module top(
  input LIOB33_SING_X0Y50_IOB_X0Y50_IPAD,
  input LIOB33_X0Y51_IOB_X0Y51_IPAD,
  input LIOB33_X0Y51_IOB_X0Y52_IPAD,
  input LIOB33_X0Y53_IOB_X0Y53_IPAD,
  input LIOB33_X0Y53_IOB_X0Y54_IPAD,
  input LIOB33_X0Y55_IOB_X0Y55_IPAD,
  input LIOB33_X0Y55_IOB_X0Y56_IPAD,
  input LIOB33_X0Y57_IOB_X0Y57_IPAD,
  input LIOB33_X0Y57_IOB_X0Y58_IPAD,
  input LIOB33_X0Y59_IOB_X0Y59_IPAD,
  input LIOB33_X0Y59_IOB_X0Y60_IPAD,
  input LIOB33_X0Y61_IOB_X0Y61_IPAD,
  input LIOB33_X0Y61_IOB_X0Y62_IPAD,
  input LIOB33_X0Y63_IOB_X0Y63_IPAD,
  input LIOB33_X0Y63_IOB_X0Y64_IPAD,
  input LIOB33_X0Y65_IOB_X0Y65_IPAD,
  input LIOB33_X0Y65_IOB_X0Y66_IPAD,
  input LIOB33_X0Y67_IOB_X0Y67_IPAD,
  input LIOB33_X0Y67_IOB_X0Y68_IPAD,
  input LIOB33_X0Y69_IOB_X0Y69_IPAD,
  input LIOB33_X0Y69_IOB_X0Y70_IPAD,
  input LIOB33_X0Y71_IOB_X0Y71_IPAD,
  input LIOB33_X0Y71_IOB_X0Y72_IPAD,
  input LIOB33_X0Y73_IOB_X0Y73_IPAD,
  input LIOB33_X0Y73_IOB_X0Y74_IPAD,
  input LIOB33_X0Y75_IOB_X0Y75_IPAD,
  input LIOB33_X0Y75_IOB_X0Y76_IPAD,
  input LIOB33_X0Y77_IOB_X0Y77_IPAD,
  input LIOB33_X0Y77_IOB_X0Y78_IPAD,
  input LIOB33_X0Y79_IOB_X0Y79_IPAD,
  input RIOB33_SING_X105Y100_IOB_X1Y100_IPAD,
  input RIOB33_SING_X105Y149_IOB_X1Y149_IPAD,
  input RIOB33_X105Y101_IOB_X1Y101_IPAD,
  input RIOB33_X105Y101_IOB_X1Y102_IPAD,
  input RIOB33_X105Y103_IOB_X1Y103_IPAD,
  input RIOB33_X105Y103_IOB_X1Y104_IPAD,
  input RIOB33_X105Y105_IOB_X1Y105_IPAD,
  input RIOB33_X105Y105_IOB_X1Y106_IPAD,
  input RIOB33_X105Y107_IOB_X1Y107_IPAD,
  input RIOB33_X105Y107_IOB_X1Y108_IPAD,
  input RIOB33_X105Y109_IOB_X1Y109_IPAD,
  input RIOB33_X105Y109_IOB_X1Y110_IPAD,
  input RIOB33_X105Y111_IOB_X1Y111_IPAD,
  input RIOB33_X105Y111_IOB_X1Y112_IPAD,
  input RIOB33_X105Y113_IOB_X1Y113_IPAD,
  input RIOB33_X105Y113_IOB_X1Y114_IPAD,
  input RIOB33_X105Y115_IOB_X1Y115_IPAD,
  input RIOB33_X105Y115_IOB_X1Y116_IPAD,
  input RIOB33_X105Y117_IOB_X1Y117_IPAD,
  input RIOB33_X105Y117_IOB_X1Y118_IPAD,
  input RIOB33_X105Y119_IOB_X1Y119_IPAD,
  input RIOB33_X105Y119_IOB_X1Y120_IPAD,
  input RIOB33_X105Y121_IOB_X1Y121_IPAD,
  input RIOB33_X105Y121_IOB_X1Y122_IPAD,
  input RIOB33_X105Y123_IOB_X1Y123_IPAD,
  input RIOB33_X105Y123_IOB_X1Y124_IPAD,
  input RIOB33_X105Y125_IOB_X1Y125_IPAD,
  input RIOB33_X105Y125_IOB_X1Y126_IPAD,
  input RIOB33_X105Y127_IOB_X1Y127_IPAD,
  input RIOB33_X105Y127_IOB_X1Y128_IPAD,
  input RIOB33_X105Y129_IOB_X1Y129_IPAD,
  input RIOB33_X105Y129_IOB_X1Y130_IPAD,
  input RIOB33_X105Y131_IOB_X1Y131_IPAD,
  input RIOB33_X105Y131_IOB_X1Y132_IPAD,
  input RIOB33_X105Y133_IOB_X1Y133_IPAD,
  input RIOB33_X105Y133_IOB_X1Y134_IPAD,
  input RIOB33_X105Y135_IOB_X1Y135_IPAD,
  input RIOB33_X105Y135_IOB_X1Y136_IPAD,
  input RIOB33_X105Y137_IOB_X1Y137_IPAD,
  input RIOB33_X105Y137_IOB_X1Y138_IPAD,
  input RIOB33_X105Y139_IOB_X1Y139_IPAD,
  input RIOB33_X105Y139_IOB_X1Y140_IPAD,
  input RIOB33_X105Y141_IOB_X1Y141_IPAD,
  input RIOB33_X105Y141_IOB_X1Y142_IPAD,
  input RIOB33_X105Y143_IOB_X1Y143_IPAD,
  input RIOB33_X105Y143_IOB_X1Y144_IPAD,
  input RIOB33_X105Y145_IOB_X1Y145_IPAD,
  input RIOB33_X105Y145_IOB_X1Y146_IPAD,
  input RIOB33_X105Y147_IOB_X1Y147_IPAD,
  input RIOB33_X105Y147_IOB_X1Y148_IPAD,
  output LIOB33_SING_X0Y100_IOB_X0Y100_OPAD,
  output LIOB33_SING_X0Y149_IOB_X0Y149_OPAD,
  output LIOB33_SING_X0Y150_IOB_X0Y150_OPAD,
  output LIOB33_SING_X0Y199_IOB_X0Y199_OPAD,
  output LIOB33_X0Y101_IOB_X0Y101_OPAD,
  output LIOB33_X0Y101_IOB_X0Y102_OPAD,
  output LIOB33_X0Y103_IOB_X0Y103_OPAD,
  output LIOB33_X0Y103_IOB_X0Y104_OPAD,
  output LIOB33_X0Y105_IOB_X0Y105_OPAD,
  output LIOB33_X0Y105_IOB_X0Y106_OPAD,
  output LIOB33_X0Y107_IOB_X0Y107_OPAD,
  output LIOB33_X0Y107_IOB_X0Y108_OPAD,
  output LIOB33_X0Y109_IOB_X0Y109_OPAD,
  output LIOB33_X0Y109_IOB_X0Y110_OPAD,
  output LIOB33_X0Y111_IOB_X0Y111_OPAD,
  output LIOB33_X0Y111_IOB_X0Y112_OPAD,
  output LIOB33_X0Y113_IOB_X0Y113_OPAD,
  output LIOB33_X0Y113_IOB_X0Y114_OPAD,
  output LIOB33_X0Y115_IOB_X0Y115_OPAD,
  output LIOB33_X0Y115_IOB_X0Y116_OPAD,
  output LIOB33_X0Y117_IOB_X0Y117_OPAD,
  output LIOB33_X0Y117_IOB_X0Y118_OPAD,
  output LIOB33_X0Y119_IOB_X0Y119_OPAD,
  output LIOB33_X0Y119_IOB_X0Y120_OPAD,
  output LIOB33_X0Y121_IOB_X0Y121_OPAD,
  output LIOB33_X0Y121_IOB_X0Y122_OPAD,
  output LIOB33_X0Y123_IOB_X0Y123_OPAD,
  output LIOB33_X0Y123_IOB_X0Y124_OPAD,
  output LIOB33_X0Y125_IOB_X0Y125_OPAD,
  output LIOB33_X0Y125_IOB_X0Y126_OPAD,
  output LIOB33_X0Y127_IOB_X0Y127_OPAD,
  output LIOB33_X0Y127_IOB_X0Y128_OPAD,
  output LIOB33_X0Y129_IOB_X0Y129_OPAD,
  output LIOB33_X0Y129_IOB_X0Y130_OPAD,
  output LIOB33_X0Y131_IOB_X0Y131_OPAD,
  output LIOB33_X0Y131_IOB_X0Y132_OPAD,
  output LIOB33_X0Y133_IOB_X0Y133_OPAD,
  output LIOB33_X0Y133_IOB_X0Y134_OPAD,
  output LIOB33_X0Y135_IOB_X0Y135_OPAD,
  output LIOB33_X0Y135_IOB_X0Y136_OPAD,
  output LIOB33_X0Y137_IOB_X0Y137_OPAD,
  output LIOB33_X0Y137_IOB_X0Y138_OPAD,
  output LIOB33_X0Y139_IOB_X0Y139_OPAD,
  output LIOB33_X0Y139_IOB_X0Y140_OPAD,
  output LIOB33_X0Y141_IOB_X0Y141_OPAD,
  output LIOB33_X0Y141_IOB_X0Y142_OPAD,
  output LIOB33_X0Y143_IOB_X0Y143_OPAD,
  output LIOB33_X0Y145_IOB_X0Y145_OPAD,
  output LIOB33_X0Y145_IOB_X0Y146_OPAD,
  output LIOB33_X0Y147_IOB_X0Y147_OPAD,
  output LIOB33_X0Y147_IOB_X0Y148_OPAD,
  output LIOB33_X0Y151_IOB_X0Y151_OPAD,
  output LIOB33_X0Y151_IOB_X0Y152_OPAD,
  output LIOB33_X0Y153_IOB_X0Y153_OPAD,
  output LIOB33_X0Y153_IOB_X0Y154_OPAD,
  output LIOB33_X0Y155_IOB_X0Y155_OPAD,
  output LIOB33_X0Y155_IOB_X0Y156_OPAD,
  output LIOB33_X0Y157_IOB_X0Y157_OPAD,
  output LIOB33_X0Y157_IOB_X0Y158_OPAD,
  output LIOB33_X0Y159_IOB_X0Y159_OPAD,
  output LIOB33_X0Y159_IOB_X0Y160_OPAD,
  output LIOB33_X0Y161_IOB_X0Y161_OPAD,
  output LIOB33_X0Y161_IOB_X0Y162_OPAD,
  output LIOB33_X0Y163_IOB_X0Y163_OPAD,
  output LIOB33_X0Y163_IOB_X0Y164_OPAD,
  output LIOB33_X0Y165_IOB_X0Y165_OPAD,
  output LIOB33_X0Y165_IOB_X0Y166_OPAD,
  output LIOB33_X0Y167_IOB_X0Y167_OPAD,
  output LIOB33_X0Y167_IOB_X0Y168_OPAD,
  output LIOB33_X0Y169_IOB_X0Y169_OPAD,
  output LIOB33_X0Y169_IOB_X0Y170_OPAD,
  output LIOB33_X0Y171_IOB_X0Y171_OPAD,
  output LIOB33_X0Y171_IOB_X0Y172_OPAD,
  output LIOB33_X0Y173_IOB_X0Y173_OPAD,
  output LIOB33_X0Y173_IOB_X0Y174_OPAD,
  output LIOB33_X0Y175_IOB_X0Y175_OPAD,
  output LIOB33_X0Y175_IOB_X0Y176_OPAD,
  output LIOB33_X0Y177_IOB_X0Y177_OPAD,
  output LIOB33_X0Y177_IOB_X0Y178_OPAD,
  output LIOB33_X0Y179_IOB_X0Y179_OPAD,
  output LIOB33_X0Y179_IOB_X0Y180_OPAD,
  output LIOB33_X0Y181_IOB_X0Y181_OPAD,
  output LIOB33_X0Y181_IOB_X0Y182_OPAD,
  output LIOB33_X0Y183_IOB_X0Y183_OPAD,
  output LIOB33_X0Y183_IOB_X0Y184_OPAD,
  output LIOB33_X0Y185_IOB_X0Y185_OPAD,
  output LIOB33_X0Y185_IOB_X0Y186_OPAD,
  output LIOB33_X0Y187_IOB_X0Y187_OPAD,
  output LIOB33_X0Y187_IOB_X0Y188_OPAD,
  output LIOB33_X0Y189_IOB_X0Y189_OPAD,
  output LIOB33_X0Y189_IOB_X0Y190_OPAD,
  output LIOB33_X0Y191_IOB_X0Y191_OPAD,
  output LIOB33_X0Y191_IOB_X0Y192_OPAD,
  output LIOB33_X0Y193_IOB_X0Y193_OPAD,
  output LIOB33_X0Y193_IOB_X0Y194_OPAD,
  output LIOB33_X0Y195_IOB_X0Y195_OPAD,
  output LIOB33_X0Y195_IOB_X0Y196_OPAD,
  output LIOB33_X0Y197_IOB_X0Y197_OPAD,
  output LIOB33_X0Y197_IOB_X0Y198_OPAD,
  output LIOB33_X0Y79_IOB_X0Y80_OPAD,
  output RIOB33_SING_X105Y150_IOB_X1Y150_OPAD,
  output RIOB33_SING_X105Y199_IOB_X1Y199_OPAD,
  output RIOB33_X105Y151_IOB_X1Y151_OPAD,
  output RIOB33_X105Y151_IOB_X1Y152_OPAD,
  output RIOB33_X105Y153_IOB_X1Y153_OPAD,
  output RIOB33_X105Y153_IOB_X1Y154_OPAD,
  output RIOB33_X105Y155_IOB_X1Y155_OPAD,
  output RIOB33_X105Y155_IOB_X1Y156_OPAD,
  output RIOB33_X105Y157_IOB_X1Y157_OPAD,
  output RIOB33_X105Y157_IOB_X1Y158_OPAD,
  output RIOB33_X105Y159_IOB_X1Y159_OPAD,
  output RIOB33_X105Y159_IOB_X1Y160_OPAD,
  output RIOB33_X105Y161_IOB_X1Y161_OPAD,
  output RIOB33_X105Y161_IOB_X1Y162_OPAD,
  output RIOB33_X105Y163_IOB_X1Y163_OPAD,
  output RIOB33_X105Y163_IOB_X1Y164_OPAD,
  output RIOB33_X105Y165_IOB_X1Y165_OPAD,
  output RIOB33_X105Y165_IOB_X1Y166_OPAD,
  output RIOB33_X105Y167_IOB_X1Y167_OPAD,
  output RIOB33_X105Y167_IOB_X1Y168_OPAD,
  output RIOB33_X105Y169_IOB_X1Y169_OPAD,
  output RIOB33_X105Y169_IOB_X1Y170_OPAD,
  output RIOB33_X105Y171_IOB_X1Y171_OPAD,
  output RIOB33_X105Y171_IOB_X1Y172_OPAD,
  output RIOB33_X105Y173_IOB_X1Y173_OPAD,
  output RIOB33_X105Y173_IOB_X1Y174_OPAD,
  output RIOB33_X105Y175_IOB_X1Y175_OPAD,
  output RIOB33_X105Y175_IOB_X1Y176_OPAD,
  output RIOB33_X105Y177_IOB_X1Y177_OPAD,
  output RIOB33_X105Y177_IOB_X1Y178_OPAD,
  output RIOB33_X105Y179_IOB_X1Y179_OPAD,
  output RIOB33_X105Y179_IOB_X1Y180_OPAD,
  output RIOB33_X105Y181_IOB_X1Y181_OPAD,
  output RIOB33_X105Y181_IOB_X1Y182_OPAD,
  output RIOB33_X105Y183_IOB_X1Y183_OPAD,
  output RIOB33_X105Y183_IOB_X1Y184_OPAD,
  output RIOB33_X105Y185_IOB_X1Y185_OPAD,
  output RIOB33_X105Y185_IOB_X1Y186_OPAD,
  output RIOB33_X105Y187_IOB_X1Y187_OPAD,
  output RIOB33_X105Y187_IOB_X1Y188_OPAD,
  output RIOB33_X105Y189_IOB_X1Y189_OPAD,
  output RIOB33_X105Y189_IOB_X1Y190_OPAD,
  output RIOB33_X105Y191_IOB_X1Y191_OPAD,
  output RIOB33_X105Y191_IOB_X1Y192_OPAD,
  output RIOB33_X105Y193_IOB_X1Y193_OPAD,
  output RIOB33_X105Y193_IOB_X1Y194_OPAD,
  output RIOB33_X105Y195_IOB_X1Y195_OPAD,
  output RIOB33_X105Y195_IOB_X1Y196_OPAD,
  output RIOB33_X105Y197_IOB_X1Y197_OPAD,
  output RIOB33_X105Y197_IOB_X1Y198_OPAD
  );
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_A;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_A1;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_A2;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_A3;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_A4;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_A5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_A6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_AO5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_AO6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_A_CY;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_A_XOR;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_B;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_B1;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_B2;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_B3;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_B4;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_B5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_B6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_BO5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_BO6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_B_CY;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_B_XOR;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_C;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_C1;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_C2;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_C3;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_C4;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_C5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_C6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_CO5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_CO6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_C_CY;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_C_XOR;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_D;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_D1;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_D2;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_D3;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_D4;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_D5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_D6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_DO5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_DO6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_D_CY;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_D_XOR;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_A;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_A1;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_A2;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_A3;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_A4;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_A5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_A6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_AO5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_AO6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_A_CY;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_A_XOR;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_B;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_B1;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_B2;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_B3;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_B4;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_B5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_B6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_BO5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_BO6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_B_CY;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_B_XOR;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_C;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_C1;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_C2;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_C3;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_C4;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_C5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_C6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_CO5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_CO6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_C_CY;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_C_XOR;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_D;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_D1;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_D2;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_D3;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_D4;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_D5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_D6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_DO5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_DO6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_D_CY;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_D_XOR;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_A;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_A1;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_A2;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_A3;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_A4;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_A5;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_A6;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_AMUX;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_AO5;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_AO6;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_A_CY;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_A_XOR;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_B;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_B1;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_B2;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_B3;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_B4;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_B5;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_B6;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_BO5;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_BO6;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_B_CY;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_B_XOR;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_C;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_C1;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_C2;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_C3;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_C4;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_C5;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_C6;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_CO5;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_CO6;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_C_CY;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_C_XOR;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_D;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_D1;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_D2;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_D3;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_D4;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_D5;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_D6;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_DO5;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_DO6;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_D_CY;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_D_XOR;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_A;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_A1;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_A2;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_A3;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_A4;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_A5;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_A6;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_AO5;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_AO6;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_A_CY;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_A_XOR;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_B;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_B1;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_B2;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_B3;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_B4;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_B5;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_B6;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_BO5;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_BO6;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_B_CY;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_B_XOR;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_C;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_C1;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_C2;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_C3;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_C4;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_C5;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_C6;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_CO5;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_CO6;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_C_CY;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_C_XOR;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_D;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_D1;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_D2;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_D3;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_D4;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_D5;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_D6;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_DO5;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_DO6;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_D_CY;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_D_XOR;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_A;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_A1;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_A2;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_A3;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_A4;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_A5;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_A6;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_AMUX;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_AO5;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_AO6;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_A_CY;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_A_XOR;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_B;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_B1;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_B2;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_B3;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_B4;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_B5;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_B6;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_BMUX;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_BO5;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_BO6;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_B_CY;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_B_XOR;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_C;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_C1;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_C2;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_C3;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_C4;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_C5;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_C6;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_CMUX;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_CO5;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_CO6;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_C_CY;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_C_XOR;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_D;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_D1;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_D2;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_D3;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_D4;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_D5;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_D6;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_DO5;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_DO6;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_D_CY;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_D_XOR;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_A;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_A1;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_A2;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_A3;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_A4;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_A5;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_A6;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_AO5;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_AO6;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_A_CY;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_A_XOR;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_B;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_B1;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_B2;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_B3;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_B4;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_B5;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_B6;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_BO5;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_BO6;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_B_CY;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_B_XOR;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_C;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_C1;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_C2;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_C3;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_C4;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_C5;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_C6;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_CO5;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_CO6;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_C_CY;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_C_XOR;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_D;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_D1;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_D2;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_D3;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_D4;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_D5;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_D6;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_DO5;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_DO6;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_D_CY;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_D_XOR;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_A;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_A1;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_A2;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_A3;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_A4;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_A5;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_A6;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_AO5;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_AO6;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_A_CY;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_A_XOR;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_B;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_B1;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_B2;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_B3;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_B4;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_B5;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_B6;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_BO5;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_BO6;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_B_CY;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_B_XOR;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_C;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_C1;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_C2;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_C3;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_C4;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_C5;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_C6;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_CO5;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_CO6;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_C_CY;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_C_XOR;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_D;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_D1;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_D2;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_D3;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_D4;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_D5;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_D6;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_DO5;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_DO6;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_D_CY;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_D_XOR;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_A;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_A1;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_A2;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_A3;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_A4;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_A5;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_A6;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_AMUX;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_AO5;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_AO6;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_A_CY;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_A_XOR;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_B;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_B1;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_B2;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_B3;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_B4;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_B5;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_B6;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_BO5;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_BO6;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_B_CY;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_B_XOR;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_C;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_C1;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_C2;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_C3;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_C4;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_C5;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_C6;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_CO5;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_CO6;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_C_CY;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_C_XOR;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_D;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_D1;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_D2;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_D3;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_D4;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_D5;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_D6;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_DO5;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_DO6;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_D_CY;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_D_XOR;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_A;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_A1;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_A2;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_A3;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_A4;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_A5;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_A6;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_AMUX;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_AO5;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_AO6;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_A_CY;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_A_XOR;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_B;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_B1;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_B2;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_B3;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_B4;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_B5;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_B6;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_BO5;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_BO6;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_B_CY;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_B_XOR;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_C;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_C1;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_C2;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_C3;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_C4;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_C5;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_C6;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_CO5;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_CO6;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_C_CY;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_C_XOR;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_D;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_D1;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_D2;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_D3;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_D4;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_D5;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_D6;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_DO5;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_DO6;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_D_CY;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_D_XOR;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_A;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_A1;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_A2;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_A3;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_A4;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_A5;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_A6;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_AMUX;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_AO5;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_AO6;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_A_CY;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_A_XOR;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_B;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_B1;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_B2;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_B3;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_B4;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_B5;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_B6;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_BMUX;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_BO5;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_BO6;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_B_CY;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_B_XOR;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_C;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_C1;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_C2;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_C3;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_C4;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_C5;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_C6;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_CO5;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_CO6;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_C_CY;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_C_XOR;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_D;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_D1;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_D2;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_D3;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_D4;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_D5;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_D6;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_DO5;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_DO6;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_D_CY;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_D_XOR;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_A;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_A1;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_A2;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_A3;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_A4;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_A5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_A6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_AO5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_AO6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_A_CY;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_A_XOR;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_B;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_B1;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_B2;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_B3;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_B4;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_B5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_B6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_BO5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_BO6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_B_CY;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_B_XOR;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_C;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_C1;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_C2;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_C3;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_C4;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_C5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_C6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_CO5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_CO6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_C_CY;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_C_XOR;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_D;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_D1;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_D2;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_D3;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_D4;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_D5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_D6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_DO5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_DO6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_D_CY;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_D_XOR;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_A;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_A1;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_A2;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_A3;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_A4;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_A5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_A6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_AO5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_AO6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_AQ;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_A_CY;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_A_XOR;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_B;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_B1;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_B2;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_B3;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_B4;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_B5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_B6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_BO5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_BO6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_B_CY;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_B_XOR;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_C;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_C1;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_C2;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_C3;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_C4;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_C5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_C6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_CLK;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_CO5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_CO6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_C_CY;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_C_XOR;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_D;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_D1;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_D2;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_D3;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_D4;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_D5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_D6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_DO5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_DO6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_D_CY;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_D_XOR;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_A;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_A1;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_A2;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_A3;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_A4;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_A5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_A6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_AO5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_AO6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_AQ;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_A_CY;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_A_XOR;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_B;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_B1;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_B2;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_B3;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_B4;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_B5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_B6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_BMUX;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_BO5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_BO6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_B_CY;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_B_XOR;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_C;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_C1;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_C2;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_C3;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_C4;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_C5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_C6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_CLK;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_CO5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_CO6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_C_CY;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_C_XOR;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_D;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_D1;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_D2;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_D3;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_D4;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_D5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_D6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_DO5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_DO6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_D_CY;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_D_XOR;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_A;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_A1;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_A2;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_A3;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_A4;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_A5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_A5Q;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_A6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_AMUX;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_AO5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_AO6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_AQ;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_AX;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_A_CY;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_A_XOR;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_B;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_B1;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_B2;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_B3;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_B4;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_B5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_B6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_BO5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_BO6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_B_CY;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_B_XOR;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_C;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_C1;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_C2;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_C3;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_C4;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_C5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_C6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_CLK;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_CO5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_CO6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_C_CY;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_C_XOR;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_D;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_D1;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_D2;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_D3;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_D4;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_D5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_D6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_DO5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_DO6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_D_CY;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_D_XOR;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_A;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_A1;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_A2;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_A3;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_A4;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_A5;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_A6;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_AO5;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_AO6;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_AQ;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_A_CY;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_A_XOR;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_B;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_B1;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_B2;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_B3;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_B4;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_B5;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_B5Q;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_B6;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_BMUX;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_BO5;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_BO6;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_BQ;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_B_CY;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_B_XOR;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_C;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_C1;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_C2;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_C3;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_C4;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_C5;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_C6;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_CLK;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_CO5;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_CO6;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_C_CY;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_C_XOR;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_D;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_D1;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_D2;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_D3;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_D4;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_D5;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_D6;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_DO5;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_DO6;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_D_CY;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_D_XOR;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_A;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_A1;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_A2;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_A3;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_A4;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_A5;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_A5Q;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_A6;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_AMUX;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_AO5;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_AO6;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_AQ;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_AX;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_A_CY;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_A_XOR;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_B;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_B1;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_B2;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_B3;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_B4;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_B5;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_B6;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_BO5;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_BO6;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_BQ;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_B_CY;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_B_XOR;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_C;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_C1;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_C2;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_C3;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_C4;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_C5;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_C6;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_CLK;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_CO5;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_CO6;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_CQ;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_C_CY;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_C_XOR;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_D;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_D1;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_D2;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_D3;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_D4;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_D5;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_D6;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_DMUX;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_DO5;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_DO6;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_D_CY;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_D_XOR;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_A;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_A1;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_A2;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_A3;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_A4;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_A5;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_A5Q;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_A6;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_AMUX;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_AO5;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_AO6;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_AQ;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_AX;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_A_CY;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_A_XOR;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_B;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_B1;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_B2;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_B3;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_B4;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_B5;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_B6;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_BO5;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_BO6;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_BQ;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_B_CY;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_B_XOR;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_C;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_C1;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_C2;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_C3;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_C4;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_C5;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_C6;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_CLK;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_CO5;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_CO6;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_CQ;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_C_CY;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_C_XOR;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_D;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_D1;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_D2;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_D3;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_D4;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_D5;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_D6;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_DMUX;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_DO5;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_DO6;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_D_CY;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_D_XOR;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_A;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_A1;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_A2;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_A3;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_A4;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_A5;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_A6;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_AO5;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_AO6;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_AQ;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_A_CY;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_A_XOR;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_B;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_B1;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_B2;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_B3;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_B4;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_B5;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_B6;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_BO5;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_BO6;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_BQ;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_B_CY;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_B_XOR;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_C;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_C1;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_C2;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_C3;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_C4;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_C5;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_C5Q;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_C6;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_CLK;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_CMUX;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_CO5;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_CO6;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_CQ;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_C_CY;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_C_XOR;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_D;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_D1;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_D2;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_D3;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_D4;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_D5;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_D5Q;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_D6;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_DMUX;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_DO5;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_DO6;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_DQ;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_D_CY;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_D_XOR;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_A;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_A1;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_A2;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_A3;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_A4;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_A5;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_A6;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_AMUX;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_AO5;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_AO6;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_AQ;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_A_CY;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_A_XOR;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_B;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_B1;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_B2;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_B3;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_B4;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_B5;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_B6;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_BO5;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_BO6;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_BQ;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_B_CY;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_B_XOR;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_C;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_C1;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_C2;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_C3;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_C4;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_C5;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_C6;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_CLK;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_CO5;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_CO6;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_CQ;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_C_CY;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_C_XOR;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_D;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_D1;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_D2;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_D3;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_D4;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_D5;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_D5Q;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_D6;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_DMUX;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_DO5;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_DO6;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_DQ;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_D_CY;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_D_XOR;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_A;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_A1;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_A2;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_A3;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_A4;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_A5;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_A5Q;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_A6;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_AMUX;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_AO5;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_AO6;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_AQ;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_AX;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_A_CY;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_A_XOR;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_B;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_B1;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_B2;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_B3;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_B4;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_B5;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_B6;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_BO5;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_BO6;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_BQ;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_B_CY;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_B_XOR;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_C;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_C1;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_C2;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_C3;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_C4;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_C5;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_C6;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_CLK;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_CO5;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_CO6;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_CQ;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_C_CY;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_C_XOR;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_D;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_D1;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_D2;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_D3;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_D4;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_D5;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_D6;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_DMUX;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_DO5;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_DO6;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_D_CY;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_D_XOR;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_A;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_A1;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_A2;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_A3;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_A4;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_A5;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_A5Q;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_A6;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_AMUX;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_AO5;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_AO6;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_AQ;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_A_CY;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_A_XOR;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_B;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_B1;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_B2;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_B3;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_B4;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_B5;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_B6;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_BO5;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_BO6;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_BQ;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_B_CY;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_B_XOR;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_C;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_C1;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_C2;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_C3;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_C4;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_C5;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_C6;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_CLK;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_CO5;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_CO6;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_CQ;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_C_CY;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_C_XOR;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_D;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_D1;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_D2;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_D3;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_D4;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_D5;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_D5Q;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_D6;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_DMUX;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_DO5;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_DO6;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_DQ;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_D_CY;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_D_XOR;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_A;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_A1;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_A2;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_A3;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_A4;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_A5;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_A6;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_AMUX;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_AO5;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_AO6;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_A_CY;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_A_XOR;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_B;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_B1;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_B2;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_B3;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_B4;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_B5;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_B6;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_BO5;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_BO6;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_BQ;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_B_CY;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_B_XOR;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_C;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_C1;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_C2;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_C3;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_C4;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_C5;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_C6;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_CLK;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_CO5;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_CO6;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_C_CY;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_C_XOR;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_D;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_D1;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_D2;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_D3;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_D4;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_D5;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_D6;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_DO5;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_DO6;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_D_CY;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_D_XOR;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_SR;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_A;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_A1;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_A2;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_A3;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_A4;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_A5;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_A6;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_AO5;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_AO6;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_AQ;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_A_CY;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_A_XOR;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_B;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_B1;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_B2;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_B3;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_B4;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_B5;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_B6;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_BO5;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_BO6;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_BQ;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_B_CY;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_B_XOR;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_C;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_C1;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_C2;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_C3;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_C4;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_C5;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_C6;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_CLK;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_CO5;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_CO6;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_C_CY;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_C_XOR;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_D;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_D1;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_D2;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_D3;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_D4;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_D5;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_D6;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_DO5;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_DO6;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_D_CY;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_D_XOR;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_SR;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_A;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_A1;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_A2;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_A3;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_A4;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_A5;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_A5Q;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_A6;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_AMUX;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_AO5;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_AO6;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_AQ;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_A_CY;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_A_XOR;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_B;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_B1;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_B2;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_B3;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_B4;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_B5;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_B5Q;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_B6;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_BMUX;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_BO5;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_BO6;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_BQ;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_BX;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_B_CY;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_B_XOR;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_C;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_C1;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_C2;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_C3;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_C4;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_C5;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_C6;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_CLK;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_CMUX;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_CO5;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_CO6;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_C_CY;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_C_XOR;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_D;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_D1;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_D2;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_D3;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_D4;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_D5;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_D6;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_DMUX;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_DO5;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_DO6;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_D_CY;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_D_XOR;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_A;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_A1;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_A2;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_A3;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_A4;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_A5;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_A6;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_AO5;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_AO6;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_AQ;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_A_CY;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_A_XOR;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_B;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_B1;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_B2;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_B3;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_B4;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_B5;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_B6;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_BO5;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_BO6;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_B_CY;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_B_XOR;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_C;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_C1;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_C2;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_C3;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_C4;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_C5;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_C6;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_CLK;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_CO5;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_CO6;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_C_CY;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_C_XOR;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_D;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_D1;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_D2;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_D3;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_D4;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_D5;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_D6;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_DO5;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_DO6;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_D_CY;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_D_XOR;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_A;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_A1;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_A2;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_A3;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_A4;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_A5;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_A6;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_AO5;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_AO6;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_AQ;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_A_CY;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_A_XOR;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_B;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_B1;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_B2;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_B3;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_B4;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_B5;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_B6;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_BO5;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_BO6;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_BQ;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_B_CY;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_B_XOR;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_C;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_C1;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_C2;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_C3;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_C4;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_C5;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_C6;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_CLK;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_CO5;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_CO6;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_C_CY;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_C_XOR;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_D;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_D1;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_D2;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_D3;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_D4;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_D5;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_D6;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_DO5;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_DO6;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_D_CY;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_D_XOR;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_A;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_A1;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_A2;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_A3;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_A4;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_A5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_A6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_AO5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_AO6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_A_CY;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_A_XOR;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_B;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_B1;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_B2;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_B3;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_B4;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_B5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_B6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_BO5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_BO6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_B_CY;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_B_XOR;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_C;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_C1;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_C2;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_C3;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_C4;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_C5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_C6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_CMUX;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_CO5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_CO6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_C_CY;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_C_XOR;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_D;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_D1;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_D2;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_D3;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_D4;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_D5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_D6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_DO5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_DO6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_D_CY;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_D_XOR;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_A;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_A1;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_A2;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_A3;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_A4;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_A5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_A6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_AO5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_AO6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_A_CY;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_A_XOR;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_B;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_B1;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_B2;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_B3;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_B4;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_B5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_B6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_BO5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_BO6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_B_CY;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_B_XOR;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_C;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_C1;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_C2;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_C3;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_C4;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_C5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_C6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_CO5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_CO6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_C_CY;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_C_XOR;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_D;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_D1;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_D2;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_D3;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_D4;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_D5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_D6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_DMUX;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_DO5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_DO6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_D_CY;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_D_XOR;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_A;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_A1;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_A2;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_A3;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_A4;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_A5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_A6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_AO5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_AO6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_A_CY;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_A_XOR;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_B;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_B1;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_B2;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_B3;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_B4;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_B5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_B6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_BO5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_BO6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_B_CY;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_B_XOR;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_C;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_C1;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_C2;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_C3;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_C4;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_C5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_C6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_CO5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_CO6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_C_CY;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_C_XOR;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_D;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_D1;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_D2;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_D3;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_D4;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_D5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_D6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_DO5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_DO6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_D_CY;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_D_XOR;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_A;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_A1;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_A2;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_A3;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_A4;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_A5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_A6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_AO5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_AO6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_A_CY;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_A_XOR;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_B;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_B1;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_B2;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_B3;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_B4;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_B5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_B6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_BO5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_BO6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_B_CY;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_B_XOR;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_C;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_C1;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_C2;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_C3;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_C4;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_C5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_C6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_CO5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_CO6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_C_CY;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_C_XOR;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_D;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_D1;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_D2;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_D3;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_D4;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_D5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_D6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_DO5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_DO6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_D_CY;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_D_XOR;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_A;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_A1;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_A2;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_A3;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_A4;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_A5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_A6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_AO5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_AO6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_A_CY;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_A_XOR;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_B;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_B1;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_B2;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_B3;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_B4;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_B5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_B6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_BO5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_BO6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_B_CY;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_B_XOR;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_C;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_C1;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_C2;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_C3;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_C4;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_C5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_C6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_CO5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_CO6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_C_CY;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_C_XOR;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_D;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_D1;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_D2;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_D3;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_D4;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_D5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_D6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_DO5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_DO6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_D_CY;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_D_XOR;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_A;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_A1;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_A2;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_A3;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_A4;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_A5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_A6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_AO5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_AO6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_A_CY;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_A_XOR;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_B;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_B1;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_B2;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_B3;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_B4;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_B5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_B6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_BO5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_BO6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_B_CY;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_B_XOR;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_C;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_C1;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_C2;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_C3;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_C4;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_C5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_C6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_CO5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_CO6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_C_CY;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_C_XOR;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_D;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_D1;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_D2;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_D3;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_D4;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_D5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_D6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_DO5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_DO6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_D_CY;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_D_XOR;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_A;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_A1;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_A2;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_A3;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_A4;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_A5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_A6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_AMUX;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_AO5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_AO6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_A_CY;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_A_XOR;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_B;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_B1;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_B2;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_B3;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_B4;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_B5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_B6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_BMUX;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_BO5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_BO6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_B_CY;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_B_XOR;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_C;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_C1;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_C2;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_C3;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_C4;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_C5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_C6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_CO5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_CO6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_C_CY;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_C_XOR;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_D;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_D1;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_D2;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_D3;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_D4;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_D5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_D6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_DO5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_DO6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_D_CY;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_D_XOR;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_A;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_A1;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_A2;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_A3;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_A4;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_A5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_A6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_AMUX;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_AO5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_AO6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_A_CY;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_A_XOR;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_B;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_B1;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_B2;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_B3;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_B4;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_B5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_B6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_BMUX;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_BO5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_BO6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_B_CY;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_B_XOR;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_C;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_C1;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_C2;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_C3;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_C4;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_C5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_C6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_CMUX;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_CO5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_CO6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_C_CY;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_C_XOR;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_D;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_D1;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_D2;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_D3;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_D4;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_D5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_D6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_DO5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_DO6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_D_CY;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_D_XOR;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_A;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_A1;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_A2;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_A3;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_A4;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_A5;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_A6;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_AO5;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_AO6;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_A_CY;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_A_XOR;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_B;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_B1;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_B2;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_B3;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_B4;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_B5;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_B6;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_BO5;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_BO6;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_B_CY;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_B_XOR;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_C;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_C1;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_C2;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_C3;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_C4;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_C5;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_C6;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_CO5;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_CO6;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_C_CY;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_C_XOR;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_D;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_D1;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_D2;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_D3;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_D4;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_D5;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_D6;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_DO5;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_DO6;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_D_CY;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_D_XOR;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_A;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_A1;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_A2;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_A3;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_A4;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_A5;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_A6;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_AO5;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_AO6;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_A_CY;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_A_XOR;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_B;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_B1;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_B2;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_B3;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_B4;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_B5;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_B6;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_BO5;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_BO6;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_B_CY;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_B_XOR;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_C;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_C1;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_C2;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_C3;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_C4;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_C5;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_C6;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_CO5;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_CO6;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_C_CY;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_C_XOR;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_D;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_D1;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_D2;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_D3;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_D4;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_D5;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_D6;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_DO5;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_DO6;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_D_CY;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_D_XOR;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A1;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A2;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A3;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A4;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_AO5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_AO6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A_CY;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A_XOR;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B1;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B2;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B3;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B4;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_BO5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_BO6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B_CY;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B_XOR;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C1;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C2;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C3;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C4;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_CO5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_CO6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C_CY;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C_XOR;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D1;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D2;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D3;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D4;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_DO5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_DO6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D_CY;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D_XOR;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A1;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A2;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A3;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A4;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_AO5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_AO6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A_CY;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A_XOR;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B1;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B2;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B3;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B4;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_BO5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_BO6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B_CY;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B_XOR;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C1;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C2;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C3;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C4;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_CO5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_CO6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C_CY;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C_XOR;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D1;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D2;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D3;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D4;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_DO5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_DO6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D_CY;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D_XOR;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_A;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_A1;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_A2;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_A3;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_A4;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_A5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_A6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_AO5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_AO6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_AQ;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_A_CY;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_A_XOR;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_B;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_B1;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_B2;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_B3;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_B4;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_B5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_B6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_BMUX;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_BO5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_BO6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_B_CY;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_B_XOR;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_C;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_C1;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_C2;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_C3;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_C4;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_C5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_C6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_CLK;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_CO5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_CO6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_C_CY;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_C_XOR;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_D;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_D1;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_D2;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_D3;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_D4;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_D5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_D6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_DO5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_DO6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_D_CY;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_D_XOR;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_A;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_A1;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_A2;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_A3;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_A4;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_A5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_A6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_AMUX;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_AO5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_AO6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_A_CY;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_A_XOR;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_B;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_B1;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_B2;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_B3;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_B4;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_B5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_B6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_BO5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_BO6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_B_CY;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_B_XOR;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_C;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_C1;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_C2;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_C3;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_C4;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_C5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_C6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_CO5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_CO6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_C_CY;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_C_XOR;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_D;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_D1;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_D2;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_D3;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_D4;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_D5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_D6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_DO5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_DO6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_D_CY;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_D_XOR;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_A;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_A1;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_A2;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_A3;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_A4;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_A5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_A6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_AMUX;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_AO5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_AO6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_A_CY;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_A_XOR;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_B;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_B1;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_B2;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_B3;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_B4;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_B5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_B6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_BO5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_BO6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_BQ;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_B_CY;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_B_XOR;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_C;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_C1;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_C2;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_C3;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_C4;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_C5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_C6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_CLK;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_CMUX;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_CO5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_CO6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_C_CY;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_C_XOR;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_D;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_D1;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_D2;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_D3;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_D4;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_D5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_D6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_DO5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_DO6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_D_CY;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_D_XOR;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_A;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_A1;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_A2;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_A3;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_A4;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_A5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_A6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_AO5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_AO6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_AQ;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_A_CY;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_A_XOR;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_B;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_B1;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_B2;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_B3;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_B4;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_B5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_B6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_BO5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_BO6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_BQ;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_B_CY;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_B_XOR;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_C;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_C1;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_C2;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_C3;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_C4;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_C5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_C6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_CLK;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_CO5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_CO6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_CQ;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_C_CY;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_C_XOR;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_D;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_D1;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_D2;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_D3;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_D4;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_D5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_D6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_DO5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_DO6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_D_CY;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_D_XOR;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_A;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_A1;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_A2;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_A3;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_A4;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_A5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_A6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_AO5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_AO6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_A_CY;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_A_XOR;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_B;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_B1;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_B2;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_B3;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_B4;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_B5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_B6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_BO5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_BO6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_B_CY;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_B_XOR;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_C;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_C1;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_C2;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_C3;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_C4;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_C5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_C6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_CMUX;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_CO5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_CO6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_C_CY;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_C_XOR;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_D;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_D1;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_D2;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_D3;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_D4;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_D5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_D6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_DO5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_DO6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_D_CY;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_D_XOR;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_A;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_A1;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_A2;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_A3;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_A4;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_A5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_A6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_AO5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_AO6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_A_CY;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_A_XOR;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_B;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_B1;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_B2;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_B3;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_B4;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_B5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_B6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_BO5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_BO6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_B_CY;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_B_XOR;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_C;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_C1;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_C2;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_C3;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_C4;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_C5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_C6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_CO5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_CO6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_C_CY;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_C_XOR;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_D;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_D1;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_D2;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_D3;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_D4;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_D5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_D6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_DO5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_DO6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_D_CY;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_D_XOR;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_A;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_A1;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_A2;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_A3;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_A4;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_A5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_A6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_AO5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_AO6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_AQ;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_A_CY;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_A_XOR;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_B;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_B1;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_B2;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_B3;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_B4;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_B5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_B6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_BO5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_BO6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_BQ;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_B_CY;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_B_XOR;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_C;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_C1;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_C2;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_C3;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_C4;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_C5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_C6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_CLK;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_CO5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_CO6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_CQ;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_C_CY;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_C_XOR;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_D;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_D1;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_D2;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_D3;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_D4;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_D5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_D6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_DMUX;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_DO5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_DO6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_D_CY;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_D_XOR;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_A;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_A1;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_A2;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_A3;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_A4;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_A5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_A6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_AO5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_AO6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_AQ;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_A_CY;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_A_XOR;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_B;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_B1;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_B2;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_B3;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_B4;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_B5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_B6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_BO5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_BO6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_BQ;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_B_CY;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_B_XOR;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_C;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_C1;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_C2;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_C3;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_C4;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_C5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_C6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_CLK;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_CO5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_CO6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_C_CY;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_C_XOR;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_D;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_D1;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_D2;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_D3;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_D4;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_D5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_D6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_DO5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_DO6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_D_CY;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_D_XOR;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_A;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_A1;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_A2;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_A3;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_A4;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_A5;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_A6;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_AO5;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_AO6;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_AQ;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_A_CY;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_A_XOR;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_B;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_B1;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_B2;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_B3;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_B4;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_B5;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_B6;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_BO5;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_BO6;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_BQ;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_B_CY;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_B_XOR;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_C;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_C1;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_C2;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_C3;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_C4;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_C5;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_C6;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_CLK;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_CO5;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_CO6;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_CQ;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_C_CY;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_C_XOR;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_D;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_D1;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_D2;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_D3;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_D4;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_D5;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_D6;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_DO5;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_DO6;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_DQ;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_D_CY;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_D_XOR;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_A;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_A1;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_A2;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_A3;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_A4;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_A5;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_A5Q;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_A6;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_AMUX;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_AO5;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_AO6;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_AQ;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_AX;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_A_CY;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_A_XOR;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_B;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_B1;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_B2;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_B3;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_B4;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_B5;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_B5Q;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_B6;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_BMUX;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_BO5;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_BO6;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_BQ;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_B_CY;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_B_XOR;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_C;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_C1;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_C2;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_C3;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_C4;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_C5;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_C6;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_CLK;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_CMUX;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_CO5;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_CO6;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_C_CY;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_C_XOR;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_D;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_D1;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_D2;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_D3;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_D4;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_D5;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_D6;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_DO5;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_DO6;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_D_CY;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_D_XOR;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_A;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_A1;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_A2;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_A3;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_A4;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_A5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_A6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_AO5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_AO6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_AQ;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_A_CY;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_A_XOR;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_B;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_B1;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_B2;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_B3;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_B4;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_B5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_B5Q;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_B6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_BMUX;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_BO5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_BO6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_BQ;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_B_CY;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_B_XOR;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_C;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_C1;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_C2;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_C3;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_C4;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_C5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_C6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_CLK;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_CO5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_CO6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_C_CY;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_C_XOR;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_D;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_D1;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_D2;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_D3;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_D4;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_D5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_D6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_DO5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_DO6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_D_CY;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_D_XOR;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_A;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_A1;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_A2;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_A3;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_A4;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_A5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_A6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_AMUX;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_AO5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_AO6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_A_CY;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_A_XOR;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_B;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_B1;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_B2;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_B3;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_B4;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_B5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_B5Q;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_B6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_BMUX;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_BO5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_BO6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_BQ;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_B_CY;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_B_XOR;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_C;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_C1;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_C2;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_C3;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_C4;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_C5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_C6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_CLK;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_CO5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_CO6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_C_CY;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_C_XOR;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_D;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_D1;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_D2;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_D3;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_D4;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_D5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_D6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_DO5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_DO6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_D_CY;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_D_XOR;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_A;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_A1;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_A2;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_A3;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_A4;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_A5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_A5Q;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_A6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_AMUX;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_AO5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_AO6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_AQ;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_AX;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_A_CY;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_A_XOR;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_B;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_B1;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_B2;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_B3;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_B4;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_B5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_B6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_BO5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_BO6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_BQ;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_B_CY;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_B_XOR;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_C;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_C1;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_C2;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_C3;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_C4;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_C5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_C6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_CLK;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_CMUX;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_CO5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_CO6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_C_CY;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_C_XOR;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_D;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_D1;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_D2;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_D3;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_D4;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_D5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_D6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_DO5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_DO6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_D_CY;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_D_XOR;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_A;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_A1;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_A2;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_A3;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_A4;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_A5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_A6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_AO5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_AO6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_A_CY;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_A_XOR;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_B;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_B1;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_B2;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_B3;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_B4;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_B5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_B6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_BO5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_BO6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_B_CY;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_B_XOR;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_C;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_C1;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_C2;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_C3;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_C4;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_C5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_C6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_CO5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_CO6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_C_CY;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_C_XOR;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_D;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_D1;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_D2;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_D3;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_D4;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_D5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_D6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_DO5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_DO6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_D_CY;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_D_XOR;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_A;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_A1;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_A2;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_A3;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_A4;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_A5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_A6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_AO5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_AO6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_AQ;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_A_CY;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_A_XOR;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_B;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_B1;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_B2;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_B3;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_B4;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_B5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_B5Q;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_B6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_BMUX;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_BO5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_BO6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_BQ;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_B_CY;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_B_XOR;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_C;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_C1;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_C2;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_C3;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_C4;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_C5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_C6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_CLK;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_CO5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_CO6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_CQ;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_C_CY;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_C_XOR;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_D;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_D1;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_D2;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_D3;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_D4;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_D5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_D6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_DO5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_DO6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_D_CY;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_D_XOR;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_A;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_A1;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_A2;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_A3;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_A4;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_A5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_A6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_AO5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_AO6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_AQ;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_A_CY;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_A_XOR;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_B;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_B1;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_B2;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_B3;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_B4;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_B5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_B6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_BO5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_BO6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_BQ;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_B_CY;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_B_XOR;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_C;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_C1;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_C2;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_C3;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_C4;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_C5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_C6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_CLK;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_CO5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_CO6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_C_CY;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_C_XOR;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_D;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_D1;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_D2;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_D3;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_D4;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_D5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_D6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_DO5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_DO6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_D_CY;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_D_XOR;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_A;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_A1;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_A2;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_A3;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_A4;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_A5;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_A5Q;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_A6;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_AMUX;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_AO5;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_AO6;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_AX;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_A_CY;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_A_XOR;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_B;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_B1;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_B2;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_B3;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_B4;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_B5;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_B6;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_BMUX;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_BO5;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_BO6;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_B_CY;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_B_XOR;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_C;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_C1;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_C2;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_C3;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_C4;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_C5;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_C6;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_CLK;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_CO5;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_CO6;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_C_CY;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_C_XOR;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_D;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_D1;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_D2;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_D3;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_D4;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_D5;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_D6;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_DO5;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_DO6;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_D_CY;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_D_XOR;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_A;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_A1;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_A2;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_A3;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_A4;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_A5;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_A6;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_AO5;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_AO6;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_AQ;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_A_CY;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_A_XOR;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_B;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_B1;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_B2;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_B3;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_B4;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_B5;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_B6;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_BO5;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_BO6;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_BQ;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_B_CY;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_B_XOR;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_C;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_C1;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_C2;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_C3;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_C4;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_C5;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_C6;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_CLK;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_CO5;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_CO6;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_CQ;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_C_CY;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_C_XOR;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_D;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_D1;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_D2;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_D3;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_D4;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_D5;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_D6;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_DO5;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_DO6;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_D_CY;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_D_XOR;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_A;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_A1;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_A2;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_A3;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_A4;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_A5;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_A6;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_AO5;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_AO6;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_AQ;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_A_CY;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_A_XOR;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_B;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_B1;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_B2;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_B3;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_B4;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_B5;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_B6;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_BO5;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_BO6;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_BQ;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_B_CY;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_B_XOR;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_C;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_C1;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_C2;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_C3;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_C4;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_C5;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_C6;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_CLK;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_CO5;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_CO6;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_C_CY;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_C_XOR;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_D;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_D1;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_D2;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_D3;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_D4;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_D5;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_D6;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_DO5;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_DO6;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_D_CY;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_D_XOR;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_A;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_A1;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_A2;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_A3;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_A4;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_A5;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_A6;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_AO5;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_AO6;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_AQ;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_A_CY;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_A_XOR;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_B;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_B1;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_B2;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_B3;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_B4;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_B5;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_B5Q;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_B6;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_BMUX;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_BO5;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_BO6;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_BQ;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_B_CY;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_B_XOR;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_C;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_C1;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_C2;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_C3;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_C4;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_C5;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_C6;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_CLK;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_CO5;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_CO6;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_CQ;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_C_CY;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_C_XOR;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_D;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_D1;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_D2;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_D3;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_D4;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_D5;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_D6;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_DO5;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_DO6;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_D_CY;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_D_XOR;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_A;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_A1;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_A2;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_A3;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_A4;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_A5;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_A5Q;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_A6;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_AMUX;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_AO5;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_AO6;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_AQ;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_AX;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_A_CY;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_A_XOR;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_B;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_B1;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_B2;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_B3;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_B4;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_B5;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_B6;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_BMUX;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_BO5;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_BO6;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_BQ;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_B_CY;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_B_XOR;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_C;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_C1;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_C2;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_C3;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_C4;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_C5;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_C6;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_CLK;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_CO5;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_CO6;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_CQ;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_C_CY;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_C_XOR;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_D;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_D1;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_D2;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_D3;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_D4;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_D5;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_D6;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_DO5;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_DO6;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_D_CY;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_D_XOR;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_A;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_A1;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_A2;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_A3;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_A4;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_A5;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_A6;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_AMUX;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_AO5;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_AO6;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_A_CY;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_A_XOR;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_B;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_B1;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_B2;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_B3;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_B4;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_B5;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_B6;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_BO5;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_BO6;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_BQ;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_B_CY;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_B_XOR;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_C;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_C1;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_C2;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_C3;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_C4;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_C5;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_C5Q;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_C6;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_CLK;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_CMUX;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_CO5;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_CO6;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_CQ;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_C_CY;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_C_XOR;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_D;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_D1;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_D2;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_D3;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_D4;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_D5;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_D6;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_DO5;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_DO6;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_DQ;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_D_CY;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_D_XOR;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_A;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_A1;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_A2;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_A3;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_A4;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_A5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_A6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_AO5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_AO6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_AQ;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_A_CY;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_A_XOR;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_B;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_B1;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_B2;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_B3;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_B4;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_B5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_B6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_BMUX;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_BO5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_BO6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_B_CY;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_B_XOR;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_C;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_C1;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_C2;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_C3;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_C4;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_C5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_C5Q;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_C6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_CLK;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_CMUX;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_CO5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_CO6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_CQ;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_C_CY;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_C_XOR;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_D;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_D1;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_D2;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_D3;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_D4;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_D5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_D6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_DO5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_DO6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_D_CY;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_D_XOR;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_A;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_A1;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_A2;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_A3;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_A4;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_A5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_A5Q;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_A6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_AMUX;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_AO5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_AO6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_AQ;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_A_CY;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_A_XOR;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_B;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_B1;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_B2;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_B3;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_B4;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_B5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_B6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_BO5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_BO6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_BQ;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_B_CY;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_B_XOR;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_C;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_C1;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_C2;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_C3;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_C4;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_C5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_C6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_CLK;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_CO5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_CO6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_CQ;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_C_CY;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_C_XOR;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_D;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_D1;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_D2;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_D3;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_D4;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_D5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_D6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_DO5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_DO6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_D_CY;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_D_XOR;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_A;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_A1;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_A2;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_A3;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_A4;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_A5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_A6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_AO5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_AO6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_AQ;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_A_CY;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_A_XOR;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_B;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_B1;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_B2;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_B3;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_B4;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_B5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_B6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_BO5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_BO6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_BQ;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_B_CY;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_B_XOR;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_C;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_C1;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_C2;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_C3;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_C4;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_C5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_C6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_CLK;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_CO5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_CO6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_CQ;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_C_CY;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_C_XOR;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_D;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_D1;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_D2;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_D3;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_D4;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_D5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_D6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_DO5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_DO6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_DQ;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_D_CY;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_D_XOR;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_A;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_A1;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_A2;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_A3;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_A4;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_A5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_A6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_AO5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_AO6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_AQ;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_A_CY;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_A_XOR;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_B;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_B1;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_B2;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_B3;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_B4;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_B5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_B6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_BO5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_BO6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_BQ;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_B_CY;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_B_XOR;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_C;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_C1;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_C2;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_C3;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_C4;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_C5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_C6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_CLK;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_CO5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_CO6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_CQ;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_C_CY;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_C_XOR;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_D;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_D1;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_D2;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_D3;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_D4;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_D5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_D6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_DO5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_DO6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_D_CY;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_D_XOR;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_A;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_A1;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_A2;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_A3;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_A4;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_A5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_A6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_AO5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_AO6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_AQ;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_A_CY;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_A_XOR;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_B;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_B1;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_B2;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_B3;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_B4;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_B5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_B6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_BO5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_BO6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_BQ;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_B_CY;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_B_XOR;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_C;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_C1;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_C2;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_C3;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_C4;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_C5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_C6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_CLK;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_CO5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_CO6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_CQ;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_C_CY;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_C_XOR;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_D;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_D1;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_D2;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_D3;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_D4;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_D5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_D6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_DO5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_DO6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_D_CY;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_D_XOR;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_A;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_A1;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_A2;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_A3;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_A4;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_A5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_A6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_AO5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_AO6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_AQ;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_AX;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_A_CY;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_A_XOR;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_B;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_B1;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_B2;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_B3;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_B4;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_B5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_B6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_BMUX;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_BO5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_BO6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_BQ;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_BX;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_B_CY;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_B_XOR;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_C;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_C1;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_C2;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_C3;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_C4;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_C5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_C6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_CE;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_CLK;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_CO5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_CO6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_C_CY;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_C_XOR;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_D;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_D1;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_D2;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_D3;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_D4;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_D5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_D6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_DO5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_DO6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_D_CY;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_D_XOR;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_SR;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_A;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_A1;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_A2;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_A3;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_A4;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_A5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_A6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_AMUX;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_AO5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_AO6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_AQ;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_AX;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_A_CY;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_A_XOR;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_B;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_B1;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_B2;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_B3;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_B4;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_B5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_B6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_BO5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_BO6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_B_CY;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_B_XOR;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_C;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_C1;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_C2;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_C3;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_C4;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_C5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_C6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_CLK;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_CO5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_CO6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_C_CY;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_C_XOR;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_D;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_D1;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_D2;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_D3;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_D4;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_D5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_D6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_DO5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_DO6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_D_CY;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_D_XOR;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_SR;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_A;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_A1;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_A2;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_A3;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_A4;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_A5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_A6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_AO5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_AO6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_AQ;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_A_CY;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_A_XOR;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_B;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_B1;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_B2;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_B3;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_B4;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_B5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_B6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_BO5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_BO6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_B_CY;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_B_XOR;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_C;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_C1;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_C2;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_C3;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_C4;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_C5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_C6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_CLK;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_CO5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_CO6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_C_CY;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_C_XOR;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_D;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_D1;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_D2;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_D3;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_D4;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_D5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_D6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_DO5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_DO6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_D_CY;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_D_XOR;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_A;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_A1;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_A2;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_A3;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_A4;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_A5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_A6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_AMUX;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_AO5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_AO6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_AQ;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_A_CY;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_A_XOR;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_B;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_B1;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_B2;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_B3;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_B4;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_B5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_B6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_BMUX;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_BO5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_BO6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_B_CY;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_B_XOR;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_C;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_C1;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_C2;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_C3;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_C4;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_C5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_C6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_CLK;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_CO5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_CO6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_C_CY;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_C_XOR;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_D;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_D1;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_D2;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_D3;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_D4;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_D5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_D6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_DO5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_DO6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_D_CY;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_D_XOR;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_A;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_A1;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_A2;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_A3;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_A4;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_A5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_A6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_AO5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_AO6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_AQ;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_A_CY;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_A_XOR;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_B;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_B1;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_B2;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_B3;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_B4;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_B5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_B6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_BMUX;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_BO5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_BO6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_B_CY;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_B_XOR;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_C;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_C1;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_C2;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_C3;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_C4;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_C5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_C6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_CLK;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_CO5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_CO6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_C_CY;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_C_XOR;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_D;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_D1;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_D2;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_D3;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_D4;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_D5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_D6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_DO5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_DO6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_D_CY;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_D_XOR;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_A;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_A1;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_A2;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_A3;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_A4;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_A5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_A6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_AMUX;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_AO5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_AO6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_A_CY;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_A_XOR;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_B;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_B1;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_B2;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_B3;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_B4;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_B5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_B6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_BO5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_BO6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_B_CY;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_B_XOR;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_C;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_C1;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_C2;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_C3;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_C4;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_C5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_C6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_CO5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_CO6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_C_CY;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_C_XOR;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_D;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_D1;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_D2;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_D3;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_D4;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_D5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_D6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_DO5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_DO6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_D_CY;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_D_XOR;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_A;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_A1;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_A2;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_A3;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_A4;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_A5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_A6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_AO5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_AO6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_A_CY;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_A_XOR;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_B;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_B1;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_B2;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_B3;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_B4;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_B5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_B6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_BO5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_BO6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_B_CY;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_B_XOR;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_C;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_C1;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_C2;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_C3;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_C4;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_C5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_C6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_CO5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_CO6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_C_CY;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_C_XOR;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_D;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_D1;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_D2;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_D3;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_D4;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_D5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_D6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_DO5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_DO6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_D_CY;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_D_XOR;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_A;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_A1;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_A2;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_A3;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_A4;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_A5;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_A6;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_AO5;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_AO6;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_AQ;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_A_CY;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_A_XOR;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_B;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_B1;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_B2;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_B3;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_B4;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_B5;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_B6;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_BO5;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_BO6;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_BQ;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_B_CY;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_B_XOR;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_C;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_C1;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_C2;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_C3;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_C4;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_C5;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_C6;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_CLK;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_CO5;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_CO6;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_CQ;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_C_CY;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_C_XOR;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_D;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_D1;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_D2;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_D3;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_D4;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_D5;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_D6;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_DMUX;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_DO5;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_DO6;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_D_CY;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_D_XOR;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_A;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_A1;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_A2;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_A3;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_A4;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_A5;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_A6;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_AO5;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_AO6;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_AQ;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_A_CY;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_A_XOR;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_B;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_B1;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_B2;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_B3;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_B4;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_B5;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_B6;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_BO5;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_BO6;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_B_CY;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_B_XOR;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_C;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_C1;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_C2;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_C3;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_C4;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_C5;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_C6;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_CLK;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_CO5;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_CO6;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_C_CY;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_C_XOR;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_D;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_D1;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_D2;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_D3;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_D4;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_D5;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_D6;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_DO5;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_DO6;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_D_CY;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_D_XOR;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_A;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_A1;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_A2;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_A3;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_A4;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_A5;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_A6;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_AO5;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_AO6;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_AQ;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_A_CY;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_A_XOR;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_B;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_B1;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_B2;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_B3;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_B4;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_B5;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_B6;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_BO5;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_BO6;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_BQ;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_B_CY;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_B_XOR;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_C;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_C1;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_C2;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_C3;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_C4;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_C5;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_C5Q;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_C6;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_CLK;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_CMUX;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_CO5;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_CO6;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_CQ;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_C_CY;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_C_XOR;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_D;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_D1;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_D2;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_D3;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_D4;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_D5;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_D6;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_DMUX;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_DO5;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_DO6;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_D_CY;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_D_XOR;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_A;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_A1;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_A2;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_A3;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_A4;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_A5;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_A6;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_AO5;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_AO6;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_AQ;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_A_CY;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_A_XOR;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_B;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_B1;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_B2;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_B3;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_B4;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_B5;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_B6;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_BO5;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_BO6;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_BQ;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_B_CY;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_B_XOR;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_C;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_C1;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_C2;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_C3;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_C4;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_C5;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_C6;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_CLK;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_CO5;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_CO6;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_C_CY;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_C_XOR;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_D;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_D1;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_D2;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_D3;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_D4;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_D5;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_D6;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_DO5;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_DO6;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_D_CY;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_D_XOR;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_A;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_A1;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_A2;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_A3;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_A4;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_A5;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_A6;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_AO5;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_AO6;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_AQ;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_AX;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_A_CY;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_A_XOR;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_B;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_B1;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_B2;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_B3;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_B4;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_B5;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_B6;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_BO5;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_BO6;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_B_CY;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_B_XOR;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_C;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_C1;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_C2;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_C3;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_C4;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_C5;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_C6;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_CE;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_CLK;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_CO5;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_CO6;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_C_CY;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_C_XOR;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_D;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_D1;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_D2;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_D3;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_D4;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_D5;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_D6;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_DO5;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_DO6;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_D_CY;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_D_XOR;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_SR;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_A;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_A1;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_A2;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_A3;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_A4;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_A5;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_A6;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_AO5;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_AO6;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_AQ;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_AX;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_A_CY;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_A_XOR;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_B;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_B1;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_B2;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_B3;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_B4;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_B5;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_B6;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_BO5;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_BO6;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_B_CY;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_B_XOR;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_C;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_C1;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_C2;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_C3;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_C4;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_C5;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_C6;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_CLK;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_CO5;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_CO6;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_C_CY;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_C_XOR;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_D;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_D1;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_D2;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_D3;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_D4;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_D5;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_D6;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_DMUX;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_DO5;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_DO6;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_D_CY;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_D_XOR;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_A;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_A1;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_A2;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_A3;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_A4;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_A5;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_A6;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_AO5;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_AO6;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_AQ;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_A_CY;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_A_XOR;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_B;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_B1;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_B2;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_B3;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_B4;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_B5;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_B6;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_BO5;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_BO6;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_BQ;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_B_CY;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_B_XOR;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_C;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_C1;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_C2;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_C3;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_C4;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_C5;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_C6;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_CLK;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_CO5;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_CO6;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_CQ;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_C_CY;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_C_XOR;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_D;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_D1;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_D2;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_D3;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_D4;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_D5;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_D6;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_DO5;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_DO6;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_DQ;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_D_CY;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_D_XOR;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_A;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_A1;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_A2;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_A3;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_A4;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_A5;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_A5Q;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_A6;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_AMUX;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_AO5;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_AO6;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_AQ;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_AX;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_A_CY;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_A_XOR;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_B;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_B1;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_B2;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_B3;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_B4;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_B5;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_B6;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_BMUX;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_BO5;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_BO6;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_B_CY;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_B_XOR;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_C;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_C1;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_C2;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_C3;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_C4;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_C5;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_C6;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_CLK;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_CO5;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_CO6;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_CQ;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_C_CY;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_C_XOR;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_D;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_D1;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_D2;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_D3;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_D4;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_D5;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_D6;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_DO5;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_DO6;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_D_CY;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_D_XOR;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_A;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_A1;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_A2;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_A3;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_A4;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_A5;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_A6;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_AO5;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_AO6;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_AQ;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_A_CY;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_A_XOR;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_B;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_B1;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_B2;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_B3;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_B4;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_B5;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_B5Q;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_B6;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_BMUX;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_BO5;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_BO6;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_BQ;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_B_CY;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_B_XOR;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_C;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_C1;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_C2;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_C3;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_C4;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_C5;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_C5Q;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_C6;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_CLK;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_CMUX;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_CO5;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_CO6;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_CQ;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_C_CY;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_C_XOR;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_D;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_D1;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_D2;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_D3;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_D4;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_D5;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_D6;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_DO5;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_DO6;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_DQ;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_D_CY;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_D_XOR;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_A;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_A1;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_A2;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_A3;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_A4;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_A5;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_A5Q;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_A6;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_AMUX;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_AO5;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_AO6;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_AQ;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_AX;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_A_CY;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_A_XOR;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_B;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_B1;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_B2;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_B3;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_B4;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_B5;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_B6;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_BMUX;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_BO5;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_BO6;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_B_CY;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_B_XOR;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_C;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_C1;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_C2;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_C3;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_C4;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_C5;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_C6;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_CLK;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_CO5;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_CO6;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_CQ;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_C_CY;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_C_XOR;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_D;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_D1;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_D2;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_D3;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_D4;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_D5;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_D6;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_DO5;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_DO6;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_DQ;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_D_CY;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_D_XOR;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_A;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_A1;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_A2;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_A3;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_A4;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_A5;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_A5Q;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_A6;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_AMUX;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_AO5;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_AO6;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_AQ;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_AX;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_A_CY;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_A_XOR;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_B;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_B1;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_B2;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_B3;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_B4;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_B5;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_B6;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_BMUX;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_BO5;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_BO6;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_B_CY;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_B_XOR;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_C;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_C1;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_C2;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_C3;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_C4;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_C5;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_C6;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_CLK;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_CO5;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_CO6;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_CQ;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_C_CY;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_C_XOR;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_D;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_D1;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_D2;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_D3;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_D4;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_D5;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_D6;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_DO5;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_DO6;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_DQ;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_D_CY;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_D_XOR;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_A;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_A1;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_A2;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_A3;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_A4;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_A5;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_A5Q;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_A6;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_AMUX;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_AO5;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_AO6;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_AQ;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_AX;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_A_CY;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_A_XOR;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_B;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_B1;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_B2;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_B3;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_B4;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_B5;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_B6;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_BMUX;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_BO5;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_BO6;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_B_CY;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_B_XOR;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_C;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_C1;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_C2;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_C3;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_C4;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_C5;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_C6;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_CLK;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_CO5;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_CO6;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_CQ;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_C_CY;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_C_XOR;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_D;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_D1;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_D2;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_D3;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_D4;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_D5;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_D6;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_DO5;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_DO6;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_D_CY;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_D_XOR;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_A;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_A1;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_A2;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_A3;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_A4;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_A5;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_A6;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_AO5;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_AO6;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_AQ;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_A_CY;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_A_XOR;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_B;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_B1;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_B2;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_B3;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_B4;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_B5;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_B6;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_BO5;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_BO6;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_BQ;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_B_CY;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_B_XOR;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_C;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_C1;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_C2;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_C3;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_C4;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_C5;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_C6;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_CLK;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_CO5;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_CO6;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_CQ;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_C_CY;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_C_XOR;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_D;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_D1;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_D2;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_D3;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_D4;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_D5;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_D6;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_DO5;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_DO6;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_DQ;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_D_CY;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_D_XOR;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_A;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_A1;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_A2;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_A3;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_A4;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_A5;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_A5Q;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_A6;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_AMUX;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_AO5;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_AO6;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_AQ;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_AX;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_A_CY;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_A_XOR;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_B;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_B1;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_B2;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_B3;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_B4;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_B5;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_B6;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_BMUX;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_BO5;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_BO6;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_BQ;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_BX;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_B_CY;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_B_XOR;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_C;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_C1;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_C2;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_C3;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_C4;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_C5;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_C6;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_CLK;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_CMUX;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_CO5;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_CO6;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_C_CY;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_C_XOR;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_D;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_D1;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_D2;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_D3;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_D4;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_D5;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_D6;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_DMUX;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_DO5;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_DO6;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_D_CY;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_D_XOR;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_A;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_A1;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_A2;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_A3;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_A4;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_A5;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_A5Q;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_A6;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_AMUX;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_AO5;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_AO6;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_AQ;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_AX;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_A_CY;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_A_XOR;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_B;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_B1;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_B2;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_B3;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_B4;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_B5;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_B6;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_BMUX;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_BO5;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_BO6;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_B_CY;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_B_XOR;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_C;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_C1;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_C2;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_C3;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_C4;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_C5;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_C6;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_CLK;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_CO5;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_CO6;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_CQ;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_C_CY;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_C_XOR;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_D;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_D1;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_D2;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_D3;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_D4;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_D5;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_D6;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_DMUX;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_DO5;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_DO6;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_D_CY;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_D_XOR;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_A;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_A1;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_A2;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_A3;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_A4;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_A5;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_A6;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_AO5;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_AO6;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_AQ;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_A_CY;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_A_XOR;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_B;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_B1;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_B2;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_B3;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_B4;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_B5;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_B6;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_BMUX;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_BO5;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_BO6;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_B_CY;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_B_XOR;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_C;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_C1;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_C2;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_C3;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_C4;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_C5;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_C6;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_CLK;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_CO5;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_CO6;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_CQ;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_C_CY;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_C_XOR;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_D;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_D1;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_D2;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_D3;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_D4;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_D5;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_D6;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_DMUX;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_DO5;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_DO6;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_D_CY;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_D_XOR;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_A;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_A1;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_A2;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_A3;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_A4;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_A5;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_A6;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_AO5;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_AO6;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_AQ;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_A_CY;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_A_XOR;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_B;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_B1;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_B2;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_B3;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_B4;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_B5;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_B6;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_BO5;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_BO6;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_BQ;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_B_CY;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_B_XOR;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_C;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_C1;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_C2;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_C3;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_C4;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_C5;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_C6;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_CLK;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_CO5;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_CO6;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_CQ;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_C_CY;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_C_XOR;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_D;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_D1;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_D2;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_D3;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_D4;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_D5;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_D6;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_DO5;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_DO6;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_DQ;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_D_CY;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_D_XOR;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_A;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_A1;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_A2;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_A3;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_A4;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_A5;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_A6;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_AO5;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_AO6;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_AQ;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_A_CY;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_A_XOR;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_B;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_B1;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_B2;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_B3;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_B4;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_B5;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_B6;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_BO5;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_BO6;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_BQ;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_B_CY;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_B_XOR;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_C;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_C1;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_C2;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_C3;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_C4;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_C5;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_C6;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_CLK;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_CO5;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_CO6;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_CQ;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_C_CY;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_C_XOR;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_D;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_D1;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_D2;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_D3;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_D4;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_D5;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_D6;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_DO5;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_DO6;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_D_CY;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_D_XOR;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_A;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_A1;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_A2;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_A3;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_A4;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_A5;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_A6;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_AO5;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_AO6;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_AQ;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_A_CY;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_A_XOR;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_B;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_B1;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_B2;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_B3;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_B4;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_B5;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_B6;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_BO5;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_BO6;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_BQ;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_B_CY;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_B_XOR;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_C;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_C1;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_C2;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_C3;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_C4;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_C5;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_C6;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_CLK;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_CO5;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_CO6;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_C_CY;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_C_XOR;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_D;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_D1;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_D2;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_D3;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_D4;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_D5;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_D6;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_DO5;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_DO6;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_D_CY;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_D_XOR;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_A;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_A1;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_A2;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_A3;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_A4;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_A5;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_A6;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_AO5;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_AO6;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_AQ;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_A_CY;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_A_XOR;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_B;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_B1;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_B2;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_B3;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_B4;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_B5;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_B6;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_BMUX;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_BO5;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_BO6;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_B_CY;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_B_XOR;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_C;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_C1;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_C2;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_C3;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_C4;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_C5;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_C6;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_CLK;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_CO5;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_CO6;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_C_CY;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_C_XOR;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_D;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_D1;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_D2;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_D3;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_D4;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_D5;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_D6;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_DMUX;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_DO5;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_DO6;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_D_CY;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_D_XOR;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_A;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_A1;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_A2;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_A3;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_A4;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_A5;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_A5Q;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_A6;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_AMUX;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_AO5;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_AO6;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_AQ;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_AX;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_A_CY;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_A_XOR;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_B;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_B1;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_B2;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_B3;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_B4;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_B5;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_B6;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_BO5;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_BO6;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_BQ;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_B_CY;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_B_XOR;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_C;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_C1;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_C2;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_C3;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_C4;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_C5;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_C6;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_CLK;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_CO5;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_CO6;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_CQ;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_C_CY;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_C_XOR;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_D;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_D1;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_D2;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_D3;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_D4;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_D5;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_D6;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_DO5;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_DO6;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_D_CY;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_D_XOR;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_A;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_A1;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_A2;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_A3;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_A4;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_A5;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_A6;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_AO5;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_AO6;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_AQ;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_A_CY;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_A_XOR;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_B;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_B1;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_B2;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_B3;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_B4;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_B5;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_B6;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_BO5;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_BO6;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_BQ;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_B_CY;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_B_XOR;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_C;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_C1;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_C2;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_C3;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_C4;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_C5;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_C6;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_CLK;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_CMUX;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_CO5;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_CO6;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_C_CY;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_C_XOR;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_D;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_D1;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_D2;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_D3;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_D4;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_D5;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_D6;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_DMUX;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_DO5;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_DO6;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_D_CY;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_D_XOR;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_A;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_A1;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_A2;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_A3;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_A4;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_A5;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_A6;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_AO5;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_AO6;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_AQ;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_A_CY;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_A_XOR;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_B;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_B1;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_B2;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_B3;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_B4;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_B5;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_B6;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_BO5;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_BO6;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_BQ;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_B_CY;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_B_XOR;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_C;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_C1;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_C2;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_C3;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_C4;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_C5;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_C6;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_CLK;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_CO5;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_CO6;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_CQ;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_C_CY;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_C_XOR;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_D;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_D1;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_D2;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_D3;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_D4;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_D5;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_D6;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_DO5;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_DO6;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_D_CY;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_D_XOR;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_A;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_A1;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_A2;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_A3;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_A4;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_A5;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_A6;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_AO5;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_AO6;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_AQ;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_A_CY;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_A_XOR;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_B;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_B1;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_B2;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_B3;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_B4;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_B5;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_B6;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_BO5;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_BO6;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_BQ;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_B_CY;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_B_XOR;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_C;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_C1;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_C2;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_C3;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_C4;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_C5;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_C6;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_CLK;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_CMUX;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_CO5;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_CO6;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_C_CY;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_C_XOR;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_D;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_D1;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_D2;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_D3;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_D4;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_D5;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_D6;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_DO5;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_DO6;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_D_CY;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_D_XOR;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_A;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_A1;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_A2;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_A3;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_A4;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_A5;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_A6;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_AO5;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_AO6;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_AQ;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_AX;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_A_CY;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_A_XOR;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_B;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_B1;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_B2;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_B3;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_B4;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_B5;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_B6;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_BO5;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_BO6;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_B_CY;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_B_XOR;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_C;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_C1;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_C2;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_C3;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_C4;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_C5;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_C6;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_CE;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_CLK;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_CO5;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_CO6;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_C_CY;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_C_XOR;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_D;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_D1;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_D2;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_D3;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_D4;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_D5;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_D6;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_DO5;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_DO6;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_D_CY;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_D_XOR;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_SR;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_A;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_A1;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_A2;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_A3;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_A4;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_A5;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_A6;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_AMUX;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_AO5;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_AO6;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_AQ;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_A_CY;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_A_XOR;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_B;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_B1;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_B2;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_B3;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_B4;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_B5;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_B6;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_BO5;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_BO6;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_B_CY;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_B_XOR;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_C;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_C1;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_C2;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_C3;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_C4;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_C5;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_C6;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_CLK;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_CO5;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_CO6;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_C_CY;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_C_XOR;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_D;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_D1;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_D2;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_D3;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_D4;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_D5;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_D6;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_DO5;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_DO6;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_D_CY;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_D_XOR;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_A;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_A1;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_A2;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_A3;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_A4;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_A5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_A6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_AMUX;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_AO5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_AO6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_A_CY;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_A_XOR;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_B;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_B1;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_B2;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_B3;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_B4;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_B5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_B6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_BO5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_BO6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_B_CY;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_B_XOR;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_C;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_C1;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_C2;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_C3;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_C4;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_C5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_C6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_CO5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_CO6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_C_CY;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_C_XOR;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_D;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_D1;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_D2;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_D3;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_D4;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_D5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_D6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_DO5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_DO6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_D_CY;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_D_XOR;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_A;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_A1;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_A2;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_A3;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_A4;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_A5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_A6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_AO5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_AO6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_A_CY;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_A_XOR;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_B;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_B1;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_B2;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_B3;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_B4;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_B5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_B6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_BO5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_BO6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_B_CY;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_B_XOR;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_C;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_C1;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_C2;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_C3;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_C4;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_C5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_C6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_CO5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_CO6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_C_CY;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_C_XOR;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_D;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_D1;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_D2;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_D3;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_D4;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_D5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_D6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_DO5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_DO6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_D_CY;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_D_XOR;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_A;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_A1;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_A2;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_A3;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_A4;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_A5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_A5Q;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_A6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_AMUX;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_AO5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_AO6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_AQ;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_AX;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_A_CY;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_A_XOR;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_B;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_B1;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_B2;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_B3;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_B4;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_B5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_B6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_BMUX;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_BO5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_BO6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_B_CY;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_B_XOR;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_C;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_C1;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_C2;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_C3;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_C4;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_C5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_C6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_CLK;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_CO5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_CO6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_C_CY;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_C_XOR;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_D;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_D1;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_D2;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_D3;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_D4;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_D5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_D6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_DO5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_DO6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_D_CY;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_D_XOR;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_A;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_A1;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_A2;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_A3;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_A4;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_A5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_A6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_AO5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_AO6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_AQ;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_A_CY;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_A_XOR;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_B;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_B1;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_B2;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_B3;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_B4;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_B5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_B6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_BO5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_BO6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_BQ;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_B_CY;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_B_XOR;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_C;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_C1;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_C2;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_C3;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_C4;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_C5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_C6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_CLK;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_CO5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_CO6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_C_CY;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_C_XOR;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_D;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_D1;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_D2;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_D3;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_D4;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_D5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_D6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_DO5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_DO6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_D_CY;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_D_XOR;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_A;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_A1;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_A2;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_A3;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_A4;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_A5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_A6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_AO5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_AO6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_AQ;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_A_CY;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_A_XOR;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_B;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_B1;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_B2;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_B3;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_B4;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_B5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_B6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_BO5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_BO6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_BQ;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_B_CY;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_B_XOR;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_C;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_C1;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_C2;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_C3;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_C4;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_C5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_C6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_CLK;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_CMUX;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_CO5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_CO6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_C_CY;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_C_XOR;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_D;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_D1;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_D2;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_D3;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_D4;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_D5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_D6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_DO5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_DO6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_D_CY;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_D_XOR;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_A;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_A1;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_A2;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_A3;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_A4;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_A5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_A6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_AO5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_AO6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_AQ;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_A_CY;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_A_XOR;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_B;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_B1;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_B2;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_B3;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_B4;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_B5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_B6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_BO5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_BO6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_BQ;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_B_CY;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_B_XOR;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_C;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_C1;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_C2;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_C3;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_C4;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_C5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_C6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_CLK;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_CO5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_CO6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_CQ;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_C_CY;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_C_XOR;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_D;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_D1;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_D2;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_D3;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_D4;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_D5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_D6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_DMUX;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_DO5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_DO6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_D_CY;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_D_XOR;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_A;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_A1;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_A2;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_A3;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_A4;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_A5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_A6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_AO5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_AO6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_AQ;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_A_CY;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_A_XOR;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_B;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_B1;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_B2;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_B3;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_B4;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_B5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_B6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_BO5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_BO6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_BQ;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_B_CY;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_B_XOR;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_C;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_C1;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_C2;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_C3;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_C4;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_C5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_C6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_CLK;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_CO5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_CO6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_CQ;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_C_CY;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_C_XOR;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_D;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_D1;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_D2;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_D3;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_D4;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_D5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_D6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_DO5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_DO6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_D_CY;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_D_XOR;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_A;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_A1;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_A2;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_A3;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_A4;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_A5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_A6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_AO5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_AO6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_AQ;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_A_CY;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_A_XOR;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_B;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_B1;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_B2;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_B3;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_B4;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_B5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_B6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_BO5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_BO6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_BQ;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_B_CY;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_B_XOR;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_C;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_C1;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_C2;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_C3;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_C4;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_C5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_C6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_CLK;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_CO5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_CO6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_CQ;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_C_CY;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_C_XOR;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_D;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_D1;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_D2;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_D3;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_D4;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_D5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_D6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_DO5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_DO6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_D_CY;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_D_XOR;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_A;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_A1;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_A2;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_A3;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_A4;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_A5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_A5Q;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_A6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_AMUX;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_AO5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_AO6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_AQ;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_AX;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_A_CY;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_A_XOR;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_B;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_B1;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_B2;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_B3;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_B4;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_B5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_B6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_BMUX;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_BO5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_BO6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_B_CY;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_B_XOR;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_C;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_C1;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_C2;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_C3;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_C4;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_C5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_C6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_CLK;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_CO5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_CO6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_C_CY;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_C_XOR;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_D;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_D1;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_D2;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_D3;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_D4;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_D5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_D6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_DO5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_DO6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_D_CY;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_D_XOR;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_A;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_A1;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_A2;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_A3;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_A4;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_A5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_A6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_AO5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_AO6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_AQ;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_A_CY;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_A_XOR;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_B;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_B1;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_B2;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_B3;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_B4;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_B5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_B6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_BO5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_BO6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_BQ;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_B_CY;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_B_XOR;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_C;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_C1;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_C2;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_C3;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_C4;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_C5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_C6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_CLK;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_CO5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_CO6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_CQ;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_C_CY;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_C_XOR;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_D;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_D1;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_D2;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_D3;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_D4;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_D5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_D6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_DO5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_DO6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_DQ;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_D_CY;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_D_XOR;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_A;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_A1;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_A2;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_A3;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_A4;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_A5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_A5Q;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_A6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_AMUX;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_AO5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_AO6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_AQ;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_AX;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_A_CY;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_A_XOR;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_B;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_B1;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_B2;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_B3;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_B4;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_B5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_B6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_BO5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_BO6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_BQ;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_B_CY;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_B_XOR;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_C;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_C1;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_C2;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_C3;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_C4;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_C5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_C6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_CLK;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_CMUX;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_CO5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_CO6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_C_CY;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_C_XOR;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_D;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_D1;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_D2;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_D3;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_D4;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_D5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_D6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_DO5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_DO6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_D_CY;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_D_XOR;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_A;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_A1;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_A2;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_A3;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_A4;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_A5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_A5Q;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_A6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_AMUX;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_AO5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_AO6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_AQ;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_A_CY;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_A_XOR;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_B;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_B1;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_B2;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_B3;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_B4;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_B5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_B5Q;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_B6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_BMUX;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_BO5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_BO6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_BQ;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_B_CY;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_B_XOR;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_C;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_C1;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_C2;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_C3;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_C4;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_C5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_C6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_CLK;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_CO5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_CO6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_CQ;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_C_CY;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_C_XOR;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_D;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_D1;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_D2;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_D3;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_D4;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_D5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_D6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_DMUX;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_DO5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_DO6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_D_CY;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_D_XOR;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_A;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_A1;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_A2;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_A3;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_A4;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_A5;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_A6;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_AO5;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_AO6;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_AQ;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_A_CY;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_A_XOR;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_B;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_B1;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_B2;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_B3;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_B4;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_B5;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_B6;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_BO5;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_BO6;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_BQ;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_B_CY;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_B_XOR;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_C;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_C1;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_C2;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_C3;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_C4;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_C5;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_C6;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_CLK;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_CO5;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_CO6;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_CQ;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_C_CY;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_C_XOR;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_D;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_D1;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_D2;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_D3;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_D4;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_D5;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_D6;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_DO5;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_DO6;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_DQ;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_D_CY;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_D_XOR;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_A;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_A1;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_A2;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_A3;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_A4;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_A5;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_A6;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_AO5;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_AO6;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_AQ;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_A_CY;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_A_XOR;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_B;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_B1;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_B2;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_B3;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_B4;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_B5;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_B6;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_BO5;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_BO6;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_BQ;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_B_CY;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_B_XOR;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_C;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_C1;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_C2;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_C3;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_C4;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_C5;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_C6;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_CLK;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_CO5;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_CO6;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_CQ;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_C_CY;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_C_XOR;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_D;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_D1;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_D2;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_D3;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_D4;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_D5;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_D6;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_DMUX;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_DO5;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_DO6;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_D_CY;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_D_XOR;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_A;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_A1;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_A2;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_A3;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_A4;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_A5;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_A6;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_AO5;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_AO6;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_AQ;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_A_CY;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_A_XOR;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_B;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_B1;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_B2;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_B3;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_B4;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_B5;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_B6;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_BMUX;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_BO5;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_BO6;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_B_CY;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_B_XOR;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_C;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_C1;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_C2;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_C3;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_C4;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_C5;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_C6;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_CLK;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_CO5;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_CO6;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_C_CY;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_C_XOR;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_D;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_D1;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_D2;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_D3;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_D4;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_D5;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_D6;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_DO5;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_DO6;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_D_CY;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_D_XOR;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_A;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_A1;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_A2;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_A3;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_A4;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_A5;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_A6;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_AO5;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_AO6;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_AQ;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_A_CY;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_A_XOR;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_B;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_B1;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_B2;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_B3;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_B4;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_B5;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_B6;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_BO5;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_BO6;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_BQ;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_B_CY;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_B_XOR;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_C;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_C1;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_C2;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_C3;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_C4;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_C5;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_C6;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_CLK;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_CMUX;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_CO5;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_CO6;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_C_CY;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_C_XOR;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_D;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_D1;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_D2;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_D3;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_D4;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_D5;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_D6;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_DO5;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_DO6;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_D_CY;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_D_XOR;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_A;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_A1;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_A2;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_A3;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_A4;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_A5;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_A6;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_AO5;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_AO6;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_AQ;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_A_CY;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_A_XOR;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_B;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_B1;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_B2;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_B3;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_B4;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_B5;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_B6;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_BO5;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_BO6;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_BQ;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_B_CY;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_B_XOR;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_C;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_C1;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_C2;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_C3;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_C4;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_C5;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_C6;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_CLK;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_CO5;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_CO6;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_CQ;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_C_CY;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_C_XOR;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_D;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_D1;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_D2;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_D3;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_D4;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_D5;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_D5Q;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_D6;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_DMUX;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_DO5;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_DO6;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_DQ;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_D_CY;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_D_XOR;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_A;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_A1;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_A2;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_A3;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_A4;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_A5;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_A6;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_AO5;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_AO6;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_AQ;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_A_CY;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_A_XOR;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_B;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_B1;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_B2;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_B3;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_B4;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_B5;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_B6;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_BO5;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_BO6;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_BQ;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_B_CY;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_B_XOR;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_C;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_C1;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_C2;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_C3;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_C4;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_C5;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_C6;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_CLK;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_CMUX;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_CO5;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_CO6;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_C_CY;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_C_XOR;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_D;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_D1;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_D2;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_D3;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_D4;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_D5;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_D6;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_DO5;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_DO6;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_D_CY;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_D_XOR;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_A;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_A1;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_A2;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_A3;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_A4;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_A5;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_A6;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_AO5;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_AO6;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_A_CY;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_A_XOR;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_B;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_B1;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_B2;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_B3;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_B4;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_B5;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_B6;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_BO5;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_BO6;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_BQ;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_B_CY;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_B_XOR;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_C;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_C1;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_C2;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_C3;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_C4;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_C5;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_C6;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_CLK;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_CO5;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_CO6;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_CQ;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_C_CY;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_C_XOR;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_D;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_D1;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_D2;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_D3;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_D4;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_D5;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_D6;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_DO5;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_DO6;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_DQ;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_D_CY;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_D_XOR;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_A;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_A1;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_A2;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_A3;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_A4;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_A5;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_A6;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_AO5;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_AO6;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_AQ;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_A_CY;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_A_XOR;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_B;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_B1;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_B2;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_B3;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_B4;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_B5;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_B6;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_BO5;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_BO6;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_BQ;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_B_CY;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_B_XOR;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_C;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_C1;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_C2;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_C3;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_C4;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_C5;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_C6;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_CLK;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_CMUX;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_CO5;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_CO6;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_C_CY;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_C_XOR;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_D;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_D1;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_D2;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_D3;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_D4;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_D5;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_D6;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_DO5;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_DO6;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_D_CY;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_D_XOR;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_A;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_A1;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_A2;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_A3;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_A4;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_A5;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_A5Q;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_A6;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_AMUX;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_AO5;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_AO6;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_AQ;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_A_CY;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_A_XOR;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_B;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_B1;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_B2;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_B3;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_B4;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_B5;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_B6;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_BO5;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_BO6;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_BQ;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_B_CY;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_B_XOR;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_C;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_C1;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_C2;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_C3;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_C4;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_C5;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_C6;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_CLK;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_CO5;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_CO6;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_CQ;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_C_CY;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_C_XOR;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_D;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_D1;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_D2;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_D3;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_D4;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_D5;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_D6;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_DO5;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_DO6;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_DQ;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_D_CY;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_D_XOR;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_A;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_A1;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_A2;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_A3;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_A4;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_A5;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_A5Q;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_A6;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_AMUX;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_AO5;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_AO6;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_AQ;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_A_CY;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_A_XOR;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_B;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_B1;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_B2;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_B3;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_B4;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_B5;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_B6;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_BO5;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_BO6;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_BQ;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_B_CY;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_B_XOR;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_C;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_C1;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_C2;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_C3;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_C4;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_C5;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_C6;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_CLK;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_CMUX;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_CO5;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_CO6;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_C_CY;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_C_XOR;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_D;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_D1;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_D2;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_D3;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_D4;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_D5;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_D6;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_DO5;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_DO6;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_D_CY;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_D_XOR;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_A;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_A1;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_A2;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_A3;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_A4;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_A5;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_A6;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_AO5;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_AO6;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_A_CY;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_A_XOR;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_B;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_B1;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_B2;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_B3;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_B4;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_B5;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_B6;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_BO5;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_BO6;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_BQ;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_B_CY;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_B_XOR;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_C;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_C1;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_C2;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_C3;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_C4;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_C5;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_C6;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_CLK;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_CO5;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_CO6;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_CQ;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_C_CY;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_C_XOR;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_D;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_D1;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_D2;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_D3;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_D4;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_D5;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_D6;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_DO5;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_DO6;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_DQ;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_D_CY;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_D_XOR;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_A;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_A1;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_A2;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_A3;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_A4;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_A5;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_A6;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_AO5;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_AO6;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_AQ;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_A_CY;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_A_XOR;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_B;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_B1;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_B2;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_B3;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_B4;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_B5;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_B6;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_BO5;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_BO6;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_BQ;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_B_CY;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_B_XOR;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_C;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_C1;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_C2;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_C3;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_C4;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_C5;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_C6;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_CLK;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_CO5;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_CO6;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_CQ;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_C_CY;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_C_XOR;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_D;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_D1;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_D2;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_D3;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_D4;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_D5;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_D6;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_DMUX;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_DO5;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_DO6;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_D_CY;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_D_XOR;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_A;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_A1;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_A2;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_A3;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_A4;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_A5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_A6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_AO5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_AO6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_AQ;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_A_CY;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_A_XOR;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_B;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_B1;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_B2;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_B3;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_B4;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_B5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_B6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_BO5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_BO6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_BQ;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_B_CY;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_B_XOR;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_C;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_C1;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_C2;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_C3;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_C4;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_C5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_C6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_CLK;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_CO5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_CO6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_CQ;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_C_CY;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_C_XOR;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_D;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_D1;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_D2;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_D3;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_D4;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_D5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_D5Q;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_D6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_DMUX;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_DO5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_DO6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_DQ;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_D_CY;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_D_XOR;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_A;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_A1;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_A2;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_A3;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_A4;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_A5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_A6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_AO5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_AO6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_AQ;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_A_CY;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_A_XOR;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_B;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_B1;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_B2;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_B3;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_B4;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_B5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_B6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_BO5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_BO6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_BQ;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_B_CY;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_B_XOR;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_C;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_C1;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_C2;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_C3;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_C4;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_C5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_C6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_CLK;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_CO5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_CO6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_CQ;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_C_CY;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_C_XOR;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_D;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_D1;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_D2;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_D3;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_D4;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_D5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_D6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_DO5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_DO6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_DQ;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_D_CY;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_D_XOR;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_A;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_A1;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_A2;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_A3;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_A4;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_A5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_A6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_AO5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_AO6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_A_CY;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_A_XOR;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_B;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_B1;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_B2;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_B3;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_B4;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_B5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_B6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_BO5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_BO6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_BQ;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_B_CY;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_B_XOR;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_C;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_C1;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_C2;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_C3;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_C4;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_C5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_C6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_CLK;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_CO5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_CO6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_CQ;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_C_CY;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_C_XOR;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_D;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_D1;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_D2;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_D3;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_D4;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_D5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_D6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_DMUX;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_DO5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_DO6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_D_CY;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_D_XOR;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_A;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_A1;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_A2;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_A3;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_A4;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_A5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_A6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_AO5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_AO6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_A_CY;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_A_XOR;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_B;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_B1;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_B2;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_B3;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_B4;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_B5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_B6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_BO5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_BO6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_B_CY;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_B_XOR;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_C;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_C1;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_C2;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_C3;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_C4;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_C5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_C6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_CO5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_CO6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_C_CY;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_C_XOR;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_D;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_D1;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_D2;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_D3;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_D4;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_D5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_D6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_DO5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_DO6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_D_CY;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_D_XOR;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_A;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_A1;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_A2;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_A3;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_A4;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_A5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_A6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_AO5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_AO6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_A_CY;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_A_XOR;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_B;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_B1;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_B2;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_B3;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_B4;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_B5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_B6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_BO5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_BO6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_B_CY;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_B_XOR;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_C;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_C1;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_C2;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_C3;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_C4;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_C5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_C6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_CO5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_CO6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_C_CY;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_C_XOR;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_D;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_D1;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_D2;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_D3;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_D4;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_D5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_D6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_DO5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_DO6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_D_CY;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_D_XOR;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_A;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_A1;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_A2;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_A3;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_A4;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_A5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_A6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_AO5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_AO6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_AQ;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_A_CY;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_A_XOR;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_B;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_B1;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_B2;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_B3;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_B4;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_B5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_B6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_BMUX;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_BO5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_BO6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_B_CY;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_B_XOR;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_C;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_C1;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_C2;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_C3;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_C4;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_C5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_C6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_CLK;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_CO5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_CO6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_C_CY;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_C_XOR;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_D;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_D1;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_D2;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_D3;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_D4;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_D5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_D6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_DO5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_DO6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_D_CY;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_D_XOR;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X162Y140_A;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X162Y140_A1;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X162Y140_A2;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X162Y140_A3;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X162Y140_A4;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X162Y140_A5;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X162Y140_A6;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X162Y140_AO5;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X162Y140_AO6;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X162Y140_A_CY;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X162Y140_A_XOR;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X162Y140_B;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X162Y140_B1;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X162Y140_B2;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X162Y140_B3;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X162Y140_B4;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X162Y140_B5;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X162Y140_B6;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X162Y140_BO5;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X162Y140_BO6;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X162Y140_B_CY;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X162Y140_B_XOR;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X162Y140_C;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X162Y140_C1;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X162Y140_C2;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X162Y140_C3;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X162Y140_C4;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X162Y140_C5;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X162Y140_C6;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X162Y140_CO5;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X162Y140_CO6;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X162Y140_C_CY;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X162Y140_C_XOR;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X162Y140_D;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X162Y140_D1;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X162Y140_D2;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X162Y140_D3;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X162Y140_D4;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X162Y140_D5;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X162Y140_D6;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X162Y140_DO5;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X162Y140_DO6;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X162Y140_D_CY;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X162Y140_D_XOR;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X163Y140_A;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X163Y140_A1;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X163Y140_A2;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X163Y140_A3;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X163Y140_A4;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X163Y140_A5;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X163Y140_A6;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X163Y140_AMUX;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X163Y140_AO5;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X163Y140_AO6;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X163Y140_A_CY;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X163Y140_A_XOR;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X163Y140_B;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X163Y140_B1;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X163Y140_B2;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X163Y140_B3;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X163Y140_B4;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X163Y140_B5;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X163Y140_B6;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X163Y140_BO5;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X163Y140_BO6;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X163Y140_B_CY;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X163Y140_B_XOR;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X163Y140_C;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X163Y140_C1;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X163Y140_C2;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X163Y140_C3;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X163Y140_C4;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X163Y140_C5;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X163Y140_C6;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X163Y140_CO5;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X163Y140_CO6;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X163Y140_C_CY;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X163Y140_C_XOR;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X163Y140_D;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X163Y140_D1;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X163Y140_D2;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X163Y140_D3;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X163Y140_D4;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X163Y140_D5;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X163Y140_D6;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X163Y140_DO5;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X163Y140_DO6;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X163Y140_D_CY;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X163Y140_D_XOR;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A1;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A2;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A3;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A4;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_AO5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_AO6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A_CY;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A_XOR;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B1;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B2;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B3;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B4;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_BO5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_BO6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B_CY;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B_XOR;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C1;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C2;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C3;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C4;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_CO5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_CO6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C_CY;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C_XOR;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D1;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D2;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D3;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D4;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_DO5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_DO6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D_CY;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D_XOR;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A1;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A2;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A3;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A4;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_AO5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_AO6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A_CY;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A_XOR;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B1;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B2;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B3;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B4;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_BO5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_BO6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B_CY;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B_XOR;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C1;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C2;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C3;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C4;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_CO5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_CO6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C_CY;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C_XOR;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D1;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D2;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D3;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D4;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_DO5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_DO6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D_CY;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D_XOR;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_A;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_A1;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_A2;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_A3;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_A4;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_A5;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_A6;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_AO5;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_AO6;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_A_CY;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_A_XOR;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_B;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_B1;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_B2;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_B3;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_B4;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_B5;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_B6;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_BO5;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_BO6;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_B_CY;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_B_XOR;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_C;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_C1;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_C2;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_C3;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_C4;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_C5;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_C6;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_CO5;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_CO6;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_C_CY;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_C_XOR;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_D;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_D1;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_D2;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_D3;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_D4;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_D5;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_D6;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_DO5;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_DO6;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_D_CY;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_D_XOR;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_A;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_A1;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_A2;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_A3;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_A4;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_A5;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_A6;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_AMUX;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_AO5;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_AO6;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_A_CY;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_A_XOR;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_B;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_B1;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_B2;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_B3;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_B4;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_B5;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_B6;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_BO5;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_BO6;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_B_CY;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_B_XOR;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_C;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_C1;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_C2;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_C3;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_C4;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_C5;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_C6;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_CO5;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_CO6;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_C_CY;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_C_XOR;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_D;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_D1;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_D2;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_D3;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_D4;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_D5;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_D6;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_DO5;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_DO6;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_D_CY;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_D_XOR;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_A;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_A1;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_A2;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_A3;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_A4;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_A5;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_A6;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_AO5;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_AO6;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_A_CY;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_A_XOR;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_B;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_B1;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_B2;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_B3;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_B4;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_B5;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_B6;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_BO5;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_BO6;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_B_CY;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_B_XOR;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_C;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_C1;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_C2;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_C3;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_C4;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_C5;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_C6;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_CO5;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_CO6;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_C_CY;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_C_XOR;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_D;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_D1;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_D2;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_D3;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_D4;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_D5;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_D6;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_DO5;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_DO6;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_D_CY;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_D_XOR;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_A;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_A1;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_A2;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_A3;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_A4;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_A5;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_A6;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_AMUX;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_AO5;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_AO6;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_A_CY;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_A_XOR;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_B;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_B1;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_B2;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_B3;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_B4;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_B5;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_B6;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_BO5;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_BO6;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_B_CY;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_B_XOR;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_C;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_C1;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_C2;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_C3;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_C4;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_C5;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_C6;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_CO5;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_CO6;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_C_CY;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_C_XOR;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_D;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_D1;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_D2;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_D3;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_D4;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_D5;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_D6;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_DO5;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_DO6;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_D_CY;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_D_XOR;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X162Y175_A;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X162Y175_A1;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X162Y175_A2;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X162Y175_A3;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X162Y175_A4;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X162Y175_A5;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X162Y175_A6;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X162Y175_AO5;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X162Y175_AO6;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X162Y175_A_CY;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X162Y175_A_XOR;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X162Y175_B;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X162Y175_B1;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X162Y175_B2;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X162Y175_B3;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X162Y175_B4;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X162Y175_B5;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X162Y175_B6;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X162Y175_BO5;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X162Y175_BO6;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X162Y175_B_CY;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X162Y175_B_XOR;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X162Y175_C;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X162Y175_C1;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X162Y175_C2;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X162Y175_C3;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X162Y175_C4;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X162Y175_C5;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X162Y175_C6;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X162Y175_CO5;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X162Y175_CO6;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X162Y175_C_CY;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X162Y175_C_XOR;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X162Y175_D;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X162Y175_D1;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X162Y175_D2;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X162Y175_D3;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X162Y175_D4;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X162Y175_D5;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X162Y175_D6;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X162Y175_DO5;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X162Y175_DO6;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X162Y175_D_CY;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X162Y175_D_XOR;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X163Y175_A;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X163Y175_A1;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X163Y175_A2;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X163Y175_A3;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X163Y175_A4;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X163Y175_A5;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X163Y175_A6;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X163Y175_AO5;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X163Y175_AO6;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X163Y175_A_CY;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X163Y175_A_XOR;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X163Y175_B;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X163Y175_B1;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X163Y175_B2;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X163Y175_B3;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X163Y175_B4;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X163Y175_B5;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X163Y175_B6;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X163Y175_BO5;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X163Y175_BO6;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X163Y175_B_CY;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X163Y175_B_XOR;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X163Y175_C;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X163Y175_C1;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X163Y175_C2;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X163Y175_C3;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X163Y175_C4;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X163Y175_C5;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X163Y175_C6;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X163Y175_CO5;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X163Y175_CO6;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X163Y175_C_CY;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X163Y175_C_XOR;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X163Y175_D;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X163Y175_D1;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X163Y175_D2;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X163Y175_D3;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X163Y175_D4;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X163Y175_D5;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X163Y175_D6;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X163Y175_DO5;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X163Y175_DO6;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X163Y175_D_CY;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X163Y175_D_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_AO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_AO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_BO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_BO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_CO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_CO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_DO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_DO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_AMUX;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_AO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_AO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_BO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_BO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_CO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_CO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_DO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_DO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D_XOR;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_A;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_A1;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_A2;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_A3;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_A4;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_A5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_A6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_AMUX;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_AO5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_AO6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_A_CY;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_A_XOR;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_B;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_B1;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_B2;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_B3;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_B4;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_B5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_B6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_BO5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_BO6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_BQ;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_B_CY;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_B_XOR;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_C;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_C1;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_C2;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_C3;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_C4;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_C5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_C6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_CLK;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_CO5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_CO6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_C_CY;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_C_XOR;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_D;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_D1;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_D2;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_D3;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_D4;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_D5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_D6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_DO5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_DO6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_D_CY;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_D_XOR;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_A;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_A1;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_A2;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_A3;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_A4;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_A5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_A6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_AMUX;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_AO5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_AO6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_A_CY;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_A_XOR;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_B;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_B1;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_B2;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_B3;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_B4;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_B5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_B6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_BO5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_BO6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_BQ;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_B_CY;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_B_XOR;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_C;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_C1;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_C2;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_C3;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_C4;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_C5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_C6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_CLK;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_CO5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_CO6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_C_CY;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_C_XOR;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_D;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_D1;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_D2;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_D3;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_D4;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_D5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_D6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_DO5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_DO6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_D_CY;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_D_XOR;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_A;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_A1;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_A2;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_A3;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_A4;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_A5;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_A6;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_AO5;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_AO6;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_AQ;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_A_CY;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_A_XOR;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_B;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_B1;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_B2;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_B3;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_B4;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_B5;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_B6;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_BO5;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_BO6;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_BQ;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_B_CY;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_B_XOR;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_C;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_C1;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_C2;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_C3;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_C4;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_C5;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_C6;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_CLK;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_CO5;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_CO6;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_C_CY;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_C_XOR;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_D;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_D1;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_D2;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_D3;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_D4;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_D5;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_D6;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_DO5;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_DO6;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_D_CY;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_D_XOR;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_A;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_A1;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_A2;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_A3;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_A4;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_A5;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_A6;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_AMUX;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_AO5;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_AO6;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_A_CY;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_A_XOR;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_B;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_B1;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_B2;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_B3;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_B4;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_B5;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_B6;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_BO5;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_BO6;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_B_CY;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_B_XOR;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_C;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_C1;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_C2;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_C3;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_C4;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_C5;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_C6;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_CMUX;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_CO5;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_CO6;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_C_CY;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_C_XOR;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_D;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_D1;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_D2;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_D3;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_D4;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_D5;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_D6;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_DO5;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_DO6;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_D_CY;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_D_XOR;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_A;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_A1;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_A2;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_A3;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_A4;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_A5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_A6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_AO5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_AO6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_AQ;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_A_CY;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_A_XOR;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_B;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_B1;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_B2;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_B3;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_B4;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_B5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_B6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_BO5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_BO6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_BQ;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_B_CY;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_B_XOR;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_C;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_C1;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_C2;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_C3;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_C4;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_C5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_C6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_CLK;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_CO5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_CO6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_CQ;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_C_CY;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_C_XOR;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_D;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_D1;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_D2;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_D3;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_D4;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_D5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_D6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_DO5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_DO6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_D_CY;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_D_XOR;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_A;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_A1;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_A2;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_A3;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_A4;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_A5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_A6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_AO5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_AO6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_AQ;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_A_CY;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_A_XOR;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_B;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_B1;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_B2;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_B3;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_B4;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_B5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_B6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_BO5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_BO6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_BQ;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_B_CY;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_B_XOR;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_C;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_C1;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_C2;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_C3;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_C4;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_C5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_C6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_CLK;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_CO5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_CO6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_CQ;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_C_CY;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_C_XOR;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_D;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_D1;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_D2;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_D3;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_D4;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_D5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_D6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_DO5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_DO6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_DQ;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_D_CY;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_D_XOR;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_A;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_A1;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_A2;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_A3;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_A4;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_A5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_A6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_AO5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_AO6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_AQ;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_A_CY;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_A_XOR;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_B;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_B1;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_B2;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_B3;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_B4;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_B5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_B6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_BO5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_BO6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_BQ;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_B_CY;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_B_XOR;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_C;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_C1;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_C2;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_C3;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_C4;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_C5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_C6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_CLK;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_CO5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_CO6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_CQ;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_C_CY;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_C_XOR;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_D;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_D1;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_D2;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_D3;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_D4;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_D5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_D6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_DO5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_DO6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_DQ;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_D_CY;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_D_XOR;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_A;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_A1;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_A2;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_A3;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_A4;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_A5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_A6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_AO5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_AO6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_AQ;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_A_CY;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_A_XOR;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_B;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_B1;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_B2;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_B3;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_B4;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_B5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_B6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_BO5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_BO6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_BQ;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_B_CY;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_B_XOR;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_C;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_C1;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_C2;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_C3;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_C4;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_C5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_C6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_CLK;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_CO5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_CO6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_CQ;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_C_CY;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_C_XOR;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_D;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_D1;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_D2;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_D3;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_D4;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_D5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_D6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_DO5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_DO6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_D_CY;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_D_XOR;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_A;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_A1;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_A2;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_A3;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_A4;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_A5;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_A6;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_AO5;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_AO6;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_AQ;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_A_CY;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_A_XOR;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_B;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_B1;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_B2;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_B3;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_B4;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_B5;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_B6;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_BO5;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_BO6;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_BQ;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_B_CY;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_B_XOR;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_C;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_C1;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_C2;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_C3;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_C4;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_C5;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_C6;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_CLK;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_CO5;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_CO6;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_CQ;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_C_CY;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_C_XOR;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_D;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_D1;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_D2;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_D3;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_D4;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_D5;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_D6;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_DO5;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_DO6;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_DQ;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_D_CY;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_D_XOR;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_A;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_A1;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_A2;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_A3;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_A4;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_A5;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_A6;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_AO5;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_AO6;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_AQ;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_A_CY;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_A_XOR;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_B;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_B1;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_B2;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_B3;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_B4;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_B5;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_B6;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_BO5;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_BO6;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_BQ;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_B_CY;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_B_XOR;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_C;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_C1;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_C2;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_C3;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_C4;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_C5;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_C6;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_CLK;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_CMUX;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_CO5;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_CO6;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_C_CY;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_C_XOR;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_D;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_D1;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_D2;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_D3;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_D4;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_D5;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_D6;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_DO5;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_DO6;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_D_CY;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_D_XOR;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_A;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_A1;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_A2;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_A3;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_A4;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_A5;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_A6;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_AO5;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_AO6;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_AQ;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_A_CY;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_A_XOR;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_B;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_B1;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_B2;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_B3;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_B4;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_B5;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_B6;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_BO5;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_BO6;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_BQ;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_B_CY;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_B_XOR;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_C;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_C1;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_C2;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_C3;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_C4;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_C5;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_C6;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_CLK;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_CMUX;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_CO5;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_CO6;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_C_CY;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_C_XOR;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_D;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_D1;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_D2;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_D3;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_D4;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_D5;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_D6;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_DO5;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_DO6;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_DQ;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_D_CY;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_D_XOR;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_A;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_A1;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_A2;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_A3;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_A4;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_A5;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_A5Q;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_A6;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_AMUX;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_AO5;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_AO6;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_AQ;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_A_CY;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_A_XOR;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_B;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_B1;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_B2;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_B3;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_B4;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_B5;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_B5Q;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_B6;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_BMUX;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_BO5;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_BO6;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_BQ;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_B_CY;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_B_XOR;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_C;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_C1;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_C2;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_C3;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_C4;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_C5;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_C6;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_CLK;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_CO5;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_CO6;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_C_CY;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_C_XOR;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_D;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_D1;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_D2;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_D3;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_D4;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_D5;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_D6;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_DO5;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_DO6;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_D_CY;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_D_XOR;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_A;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_A1;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_A2;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_A3;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_A4;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_A5;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_A6;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_AO5;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_AO6;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_AQ;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_A_CY;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_A_XOR;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_B;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_B1;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_B2;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_B3;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_B4;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_B5;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_B6;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_BMUX;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_BO5;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_BO6;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_B_CY;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_B_XOR;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_C;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_C1;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_C2;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_C3;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_C4;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_C5;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_C6;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_CLK;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_CMUX;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_CO5;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_CO6;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_C_CY;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_C_XOR;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_D;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_D1;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_D2;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_D3;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_D4;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_D5;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_D6;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_DO5;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_DO6;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_D_CY;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_D_XOR;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_A;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_A1;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_A2;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_A3;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_A4;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_A5;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_A6;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_AO5;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_AO6;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_AQ;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_A_CY;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_A_XOR;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_B;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_B1;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_B2;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_B3;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_B4;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_B5;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_B6;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_BO5;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_BO6;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_B_CY;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_B_XOR;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_C;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_C1;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_C2;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_C3;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_C4;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_C5;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_C6;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_CLK;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_CO5;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_CO6;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_C_CY;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_C_XOR;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_D;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_D1;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_D2;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_D3;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_D4;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_D5;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_D6;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_DMUX;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_DO5;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_DO6;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_D_CY;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_D_XOR;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_A;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_A1;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_A2;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_A3;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_A4;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_A5;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_A6;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_AO5;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_AO6;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_AQ;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_A_CY;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_A_XOR;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_B;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_B1;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_B2;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_B3;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_B4;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_B5;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_B6;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_BO5;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_BO6;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_BQ;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_B_CY;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_B_XOR;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_C;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_C1;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_C2;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_C3;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_C4;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_C5;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_C6;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_CLK;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_CO5;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_CO6;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_CQ;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_C_CY;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_C_XOR;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_D;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_D1;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_D2;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_D3;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_D4;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_D5;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_D5Q;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_D6;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_DMUX;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_DO5;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_DO6;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_DQ;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_D_CY;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_D_XOR;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_A;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_A1;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_A2;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_A3;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_A4;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_A5;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_A6;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_AO5;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_AO6;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_AQ;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_A_CY;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_A_XOR;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_B;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_B1;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_B2;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_B3;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_B4;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_B5;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_B5Q;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_B6;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_BMUX;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_BO5;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_BO6;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_BQ;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_B_CY;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_B_XOR;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_C;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_C1;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_C2;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_C3;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_C4;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_C5;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_C6;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_CLK;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_CO5;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_CO6;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_CQ;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_C_CY;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_C_XOR;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_D;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_D1;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_D2;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_D3;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_D4;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_D5;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_D5Q;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_D6;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_DMUX;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_DO5;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_DO6;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_DQ;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_D_CY;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_D_XOR;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_A;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_A1;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_A2;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_A3;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_A4;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_A5;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_A6;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_AO5;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_AO6;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_AQ;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_A_CY;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_A_XOR;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_B;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_B1;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_B2;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_B3;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_B4;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_B5;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_B5Q;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_B6;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_BMUX;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_BO5;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_BO6;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_BQ;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_B_CY;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_B_XOR;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_C;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_C1;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_C2;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_C3;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_C4;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_C5;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_C6;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_CLK;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_CO5;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_CO6;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_CQ;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_C_CY;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_C_XOR;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_D;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_D1;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_D2;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_D3;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_D4;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_D5;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_D6;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_DO5;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_DO6;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_D_CY;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_D_XOR;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_A;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_A1;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_A2;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_A3;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_A4;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_A5;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_A5Q;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_A6;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_AMUX;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_AO5;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_AO6;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_AQ;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_A_CY;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_A_XOR;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_B;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_B1;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_B2;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_B3;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_B4;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_B5;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_B6;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_BO5;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_BO6;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_BQ;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_B_CY;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_B_XOR;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_C;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_C1;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_C2;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_C3;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_C4;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_C5;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_C6;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_CLK;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_CO5;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_CO6;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_CQ;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_C_CY;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_C_XOR;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_D;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_D1;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_D2;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_D3;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_D4;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_D5;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_D6;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_DO5;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_DO6;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_DQ;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_D_CY;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_D_XOR;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_A;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_A1;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_A2;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_A3;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_A4;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_A5;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_A6;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_AO5;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_AO6;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_AQ;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_A_CY;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_A_XOR;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_B;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_B1;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_B2;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_B3;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_B4;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_B5;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_B6;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_BO5;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_BO6;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_BQ;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_B_CY;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_B_XOR;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_C;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_C1;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_C2;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_C3;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_C4;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_C5;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_C6;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_CLK;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_CO5;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_CO6;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_CQ;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_C_CY;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_C_XOR;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_D;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_D1;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_D2;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_D3;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_D4;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_D5;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_D6;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_DO5;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_DO6;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_D_CY;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_D_XOR;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_A;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_A1;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_A2;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_A3;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_A4;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_A5;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_A6;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_AMUX;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_AO5;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_AO6;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_A_CY;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_A_XOR;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_B;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_B1;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_B2;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_B3;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_B4;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_B5;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_B6;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_BO5;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_BO6;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_BQ;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_B_CY;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_B_XOR;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_C;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_C1;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_C2;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_C3;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_C4;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_C5;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_C5Q;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_C6;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_CLK;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_CMUX;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_CO5;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_CO6;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_CQ;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_C_CY;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_C_XOR;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_D;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_D1;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_D2;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_D3;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_D4;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_D5;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_D6;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_DO5;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_DO6;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_DQ;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_D_CY;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_D_XOR;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_A;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_A1;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_A2;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_A3;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_A4;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_A5;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_A6;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_AO5;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_AO6;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_AQ;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_A_CY;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_A_XOR;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_B;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_B1;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_B2;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_B3;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_B4;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_B5;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_B6;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_BO5;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_BO6;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_BQ;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_B_CY;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_B_XOR;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_C;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_C1;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_C2;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_C3;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_C4;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_C5;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_C6;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_CLK;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_CMUX;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_CO5;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_CO6;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_C_CY;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_C_XOR;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_D;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_D1;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_D2;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_D3;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_D4;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_D5;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_D6;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_DMUX;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_DO5;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_DO6;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_D_CY;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_D_XOR;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_A;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_A1;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_A2;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_A3;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_A4;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_A5;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_A6;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_AO5;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_AO6;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_AQ;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_A_CY;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_A_XOR;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_B;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_B1;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_B2;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_B3;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_B4;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_B5;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_B6;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_BO5;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_BO6;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_BQ;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_B_CY;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_B_XOR;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_C;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_C1;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_C2;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_C3;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_C4;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_C5;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_C6;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_CLK;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_CO5;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_CO6;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_CQ;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_C_CY;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_C_XOR;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_D;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_D1;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_D2;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_D3;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_D4;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_D5;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_D6;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_DO5;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_DO6;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_DQ;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_D_CY;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_D_XOR;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_A;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_A1;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_A2;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_A3;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_A4;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_A5;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_A6;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_AO5;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_AO6;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_AQ;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_A_CY;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_A_XOR;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_B;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_B1;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_B2;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_B3;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_B4;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_B5;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_B6;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_BO5;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_BO6;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_BQ;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_B_CY;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_B_XOR;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_C;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_C1;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_C2;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_C3;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_C4;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_C5;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_C6;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_CLK;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_CO5;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_CO6;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_C_CY;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_C_XOR;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_D;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_D1;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_D2;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_D3;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_D4;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_D5;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_D6;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_DO5;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_DO6;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_D_CY;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_D_XOR;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_A;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_A1;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_A2;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_A3;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_A4;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_A5;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_A6;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_AO5;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_AO6;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_AQ;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_A_CY;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_A_XOR;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_B;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_B1;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_B2;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_B3;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_B4;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_B5;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_B6;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_BO5;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_BO6;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_BQ;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_B_CY;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_B_XOR;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_C;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_C1;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_C2;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_C3;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_C4;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_C5;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_C6;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_CLK;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_CO5;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_CO6;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_CQ;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_C_CY;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_C_XOR;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_D;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_D1;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_D2;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_D3;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_D4;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_D5;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_D6;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_DO5;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_DO6;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_DQ;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_D_CY;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_D_XOR;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_A;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_A1;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_A2;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_A3;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_A4;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_A5;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_A6;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_AO5;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_AO6;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_AQ;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_A_CY;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_A_XOR;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_B;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_B1;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_B2;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_B3;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_B4;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_B5;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_B6;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_BMUX;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_BO5;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_BO6;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_B_CY;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_B_XOR;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_C;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_C1;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_C2;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_C3;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_C4;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_C5;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_C6;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_CLK;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_CMUX;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_CO5;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_CO6;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_C_CY;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_C_XOR;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_D;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_D1;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_D2;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_D3;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_D4;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_D5;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_D6;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_DO5;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_DO6;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_D_CY;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_D_XOR;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_A;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_A1;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_A2;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_A3;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_A4;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_A5;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_A6;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_AO5;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_AO6;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_AQ;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_A_CY;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_A_XOR;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_B;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_B1;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_B2;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_B3;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_B4;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_B5;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_B6;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_BO5;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_BO6;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_BQ;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_B_CY;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_B_XOR;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_C;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_C1;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_C2;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_C3;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_C4;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_C5;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_C6;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_CLK;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_CMUX;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_CO5;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_CO6;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_C_CY;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_C_XOR;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_D;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_D1;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_D2;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_D3;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_D4;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_D5;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_D6;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_DO5;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_DO6;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_D_CY;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_D_XOR;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_A;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_A1;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_A2;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_A3;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_A4;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_A5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_A6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_AO5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_AO6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_AQ;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_A_CY;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_A_XOR;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_B;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_B1;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_B2;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_B3;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_B4;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_B5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_B6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_BMUX;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_BO5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_BO6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_B_CY;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_B_XOR;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_C;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_C1;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_C2;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_C3;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_C4;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_C5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_C6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_CLK;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_CO5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_CO6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_C_CY;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_C_XOR;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_D;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_D1;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_D2;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_D3;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_D4;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_D5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_D6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_DO5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_DO6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_D_CY;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_D_XOR;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_A;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_A1;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_A2;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_A3;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_A4;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_A5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_A6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_AO5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_AO6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_AQ;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_A_CY;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_A_XOR;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_B;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_B1;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_B2;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_B3;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_B4;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_B5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_B6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_BO5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_BO6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_BQ;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_B_CY;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_B_XOR;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_C;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_C1;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_C2;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_C3;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_C4;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_C5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_C6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_CLK;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_CMUX;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_CO5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_CO6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_C_CY;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_C_XOR;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_D;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_D1;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_D2;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_D3;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_D4;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_D5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_D6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_DO5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_DO6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_D_CY;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_D_XOR;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_A;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_A1;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_A2;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_A3;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_A4;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_A5;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_A6;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_AMUX;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_AO5;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_AO6;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_A_CY;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_A_XOR;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_B;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_B1;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_B2;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_B3;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_B4;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_B5;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_B6;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_BO5;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_BO6;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_B_CY;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_B_XOR;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_C;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_C1;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_C2;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_C3;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_C4;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_C5;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_C6;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_CO5;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_CO6;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_C_CY;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_C_XOR;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_D;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_D1;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_D2;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_D3;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_D4;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_D5;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_D6;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_DO5;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_DO6;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_D_CY;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_D_XOR;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_A;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_A1;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_A2;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_A3;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_A4;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_A5;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_A6;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_AO5;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_AO6;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_A_CY;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_A_XOR;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_B;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_B1;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_B2;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_B3;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_B4;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_B5;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_B6;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_BO5;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_BO6;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_B_CY;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_B_XOR;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_C;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_C1;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_C2;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_C3;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_C4;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_C5;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_C6;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_CO5;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_CO6;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_C_CY;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_C_XOR;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_D;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_D1;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_D2;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_D3;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_D4;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_D5;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_D6;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_DO5;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_DO6;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_D_CY;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_D_XOR;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_A;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_A1;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_A2;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_A3;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_A4;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_A5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_A6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_AO5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_AO6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_AQ;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_AX;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_A_CY;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_A_XOR;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_B;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_B1;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_B2;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_B3;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_B4;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_B5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_B6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_BO5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_BO6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_B_CY;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_B_XOR;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_C;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_C1;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_C2;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_C3;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_C4;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_C5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_C6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_CLK;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_CO5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_CO6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_C_CY;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_C_XOR;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_D;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_D1;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_D2;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_D3;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_D4;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_D5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_D6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_DO5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_DO6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_D_CY;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_D_XOR;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_A;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_A1;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_A2;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_A3;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_A4;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_A5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_A6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_AO5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_AO6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_A_CY;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_A_XOR;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_B;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_B1;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_B2;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_B3;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_B4;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_B5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_B6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_BO5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_BO6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_B_CY;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_B_XOR;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_C;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_C1;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_C2;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_C3;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_C4;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_C5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_C6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_CO5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_CO6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_C_CY;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_C_XOR;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_D;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_D1;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_D2;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_D3;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_D4;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_D5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_D6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_DO5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_DO6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_D_CY;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_D_XOR;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_A;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_A1;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_A2;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_A3;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_A4;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_A5;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_A6;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_AO5;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_AO6;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_A_CY;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_A_XOR;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_B;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_B1;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_B2;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_B3;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_B4;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_B5;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_B6;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_BO5;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_BO6;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_B_CY;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_B_XOR;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_C;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_C1;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_C2;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_C3;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_C4;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_C5;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_C6;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_CO5;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_CO6;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_C_CY;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_C_XOR;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_D;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_D1;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_D2;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_D3;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_D4;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_D5;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_D6;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_DO5;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_DO6;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_D_CY;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_D_XOR;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_A;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_A1;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_A2;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_A3;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_A4;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_A5;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_A6;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_AO5;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_AO6;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_A_CY;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_A_XOR;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_B;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_B1;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_B2;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_B3;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_B4;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_B5;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_B6;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_BO5;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_BO6;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_B_CY;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_B_XOR;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_C;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_C1;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_C2;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_C3;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_C4;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_C5;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_C6;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_CO5;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_CO6;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_C_CY;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_C_XOR;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_D;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_D1;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_D2;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_D3;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_D4;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_D5;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_D6;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_DO5;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_DO6;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_D_CY;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_D_XOR;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_A;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_A1;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_A2;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_A3;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_A4;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_A5;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_A6;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_AO5;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_AO6;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_AQ;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_A_CY;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_A_XOR;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_B;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_B1;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_B2;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_B3;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_B4;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_B5;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_B6;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_BO5;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_BO6;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_BQ;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_B_CY;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_B_XOR;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_C;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_C1;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_C2;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_C3;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_C4;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_C5;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_C6;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_CLK;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_CO5;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_CO6;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_C_CY;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_C_XOR;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_D;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_D1;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_D2;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_D3;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_D4;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_D5;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_D6;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_DO5;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_DO6;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_D_CY;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X18Y133_D_XOR;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_A;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_A1;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_A2;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_A3;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_A4;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_A5;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_A6;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_AO5;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_AO6;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_A_CY;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_A_XOR;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_B;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_B1;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_B2;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_B3;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_B4;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_B5;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_B6;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_BO5;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_BO6;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_B_CY;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_B_XOR;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_C;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_C1;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_C2;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_C3;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_C4;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_C5;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_C6;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_CO5;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_CO6;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_C_CY;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_C_XOR;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_D;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_D1;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_D2;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_D3;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_D4;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_D5;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_D6;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_DO5;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_DO6;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_D_CY;
  wire [0:0] CLBLM_R_X13Y133_SLICE_X19Y133_D_XOR;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_A;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_A1;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_A2;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_A3;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_A4;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_A5;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_A6;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_AMUX;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_AO5;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_AO6;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_A_CY;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_A_XOR;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_B;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_B1;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_B2;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_B3;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_B4;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_B5;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_B6;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_BO5;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_BO6;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_B_CY;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_B_XOR;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_C;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_C1;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_C2;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_C3;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_C4;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_C5;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_C6;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_CMUX;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_CO5;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_CO6;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_C_CY;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_C_XOR;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_D;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_D1;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_D2;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_D3;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_D4;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_D5;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_D6;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_DO5;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_DO6;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_D_CY;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_D_XOR;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_A;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_A1;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_A2;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_A3;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_A4;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_A5;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_A6;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_AO5;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_AO6;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_AQ;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_A_CY;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_A_XOR;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_B;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_B1;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_B2;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_B3;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_B4;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_B5;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_B6;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_BO5;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_BO6;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_BQ;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_B_CY;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_B_XOR;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_C;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_C1;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_C2;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_C3;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_C4;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_C5;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_C6;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_CLK;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_CO5;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_CO6;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_CQ;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_C_CY;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_C_XOR;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_D;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_D1;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_D2;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_D3;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_D4;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_D5;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_D6;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_DO5;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_DO6;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_DQ;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_D_CY;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_D_XOR;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_A;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_A1;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_A2;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_A3;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_A4;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_A5;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_A6;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_AO5;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_AO6;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_AQ;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_A_CY;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_A_XOR;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_B;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_B1;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_B2;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_B3;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_B4;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_B5;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_B6;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_BO5;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_BO6;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_BQ;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_B_CY;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_B_XOR;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_C;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_C1;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_C2;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_C3;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_C4;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_C5;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_C6;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_CLK;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_CO5;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_CO6;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_C_CY;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_C_XOR;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_D;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_D1;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_D2;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_D3;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_D4;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_D5;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_D6;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_DO5;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_DO6;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_D_CY;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X18Y135_D_XOR;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_A;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_A1;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_A2;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_A3;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_A4;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_A5;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_A6;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_AO5;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_AO6;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_A_CY;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_A_XOR;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_B;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_B1;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_B2;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_B3;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_B4;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_B5;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_B6;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_BO5;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_BO6;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_B_CY;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_B_XOR;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_C;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_C1;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_C2;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_C3;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_C4;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_C5;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_C6;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_CO5;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_CO6;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_C_CY;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_C_XOR;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_D;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_D1;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_D2;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_D3;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_D4;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_D5;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_D6;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_DO5;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_DO6;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_D_CY;
  wire [0:0] CLBLM_R_X13Y135_SLICE_X19Y135_D_XOR;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_A;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_A1;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_A2;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_A3;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_A4;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_A5;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_A6;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_AO5;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_AO6;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_AQ;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_A_CY;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_A_XOR;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_B;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_B1;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_B2;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_B3;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_B4;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_B5;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_B6;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_BO5;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_BO6;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_BQ;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_B_CY;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_B_XOR;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_C;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_C1;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_C2;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_C3;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_C4;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_C5;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_C6;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_CLK;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_CO5;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_CO6;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_CQ;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_C_CY;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_C_XOR;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_D;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_D1;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_D2;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_D3;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_D4;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_D5;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_D6;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_DO5;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_DO6;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_D_CY;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X18Y136_D_XOR;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_A;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_A1;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_A2;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_A3;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_A4;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_A5;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_A6;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_AO5;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_AO6;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_A_CY;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_A_XOR;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_B;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_B1;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_B2;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_B3;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_B4;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_B5;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_B6;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_BO5;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_BO6;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_B_CY;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_B_XOR;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_C;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_C1;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_C2;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_C3;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_C4;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_C5;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_C6;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_CO5;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_CO6;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_C_CY;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_C_XOR;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_D;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_D1;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_D2;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_D3;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_D4;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_D5;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_D6;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_DO5;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_DO6;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_D_CY;
  wire [0:0] CLBLM_R_X13Y136_SLICE_X19Y136_D_XOR;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_A;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_A1;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_A2;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_A3;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_A4;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_A5;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_A5Q;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_A6;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_AMUX;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_AO5;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_AO6;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_AQ;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_AX;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_A_CY;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_A_XOR;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_B;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_B1;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_B2;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_B3;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_B4;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_B5;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_B6;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_BMUX;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_BO5;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_BO6;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_B_CY;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_B_XOR;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_C;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_C1;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_C2;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_C3;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_C4;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_C5;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_C6;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_CLK;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_CMUX;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_CO5;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_CO6;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_C_CY;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_C_XOR;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_D;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_D1;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_D2;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_D3;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_D4;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_D5;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_D6;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_DO5;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_DO6;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_D_CY;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_D_XOR;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_A;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_A1;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_A2;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_A3;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_A4;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_A5;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_A6;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_AO5;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_AO6;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_AQ;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_A_CY;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_A_XOR;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_B;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_B1;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_B2;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_B3;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_B4;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_B5;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_B6;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_BO5;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_BO6;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_BQ;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_B_CY;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_B_XOR;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_C;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_C1;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_C2;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_C3;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_C4;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_C5;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_C6;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_CLK;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_CO5;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_CO6;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_CQ;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_C_CY;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_C_XOR;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_D;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_D1;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_D2;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_D3;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_D4;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_D5;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_D6;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_DO5;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_DO6;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_D_CY;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_D_XOR;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_A;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_A1;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_A2;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_A3;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_A4;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_A5;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_A6;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_AO5;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_AO6;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_AQ;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_A_CY;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_A_XOR;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_B;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_B1;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_B2;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_B3;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_B4;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_B5;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_B6;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_BO5;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_BO6;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_B_CY;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_B_XOR;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_C;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_C1;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_C2;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_C3;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_C4;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_C5;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_C6;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_CLK;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_CO5;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_CO6;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_C_CY;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_C_XOR;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_D;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_D1;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_D2;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_D3;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_D4;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_D5;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_D6;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_DO5;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_DO6;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_D_CY;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_D_XOR;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_A;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_A1;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_A2;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_A3;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_A4;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_A5;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_A6;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_AO5;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_AO6;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_A_CY;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_A_XOR;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_B;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_B1;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_B2;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_B3;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_B4;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_B5;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_B6;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_BO5;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_BO6;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_B_CY;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_B_XOR;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_C;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_C1;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_C2;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_C3;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_C4;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_C5;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_C6;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_CO5;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_CO6;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_C_CY;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_C_XOR;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_D;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_D1;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_D2;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_D3;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_D4;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_D5;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_D6;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_DO5;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_DO6;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_D_CY;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_D_XOR;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_A;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_A1;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_A2;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_A3;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_A4;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_A5;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_A6;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_AO5;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_AO6;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_AQ;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_A_CY;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_A_XOR;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_B;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_B1;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_B2;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_B3;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_B4;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_B5;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_B6;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_BO5;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_BO6;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_B_CY;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_B_XOR;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_C;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_C1;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_C2;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_C3;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_C4;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_C5;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_C6;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_CLK;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_CO5;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_CO6;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_C_CY;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_C_XOR;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_D;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_D1;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_D2;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_D3;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_D4;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_D5;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_D6;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_DO5;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_DO6;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_D_CY;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X18Y139_D_XOR;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_A;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_A1;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_A2;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_A3;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_A4;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_A5;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_A6;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_AO5;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_AO6;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_AQ;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_A_CY;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_A_XOR;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_B;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_B1;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_B2;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_B3;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_B4;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_B5;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_B6;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_BO5;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_BO6;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_B_CY;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_B_XOR;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_C;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_C1;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_C2;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_C3;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_C4;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_C5;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_C6;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_CLK;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_CO5;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_CO6;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_C_CY;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_C_XOR;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_D;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_D1;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_D2;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_D3;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_D4;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_D5;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_D6;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_DO5;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_DO6;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_D_CY;
  wire [0:0] CLBLM_R_X13Y139_SLICE_X19Y139_D_XOR;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_A;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_A1;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_A2;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_A3;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_A4;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_A5;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_A6;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_AO5;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_AO6;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_AQ;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_A_CY;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_A_XOR;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_B;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_B1;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_B2;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_B3;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_B4;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_B5;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_B6;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_BO5;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_BO6;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_BQ;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_B_CY;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_B_XOR;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_C;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_C1;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_C2;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_C3;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_C4;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_C5;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_C6;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_CLK;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_CO5;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_CO6;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_CQ;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_C_CY;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_C_XOR;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_D;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_D1;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_D2;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_D3;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_D4;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_D5;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_D6;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_DO5;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_DO6;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_D_CY;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X18Y140_D_XOR;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_A;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_A1;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_A2;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_A3;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_A4;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_A5;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_A6;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_AO5;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_AO6;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_AQ;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_A_CY;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_A_XOR;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_B;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_B1;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_B2;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_B3;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_B4;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_B5;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_B6;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_BO5;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_BO6;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_BQ;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_B_CY;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_B_XOR;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_C;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_C1;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_C2;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_C3;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_C4;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_C5;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_C6;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_CLK;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_CO5;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_CO6;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_C_CY;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_C_XOR;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_D;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_D1;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_D2;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_D3;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_D4;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_D5;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_D6;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_DO5;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_DO6;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_D_CY;
  wire [0:0] CLBLM_R_X13Y140_SLICE_X19Y140_D_XOR;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_A;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_A1;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_A2;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_A3;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_A4;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_A5;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_A6;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_AMUX;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_AO5;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_AO6;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_A_CY;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_A_XOR;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_B;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_B1;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_B2;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_B3;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_B4;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_B5;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_B6;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_BMUX;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_BO5;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_BO6;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_B_CY;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_B_XOR;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_C;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_C1;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_C2;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_C3;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_C4;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_C5;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_C6;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_CMUX;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_CO5;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_CO6;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_C_CY;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_C_XOR;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_D;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_D1;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_D2;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_D3;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_D4;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_D5;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_D6;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_DMUX;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_DO5;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_DO6;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_D_CY;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X18Y141_D_XOR;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_A;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_A1;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_A2;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_A3;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_A4;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_A5;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_A6;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_AO5;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_AO6;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_AQ;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_A_CY;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_A_XOR;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_B;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_B1;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_B2;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_B3;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_B4;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_B5;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_B6;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_BO5;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_BO6;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_BQ;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_B_CY;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_B_XOR;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_C;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_C1;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_C2;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_C3;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_C4;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_C5;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_C6;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_CLK;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_CMUX;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_CO5;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_CO6;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_C_CY;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_C_XOR;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_D;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_D1;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_D2;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_D3;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_D4;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_D5;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_D6;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_DO5;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_DO6;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_D_CY;
  wire [0:0] CLBLM_R_X13Y141_SLICE_X19Y141_D_XOR;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_A;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_A1;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_A2;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_A3;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_A4;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_A5;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_A6;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_AO5;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_AO6;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_A_CY;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_A_XOR;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_B;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_B1;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_B2;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_B3;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_B4;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_B5;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_B6;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_BO5;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_BO6;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_B_CY;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_B_XOR;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_C;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_C1;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_C2;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_C3;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_C4;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_C5;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_C6;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_CO5;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_CO6;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_C_CY;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_C_XOR;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_D;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_D1;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_D2;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_D3;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_D4;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_D5;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_D6;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_DO5;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_DO6;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_D_CY;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X18Y142_D_XOR;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_A;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_A1;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_A2;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_A3;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_A4;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_A5;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_A6;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_AO5;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_AO6;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_AQ;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_A_CY;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_A_XOR;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_B;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_B1;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_B2;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_B3;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_B4;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_B5;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_B6;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_BO5;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_BO6;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_B_CY;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_B_XOR;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_C;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_C1;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_C2;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_C3;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_C4;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_C5;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_C6;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_CLK;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_CO5;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_CO6;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_C_CY;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_C_XOR;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_D;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_D1;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_D2;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_D3;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_D4;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_D5;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_D6;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_DO5;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_DO6;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_D_CY;
  wire [0:0] CLBLM_R_X13Y142_SLICE_X19Y142_D_XOR;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_A;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_A1;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_A2;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_A3;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_A4;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_A5;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_A6;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_AMUX;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_AO5;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_AO6;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_AQ;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_AX;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_A_CY;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_A_XOR;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_B;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_B1;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_B2;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_B3;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_B4;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_B5;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_B6;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_BO5;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_BO6;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_BQ;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_BX;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_B_CY;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_B_XOR;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_C;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_C1;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_C2;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_C3;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_C4;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_C5;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_C6;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_CE;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_CLK;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_CMUX;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_CO5;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_CO6;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_C_CY;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_C_XOR;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_D;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_D1;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_D2;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_D3;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_D4;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_D5;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_D6;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_DO5;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_DO6;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_D_CY;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_D_XOR;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X18Y143_SR;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X19Y143_A;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X19Y143_A1;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X19Y143_A2;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X19Y143_A3;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X19Y143_A4;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X19Y143_A5;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X19Y143_A6;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X19Y143_AO5;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X19Y143_AO6;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X19Y143_A_CY;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X19Y143_A_XOR;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X19Y143_B;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X19Y143_B1;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X19Y143_B2;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X19Y143_B3;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X19Y143_B4;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X19Y143_B5;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X19Y143_B6;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X19Y143_BO5;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X19Y143_BO6;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X19Y143_B_CY;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X19Y143_B_XOR;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X19Y143_C;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X19Y143_C1;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X19Y143_C2;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X19Y143_C3;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X19Y143_C4;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X19Y143_C5;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X19Y143_C6;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X19Y143_CO5;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X19Y143_CO6;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X19Y143_C_CY;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X19Y143_C_XOR;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X19Y143_D;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X19Y143_D1;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X19Y143_D2;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X19Y143_D3;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X19Y143_D4;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X19Y143_D5;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X19Y143_D6;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X19Y143_DO5;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X19Y143_DO6;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X19Y143_D_CY;
  wire [0:0] CLBLM_R_X13Y143_SLICE_X19Y143_D_XOR;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_A;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_A1;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_A2;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_A3;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_A4;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_A5;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_A6;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_AO5;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_AO6;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_AQ;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_A_CY;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_A_XOR;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_B;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_B1;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_B2;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_B3;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_B4;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_B5;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_B6;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_BMUX;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_BO5;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_BO6;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_B_CY;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_B_XOR;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_C;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_C1;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_C2;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_C3;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_C4;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_C5;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_C6;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_CLK;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_CO5;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_CO6;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_C_CY;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_C_XOR;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_D;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_D1;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_D2;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_D3;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_D4;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_D5;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_D6;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_DO5;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_DO6;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_D_CY;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X18Y144_D_XOR;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_A;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_A1;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_A2;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_A3;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_A4;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_A5;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_A6;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_AO5;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_AO6;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_AQ;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_A_CY;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_A_XOR;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_B;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_B1;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_B2;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_B3;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_B4;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_B5;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_B6;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_BO5;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_BO6;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_B_CY;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_B_XOR;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_C;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_C1;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_C2;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_C3;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_C4;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_C5;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_C6;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_CLK;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_CO5;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_CO6;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_C_CY;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_C_XOR;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_D;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_D1;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_D2;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_D3;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_D4;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_D5;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_D6;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_DO5;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_DO6;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_D_CY;
  wire [0:0] CLBLM_R_X13Y144_SLICE_X19Y144_D_XOR;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_A;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_A1;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_A2;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_A3;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_A4;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_A5;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_A6;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_AO5;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_AO6;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_AQ;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_A_CY;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_A_XOR;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_B;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_B1;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_B2;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_B3;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_B4;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_B5;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_B6;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_BO5;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_BO6;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_B_CY;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_B_XOR;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_C;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_C1;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_C2;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_C3;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_C4;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_C5;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_C6;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_CLK;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_CO5;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_CO6;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_C_CY;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_C_XOR;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_D;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_D1;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_D2;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_D3;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_D4;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_D5;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_D6;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_DO5;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_DO6;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_D_CY;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X20Y142_D_XOR;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_A;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_A1;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_A2;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_A3;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_A4;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_A5;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_A6;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_AO5;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_AO6;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_A_CY;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_A_XOR;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_B;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_B1;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_B2;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_B3;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_B4;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_B5;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_B6;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_BO5;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_BO6;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_B_CY;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_B_XOR;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_C;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_C1;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_C2;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_C3;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_C4;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_C5;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_C6;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_CO5;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_CO6;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_C_CY;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_C_XOR;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_D;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_D1;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_D2;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_D3;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_D4;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_D5;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_D6;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_DO5;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_DO6;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_D_CY;
  wire [0:0] CLBLM_R_X15Y142_SLICE_X21Y142_D_XOR;
  wire [0:0] CLBLM_R_X37Y138_SLICE_X56Y138_A;
  wire [0:0] CLBLM_R_X37Y138_SLICE_X56Y138_A1;
  wire [0:0] CLBLM_R_X37Y138_SLICE_X56Y138_A2;
  wire [0:0] CLBLM_R_X37Y138_SLICE_X56Y138_A3;
  wire [0:0] CLBLM_R_X37Y138_SLICE_X56Y138_A4;
  wire [0:0] CLBLM_R_X37Y138_SLICE_X56Y138_A5;
  wire [0:0] CLBLM_R_X37Y138_SLICE_X56Y138_A6;
  wire [0:0] CLBLM_R_X37Y138_SLICE_X56Y138_AO5;
  wire [0:0] CLBLM_R_X37Y138_SLICE_X56Y138_AO6;
  wire [0:0] CLBLM_R_X37Y138_SLICE_X56Y138_A_CY;
  wire [0:0] CLBLM_R_X37Y138_SLICE_X56Y138_A_XOR;
  wire [0:0] CLBLM_R_X37Y138_SLICE_X56Y138_B;
  wire [0:0] CLBLM_R_X37Y138_SLICE_X56Y138_B1;
  wire [0:0] CLBLM_R_X37Y138_SLICE_X56Y138_B2;
  wire [0:0] CLBLM_R_X37Y138_SLICE_X56Y138_B3;
  wire [0:0] CLBLM_R_X37Y138_SLICE_X56Y138_B4;
  wire [0:0] CLBLM_R_X37Y138_SLICE_X56Y138_B5;
  wire [0:0] CLBLM_R_X37Y138_SLICE_X56Y138_B6;
  wire [0:0] CLBLM_R_X37Y138_SLICE_X56Y138_BO5;
  wire [0:0] CLBLM_R_X37Y138_SLICE_X56Y138_BO6;
  wire [0:0] CLBLM_R_X37Y138_SLICE_X56Y138_B_CY;
  wire [0:0] CLBLM_R_X37Y138_SLICE_X56Y138_B_XOR;
  wire [0:0] CLBLM_R_X37Y138_SLICE_X56Y138_C;
  wire [0:0] CLBLM_R_X37Y138_SLICE_X56Y138_C1;
  wire [0:0] CLBLM_R_X37Y138_SLICE_X56Y138_C2;
  wire [0:0] CLBLM_R_X37Y138_SLICE_X56Y138_C3;
  wire [0:0] CLBLM_R_X37Y138_SLICE_X56Y138_C4;
  wire [0:0] CLBLM_R_X37Y138_SLICE_X56Y138_C5;
  wire [0:0] CLBLM_R_X37Y138_SLICE_X56Y138_C6;
  wire [0:0] CLBLM_R_X37Y138_SLICE_X56Y138_CO5;
  wire [0:0] CLBLM_R_X37Y138_SLICE_X56Y138_CO6;
  wire [0:0] CLBLM_R_X37Y138_SLICE_X56Y138_C_CY;
  wire [0:0] CLBLM_R_X37Y138_SLICE_X56Y138_C_XOR;
  wire [0:0] CLBLM_R_X37Y138_SLICE_X56Y138_D;
  wire [0:0] CLBLM_R_X37Y138_SLICE_X56Y138_D1;
  wire [0:0] CLBLM_R_X37Y138_SLICE_X56Y138_D2;
  wire [0:0] CLBLM_R_X37Y138_SLICE_X56Y138_D3;
  wire [0:0] CLBLM_R_X37Y138_SLICE_X56Y138_D4;
  wire [0:0] CLBLM_R_X37Y138_SLICE_X56Y138_D5;
  wire [0:0] CLBLM_R_X37Y138_SLICE_X56Y138_D6;
  wire [0:0] CLBLM_R_X37Y138_SLICE_X56Y138_DO5;
  wire [0:0] CLBLM_R_X37Y138_SLICE_X56Y138_DO6;
  wire [0:0] CLBLM_R_X37Y138_SLICE_X56Y138_D_CY;
  wire [0:0] CLBLM_R_X37Y138_SLICE_X56Y138_D_XOR;
  wire [0:0] CLBLM_R_X37Y138_SLICE_X57Y138_A;
  wire [0:0] CLBLM_R_X37Y138_SLICE_X57Y138_A1;
  wire [0:0] CLBLM_R_X37Y138_SLICE_X57Y138_A2;
  wire [0:0] CLBLM_R_X37Y138_SLICE_X57Y138_A3;
  wire [0:0] CLBLM_R_X37Y138_SLICE_X57Y138_A4;
  wire [0:0] CLBLM_R_X37Y138_SLICE_X57Y138_A5;
  wire [0:0] CLBLM_R_X37Y138_SLICE_X57Y138_A6;
  wire [0:0] CLBLM_R_X37Y138_SLICE_X57Y138_AO5;
  wire [0:0] CLBLM_R_X37Y138_SLICE_X57Y138_AO6;
  wire [0:0] CLBLM_R_X37Y138_SLICE_X57Y138_A_CY;
  wire [0:0] CLBLM_R_X37Y138_SLICE_X57Y138_A_XOR;
  wire [0:0] CLBLM_R_X37Y138_SLICE_X57Y138_B;
  wire [0:0] CLBLM_R_X37Y138_SLICE_X57Y138_B1;
  wire [0:0] CLBLM_R_X37Y138_SLICE_X57Y138_B2;
  wire [0:0] CLBLM_R_X37Y138_SLICE_X57Y138_B3;
  wire [0:0] CLBLM_R_X37Y138_SLICE_X57Y138_B4;
  wire [0:0] CLBLM_R_X37Y138_SLICE_X57Y138_B5;
  wire [0:0] CLBLM_R_X37Y138_SLICE_X57Y138_B6;
  wire [0:0] CLBLM_R_X37Y138_SLICE_X57Y138_BO5;
  wire [0:0] CLBLM_R_X37Y138_SLICE_X57Y138_BO6;
  wire [0:0] CLBLM_R_X37Y138_SLICE_X57Y138_B_CY;
  wire [0:0] CLBLM_R_X37Y138_SLICE_X57Y138_B_XOR;
  wire [0:0] CLBLM_R_X37Y138_SLICE_X57Y138_C;
  wire [0:0] CLBLM_R_X37Y138_SLICE_X57Y138_C1;
  wire [0:0] CLBLM_R_X37Y138_SLICE_X57Y138_C2;
  wire [0:0] CLBLM_R_X37Y138_SLICE_X57Y138_C3;
  wire [0:0] CLBLM_R_X37Y138_SLICE_X57Y138_C4;
  wire [0:0] CLBLM_R_X37Y138_SLICE_X57Y138_C5;
  wire [0:0] CLBLM_R_X37Y138_SLICE_X57Y138_C6;
  wire [0:0] CLBLM_R_X37Y138_SLICE_X57Y138_CO5;
  wire [0:0] CLBLM_R_X37Y138_SLICE_X57Y138_CO6;
  wire [0:0] CLBLM_R_X37Y138_SLICE_X57Y138_C_CY;
  wire [0:0] CLBLM_R_X37Y138_SLICE_X57Y138_C_XOR;
  wire [0:0] CLBLM_R_X37Y138_SLICE_X57Y138_D;
  wire [0:0] CLBLM_R_X37Y138_SLICE_X57Y138_D1;
  wire [0:0] CLBLM_R_X37Y138_SLICE_X57Y138_D2;
  wire [0:0] CLBLM_R_X37Y138_SLICE_X57Y138_D3;
  wire [0:0] CLBLM_R_X37Y138_SLICE_X57Y138_D4;
  wire [0:0] CLBLM_R_X37Y138_SLICE_X57Y138_D5;
  wire [0:0] CLBLM_R_X37Y138_SLICE_X57Y138_D6;
  wire [0:0] CLBLM_R_X37Y138_SLICE_X57Y138_DO5;
  wire [0:0] CLBLM_R_X37Y138_SLICE_X57Y138_DO6;
  wire [0:0] CLBLM_R_X37Y138_SLICE_X57Y138_D_CY;
  wire [0:0] CLBLM_R_X37Y138_SLICE_X57Y138_D_XOR;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_A;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_A1;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_A2;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_A3;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_A4;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_A5;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_A6;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_AMUX;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_AO5;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_AO6;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_A_CY;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_A_XOR;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_B;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_B1;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_B2;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_B3;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_B4;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_B5;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_B6;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_BO5;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_BO6;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_B_CY;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_B_XOR;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_C;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_C1;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_C2;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_C3;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_C4;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_C5;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_C6;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_CMUX;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_CO5;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_CO6;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_C_CY;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_C_XOR;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_D;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_D1;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_D2;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_D3;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_D4;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_D5;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_D6;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_DO5;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_DO6;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_D_CY;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_D_XOR;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_A;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_A1;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_A2;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_A3;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_A4;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_A5;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_A6;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_AO5;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_AO6;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_AQ;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_A_CY;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_A_XOR;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_B;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_B1;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_B2;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_B3;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_B4;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_B5;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_B6;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_BO5;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_BO6;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_B_CY;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_B_XOR;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_C;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_C1;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_C2;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_C3;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_C4;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_C5;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_C6;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_CLK;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_CO5;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_CO6;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_C_CY;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_C_XOR;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_D;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_D1;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_D2;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_D3;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_D4;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_D5;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_D6;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_DO5;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_DO6;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_D_CY;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_D_XOR;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_A;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_A1;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_A2;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_A3;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_A4;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_A5;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_A6;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_AO5;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_AO6;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_A_CY;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_A_XOR;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_B;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_B1;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_B2;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_B3;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_B4;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_B5;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_B6;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_BO5;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_BO6;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_B_CY;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_B_XOR;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_C;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_C1;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_C2;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_C3;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_C4;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_C5;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_C6;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_CO5;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_CO6;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_C_CY;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_C_XOR;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_D;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_D1;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_D2;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_D3;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_D4;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_D5;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_D6;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_DO5;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_DO6;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_D_CY;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_D_XOR;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_A;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_A1;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_A2;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_A3;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_A4;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_A5;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_A6;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_AO5;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_AO6;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_AQ;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_A_CY;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_A_XOR;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_B;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_B1;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_B2;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_B3;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_B4;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_B5;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_B6;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_BO5;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_BO6;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_BQ;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_B_CY;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_B_XOR;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_C;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_C1;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_C2;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_C3;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_C4;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_C5;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_C6;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_CLK;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_CMUX;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_CO5;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_CO6;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_C_CY;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_C_XOR;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_D;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_D1;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_D2;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_D3;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_D4;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_D5;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_D6;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_DO5;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_DO6;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_D_CY;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_D_XOR;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_A;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_A1;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_A2;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_A3;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_A4;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_A5;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_A6;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_AO5;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_AO6;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_AQ;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_A_CY;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_A_XOR;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_B;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_B1;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_B2;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_B3;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_B4;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_B5;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_B6;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_BMUX;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_BO5;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_BO6;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_B_CY;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_B_XOR;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_C;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_C1;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_C2;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_C3;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_C4;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_C5;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_C6;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_CLK;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_CO5;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_CO6;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_C_CY;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_C_XOR;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_D;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_D1;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_D2;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_D3;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_D4;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_D5;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_D6;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_DO5;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_DO6;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_D_CY;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_D_XOR;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_A;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_A1;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_A2;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_A3;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_A4;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_A5;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_A6;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_AO5;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_AO6;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_AQ;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_A_CY;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_A_XOR;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_B;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_B1;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_B2;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_B3;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_B4;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_B5;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_B6;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_BO5;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_BO6;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_BQ;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_B_CY;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_B_XOR;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_C;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_C1;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_C2;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_C3;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_C4;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_C5;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_C6;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_CLK;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_CO5;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_CO6;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_CQ;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_C_CY;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_C_XOR;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_D;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_D1;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_D2;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_D3;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_D4;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_D5;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_D6;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_DO5;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_DO6;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_DQ;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_D_CY;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_D_XOR;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_A;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_A1;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_A2;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_A3;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_A4;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_A5;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_A6;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_AO5;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_AO6;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_AQ;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_A_CY;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_A_XOR;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_B;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_B1;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_B2;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_B3;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_B4;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_B5;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_B6;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_BO5;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_BO6;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_BQ;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_B_CY;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_B_XOR;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_C;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_C1;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_C2;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_C3;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_C4;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_C5;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_C6;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_CLK;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_CO5;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_CO6;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_C_CY;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_C_XOR;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_D;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_D1;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_D2;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_D3;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_D4;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_D5;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_D6;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_DO5;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_DO6;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_D_CY;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_D_XOR;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_A;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_A1;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_A2;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_A3;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_A4;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_A5;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_A6;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_AMUX;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_AO5;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_AO6;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_AQ;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_A_CY;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_A_XOR;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_B;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_B1;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_B2;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_B3;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_B4;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_B5;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_B6;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_BMUX;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_BO5;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_BO6;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_BQ;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_B_CY;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_B_XOR;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_C;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_C1;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_C2;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_C3;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_C4;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_C5;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_C6;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_CLK;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_CO5;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_CO6;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_CQ;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_C_CY;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_C_XOR;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_D;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_D1;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_D2;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_D3;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_D4;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_D5;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_D6;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_DO5;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_DO6;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_D_CY;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_D_XOR;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_A;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_A1;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_A2;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_A3;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_A4;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_A5;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_A6;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_AMUX;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_AO5;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_AO6;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_A_CY;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_A_XOR;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_B;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_B1;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_B2;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_B3;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_B4;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_B5;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_B6;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_BO5;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_BO6;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_B_CY;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_B_XOR;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_C;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_C1;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_C2;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_C3;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_C4;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_C5;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_C6;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_CO5;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_CO6;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_C_CY;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_C_XOR;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_D;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_D1;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_D2;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_D3;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_D4;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_D5;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_D6;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_DO5;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_DO6;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_D_CY;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_D_XOR;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_A;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_A1;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_A2;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_A3;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_A4;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_A5;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_A6;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_AO5;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_AO6;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_AQ;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_A_CY;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_A_XOR;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_B;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_B1;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_B2;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_B3;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_B4;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_B5;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_B6;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_BO5;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_BO6;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_B_CY;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_B_XOR;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_C;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_C1;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_C2;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_C3;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_C4;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_C5;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_C6;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_CLK;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_CO5;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_CO6;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_C_CY;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_C_XOR;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_D;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_D1;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_D2;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_D3;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_D4;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_D5;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_D6;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_DO5;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_DO6;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_D_CY;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_D_XOR;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_A;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_A1;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_A2;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_A3;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_A4;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_A5;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_A6;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_AMUX;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_AO5;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_AO6;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_A_CY;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_A_XOR;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_B;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_B1;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_B2;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_B3;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_B4;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_B5;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_B6;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_BO5;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_BO6;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_B_CY;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_B_XOR;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_C;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_C1;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_C2;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_C3;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_C4;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_C5;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_C6;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_CO5;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_CO6;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_C_CY;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_C_XOR;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_D;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_D1;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_D2;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_D3;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_D4;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_D5;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_D6;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_DO5;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_DO6;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_D_CY;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_D_XOR;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_A;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_A1;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_A2;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_A3;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_A4;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_A5;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_A6;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_AO5;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_AO6;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_AQ;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_A_CY;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_A_XOR;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_B;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_B1;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_B2;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_B3;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_B4;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_B5;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_B6;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_BO5;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_BO6;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_B_CY;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_B_XOR;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_C;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_C1;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_C2;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_C3;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_C4;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_C5;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_C6;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_CLK;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_CO5;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_CO6;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_C_CY;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_C_XOR;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_D;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_D1;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_D2;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_D3;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_D4;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_D5;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_D6;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_DO5;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_DO6;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_D_CY;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_D_XOR;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_A;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_A1;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_A2;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_A3;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_A4;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_A5;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_A6;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_AO5;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_AO6;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_A_CY;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_A_XOR;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_B;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_B1;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_B2;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_B3;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_B4;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_B5;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_B6;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_BO5;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_BO6;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_B_CY;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_B_XOR;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_C;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_C1;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_C2;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_C3;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_C4;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_C5;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_C6;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_CO5;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_CO6;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_C_CY;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_C_XOR;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_D;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_D1;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_D2;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_D3;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_D4;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_D5;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_D6;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_DO5;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_DO6;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_D_CY;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_D_XOR;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_A;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_A1;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_A2;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_A3;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_A4;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_A5;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_A6;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_AO5;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_AO6;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_A_CY;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_A_XOR;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_B;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_B1;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_B2;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_B3;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_B4;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_B5;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_B6;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_BO5;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_BO6;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_B_CY;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_B_XOR;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_C;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_C1;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_C2;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_C3;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_C4;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_C5;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_C6;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_CMUX;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_CO5;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_CO6;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_C_CY;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_C_XOR;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_D;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_D1;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_D2;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_D3;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_D4;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_D5;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_D6;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_DO5;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_DO6;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_D_CY;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_D_XOR;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_A;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_A1;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_A2;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_A3;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_A4;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_A5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_A6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_AMUX;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_AO5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_AO6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_A_CY;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_A_XOR;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_B;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_B1;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_B2;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_B3;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_B4;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_B5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_B6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_BO5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_BO6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_B_CY;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_B_XOR;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_C;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_C1;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_C2;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_C3;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_C4;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_C5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_C6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_CO5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_CO6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_C_CY;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_C_XOR;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_D;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_D1;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_D2;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_D3;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_D4;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_D5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_D6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_DO5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_DO6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_D_CY;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_D_XOR;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_A;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_A1;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_A2;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_A3;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_A4;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_A5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_A6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_AMUX;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_AO5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_AO6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_A_CY;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_A_XOR;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_B;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_B1;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_B2;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_B3;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_B4;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_B5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_B6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_BO5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_BO6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_B_CY;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_B_XOR;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_C;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_C1;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_C2;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_C3;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_C4;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_C5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_C6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_CO5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_CO6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_C_CY;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_C_XOR;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_D;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_D1;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_D2;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_D3;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_D4;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_D5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_D6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_DO5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_DO6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_D_CY;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_D_XOR;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_A;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_A1;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_A2;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_A3;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_A4;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_A5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_A6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_AMUX;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_AO5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_AO6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_A_CY;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_A_XOR;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_B;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_B1;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_B2;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_B3;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_B4;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_B5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_B6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_BO5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_BO6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_B_CY;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_B_XOR;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_C;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_C1;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_C2;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_C3;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_C4;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_C5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_C6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_CO5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_CO6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_C_CY;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_C_XOR;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_D;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_D1;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_D2;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_D3;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_D4;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_D5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_D6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_DO5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_DO6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_D_CY;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_D_XOR;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_A;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_A1;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_A2;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_A3;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_A4;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_A5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_A6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_AMUX;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_AO5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_AO6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_A_CY;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_A_XOR;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_B;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_B1;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_B2;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_B3;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_B4;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_B5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_B6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_BO5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_BO6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_B_CY;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_B_XOR;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_C;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_C1;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_C2;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_C3;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_C4;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_C5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_C6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_CO5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_CO6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_C_CY;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_C_XOR;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_D;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_D1;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_D2;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_D3;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_D4;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_D5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_D6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_DO5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_DO6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_D_CY;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_D_XOR;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_A;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_A1;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_A2;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_A3;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_A4;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_A5;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_A6;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_AMUX;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_AO5;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_AO6;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_A_CY;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_A_XOR;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_B;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_B1;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_B2;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_B3;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_B4;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_B5;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_B6;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_BO5;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_BO6;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_B_CY;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_B_XOR;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_C;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_C1;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_C2;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_C3;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_C4;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_C5;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_C6;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_CO5;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_CO6;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_C_CY;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_C_XOR;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_D;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_D1;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_D2;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_D3;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_D4;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_D5;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_D6;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_DO5;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_DO6;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_D_CY;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_D_XOR;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_A;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_A1;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_A2;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_A3;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_A4;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_A5;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_A6;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_AMUX;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_AO5;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_AO6;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_A_CY;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_A_XOR;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_B;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_B1;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_B2;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_B3;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_B4;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_B5;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_B6;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_BO5;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_BO6;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_B_CY;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_B_XOR;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_C;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_C1;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_C2;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_C3;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_C4;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_C5;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_C6;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_CO5;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_CO6;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_C_CY;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_C_XOR;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_D;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_D1;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_D2;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_D3;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_D4;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_D5;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_D6;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_DO5;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_DO6;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_D_CY;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_D_XOR;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_A;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_A1;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_A2;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_A3;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_A4;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_A5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_A6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_AO5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_AO6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_A_CY;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_A_XOR;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_B;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_B1;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_B2;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_B3;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_B4;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_B5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_B6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_BO5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_BO6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_B_CY;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_B_XOR;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_C;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_C1;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_C2;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_C3;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_C4;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_C5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_C6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_CO5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_CO6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_C_CY;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_C_XOR;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_D;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_D1;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_D2;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_D3;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_D4;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_D5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_D6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_DO5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_DO6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_D_CY;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_D_XOR;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_A;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_A1;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_A2;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_A3;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_A4;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_A5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_A6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_AO5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_AO6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_AQ;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_A_CY;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_A_XOR;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_B;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_B1;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_B2;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_B3;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_B4;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_B5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_B6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_BMUX;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_BO5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_BO6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_B_CY;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_B_XOR;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_C;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_C1;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_C2;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_C3;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_C4;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_C5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_C6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_CLK;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_CMUX;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_CO5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_CO6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_C_CY;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_C_XOR;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_D;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_D1;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_D2;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_D3;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_D4;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_D5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_D6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_DMUX;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_DO5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_DO6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_D_CY;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_D_XOR;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_A;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_A1;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_A2;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_A3;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_A4;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_A5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_A6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_AMUX;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_AO5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_AO6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_A_CY;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_A_XOR;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_B;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_B1;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_B2;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_B3;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_B4;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_B5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_B6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_BMUX;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_BO5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_BO6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_B_CY;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_B_XOR;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_C;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_C1;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_C2;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_C3;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_C4;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_C5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_C6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_CO5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_CO6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_C_CY;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_C_XOR;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_D;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_D1;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_D2;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_D3;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_D4;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_D5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_D6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_DMUX;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_DO5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_DO6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_D_CY;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_D_XOR;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_A;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_A1;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_A2;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_A3;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_A4;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_A5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_A6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_AO5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_AO6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_A_CY;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_A_XOR;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_B;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_B1;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_B2;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_B3;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_B4;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_B5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_B6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_BO5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_BO6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_B_CY;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_B_XOR;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_C;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_C1;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_C2;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_C3;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_C4;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_C5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_C6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_CO5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_CO6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_C_CY;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_C_XOR;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_D;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_D1;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_D2;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_D3;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_D4;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_D5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_D6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_DO5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_DO6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_D_CY;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_D_XOR;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_A;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_A1;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_A2;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_A3;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_A4;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_A5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_A5Q;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_A6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_AMUX;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_AO5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_AO6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_AQ;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_AX;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_A_CY;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_A_XOR;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_B;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_B1;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_B2;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_B3;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_B4;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_B5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_B6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_BMUX;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_BO5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_BO6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_B_CY;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_B_XOR;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_C;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_C1;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_C2;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_C3;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_C4;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_C5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_C6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_CLK;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_CMUX;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_CO5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_CO6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_C_CY;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_C_XOR;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_D;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_D1;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_D2;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_D3;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_D4;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_D5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_D6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_DO5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_DO6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_D_CY;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_D_XOR;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_A;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_A1;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_A2;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_A3;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_A4;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_A5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_A6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_AMUX;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_AO5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_AO6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_A_CY;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_A_XOR;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_B;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_B1;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_B2;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_B3;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_B4;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_B5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_B6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_BO5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_BO6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_BQ;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_B_CY;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_B_XOR;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_C;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_C1;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_C2;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_C3;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_C4;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_C5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_C6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_CLK;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_CO5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_CO6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_CQ;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_C_CY;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_C_XOR;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_D;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_D1;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_D2;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_D3;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_D4;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_D5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_D6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_DMUX;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_DO5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_DO6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_D_CY;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_D_XOR;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_A;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_A1;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_A2;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_A3;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_A4;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_A5;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_A6;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_AO5;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_AO6;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_AQ;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_A_CY;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_A_XOR;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_B;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_B1;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_B2;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_B3;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_B4;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_B5;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_B6;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_BO5;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_BO6;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_BQ;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_B_CY;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_B_XOR;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_C;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_C1;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_C2;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_C3;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_C4;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_C5;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_C6;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_CLK;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_CO5;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_CO6;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_CQ;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_C_CY;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_C_XOR;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_D;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_D1;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_D2;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_D3;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_D4;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_D5;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_D5Q;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_D6;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_DMUX;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_DO5;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_DO6;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_DQ;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_D_CY;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_D_XOR;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_A;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_A1;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_A2;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_A3;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_A4;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_A5;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_A5Q;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_A6;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_AMUX;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_AO5;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_AO6;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_AQ;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_AX;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_A_CY;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_A_XOR;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_B;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_B1;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_B2;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_B3;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_B4;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_B5;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_B6;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_BMUX;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_BO5;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_BO6;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_B_CY;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_B_XOR;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_C;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_C1;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_C2;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_C3;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_C4;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_C5;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_C6;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_CLK;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_CMUX;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_CO5;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_CO6;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_C_CY;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_C_XOR;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_D;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_D1;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_D2;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_D3;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_D4;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_D5;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_D6;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_DO5;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_DO6;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_D_CY;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_D_XOR;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_A;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_A1;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_A2;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_A3;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_A4;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_A5;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_A6;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_AO5;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_AO6;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_AQ;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_A_CY;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_A_XOR;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_B;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_B1;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_B2;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_B3;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_B4;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_B5;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_B6;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_BO5;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_BO6;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_BQ;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_B_CY;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_B_XOR;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_C;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_C1;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_C2;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_C3;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_C4;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_C5;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_C6;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_CLK;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_CO5;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_CO6;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_CQ;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_C_CY;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_C_XOR;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_D;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_D1;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_D2;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_D3;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_D4;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_D5;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_D5Q;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_D6;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_DMUX;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_DO5;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_DO6;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_DQ;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_D_CY;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_D_XOR;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_A;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_A1;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_A2;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_A3;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_A4;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_A5;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_A6;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_AO5;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_AO6;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_AQ;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_A_CY;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_A_XOR;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_B;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_B1;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_B2;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_B3;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_B4;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_B5;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_B6;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_BO5;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_BO6;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_BQ;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_B_CY;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_B_XOR;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_C;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_C1;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_C2;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_C3;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_C4;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_C5;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_C6;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_CLK;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_CO5;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_CO6;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_CQ;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_C_CY;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_C_XOR;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_D;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_D1;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_D2;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_D3;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_D4;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_D5;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_D6;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_DMUX;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_DO5;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_DO6;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_D_CY;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_D_XOR;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_A;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_A1;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_A2;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_A3;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_A4;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_A5;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_A6;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_AO5;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_AO6;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_AQ;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_A_CY;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_A_XOR;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_B;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_B1;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_B2;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_B3;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_B4;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_B5;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_B6;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_BO5;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_BO6;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_BQ;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_B_CY;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_B_XOR;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_C;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_C1;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_C2;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_C3;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_C4;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_C5;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_C6;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_CLK;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_CO5;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_CO6;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_CQ;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_C_CY;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_C_XOR;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_D;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_D1;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_D2;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_D3;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_D4;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_D5;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_D6;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_DO5;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_DO6;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_D_CY;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_D_XOR;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_A;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_A1;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_A2;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_A3;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_A4;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_A5;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_A6;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_AO5;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_AO6;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_AQ;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_A_CY;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_A_XOR;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_B;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_B1;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_B2;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_B3;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_B4;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_B5;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_B5Q;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_B6;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_BMUX;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_BO5;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_BO6;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_BQ;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_B_CY;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_B_XOR;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_C;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_C1;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_C2;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_C3;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_C4;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_C5;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_C5Q;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_C6;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_CLK;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_CMUX;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_CO5;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_CO6;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_CQ;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_C_CY;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_C_XOR;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_D;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_D1;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_D2;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_D3;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_D4;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_D5;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_D6;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_DO5;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_DO6;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_D_CY;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_D_XOR;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_A;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_A1;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_A2;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_A3;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_A4;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_A5;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_A6;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_AO5;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_AO6;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_AQ;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_A_CY;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_A_XOR;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_B;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_B1;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_B2;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_B3;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_B4;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_B5;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_B6;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_BO5;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_BO6;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_BQ;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_B_CY;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_B_XOR;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_C;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_C1;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_C2;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_C3;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_C4;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_C5;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_C6;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_CLK;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_CO5;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_CO6;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_CQ;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_C_CY;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_C_XOR;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_D;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_D1;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_D2;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_D3;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_D4;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_D5;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_D6;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_DMUX;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_DO5;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_DO6;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_D_CY;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_D_XOR;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_A;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_A1;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_A2;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_A3;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_A4;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_A5;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_A6;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_AO5;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_AO6;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_AQ;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_A_CY;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_A_XOR;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_B;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_B1;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_B2;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_B3;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_B4;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_B5;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_B6;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_BO5;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_BO6;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_BQ;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_B_CY;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_B_XOR;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_C;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_C1;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_C2;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_C3;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_C4;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_C5;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_C6;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_CLK;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_CO5;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_CO6;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_CQ;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_C_CY;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_C_XOR;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_D;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_D1;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_D2;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_D3;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_D4;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_D5;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_D6;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_DO5;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_DO6;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_D_CY;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_D_XOR;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_A;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_A1;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_A2;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_A3;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_A4;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_A5;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_A6;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_AO5;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_AO6;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_AQ;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_A_CY;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_A_XOR;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_B;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_B1;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_B2;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_B3;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_B4;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_B5;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_B6;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_BO5;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_BO6;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_BQ;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_B_CY;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_B_XOR;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_C;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_C1;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_C2;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_C3;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_C4;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_C5;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_C6;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_CLK;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_CO5;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_CO6;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_C_CY;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_C_XOR;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_D;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_D1;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_D2;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_D3;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_D4;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_D5;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_D6;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_DO5;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_DO6;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_D_CY;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_D_XOR;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_A;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_A1;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_A2;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_A3;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_A4;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_A5;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_A6;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_AO5;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_AO6;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_AQ;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_A_CY;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_A_XOR;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_B;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_B1;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_B2;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_B3;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_B4;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_B5;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_B6;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_BO5;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_BO6;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_BQ;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_B_CY;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_B_XOR;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_C;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_C1;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_C2;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_C3;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_C4;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_C5;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_C6;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_CLK;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_CO5;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_CO6;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_CQ;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_C_CY;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_C_XOR;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_D;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_D1;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_D2;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_D3;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_D4;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_D5;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_D6;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_DO5;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_DO6;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_D_CY;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_D_XOR;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_A;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_A1;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_A2;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_A3;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_A4;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_A5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_A6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_AO5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_AO6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_A_CY;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_A_XOR;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_B;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_B1;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_B2;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_B3;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_B4;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_B5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_B6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_BO5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_BO6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_B_CY;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_B_XOR;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_C;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_C1;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_C2;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_C3;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_C4;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_C5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_C6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_CMUX;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_CO5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_CO6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_C_CY;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_C_XOR;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_D;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_D1;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_D2;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_D3;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_D4;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_D5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_D6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_DO5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_DO6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_D_CY;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_D_XOR;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_A;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_A1;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_A2;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_A3;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_A4;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_A5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_A6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_AO5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_AO6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_AQ;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_A_CY;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_A_XOR;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_B;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_B1;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_B2;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_B3;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_B4;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_B5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_B6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_BO5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_BO6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_BQ;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_B_CY;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_B_XOR;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_C;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_C1;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_C2;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_C3;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_C4;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_C5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_C6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_CLK;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_CMUX;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_CO5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_CO6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_C_CY;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_C_XOR;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_D;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_D1;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_D2;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_D3;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_D4;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_D5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_D6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_DO5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_DO6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_D_CY;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_D_XOR;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_A;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_A1;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_A2;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_A3;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_A4;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_A5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_A5Q;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_A6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_AMUX;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_AO5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_AO6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_AQ;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_AX;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_A_CY;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_A_XOR;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_B;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_B1;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_B2;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_B3;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_B4;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_B5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_B6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_BO5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_BO6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_BQ;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_B_CY;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_B_XOR;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_C;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_C1;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_C2;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_C3;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_C4;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_C5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_C6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_CLK;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_CO5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_CO6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_CQ;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_C_CY;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_C_XOR;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_D;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_D1;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_D2;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_D3;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_D4;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_D5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_D6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_DO5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_DO6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_D_CY;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_D_XOR;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_A;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_A1;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_A2;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_A3;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_A4;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_A5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_A6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_AO5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_AO6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_AQ;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_A_CY;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_A_XOR;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_B;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_B1;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_B2;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_B3;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_B4;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_B5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_B6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_BO5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_BO6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_BQ;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_B_CY;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_B_XOR;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_C;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_C1;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_C2;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_C3;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_C4;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_C5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_C6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_CLK;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_CO5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_CO6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_C_CY;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_C_XOR;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_D;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_D1;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_D2;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_D3;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_D4;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_D5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_D6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_DO5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_DO6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_D_CY;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_D_XOR;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_A;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_A1;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_A2;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_A3;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_A4;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_A5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_A6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_AO5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_AO6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_A_CY;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_A_XOR;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_B;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_B1;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_B2;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_B3;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_B4;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_B5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_B6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_BO5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_BO6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_B_CY;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_B_XOR;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_C;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_C1;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_C2;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_C3;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_C4;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_C5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_C6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_CO5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_CO6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_C_CY;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_C_XOR;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_D;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_D1;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_D2;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_D3;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_D4;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_D5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_D6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_DO5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_DO6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_D_CY;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_D_XOR;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_A;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_A1;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_A2;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_A3;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_A4;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_A5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_A6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_AO5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_AO6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_A_CY;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_A_XOR;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_B;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_B1;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_B2;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_B3;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_B4;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_B5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_B6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_BO5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_BO6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_B_CY;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_B_XOR;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_C;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_C1;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_C2;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_C3;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_C4;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_C5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_C6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_CO5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_CO6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_C_CY;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_C_XOR;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_D;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_D1;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_D2;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_D3;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_D4;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_D5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_D6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_DO5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_DO6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_D_CY;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_D_XOR;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_A;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_A1;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_A2;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_A3;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_A4;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_A5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_A6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_AMUX;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_AO5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_AO6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_A_CY;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_A_XOR;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_B;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_B1;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_B2;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_B3;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_B4;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_B5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_B6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_BMUX;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_BO5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_BO6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_B_CY;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_B_XOR;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_C;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_C1;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_C2;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_C3;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_C4;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_C5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_C6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_CO5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_CO6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_C_CY;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_C_XOR;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_D;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_D1;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_D2;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_D3;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_D4;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_D5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_D6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_DO5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_DO6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_D_CY;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_D_XOR;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_A;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_A1;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_A2;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_A3;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_A4;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_A5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_A6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_AO5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_AO6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_A_CY;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_A_XOR;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_B;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_B1;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_B2;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_B3;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_B4;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_B5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_B6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_BO5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_BO6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_B_CY;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_B_XOR;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_C;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_C1;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_C2;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_C3;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_C4;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_C5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_C6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_CO5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_CO6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_C_CY;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_C_XOR;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_D;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_D1;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_D2;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_D3;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_D4;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_D5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_D6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_DO5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_DO6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_D_CY;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_D_XOR;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_A;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_A1;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_A2;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_A3;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_A4;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_A5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_A6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_AO5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_AO6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_A_CY;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_A_XOR;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_B;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_B1;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_B2;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_B3;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_B4;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_B5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_B6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_BO5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_BO6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_B_CY;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_B_XOR;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_C;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_C1;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_C2;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_C3;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_C4;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_C5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_C6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_CO5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_CO6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_C_CY;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_C_XOR;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_D;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_D1;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_D2;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_D3;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_D4;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_D5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_D6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_DO5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_DO6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_D_CY;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_D_XOR;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_A;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_A1;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_A2;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_A3;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_A4;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_A5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_A6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_AMUX;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_AO5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_AO6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_AQ;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_A_CY;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_A_XOR;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_B;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_B1;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_B2;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_B3;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_B4;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_B5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_B6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_BO5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_BO6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_BQ;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_B_CY;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_B_XOR;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_C;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_C1;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_C2;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_C3;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_C4;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_C5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_C6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_CLK;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_CO5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_CO6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_C_CY;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_C_XOR;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_D;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_D1;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_D2;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_D3;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_D4;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_D5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_D6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_DO5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_DO6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_D_CY;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_D_XOR;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_A;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_A1;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_A2;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_A3;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_A4;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_A5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_A6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_AMUX;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_AO5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_AO6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_AQ;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_A_CY;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_A_XOR;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_B;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_B1;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_B2;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_B3;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_B4;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_B5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_B6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_BO5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_BO6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_BQ;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_B_CY;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_B_XOR;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_C;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_C1;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_C2;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_C3;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_C4;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_C5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_C6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_CLK;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_CO5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_CO6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_CQ;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_C_CY;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_C_XOR;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_D;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_D1;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_D2;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_D3;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_D4;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_D5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_D6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_DO5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_DO6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_D_CY;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_D_XOR;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_A;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_A1;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_A2;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_A3;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_A4;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_A5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_A6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_AO5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_AO6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_AQ;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_A_CY;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_A_XOR;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_B;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_B1;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_B2;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_B3;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_B4;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_B5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_B6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_BO5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_BO6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_BQ;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_B_CY;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_B_XOR;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_C;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_C1;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_C2;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_C3;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_C4;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_C5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_C6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_CLK;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_CO5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_CO6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_CQ;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_C_CY;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_C_XOR;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_D;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_D1;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_D2;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_D3;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_D4;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_D5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_D5Q;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_D6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_DMUX;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_DO5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_DO6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_DQ;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_D_CY;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_D_XOR;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_A;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_A1;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_A2;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_A3;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_A4;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_A5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_A6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_AO5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_AO6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_AQ;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_A_CY;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_A_XOR;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_B;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_B1;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_B2;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_B3;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_B4;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_B5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_B6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_BO5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_BO6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_BQ;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_B_CY;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_B_XOR;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_C;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_C1;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_C2;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_C3;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_C4;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_C5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_C6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_CLK;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_CO5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_CO6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_CQ;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_C_CY;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_C_XOR;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_D;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_D1;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_D2;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_D3;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_D4;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_D5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_D6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_DO5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_DO6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_D_CY;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_D_XOR;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_A;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_A1;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_A2;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_A3;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_A4;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_A5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_A6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_AO5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_AO6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_AQ;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_A_CY;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_A_XOR;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_B;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_B1;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_B2;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_B3;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_B4;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_B5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_B6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_BO5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_BO6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_BQ;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_B_CY;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_B_XOR;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_C;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_C1;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_C2;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_C3;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_C4;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_C5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_C6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_CLK;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_CO5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_CO6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_CQ;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_C_CY;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_C_XOR;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_D;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_D1;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_D2;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_D3;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_D4;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_D5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_D6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_DO5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_DO6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_D_CY;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_D_XOR;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_A;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_A1;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_A2;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_A3;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_A4;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_A5;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_A6;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_AO5;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_AO6;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_AQ;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_A_CY;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_A_XOR;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_B;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_B1;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_B2;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_B3;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_B4;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_B5;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_B6;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_BO5;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_BO6;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_BQ;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_B_CY;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_B_XOR;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_C;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_C1;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_C2;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_C3;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_C4;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_C5;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_C5Q;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_C6;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_CLK;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_CMUX;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_CO5;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_CO6;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_CQ;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_C_CY;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_C_XOR;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_D;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_D1;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_D2;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_D3;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_D4;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_D5;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_D6;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_DMUX;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_DO5;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_DO6;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_D_CY;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_D_XOR;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_A;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_A1;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_A2;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_A3;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_A4;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_A5;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_A6;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_AO5;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_AO6;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_AQ;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_A_CY;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_A_XOR;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_B;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_B1;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_B2;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_B3;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_B4;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_B5;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_B6;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_BO5;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_BO6;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_BQ;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_B_CY;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_B_XOR;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_C;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_C1;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_C2;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_C3;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_C4;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_C5;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_C6;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_CLK;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_CO5;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_CO6;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_C_CY;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_C_XOR;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_D;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_D1;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_D2;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_D3;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_D4;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_D5;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_D6;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_DO5;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_DO6;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_D_CY;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_D_XOR;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_A;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_A1;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_A2;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_A3;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_A4;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_A5;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_A6;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_AO5;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_AO6;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_AQ;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_A_CY;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_A_XOR;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_B;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_B1;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_B2;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_B3;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_B4;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_B5;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_B6;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_BO5;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_BO6;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_BQ;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_B_CY;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_B_XOR;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_C;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_C1;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_C2;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_C3;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_C4;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_C5;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_C6;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_CLK;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_CO5;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_CO6;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_CQ;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_C_CY;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_C_XOR;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_D;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_D1;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_D2;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_D3;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_D4;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_D5;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_D6;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_DMUX;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_DO5;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_DO6;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_D_CY;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_D_XOR;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_A;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_A1;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_A2;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_A3;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_A4;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_A5;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_A5Q;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_A6;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_AMUX;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_AO5;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_AO6;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_AQ;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_AX;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_A_CY;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_A_XOR;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_B;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_B1;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_B2;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_B3;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_B4;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_B5;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_B5Q;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_B6;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_BMUX;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_BO5;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_BO6;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_BQ;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_BX;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_B_CY;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_B_XOR;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_C;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_C1;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_C2;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_C3;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_C4;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_C5;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_C6;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_CLK;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_CMUX;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_CO5;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_CO6;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_C_CY;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_C_XOR;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_D;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_D1;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_D2;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_D3;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_D4;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_D5;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_D6;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_DO5;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_DO6;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_D_CY;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_D_XOR;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_A;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_A1;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_A2;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_A3;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_A4;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_A5;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_A6;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_AO5;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_AO6;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_AQ;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_A_CY;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_A_XOR;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_B;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_B1;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_B2;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_B3;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_B4;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_B5;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_B6;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_BO5;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_BO6;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_BQ;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_B_CY;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_B_XOR;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_C;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_C1;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_C2;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_C3;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_C4;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_C5;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_C6;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_CLK;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_CO5;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_CO6;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_CQ;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_C_CY;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_C_XOR;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_D;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_D1;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_D2;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_D3;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_D4;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_D5;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_D6;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_DMUX;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_DO5;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_DO6;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_D_CY;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_D_XOR;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_A;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_A1;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_A2;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_A3;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_A4;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_A5;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_A6;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_AO5;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_AO6;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_AQ;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_A_CY;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_A_XOR;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_B;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_B1;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_B2;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_B3;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_B4;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_B5;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_B6;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_BMUX;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_BO5;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_BO6;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_B_CY;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_B_XOR;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_C;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_C1;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_C2;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_C3;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_C4;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_C5;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_C6;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_CLK;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_CO5;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_CO6;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_CQ;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_C_CY;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_C_XOR;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_D;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_D1;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_D2;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_D3;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_D4;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_D5;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_D6;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_DO5;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_DO6;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_D_CY;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_D_XOR;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_A;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_A1;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_A2;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_A3;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_A4;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_A5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_A6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_AO5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_AO6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_AQ;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_A_CY;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_A_XOR;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_B;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_B1;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_B2;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_B3;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_B4;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_B5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_B6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_BO5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_BO6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_BQ;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_B_CY;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_B_XOR;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_C;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_C1;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_C2;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_C3;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_C4;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_C5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_C6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_CLK;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_CO5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_CO6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_CQ;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_C_CY;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_C_XOR;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_D;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_D1;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_D2;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_D3;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_D4;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_D5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_D6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_DMUX;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_DO5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_DO6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_D_CY;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_D_XOR;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_A;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_A1;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_A2;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_A3;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_A4;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_A5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_A6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_AO5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_AO6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_AQ;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_A_CY;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_A_XOR;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_B;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_B1;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_B2;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_B3;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_B4;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_B5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_B6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_BO5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_BO6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_BQ;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_B_CY;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_B_XOR;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_C;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_C1;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_C2;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_C3;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_C4;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_C5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_C6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_CLK;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_CO5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_CO6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_C_CY;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_C_XOR;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_D;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_D1;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_D2;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_D3;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_D4;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_D5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_D6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_DO5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_DO6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_D_CY;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_D_XOR;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_A;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_A1;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_A2;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_A3;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_A4;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_A5;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_A6;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_AO5;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_AO6;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_AQ;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_A_CY;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_A_XOR;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_B;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_B1;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_B2;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_B3;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_B4;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_B5;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_B6;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_BO5;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_BO6;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_BQ;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_B_CY;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_B_XOR;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_C;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_C1;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_C2;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_C3;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_C4;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_C5;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_C6;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_CLK;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_CO5;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_CO6;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_CQ;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_C_CY;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_C_XOR;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_D;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_D1;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_D2;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_D3;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_D4;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_D5;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_D6;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_DO5;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_DO6;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_D_CY;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_D_XOR;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_A;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_A1;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_A2;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_A3;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_A4;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_A5;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_A6;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_AO5;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_AO6;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_AQ;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_A_CY;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_A_XOR;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_B;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_B1;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_B2;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_B3;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_B4;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_B5;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_B6;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_BO5;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_BO6;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_B_CY;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_B_XOR;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_C;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_C1;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_C2;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_C3;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_C4;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_C5;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_C6;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_CLK;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_CO5;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_CO6;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_C_CY;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_C_XOR;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_D;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_D1;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_D2;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_D3;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_D4;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_D5;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_D6;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_DO5;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_DO6;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_D_CY;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_D_XOR;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_A;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_A1;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_A2;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_A3;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_A4;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_A5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_A5Q;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_A6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_AMUX;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_AO5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_AO6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_AQ;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_AX;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_A_CY;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_A_XOR;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_B;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_B1;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_B2;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_B3;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_B4;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_B5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_B6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_BO5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_BO6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_BQ;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_B_CY;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_B_XOR;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_C;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_C1;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_C2;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_C3;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_C4;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_C5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_C6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_CLK;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_CMUX;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_CO5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_CO6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_C_CY;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_C_XOR;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_D;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_D1;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_D2;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_D3;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_D4;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_D5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_D6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_DMUX;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_DO5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_DO6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_D_CY;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_D_XOR;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_A;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_A1;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_A2;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_A3;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_A4;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_A5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_A5Q;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_A6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_AMUX;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_AO5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_AO6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_AQ;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_A_CY;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_A_XOR;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_B;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_B1;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_B2;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_B3;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_B4;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_B5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_B6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_BMUX;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_BO5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_BO6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_B_CY;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_B_XOR;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_C;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_C1;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_C2;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_C3;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_C4;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_C5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_C6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_CLK;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_CO5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_CO6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_C_CY;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_C_XOR;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_D;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_D1;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_D2;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_D3;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_D4;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_D5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_D6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_DO5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_DO6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_D_CY;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_D_XOR;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_A;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_A1;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_A2;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_A3;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_A4;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_A5;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_A6;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_AO5;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_AO6;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_AQ;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_A_CY;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_A_XOR;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_B;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_B1;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_B2;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_B3;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_B4;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_B5;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_B6;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_BMUX;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_BO5;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_BO6;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_B_CY;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_B_XOR;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_C;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_C1;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_C2;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_C3;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_C4;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_C5;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_C6;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_CLK;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_CO5;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_CO6;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_C_CY;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_C_XOR;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_D;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_D1;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_D2;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_D3;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_D4;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_D5;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_D6;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_DO5;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_DO6;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_D_CY;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_D_XOR;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_A;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_A1;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_A2;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_A3;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_A4;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_A5;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_A6;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_AO5;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_AO6;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_AQ;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_A_CY;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_A_XOR;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_B;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_B1;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_B2;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_B3;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_B4;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_B5;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_B6;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_BO5;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_BO6;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_BQ;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_B_CY;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_B_XOR;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_C;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_C1;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_C2;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_C3;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_C4;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_C5;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_C6;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_CLK;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_CO5;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_CO6;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_CQ;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_C_CY;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_C_XOR;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_D;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_D1;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_D2;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_D3;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_D4;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_D5;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_D6;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_DO5;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_DO6;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_D_CY;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_D_XOR;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_A;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_A1;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_A2;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_A3;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_A4;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_A5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_A6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_AO5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_AO6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_AQ;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_A_CY;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_A_XOR;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_B;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_B1;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_B2;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_B3;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_B4;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_B5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_B6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_BMUX;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_BO5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_BO6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_B_CY;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_B_XOR;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_C;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_C1;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_C2;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_C3;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_C4;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_C5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_C6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_CLK;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_CO5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_CO6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_C_CY;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_C_XOR;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_D;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_D1;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_D2;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_D3;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_D4;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_D5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_D6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_DO5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_DO6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_D_CY;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_D_XOR;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_A;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_A1;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_A2;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_A3;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_A4;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_A5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_A6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_AO5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_AO6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_AQ;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_A_CY;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_A_XOR;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_B;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_B1;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_B2;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_B3;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_B4;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_B5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_B6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_BO5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_BO6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_BQ;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_B_CY;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_B_XOR;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_C;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_C1;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_C2;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_C3;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_C4;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_C5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_C6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_CLK;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_CO5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_CO6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_C_CY;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_C_XOR;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_D;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_D1;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_D2;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_D3;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_D4;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_D5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_D6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_DO5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_DO6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_D_CY;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_D_XOR;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_A;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_A1;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_A2;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_A3;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_A4;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_A5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_A6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_AO5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_AO6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_AQ;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_A_CY;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_A_XOR;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_B;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_B1;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_B2;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_B3;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_B4;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_B5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_B6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_BO5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_BO6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_B_CY;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_B_XOR;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_C;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_C1;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_C2;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_C3;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_C4;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_C5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_C6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_CLK;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_CO5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_CO6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_C_CY;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_C_XOR;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_D;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_D1;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_D2;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_D3;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_D4;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_D5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_D6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_DO5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_DO6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_D_CY;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_D_XOR;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_A;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_A1;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_A2;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_A3;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_A4;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_A5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_A6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_AO5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_AO6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_AQ;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_A_CY;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_A_XOR;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_B;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_B1;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_B2;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_B3;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_B4;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_B5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_B6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_BO5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_BO6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_BQ;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_B_CY;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_B_XOR;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_C;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_C1;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_C2;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_C3;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_C4;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_C5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_C6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_CLK;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_CMUX;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_CO5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_CO6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_C_CY;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_C_XOR;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_D;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_D1;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_D2;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_D3;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_D4;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_D5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_D6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_DMUX;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_DO5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_DO6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_D_CY;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_D_XOR;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_A;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_A1;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_A2;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_A3;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_A4;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_A5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_A5Q;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_A6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_AMUX;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_AO5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_AO6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_AQ;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_AX;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_A_CY;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_A_XOR;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_B;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_B1;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_B2;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_B3;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_B4;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_B5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_B6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_BMUX;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_BO5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_BO6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_B_CY;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_B_XOR;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_C;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_C1;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_C2;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_C3;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_C4;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_C5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_C6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_CLK;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_CO5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_CO6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_CQ;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_C_CY;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_C_XOR;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_D;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_D1;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_D2;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_D3;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_D4;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_D5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_D6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_DO5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_DO6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_D_CY;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_D_XOR;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_A;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_A1;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_A2;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_A3;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_A4;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_A5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_A6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_AO5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_AO6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_AQ;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_A_CY;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_A_XOR;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_B;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_B1;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_B2;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_B3;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_B4;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_B5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_B6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_BO5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_BO6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_BQ;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_B_CY;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_B_XOR;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_C;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_C1;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_C2;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_C3;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_C4;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_C5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_C6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_CLK;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_CO5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_CO6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_CQ;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_C_CY;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_C_XOR;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_D;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_D1;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_D2;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_D3;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_D4;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_D5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_D6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_DO5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_DO6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_D_CY;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_D_XOR;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_A;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_A1;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_A2;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_A3;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_A4;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_A5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_A6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_AO5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_AO6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_AQ;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_A_CY;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_A_XOR;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_B;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_B1;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_B2;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_B3;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_B4;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_B5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_B6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_BO5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_BO6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_BQ;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_B_CY;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_B_XOR;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_C;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_C1;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_C2;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_C3;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_C4;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_C5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_C6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_CLK;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_CO5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_CO6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_CQ;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_C_CY;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_C_XOR;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_D;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_D1;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_D2;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_D3;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_D4;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_D5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_D6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_DO5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_DO6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_D_CY;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_D_XOR;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_A;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_A1;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_A2;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_A3;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_A4;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_A5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_A6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_AO5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_AO6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_AQ;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_A_CY;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_A_XOR;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_B;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_B1;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_B2;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_B3;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_B4;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_B5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_B6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_BO5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_BO6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_B_CY;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_B_XOR;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_C;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_C1;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_C2;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_C3;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_C4;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_C5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_C6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_CLK;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_CO5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_CO6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_C_CY;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_C_XOR;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_D;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_D1;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_D2;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_D3;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_D4;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_D5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_D6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_DO5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_DO6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_D_CY;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_D_XOR;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_A;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_A1;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_A2;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_A3;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_A4;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_A5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_A6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_AO5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_AO6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_AX;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_A_CY;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_A_XOR;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_B;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_B1;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_B2;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_B3;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_B4;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_B5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_B6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_BO5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_BO6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_B_CY;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_B_XOR;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_C;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_C1;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_C2;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_C3;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_C4;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_C5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_C6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_CLK;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_CO5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_CO6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_C_CY;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_C_XOR;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_D;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_D1;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_D2;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_D3;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_D4;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_D5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_D6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_DO5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_DO6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_D_CY;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_D_XOR;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_A;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_A1;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_A2;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_A3;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_A4;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_A5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_A6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_AO5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_AO6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_A_CY;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_A_XOR;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_B;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_B1;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_B2;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_B3;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_B4;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_B5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_B6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_BO5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_BO6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_B_CY;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_B_XOR;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_C;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_C1;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_C2;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_C3;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_C4;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_C5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_C6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_CO5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_CO6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_C_CY;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_C_XOR;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_D;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_D1;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_D2;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_D3;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_D4;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_D5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_D6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_DO5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_DO6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_D_CY;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_D_XOR;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE1;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I1;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE1;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S1;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_CE;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_I;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  wire [0:0] LIOB33_SING_X0Y100_IOB_X0Y100_O;
  wire [0:0] LIOB33_SING_X0Y149_IOB_X0Y149_O;
  wire [0:0] LIOB33_SING_X0Y150_IOB_X0Y150_O;
  wire [0:0] LIOB33_SING_X0Y199_IOB_X0Y199_O;
  wire [0:0] LIOB33_SING_X0Y50_IOB_X0Y50_I;
  wire [0:0] LIOB33_X0Y101_IOB_X0Y101_O;
  wire [0:0] LIOB33_X0Y101_IOB_X0Y102_O;
  wire [0:0] LIOB33_X0Y103_IOB_X0Y103_O;
  wire [0:0] LIOB33_X0Y103_IOB_X0Y104_O;
  wire [0:0] LIOB33_X0Y105_IOB_X0Y105_O;
  wire [0:0] LIOB33_X0Y105_IOB_X0Y106_O;
  wire [0:0] LIOB33_X0Y107_IOB_X0Y107_O;
  wire [0:0] LIOB33_X0Y107_IOB_X0Y108_O;
  wire [0:0] LIOB33_X0Y109_IOB_X0Y109_O;
  wire [0:0] LIOB33_X0Y109_IOB_X0Y110_O;
  wire [0:0] LIOB33_X0Y111_IOB_X0Y111_O;
  wire [0:0] LIOB33_X0Y111_IOB_X0Y112_O;
  wire [0:0] LIOB33_X0Y113_IOB_X0Y113_O;
  wire [0:0] LIOB33_X0Y113_IOB_X0Y114_O;
  wire [0:0] LIOB33_X0Y115_IOB_X0Y115_O;
  wire [0:0] LIOB33_X0Y115_IOB_X0Y116_O;
  wire [0:0] LIOB33_X0Y117_IOB_X0Y117_O;
  wire [0:0] LIOB33_X0Y117_IOB_X0Y118_O;
  wire [0:0] LIOB33_X0Y119_IOB_X0Y119_O;
  wire [0:0] LIOB33_X0Y119_IOB_X0Y120_O;
  wire [0:0] LIOB33_X0Y121_IOB_X0Y121_O;
  wire [0:0] LIOB33_X0Y121_IOB_X0Y122_O;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y123_O;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y124_O;
  wire [0:0] LIOB33_X0Y125_IOB_X0Y125_O;
  wire [0:0] LIOB33_X0Y125_IOB_X0Y126_O;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y127_O;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y128_O;
  wire [0:0] LIOB33_X0Y129_IOB_X0Y129_O;
  wire [0:0] LIOB33_X0Y129_IOB_X0Y130_O;
  wire [0:0] LIOB33_X0Y131_IOB_X0Y131_O;
  wire [0:0] LIOB33_X0Y131_IOB_X0Y132_O;
  wire [0:0] LIOB33_X0Y133_IOB_X0Y133_O;
  wire [0:0] LIOB33_X0Y133_IOB_X0Y134_O;
  wire [0:0] LIOB33_X0Y135_IOB_X0Y135_O;
  wire [0:0] LIOB33_X0Y135_IOB_X0Y136_O;
  wire [0:0] LIOB33_X0Y137_IOB_X0Y137_O;
  wire [0:0] LIOB33_X0Y137_IOB_X0Y138_O;
  wire [0:0] LIOB33_X0Y139_IOB_X0Y139_O;
  wire [0:0] LIOB33_X0Y139_IOB_X0Y140_O;
  wire [0:0] LIOB33_X0Y141_IOB_X0Y141_O;
  wire [0:0] LIOB33_X0Y141_IOB_X0Y142_O;
  wire [0:0] LIOB33_X0Y143_IOB_X0Y143_O;
  wire [0:0] LIOB33_X0Y145_IOB_X0Y145_O;
  wire [0:0] LIOB33_X0Y145_IOB_X0Y146_O;
  wire [0:0] LIOB33_X0Y147_IOB_X0Y147_O;
  wire [0:0] LIOB33_X0Y147_IOB_X0Y148_O;
  wire [0:0] LIOB33_X0Y151_IOB_X0Y151_O;
  wire [0:0] LIOB33_X0Y151_IOB_X0Y152_O;
  wire [0:0] LIOB33_X0Y153_IOB_X0Y153_O;
  wire [0:0] LIOB33_X0Y153_IOB_X0Y154_O;
  wire [0:0] LIOB33_X0Y155_IOB_X0Y155_O;
  wire [0:0] LIOB33_X0Y155_IOB_X0Y156_O;
  wire [0:0] LIOB33_X0Y157_IOB_X0Y157_O;
  wire [0:0] LIOB33_X0Y157_IOB_X0Y158_O;
  wire [0:0] LIOB33_X0Y159_IOB_X0Y159_O;
  wire [0:0] LIOB33_X0Y159_IOB_X0Y160_O;
  wire [0:0] LIOB33_X0Y161_IOB_X0Y161_O;
  wire [0:0] LIOB33_X0Y161_IOB_X0Y162_O;
  wire [0:0] LIOB33_X0Y163_IOB_X0Y163_O;
  wire [0:0] LIOB33_X0Y163_IOB_X0Y164_O;
  wire [0:0] LIOB33_X0Y165_IOB_X0Y165_O;
  wire [0:0] LIOB33_X0Y165_IOB_X0Y166_O;
  wire [0:0] LIOB33_X0Y167_IOB_X0Y167_O;
  wire [0:0] LIOB33_X0Y167_IOB_X0Y168_O;
  wire [0:0] LIOB33_X0Y169_IOB_X0Y169_O;
  wire [0:0] LIOB33_X0Y169_IOB_X0Y170_O;
  wire [0:0] LIOB33_X0Y171_IOB_X0Y171_O;
  wire [0:0] LIOB33_X0Y171_IOB_X0Y172_O;
  wire [0:0] LIOB33_X0Y173_IOB_X0Y173_O;
  wire [0:0] LIOB33_X0Y173_IOB_X0Y174_O;
  wire [0:0] LIOB33_X0Y175_IOB_X0Y175_O;
  wire [0:0] LIOB33_X0Y175_IOB_X0Y176_O;
  wire [0:0] LIOB33_X0Y177_IOB_X0Y177_O;
  wire [0:0] LIOB33_X0Y177_IOB_X0Y178_O;
  wire [0:0] LIOB33_X0Y179_IOB_X0Y179_O;
  wire [0:0] LIOB33_X0Y179_IOB_X0Y180_O;
  wire [0:0] LIOB33_X0Y181_IOB_X0Y181_O;
  wire [0:0] LIOB33_X0Y181_IOB_X0Y182_O;
  wire [0:0] LIOB33_X0Y183_IOB_X0Y183_O;
  wire [0:0] LIOB33_X0Y183_IOB_X0Y184_O;
  wire [0:0] LIOB33_X0Y185_IOB_X0Y185_O;
  wire [0:0] LIOB33_X0Y185_IOB_X0Y186_O;
  wire [0:0] LIOB33_X0Y187_IOB_X0Y187_O;
  wire [0:0] LIOB33_X0Y187_IOB_X0Y188_O;
  wire [0:0] LIOB33_X0Y189_IOB_X0Y189_O;
  wire [0:0] LIOB33_X0Y189_IOB_X0Y190_O;
  wire [0:0] LIOB33_X0Y191_IOB_X0Y191_O;
  wire [0:0] LIOB33_X0Y191_IOB_X0Y192_O;
  wire [0:0] LIOB33_X0Y193_IOB_X0Y193_O;
  wire [0:0] LIOB33_X0Y193_IOB_X0Y194_O;
  wire [0:0] LIOB33_X0Y195_IOB_X0Y195_O;
  wire [0:0] LIOB33_X0Y195_IOB_X0Y196_O;
  wire [0:0] LIOB33_X0Y197_IOB_X0Y197_O;
  wire [0:0] LIOB33_X0Y197_IOB_X0Y198_O;
  wire [0:0] LIOB33_X0Y51_IOB_X0Y51_I;
  wire [0:0] LIOB33_X0Y51_IOB_X0Y52_I;
  wire [0:0] LIOB33_X0Y53_IOB_X0Y53_I;
  wire [0:0] LIOB33_X0Y53_IOB_X0Y54_I;
  wire [0:0] LIOB33_X0Y55_IOB_X0Y55_I;
  wire [0:0] LIOB33_X0Y55_IOB_X0Y56_I;
  wire [0:0] LIOB33_X0Y57_IOB_X0Y57_I;
  wire [0:0] LIOB33_X0Y57_IOB_X0Y58_I;
  wire [0:0] LIOB33_X0Y59_IOB_X0Y59_I;
  wire [0:0] LIOB33_X0Y59_IOB_X0Y60_I;
  wire [0:0] LIOB33_X0Y61_IOB_X0Y61_I;
  wire [0:0] LIOB33_X0Y61_IOB_X0Y62_I;
  wire [0:0] LIOB33_X0Y63_IOB_X0Y63_I;
  wire [0:0] LIOB33_X0Y63_IOB_X0Y64_I;
  wire [0:0] LIOB33_X0Y65_IOB_X0Y65_I;
  wire [0:0] LIOB33_X0Y65_IOB_X0Y66_I;
  wire [0:0] LIOB33_X0Y67_IOB_X0Y67_I;
  wire [0:0] LIOB33_X0Y67_IOB_X0Y68_I;
  wire [0:0] LIOB33_X0Y69_IOB_X0Y69_I;
  wire [0:0] LIOB33_X0Y69_IOB_X0Y70_I;
  wire [0:0] LIOB33_X0Y71_IOB_X0Y71_I;
  wire [0:0] LIOB33_X0Y71_IOB_X0Y72_I;
  wire [0:0] LIOB33_X0Y73_IOB_X0Y73_I;
  wire [0:0] LIOB33_X0Y73_IOB_X0Y74_I;
  wire [0:0] LIOB33_X0Y75_IOB_X0Y75_I;
  wire [0:0] LIOB33_X0Y75_IOB_X0Y76_I;
  wire [0:0] LIOB33_X0Y77_IOB_X0Y77_I;
  wire [0:0] LIOB33_X0Y77_IOB_X0Y78_I;
  wire [0:0] LIOB33_X0Y79_IOB_X0Y79_I;
  wire [0:0] LIOB33_X0Y79_IOB_X0Y80_O;
  wire [0:0] LIOI3_SING_X0Y100_OLOGIC_X0Y100_D1;
  wire [0:0] LIOI3_SING_X0Y100_OLOGIC_X0Y100_OQ;
  wire [0:0] LIOI3_SING_X0Y100_OLOGIC_X0Y100_T1;
  wire [0:0] LIOI3_SING_X0Y100_OLOGIC_X0Y100_TQ;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_D1;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_OQ;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_T1;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_TQ;
  wire [0:0] LIOI3_SING_X0Y150_OLOGIC_X0Y150_D1;
  wire [0:0] LIOI3_SING_X0Y150_OLOGIC_X0Y150_OQ;
  wire [0:0] LIOI3_SING_X0Y150_OLOGIC_X0Y150_T1;
  wire [0:0] LIOI3_SING_X0Y150_OLOGIC_X0Y150_TQ;
  wire [0:0] LIOI3_SING_X0Y199_OLOGIC_X0Y199_D1;
  wire [0:0] LIOI3_SING_X0Y199_OLOGIC_X0Y199_OQ;
  wire [0:0] LIOI3_SING_X0Y199_OLOGIC_X0Y199_T1;
  wire [0:0] LIOI3_SING_X0Y199_OLOGIC_X0Y199_TQ;
  wire [0:0] LIOI3_SING_X0Y50_ILOGIC_X0Y50_D;
  wire [0:0] LIOI3_SING_X0Y50_ILOGIC_X0Y50_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y57_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y57_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y58_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y58_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y69_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y69_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y70_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y70_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y63_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y63_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y64_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y64_O;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y101_D1;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y101_OQ;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y101_T1;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y101_TQ;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y102_D1;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y102_OQ;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y102_T1;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y102_TQ;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y103_D1;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y103_OQ;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y103_T1;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y103_TQ;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y104_D1;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y104_OQ;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y104_T1;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y104_TQ;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y105_D1;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y105_OQ;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y105_T1;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y105_TQ;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y106_D1;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y106_OQ;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y106_T1;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y106_TQ;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y109_D1;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y109_OQ;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y109_T1;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y109_TQ;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y110_D1;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y110_OQ;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y110_T1;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y110_TQ;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_D1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_OQ;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_T1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_TQ;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y112_D1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y112_OQ;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y112_T1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y112_TQ;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y115_D1;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y115_OQ;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y115_T1;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y115_TQ;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y116_D1;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y116_OQ;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y116_T1;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y116_TQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y117_D1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y117_OQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y117_T1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y117_TQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_D1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_OQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_T1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_TQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_D1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_OQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_T1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_TQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_D1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_OQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_T1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_TQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_D1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_OQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_T1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_TQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_D1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_OQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_T1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_TQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_D1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_OQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_T1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_TQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_D1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_OQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_T1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_TQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_D1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_OQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_T1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_TQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_D1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_OQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_T1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_TQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_D1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_OQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_T1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_TQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_D1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_OQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_T1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_TQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_D1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_OQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_T1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_TQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_D1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_OQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_T1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_TQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_D1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_OQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_T1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_TQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_D1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_OQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_T1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_TQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_D1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_OQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_T1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_TQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_D1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_OQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_T1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_TQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_D1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_OQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_T1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_TQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_D1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_OQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_T1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_TQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_D1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_OQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_T1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_TQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_D1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_OQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_T1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_TQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_D1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_OQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_T1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_TQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_D1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_OQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_T1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_TQ;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y151_D1;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y151_OQ;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y151_T1;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y151_TQ;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y152_D1;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y152_OQ;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y152_T1;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y152_TQ;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y153_D1;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y153_OQ;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y153_T1;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y153_TQ;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y154_D1;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y154_OQ;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y154_T1;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y154_TQ;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y155_D1;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y155_OQ;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y155_T1;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y155_TQ;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y156_D1;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y156_OQ;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y156_T1;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y156_TQ;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y159_D1;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y159_OQ;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y159_T1;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y159_TQ;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y160_D1;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y160_OQ;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y160_T1;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y160_TQ;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y161_D1;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y161_OQ;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y161_T1;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y161_TQ;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y162_D1;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y162_OQ;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y162_T1;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y162_TQ;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y165_D1;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y165_OQ;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y165_T1;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y165_TQ;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y166_D1;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y166_OQ;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y166_T1;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y166_TQ;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y167_D1;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y167_OQ;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y167_T1;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y167_TQ;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y168_D1;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y168_OQ;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y168_T1;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y168_TQ;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y171_D1;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y171_OQ;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y171_T1;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y171_TQ;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y172_D1;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y172_OQ;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y172_T1;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y172_TQ;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y173_D1;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y173_OQ;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y173_T1;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y173_TQ;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y174_D1;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y174_OQ;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y174_T1;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y174_TQ;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y175_D1;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y175_OQ;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y175_T1;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y175_TQ;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y176_D1;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y176_OQ;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y176_T1;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y176_TQ;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y177_D1;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y177_OQ;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y177_T1;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y177_TQ;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y178_D1;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y178_OQ;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y178_T1;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y178_TQ;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y179_D1;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y179_OQ;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y179_T1;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y179_TQ;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y180_D1;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y180_OQ;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y180_T1;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y180_TQ;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y183_D1;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y183_OQ;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y183_T1;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y183_TQ;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y184_D1;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y184_OQ;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y184_T1;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y184_TQ;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y185_D1;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y185_OQ;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y185_T1;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y185_TQ;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y186_D1;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y186_OQ;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y186_T1;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y186_TQ;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y189_D1;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y189_OQ;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y189_T1;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y189_TQ;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y190_D1;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y190_OQ;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y190_T1;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y190_TQ;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y191_D1;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y191_OQ;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y191_T1;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y191_TQ;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y192_D1;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y192_OQ;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y192_T1;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y192_TQ;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y195_D1;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y195_OQ;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y195_T1;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y195_TQ;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y196_D1;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y196_OQ;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y196_T1;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y196_TQ;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y197_D1;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y197_OQ;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y197_T1;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y197_TQ;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y198_D1;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y198_OQ;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y198_T1;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y198_TQ;
  wire [0:0] LIOI3_X0Y51_ILOGIC_X0Y51_D;
  wire [0:0] LIOI3_X0Y51_ILOGIC_X0Y51_O;
  wire [0:0] LIOI3_X0Y51_ILOGIC_X0Y52_D;
  wire [0:0] LIOI3_X0Y51_ILOGIC_X0Y52_O;
  wire [0:0] LIOI3_X0Y53_ILOGIC_X0Y53_D;
  wire [0:0] LIOI3_X0Y53_ILOGIC_X0Y53_O;
  wire [0:0] LIOI3_X0Y53_ILOGIC_X0Y54_D;
  wire [0:0] LIOI3_X0Y53_ILOGIC_X0Y54_O;
  wire [0:0] LIOI3_X0Y55_ILOGIC_X0Y55_D;
  wire [0:0] LIOI3_X0Y55_ILOGIC_X0Y55_O;
  wire [0:0] LIOI3_X0Y55_ILOGIC_X0Y56_D;
  wire [0:0] LIOI3_X0Y55_ILOGIC_X0Y56_O;
  wire [0:0] LIOI3_X0Y59_ILOGIC_X0Y59_D;
  wire [0:0] LIOI3_X0Y59_ILOGIC_X0Y59_O;
  wire [0:0] LIOI3_X0Y59_ILOGIC_X0Y60_D;
  wire [0:0] LIOI3_X0Y59_ILOGIC_X0Y60_O;
  wire [0:0] LIOI3_X0Y61_ILOGIC_X0Y61_D;
  wire [0:0] LIOI3_X0Y61_ILOGIC_X0Y61_O;
  wire [0:0] LIOI3_X0Y61_ILOGIC_X0Y62_D;
  wire [0:0] LIOI3_X0Y61_ILOGIC_X0Y62_O;
  wire [0:0] LIOI3_X0Y65_ILOGIC_X0Y65_D;
  wire [0:0] LIOI3_X0Y65_ILOGIC_X0Y65_O;
  wire [0:0] LIOI3_X0Y65_ILOGIC_X0Y66_D;
  wire [0:0] LIOI3_X0Y65_ILOGIC_X0Y66_O;
  wire [0:0] LIOI3_X0Y67_ILOGIC_X0Y67_D;
  wire [0:0] LIOI3_X0Y67_ILOGIC_X0Y67_O;
  wire [0:0] LIOI3_X0Y67_ILOGIC_X0Y68_D;
  wire [0:0] LIOI3_X0Y67_ILOGIC_X0Y68_O;
  wire [0:0] LIOI3_X0Y71_ILOGIC_X0Y71_D;
  wire [0:0] LIOI3_X0Y71_ILOGIC_X0Y71_O;
  wire [0:0] LIOI3_X0Y71_ILOGIC_X0Y72_D;
  wire [0:0] LIOI3_X0Y71_ILOGIC_X0Y72_O;
  wire [0:0] LIOI3_X0Y73_ILOGIC_X0Y73_D;
  wire [0:0] LIOI3_X0Y73_ILOGIC_X0Y73_O;
  wire [0:0] LIOI3_X0Y73_ILOGIC_X0Y74_D;
  wire [0:0] LIOI3_X0Y73_ILOGIC_X0Y74_O;
  wire [0:0] LIOI3_X0Y75_ILOGIC_X0Y75_D;
  wire [0:0] LIOI3_X0Y75_ILOGIC_X0Y75_O;
  wire [0:0] LIOI3_X0Y75_ILOGIC_X0Y76_D;
  wire [0:0] LIOI3_X0Y75_ILOGIC_X0Y76_O;
  wire [0:0] LIOI3_X0Y77_ILOGIC_X0Y77_D;
  wire [0:0] LIOI3_X0Y77_ILOGIC_X0Y77_O;
  wire [0:0] LIOI3_X0Y77_ILOGIC_X0Y78_D;
  wire [0:0] LIOI3_X0Y77_ILOGIC_X0Y78_O;
  wire [0:0] LIOI3_X0Y79_ILOGIC_X0Y79_D;
  wire [0:0] LIOI3_X0Y79_ILOGIC_X0Y79_O;
  wire [0:0] LIOI3_X0Y79_OLOGIC_X0Y80_D1;
  wire [0:0] LIOI3_X0Y79_OLOGIC_X0Y80_OQ;
  wire [0:0] LIOI3_X0Y79_OLOGIC_X0Y80_T1;
  wire [0:0] LIOI3_X0Y79_OLOGIC_X0Y80_TQ;
  wire [0:0] RIOB33_SING_X105Y100_IOB_X1Y100_I;
  wire [0:0] RIOB33_SING_X105Y149_IOB_X1Y149_I;
  wire [0:0] RIOB33_SING_X105Y150_IOB_X1Y150_O;
  wire [0:0] RIOB33_SING_X105Y199_IOB_X1Y199_O;
  wire [0:0] RIOB33_X105Y101_IOB_X1Y101_I;
  wire [0:0] RIOB33_X105Y101_IOB_X1Y102_I;
  wire [0:0] RIOB33_X105Y103_IOB_X1Y103_I;
  wire [0:0] RIOB33_X105Y103_IOB_X1Y104_I;
  wire [0:0] RIOB33_X105Y105_IOB_X1Y105_I;
  wire [0:0] RIOB33_X105Y105_IOB_X1Y106_I;
  wire [0:0] RIOB33_X105Y107_IOB_X1Y107_I;
  wire [0:0] RIOB33_X105Y107_IOB_X1Y108_I;
  wire [0:0] RIOB33_X105Y109_IOB_X1Y109_I;
  wire [0:0] RIOB33_X105Y109_IOB_X1Y110_I;
  wire [0:0] RIOB33_X105Y111_IOB_X1Y111_I;
  wire [0:0] RIOB33_X105Y111_IOB_X1Y112_I;
  wire [0:0] RIOB33_X105Y113_IOB_X1Y113_I;
  wire [0:0] RIOB33_X105Y113_IOB_X1Y114_I;
  wire [0:0] RIOB33_X105Y115_IOB_X1Y115_I;
  wire [0:0] RIOB33_X105Y115_IOB_X1Y116_I;
  wire [0:0] RIOB33_X105Y117_IOB_X1Y117_I;
  wire [0:0] RIOB33_X105Y117_IOB_X1Y118_I;
  wire [0:0] RIOB33_X105Y119_IOB_X1Y119_I;
  wire [0:0] RIOB33_X105Y119_IOB_X1Y120_I;
  wire [0:0] RIOB33_X105Y121_IOB_X1Y121_I;
  wire [0:0] RIOB33_X105Y121_IOB_X1Y122_I;
  wire [0:0] RIOB33_X105Y123_IOB_X1Y123_I;
  wire [0:0] RIOB33_X105Y123_IOB_X1Y124_I;
  wire [0:0] RIOB33_X105Y125_IOB_X1Y125_I;
  wire [0:0] RIOB33_X105Y125_IOB_X1Y126_I;
  wire [0:0] RIOB33_X105Y127_IOB_X1Y127_I;
  wire [0:0] RIOB33_X105Y127_IOB_X1Y128_I;
  wire [0:0] RIOB33_X105Y129_IOB_X1Y129_I;
  wire [0:0] RIOB33_X105Y129_IOB_X1Y130_I;
  wire [0:0] RIOB33_X105Y131_IOB_X1Y131_I;
  wire [0:0] RIOB33_X105Y131_IOB_X1Y132_I;
  wire [0:0] RIOB33_X105Y133_IOB_X1Y133_I;
  wire [0:0] RIOB33_X105Y133_IOB_X1Y134_I;
  wire [0:0] RIOB33_X105Y135_IOB_X1Y135_I;
  wire [0:0] RIOB33_X105Y135_IOB_X1Y136_I;
  wire [0:0] RIOB33_X105Y137_IOB_X1Y137_I;
  wire [0:0] RIOB33_X105Y137_IOB_X1Y138_I;
  wire [0:0] RIOB33_X105Y139_IOB_X1Y139_I;
  wire [0:0] RIOB33_X105Y139_IOB_X1Y140_I;
  wire [0:0] RIOB33_X105Y141_IOB_X1Y141_I;
  wire [0:0] RIOB33_X105Y141_IOB_X1Y142_I;
  wire [0:0] RIOB33_X105Y143_IOB_X1Y143_I;
  wire [0:0] RIOB33_X105Y143_IOB_X1Y144_I;
  wire [0:0] RIOB33_X105Y145_IOB_X1Y145_I;
  wire [0:0] RIOB33_X105Y145_IOB_X1Y146_I;
  wire [0:0] RIOB33_X105Y147_IOB_X1Y147_I;
  wire [0:0] RIOB33_X105Y147_IOB_X1Y148_I;
  wire [0:0] RIOB33_X105Y151_IOB_X1Y151_O;
  wire [0:0] RIOB33_X105Y151_IOB_X1Y152_O;
  wire [0:0] RIOB33_X105Y153_IOB_X1Y153_O;
  wire [0:0] RIOB33_X105Y153_IOB_X1Y154_O;
  wire [0:0] RIOB33_X105Y155_IOB_X1Y155_O;
  wire [0:0] RIOB33_X105Y155_IOB_X1Y156_O;
  wire [0:0] RIOB33_X105Y157_IOB_X1Y157_O;
  wire [0:0] RIOB33_X105Y157_IOB_X1Y158_O;
  wire [0:0] RIOB33_X105Y159_IOB_X1Y159_O;
  wire [0:0] RIOB33_X105Y159_IOB_X1Y160_O;
  wire [0:0] RIOB33_X105Y161_IOB_X1Y161_O;
  wire [0:0] RIOB33_X105Y161_IOB_X1Y162_O;
  wire [0:0] RIOB33_X105Y163_IOB_X1Y163_O;
  wire [0:0] RIOB33_X105Y163_IOB_X1Y164_O;
  wire [0:0] RIOB33_X105Y165_IOB_X1Y165_O;
  wire [0:0] RIOB33_X105Y165_IOB_X1Y166_O;
  wire [0:0] RIOB33_X105Y167_IOB_X1Y167_O;
  wire [0:0] RIOB33_X105Y167_IOB_X1Y168_O;
  wire [0:0] RIOB33_X105Y169_IOB_X1Y169_O;
  wire [0:0] RIOB33_X105Y169_IOB_X1Y170_O;
  wire [0:0] RIOB33_X105Y171_IOB_X1Y171_O;
  wire [0:0] RIOB33_X105Y171_IOB_X1Y172_O;
  wire [0:0] RIOB33_X105Y173_IOB_X1Y173_O;
  wire [0:0] RIOB33_X105Y173_IOB_X1Y174_O;
  wire [0:0] RIOB33_X105Y175_IOB_X1Y175_O;
  wire [0:0] RIOB33_X105Y175_IOB_X1Y176_O;
  wire [0:0] RIOB33_X105Y177_IOB_X1Y177_O;
  wire [0:0] RIOB33_X105Y177_IOB_X1Y178_O;
  wire [0:0] RIOB33_X105Y179_IOB_X1Y179_O;
  wire [0:0] RIOB33_X105Y179_IOB_X1Y180_O;
  wire [0:0] RIOB33_X105Y181_IOB_X1Y181_O;
  wire [0:0] RIOB33_X105Y181_IOB_X1Y182_O;
  wire [0:0] RIOB33_X105Y183_IOB_X1Y183_O;
  wire [0:0] RIOB33_X105Y183_IOB_X1Y184_O;
  wire [0:0] RIOB33_X105Y185_IOB_X1Y185_O;
  wire [0:0] RIOB33_X105Y185_IOB_X1Y186_O;
  wire [0:0] RIOB33_X105Y187_IOB_X1Y187_O;
  wire [0:0] RIOB33_X105Y187_IOB_X1Y188_O;
  wire [0:0] RIOB33_X105Y189_IOB_X1Y189_O;
  wire [0:0] RIOB33_X105Y189_IOB_X1Y190_O;
  wire [0:0] RIOB33_X105Y191_IOB_X1Y191_O;
  wire [0:0] RIOB33_X105Y191_IOB_X1Y192_O;
  wire [0:0] RIOB33_X105Y193_IOB_X1Y193_O;
  wire [0:0] RIOB33_X105Y193_IOB_X1Y194_O;
  wire [0:0] RIOB33_X105Y195_IOB_X1Y195_O;
  wire [0:0] RIOB33_X105Y195_IOB_X1Y196_O;
  wire [0:0] RIOB33_X105Y197_IOB_X1Y197_O;
  wire [0:0] RIOB33_X105Y197_IOB_X1Y198_O;
  wire [0:0] RIOI3_SING_X105Y100_ILOGIC_X1Y100_D;
  wire [0:0] RIOI3_SING_X105Y100_ILOGIC_X1Y100_O;
  wire [0:0] RIOI3_SING_X105Y149_ILOGIC_X1Y149_D;
  wire [0:0] RIOI3_SING_X105Y149_ILOGIC_X1Y149_O;
  wire [0:0] RIOI3_SING_X105Y150_OLOGIC_X1Y150_D1;
  wire [0:0] RIOI3_SING_X105Y150_OLOGIC_X1Y150_OQ;
  wire [0:0] RIOI3_SING_X105Y150_OLOGIC_X1Y150_T1;
  wire [0:0] RIOI3_SING_X105Y150_OLOGIC_X1Y150_TQ;
  wire [0:0] RIOI3_SING_X105Y199_OLOGIC_X1Y199_D1;
  wire [0:0] RIOI3_SING_X105Y199_OLOGIC_X1Y199_OQ;
  wire [0:0] RIOI3_SING_X105Y199_OLOGIC_X1Y199_T1;
  wire [0:0] RIOI3_SING_X105Y199_OLOGIC_X1Y199_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y131_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y131_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y132_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y132_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y143_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y143_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y144_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y144_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y114_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y114_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y137_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y137_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y138_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y138_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_TQ;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y101_D;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y101_O;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y102_D;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y102_O;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y103_D;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y103_O;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y104_D;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y104_O;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y105_D;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y105_O;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y106_D;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y106_O;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y109_D;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y109_O;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y110_D;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y110_O;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y111_D;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y111_O;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y112_D;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y112_O;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y115_D;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y115_O;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y116_D;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y116_O;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y117_D;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y117_O;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y118_D;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y118_O;
  wire [0:0] RIOI3_X105Y121_ILOGIC_X1Y121_D;
  wire [0:0] RIOI3_X105Y121_ILOGIC_X1Y121_O;
  wire [0:0] RIOI3_X105Y121_ILOGIC_X1Y122_D;
  wire [0:0] RIOI3_X105Y121_ILOGIC_X1Y122_O;
  wire [0:0] RIOI3_X105Y123_ILOGIC_X1Y123_D;
  wire [0:0] RIOI3_X105Y123_ILOGIC_X1Y123_O;
  wire [0:0] RIOI3_X105Y123_ILOGIC_X1Y124_D;
  wire [0:0] RIOI3_X105Y123_ILOGIC_X1Y124_O;
  wire [0:0] RIOI3_X105Y125_ILOGIC_X1Y125_D;
  wire [0:0] RIOI3_X105Y125_ILOGIC_X1Y125_O;
  wire [0:0] RIOI3_X105Y125_ILOGIC_X1Y126_D;
  wire [0:0] RIOI3_X105Y125_ILOGIC_X1Y126_O;
  wire [0:0] RIOI3_X105Y127_ILOGIC_X1Y127_D;
  wire [0:0] RIOI3_X105Y127_ILOGIC_X1Y127_O;
  wire [0:0] RIOI3_X105Y127_ILOGIC_X1Y128_D;
  wire [0:0] RIOI3_X105Y127_ILOGIC_X1Y128_O;
  wire [0:0] RIOI3_X105Y129_ILOGIC_X1Y129_D;
  wire [0:0] RIOI3_X105Y129_ILOGIC_X1Y129_O;
  wire [0:0] RIOI3_X105Y129_ILOGIC_X1Y130_D;
  wire [0:0] RIOI3_X105Y129_ILOGIC_X1Y130_O;
  wire [0:0] RIOI3_X105Y133_ILOGIC_X1Y133_D;
  wire [0:0] RIOI3_X105Y133_ILOGIC_X1Y133_O;
  wire [0:0] RIOI3_X105Y133_ILOGIC_X1Y134_D;
  wire [0:0] RIOI3_X105Y133_ILOGIC_X1Y134_O;
  wire [0:0] RIOI3_X105Y135_ILOGIC_X1Y135_D;
  wire [0:0] RIOI3_X105Y135_ILOGIC_X1Y135_O;
  wire [0:0] RIOI3_X105Y135_ILOGIC_X1Y136_D;
  wire [0:0] RIOI3_X105Y135_ILOGIC_X1Y136_O;
  wire [0:0] RIOI3_X105Y139_ILOGIC_X1Y139_D;
  wire [0:0] RIOI3_X105Y139_ILOGIC_X1Y139_O;
  wire [0:0] RIOI3_X105Y139_ILOGIC_X1Y140_D;
  wire [0:0] RIOI3_X105Y139_ILOGIC_X1Y140_O;
  wire [0:0] RIOI3_X105Y141_ILOGIC_X1Y141_D;
  wire [0:0] RIOI3_X105Y141_ILOGIC_X1Y141_O;
  wire [0:0] RIOI3_X105Y141_ILOGIC_X1Y142_D;
  wire [0:0] RIOI3_X105Y141_ILOGIC_X1Y142_O;
  wire [0:0] RIOI3_X105Y145_ILOGIC_X1Y145_D;
  wire [0:0] RIOI3_X105Y145_ILOGIC_X1Y145_O;
  wire [0:0] RIOI3_X105Y145_ILOGIC_X1Y146_D;
  wire [0:0] RIOI3_X105Y145_ILOGIC_X1Y146_O;
  wire [0:0] RIOI3_X105Y147_ILOGIC_X1Y147_D;
  wire [0:0] RIOI3_X105Y147_ILOGIC_X1Y147_O;
  wire [0:0] RIOI3_X105Y147_ILOGIC_X1Y148_D;
  wire [0:0] RIOI3_X105Y147_ILOGIC_X1Y148_O;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y151_D1;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y151_OQ;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y151_T1;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y151_TQ;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y152_D1;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y152_OQ;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y152_T1;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y152_TQ;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y153_D1;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y153_OQ;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y153_T1;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y153_TQ;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y154_D1;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y154_OQ;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y154_T1;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y154_TQ;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y155_D1;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y155_OQ;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y155_T1;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y155_TQ;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y156_D1;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y156_OQ;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y156_T1;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y156_TQ;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y159_D1;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y159_OQ;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y159_T1;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y159_TQ;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y160_D1;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y160_OQ;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y160_T1;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y160_TQ;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y161_D1;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y161_OQ;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y161_T1;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y161_TQ;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y162_D1;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y162_OQ;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y162_T1;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y162_TQ;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y165_D1;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y165_OQ;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y165_T1;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y165_TQ;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y166_D1;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y166_OQ;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y166_T1;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y166_TQ;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y167_D1;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y167_OQ;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y167_T1;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y167_TQ;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y168_D1;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y168_OQ;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y168_T1;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y168_TQ;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y171_D1;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y171_OQ;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y171_T1;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y171_TQ;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y172_D1;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y172_OQ;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y172_T1;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y172_TQ;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y173_D1;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y173_OQ;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y173_T1;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y173_TQ;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y174_D1;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y174_OQ;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y174_T1;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y174_TQ;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y175_D1;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y175_OQ;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y175_T1;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y175_TQ;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y176_D1;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y176_OQ;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y176_T1;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y176_TQ;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y177_D1;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y177_OQ;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y177_T1;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y177_TQ;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y178_D1;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y178_OQ;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y178_T1;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y178_TQ;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y179_D1;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y179_OQ;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y179_T1;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y179_TQ;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y180_D1;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y180_OQ;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y180_T1;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y180_TQ;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y183_D1;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y183_OQ;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y183_T1;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y183_TQ;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y184_D1;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y184_OQ;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y184_T1;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y184_TQ;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y185_D1;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y185_OQ;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y185_T1;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y185_TQ;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y186_D1;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y186_OQ;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y186_T1;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y186_TQ;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y189_D1;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y189_OQ;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y189_T1;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y189_TQ;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y190_D1;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y190_OQ;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y190_T1;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y190_TQ;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y191_D1;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y191_OQ;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y191_T1;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y191_TQ;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y192_D1;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y192_OQ;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y192_T1;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y192_TQ;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y195_D1;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y195_OQ;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y195_T1;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y195_TQ;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y196_D1;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y196_OQ;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y196_T1;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y196_TQ;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y197_D1;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y197_OQ;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y197_T1;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y197_TQ;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y198_D1;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y198_OQ;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y198_T1;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y198_TQ;


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y108_SLICE_X0Y108_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y108_SLICE_X0Y108_DO5),
.O6(CLBLL_L_X2Y108_SLICE_X0Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y108_SLICE_X0Y108_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y108_SLICE_X0Y108_CO5),
.O6(CLBLL_L_X2Y108_SLICE_X0Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y108_SLICE_X0Y108_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y108_SLICE_X0Y108_BO5),
.O6(CLBLL_L_X2Y108_SLICE_X0Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00ff00ff00ff)
  ) CLBLL_L_X2Y108_SLICE_X0Y108_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X3Y133_SLICE_X2Y133_BO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y108_SLICE_X0Y108_AO5),
.O6(CLBLL_L_X2Y108_SLICE_X0Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y108_SLICE_X1Y108_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y108_SLICE_X1Y108_DO5),
.O6(CLBLL_L_X2Y108_SLICE_X1Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y108_SLICE_X1Y108_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y108_SLICE_X1Y108_CO5),
.O6(CLBLL_L_X2Y108_SLICE_X1Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y108_SLICE_X1Y108_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y108_SLICE_X1Y108_BO5),
.O6(CLBLL_L_X2Y108_SLICE_X1Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y108_SLICE_X1Y108_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y108_SLICE_X1Y108_AO5),
.O6(CLBLL_L_X2Y108_SLICE_X1Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y127_SLICE_X0Y127_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y127_SLICE_X0Y127_DO5),
.O6(CLBLL_L_X2Y127_SLICE_X0Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y127_SLICE_X0Y127_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y127_SLICE_X0Y127_CO5),
.O6(CLBLL_L_X2Y127_SLICE_X0Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y127_SLICE_X0Y127_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y127_SLICE_X0Y127_BO5),
.O6(CLBLL_L_X2Y127_SLICE_X0Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h666666660a0a0a0a)
  ) CLBLL_L_X2Y127_SLICE_X0Y127_ALUT (
.I0(CLBLL_L_X4Y133_SLICE_X4Y133_CO6),
.I1(CLBLM_R_X5Y136_SLICE_X7Y136_DO5),
.I2(CLBLM_R_X3Y133_SLICE_X2Y133_BO6),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y127_SLICE_X0Y127_AO5),
.O6(CLBLL_L_X2Y127_SLICE_X0Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y127_SLICE_X1Y127_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y127_SLICE_X1Y127_DO5),
.O6(CLBLL_L_X2Y127_SLICE_X1Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y127_SLICE_X1Y127_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y127_SLICE_X1Y127_CO5),
.O6(CLBLL_L_X2Y127_SLICE_X1Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y127_SLICE_X1Y127_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y127_SLICE_X1Y127_BO5),
.O6(CLBLL_L_X2Y127_SLICE_X1Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y127_SLICE_X1Y127_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y127_SLICE_X1Y127_AO5),
.O6(CLBLL_L_X2Y127_SLICE_X1Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y133_SLICE_X0Y133_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y133_SLICE_X0Y133_DO5),
.O6(CLBLL_L_X2Y133_SLICE_X0Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffdfdffffffdd)
  ) CLBLL_L_X2Y133_SLICE_X0Y133_CLUT (
.I0(RIOB33_X105Y137_IOB_X1Y137_I),
.I1(RIOB33_X105Y127_IOB_X1Y128_I),
.I2(CLBLL_L_X4Y139_SLICE_X4Y139_BO6),
.I3(CLBLM_R_X5Y136_SLICE_X7Y136_DO5),
.I4(RIOB33_X105Y129_IOB_X1Y129_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y133_SLICE_X0Y133_CO5),
.O6(CLBLL_L_X2Y133_SLICE_X0Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffafffffefef)
  ) CLBLL_L_X2Y133_SLICE_X0Y133_BLUT (
.I0(RIOB33_X105Y129_IOB_X1Y129_I),
.I1(CLBLM_R_X3Y140_SLICE_X2Y140_DO6),
.I2(RIOB33_X105Y137_IOB_X1Y137_I),
.I3(CLBLM_R_X5Y142_SLICE_X6Y142_CO6),
.I4(RIOB33_X105Y127_IOB_X1Y128_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y133_SLICE_X0Y133_BO5),
.O6(CLBLL_L_X2Y133_SLICE_X0Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffefefffffffaf)
  ) CLBLL_L_X2Y133_SLICE_X0Y133_ALUT (
.I0(RIOB33_X105Y129_IOB_X1Y129_I),
.I1(CLBLL_L_X4Y142_SLICE_X4Y142_BO6),
.I2(RIOB33_X105Y137_IOB_X1Y137_I),
.I3(CLBLM_R_X5Y140_SLICE_X6Y140_AO6),
.I4(RIOB33_X105Y127_IOB_X1Y128_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y133_SLICE_X0Y133_AO5),
.O6(CLBLL_L_X2Y133_SLICE_X0Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y133_SLICE_X1Y133_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y133_SLICE_X1Y133_DO5),
.O6(CLBLL_L_X2Y133_SLICE_X1Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y133_SLICE_X1Y133_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y133_SLICE_X1Y133_CO5),
.O6(CLBLL_L_X2Y133_SLICE_X1Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y133_SLICE_X1Y133_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y133_SLICE_X1Y133_BO5),
.O6(CLBLL_L_X2Y133_SLICE_X1Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y133_SLICE_X1Y133_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y133_SLICE_X1Y133_AO5),
.O6(CLBLL_L_X2Y133_SLICE_X1Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y140_SLICE_X0Y140_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y140_SLICE_X0Y140_DO5),
.O6(CLBLL_L_X2Y140_SLICE_X0Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y140_SLICE_X0Y140_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y140_SLICE_X0Y140_CO5),
.O6(CLBLL_L_X2Y140_SLICE_X0Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y140_SLICE_X0Y140_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y140_SLICE_X0Y140_BO5),
.O6(CLBLL_L_X2Y140_SLICE_X0Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y140_SLICE_X0Y140_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y140_SLICE_X0Y140_AO5),
.O6(CLBLL_L_X2Y140_SLICE_X0Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y140_SLICE_X1Y140_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y140_SLICE_X1Y140_DO5),
.O6(CLBLL_L_X2Y140_SLICE_X1Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y140_SLICE_X1Y140_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y140_SLICE_X1Y140_CO5),
.O6(CLBLL_L_X2Y140_SLICE_X1Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y140_SLICE_X1Y140_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y140_SLICE_X1Y140_BO5),
.O6(CLBLL_L_X2Y140_SLICE_X1Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffefffef02000000)
  ) CLBLL_L_X2Y140_SLICE_X1Y140_ALUT (
.I0(RIOB33_X105Y133_IOB_X1Y133_I),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(RIOB33_X105Y133_IOB_X1Y134_I),
.I3(RIOB33_X105Y131_IOB_X1Y132_I),
.I4(RIOB33_X105Y135_IOB_X1Y136_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y140_SLICE_X1Y140_AO5),
.O6(CLBLL_L_X2Y140_SLICE_X1Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y141_SLICE_X0Y141_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y141_SLICE_X0Y141_DO5),
.O6(CLBLL_L_X2Y141_SLICE_X0Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y141_SLICE_X0Y141_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y141_SLICE_X0Y141_CO5),
.O6(CLBLL_L_X2Y141_SLICE_X0Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y141_SLICE_X0Y141_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y141_SLICE_X0Y141_BO5),
.O6(CLBLL_L_X2Y141_SLICE_X0Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0030001000200000)
  ) CLBLL_L_X2Y141_SLICE_X0Y141_ALUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(CLBLM_R_X3Y143_SLICE_X2Y143_AO6),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(CLBLM_R_X3Y138_SLICE_X2Y138_AO5),
.I4(LIOB33_X0Y61_IOB_X0Y61_I),
.I5(LIOB33_X0Y71_IOB_X0Y71_I),
.O5(CLBLL_L_X2Y141_SLICE_X0Y141_AO5),
.O6(CLBLL_L_X2Y141_SLICE_X0Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffddfffdccccfcfc)
  ) CLBLL_L_X2Y141_SLICE_X1Y141_DLUT (
.I0(RIOB33_X105Y137_IOB_X1Y137_I),
.I1(CLBLL_L_X2Y141_SLICE_X0Y141_AO6),
.I2(LIOB33_X0Y55_IOB_X0Y55_I),
.I3(RIOB33_X105Y129_IOB_X1Y129_I),
.I4(CLBLL_L_X2Y141_SLICE_X1Y141_BO5),
.I5(CLBLM_L_X10Y140_SLICE_X13Y140_C5Q),
.O5(CLBLL_L_X2Y141_SLICE_X1Y141_DO5),
.O6(CLBLL_L_X2Y141_SLICE_X1Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h000a000000ce00cc)
  ) CLBLL_L_X2Y141_SLICE_X1Y141_CLUT (
.I0(CLBLL_L_X2Y141_SLICE_X1Y141_AO6),
.I1(LIOB33_X0Y53_IOB_X0Y54_I),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(CLBLM_R_X3Y143_SLICE_X2Y143_AO6),
.I4(LIOB33_X0Y69_IOB_X0Y70_I),
.I5(CLBLL_L_X2Y141_SLICE_X1Y141_BO6),
.O5(CLBLL_L_X2Y141_SLICE_X1Y141_CO5),
.O6(CLBLL_L_X2Y141_SLICE_X1Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff5fffffffdfffff)
  ) CLBLL_L_X2Y141_SLICE_X1Y141_BLUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(CLBLM_R_X3Y143_SLICE_X2Y143_AO6),
.I2(RIOB33_X105Y133_IOB_X1Y134_I),
.I3(RIOB33_X105Y133_IOB_X1Y133_I),
.I4(RIOB33_X105Y131_IOB_X1Y132_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y141_SLICE_X1Y141_BO5),
.O6(CLBLL_L_X2Y141_SLICE_X1Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00cc0000ffffccff)
  ) CLBLL_L_X2Y141_SLICE_X1Y141_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y133_IOB_X1Y133_I),
.I2(1'b1),
.I3(RIOB33_X105Y133_IOB_X1Y134_I),
.I4(RIOB33_X105Y131_IOB_X1Y132_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y141_SLICE_X1Y141_AO5),
.O6(CLBLL_L_X2Y141_SLICE_X1Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y132_SLICE_X4Y132_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y132_SLICE_X4Y132_DO5),
.O6(CLBLL_L_X4Y132_SLICE_X4Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y132_SLICE_X4Y132_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y132_SLICE_X4Y132_CO5),
.O6(CLBLL_L_X4Y132_SLICE_X4Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y132_SLICE_X4Y132_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y132_SLICE_X4Y132_BO5),
.O6(CLBLL_L_X4Y132_SLICE_X4Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y132_SLICE_X4Y132_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y132_SLICE_X4Y132_AO5),
.O6(CLBLL_L_X4Y132_SLICE_X4Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y132_SLICE_X5Y132_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y132_SLICE_X5Y132_AO6),
.Q(CLBLL_L_X4Y132_SLICE_X5Y132_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y132_SLICE_X5Y132_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y132_SLICE_X5Y132_DO5),
.O6(CLBLL_L_X4Y132_SLICE_X5Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y132_SLICE_X5Y132_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y132_SLICE_X5Y132_CO5),
.O6(CLBLL_L_X4Y132_SLICE_X5Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y132_SLICE_X5Y132_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y132_SLICE_X5Y132_BO5),
.O6(CLBLL_L_X4Y132_SLICE_X5Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00ff55aa00fa50)
  ) CLBLL_L_X4Y132_SLICE_X5Y132_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(1'b1),
.I2(CLBLM_L_X10Y131_SLICE_X13Y131_AQ),
.I3(CLBLM_R_X5Y136_SLICE_X6Y136_DQ),
.I4(CLBLM_R_X5Y133_SLICE_X7Y133_DO6),
.I5(CLBLL_L_X4Y132_SLICE_X5Y132_AQ),
.O5(CLBLL_L_X4Y132_SLICE_X5Y132_AO5),
.O6(CLBLL_L_X4Y132_SLICE_X5Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y133_SLICE_X4Y133_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y133_SLICE_X4Y133_AO6),
.Q(CLBLL_L_X4Y133_SLICE_X4Y133_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y133_SLICE_X4Y133_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y133_SLICE_X4Y133_DO5),
.O6(CLBLL_L_X4Y133_SLICE_X4Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h550555057727ffaf)
  ) CLBLL_L_X4Y133_SLICE_X4Y133_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLL_L_X4Y139_SLICE_X4Y139_BO6),
.I2(CLBLL_L_X4Y142_SLICE_X4Y142_BO6),
.I3(CLBLL_L_X4Y136_SLICE_X4Y136_AO5),
.I4(CLBLM_L_X12Y134_SLICE_X17Y134_AQ),
.I5(CLBLM_R_X5Y133_SLICE_X6Y133_CO6),
.O5(CLBLL_L_X4Y133_SLICE_X4Y133_CO5),
.O6(CLBLL_L_X4Y133_SLICE_X4Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0ccc8cc0000aaaa)
  ) CLBLL_L_X4Y133_SLICE_X4Y133_BLUT (
.I0(CLBLL_L_X4Y134_SLICE_X5Y134_A5Q),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLL_L_X4Y135_SLICE_X5Y135_C5Q),
.I3(CLBLM_R_X11Y138_SLICE_X15Y138_BQ),
.I4(CLBLL_L_X4Y134_SLICE_X4Y134_B5Q),
.I5(1'b1),
.O5(CLBLL_L_X4Y133_SLICE_X4Y133_BO5),
.O6(CLBLL_L_X4Y133_SLICE_X4Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00ea40ae04)
  ) CLBLL_L_X4Y133_SLICE_X4Y133_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLL_L_X4Y133_SLICE_X4Y133_AQ),
.I3(CLBLM_R_X3Y135_SLICE_X3Y135_BQ),
.I4(CLBLM_R_X5Y132_SLICE_X7Y132_CO5),
.I5(CLBLM_R_X11Y138_SLICE_X15Y138_BQ),
.O5(CLBLL_L_X4Y133_SLICE_X4Y133_AO5),
.O6(CLBLL_L_X4Y133_SLICE_X4Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y133_SLICE_X5Y133_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y136_SLICE_X5Y136_DO6),
.Q(CLBLL_L_X4Y133_SLICE_X5Y133_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y133_SLICE_X5Y133_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y133_SLICE_X5Y133_AO6),
.Q(CLBLL_L_X4Y133_SLICE_X5Y133_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbffbbffffffffff)
  ) CLBLL_L_X4Y133_SLICE_X5Y133_DLUT (
.I0(CLBLM_L_X10Y132_SLICE_X12Y132_AO6),
.I1(CLBLL_L_X4Y134_SLICE_X5Y134_AQ),
.I2(1'b1),
.I3(CLBLM_R_X5Y132_SLICE_X7Y132_BO5),
.I4(1'b1),
.I5(CLBLM_R_X5Y132_SLICE_X7Y132_DO6),
.O5(CLBLL_L_X4Y133_SLICE_X5Y133_DO5),
.O6(CLBLL_L_X4Y133_SLICE_X5Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hbfffffffffffffff)
  ) CLBLL_L_X4Y133_SLICE_X5Y133_CLUT (
.I0(CLBLM_L_X10Y132_SLICE_X12Y132_AO6),
.I1(CLBLL_L_X4Y134_SLICE_X5Y134_CQ),
.I2(CLBLL_L_X4Y134_SLICE_X5Y134_AQ),
.I3(CLBLM_R_X5Y132_SLICE_X7Y132_BO5),
.I4(CLBLL_L_X4Y133_SLICE_X5Y133_AQ),
.I5(CLBLM_R_X5Y132_SLICE_X7Y132_DO6),
.O5(CLBLL_L_X4Y133_SLICE_X5Y133_CO5),
.O6(CLBLL_L_X4Y133_SLICE_X5Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h000a002a00000000)
  ) CLBLL_L_X4Y133_SLICE_X5Y133_BLUT (
.I0(CLBLM_R_X5Y132_SLICE_X7Y132_DO6),
.I1(CLBLL_L_X4Y133_SLICE_X4Y133_BO5),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_L_X10Y132_SLICE_X12Y132_AO6),
.I4(CLBLL_L_X4Y135_SLICE_X5Y135_C5Q),
.I5(CLBLM_R_X5Y132_SLICE_X7Y132_BO5),
.O5(CLBLL_L_X4Y133_SLICE_X5Y133_BO5),
.O6(CLBLL_L_X4Y133_SLICE_X5Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcca5cc00ccf0cc00)
  ) CLBLL_L_X4Y133_SLICE_X5Y133_ALUT (
.I0(CLBLL_L_X4Y133_SLICE_X5Y133_DO6),
.I1(CLBLM_R_X11Y133_SLICE_X15Y133_BQ),
.I2(CLBLL_L_X4Y133_SLICE_X5Y133_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLL_L_X4Y133_SLICE_X4Y133_BO6),
.I5(CLBLL_L_X4Y134_SLICE_X5Y134_CQ),
.O5(CLBLL_L_X4Y133_SLICE_X5Y133_AO5),
.O6(CLBLL_L_X4Y133_SLICE_X5Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y134_SLICE_X4Y134_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y134_SLICE_X4Y134_BO5),
.Q(CLBLL_L_X4Y134_SLICE_X4Y134_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y134_SLICE_X4Y134_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y134_SLICE_X4Y134_AO6),
.Q(CLBLL_L_X4Y134_SLICE_X4Y134_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y134_SLICE_X4Y134_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y134_SLICE_X4Y134_BO6),
.Q(CLBLL_L_X4Y134_SLICE_X4Y134_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y134_SLICE_X4Y134_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y134_SLICE_X4Y134_DO5),
.O6(CLBLL_L_X4Y134_SLICE_X4Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y134_SLICE_X4Y134_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y134_SLICE_X4Y134_CO5),
.O6(CLBLL_L_X4Y134_SLICE_X4Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaa5500dddd8888)
  ) CLBLL_L_X4Y134_SLICE_X4Y134_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.I2(1'b1),
.I3(CLBLM_R_X11Y135_SLICE_X14Y135_AQ),
.I4(CLBLL_L_X4Y134_SLICE_X5Y134_A5Q),
.I5(1'b1),
.O5(CLBLL_L_X4Y134_SLICE_X4Y134_BO5),
.O6(CLBLL_L_X4Y134_SLICE_X4Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaa5500feba5410)
  ) CLBLL_L_X4Y134_SLICE_X4Y134_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y138_SLICE_X10Y138_AQ),
.I2(CLBLL_L_X4Y134_SLICE_X4Y134_AQ),
.I3(CLBLM_R_X11Y135_SLICE_X14Y135_AQ),
.I4(CLBLM_R_X3Y137_SLICE_X3Y137_AQ),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLL_L_X4Y134_SLICE_X4Y134_AO5),
.O6(CLBLL_L_X4Y134_SLICE_X4Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y134_SLICE_X5Y134_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y134_SLICE_X5Y134_DO5),
.Q(CLBLL_L_X4Y134_SLICE_X5Y134_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y134_SLICE_X5Y134_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y134_SLICE_X5Y134_AO6),
.Q(CLBLL_L_X4Y134_SLICE_X5Y134_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y134_SLICE_X5Y134_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y134_SLICE_X5Y134_BO6),
.Q(CLBLL_L_X4Y134_SLICE_X5Y134_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y134_SLICE_X5Y134_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y134_SLICE_X5Y134_CO6),
.Q(CLBLL_L_X4Y134_SLICE_X5Y134_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h88000000f8f00000)
  ) CLBLL_L_X4Y134_SLICE_X5Y134_DLUT (
.I0(CLBLL_L_X4Y134_SLICE_X5Y134_BQ),
.I1(CLBLL_L_X4Y134_SLICE_X5Y134_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLL_L_X4Y134_SLICE_X5Y134_AQ),
.I4(CLBLL_L_X4Y133_SLICE_X5Y133_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y134_SLICE_X5Y134_DO5),
.O6(CLBLL_L_X4Y134_SLICE_X5Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf909fc0cf000f000)
  ) CLBLL_L_X4Y134_SLICE_X5Y134_CLUT (
.I0(CLBLM_R_X5Y132_SLICE_X6Y132_AO6),
.I1(CLBLL_L_X4Y134_SLICE_X5Y134_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y133_SLICE_X8Y133_CQ),
.I4(CLBLL_L_X4Y134_SLICE_X5Y134_AQ),
.I5(CLBLL_L_X4Y133_SLICE_X4Y133_BO6),
.O5(CLBLL_L_X4Y134_SLICE_X5Y134_CO5),
.O6(CLBLL_L_X4Y134_SLICE_X5Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcdcccdc30100010)
  ) CLBLL_L_X4Y134_SLICE_X5Y134_BLUT (
.I0(CLBLL_L_X4Y134_SLICE_X5Y134_DO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLL_L_X4Y133_SLICE_X4Y133_BO6),
.I3(CLBLL_L_X4Y133_SLICE_X5Y133_CO6),
.I4(CLBLL_L_X4Y134_SLICE_X5Y134_BQ),
.I5(CLBLM_L_X8Y134_SLICE_X11Y134_CQ),
.O5(CLBLL_L_X4Y134_SLICE_X5Y134_BO5),
.O6(CLBLL_L_X4Y134_SLICE_X5Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hd888d88888d888d8)
  ) CLBLL_L_X4Y134_SLICE_X5Y134_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLL_L_X4Y134_SLICE_X5Y134_BQ),
.I2(CLBLL_L_X4Y133_SLICE_X4Y133_BO6),
.I3(CLBLM_R_X5Y132_SLICE_X6Y132_AO6),
.I4(1'b1),
.I5(CLBLL_L_X4Y134_SLICE_X5Y134_AQ),
.O5(CLBLL_L_X4Y134_SLICE_X5Y134_AO5),
.O6(CLBLL_L_X4Y134_SLICE_X5Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y135_SLICE_X4Y135_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y135_SLICE_X4Y135_DO6),
.Q(CLBLL_L_X4Y135_SLICE_X4Y135_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y135_SLICE_X4Y135_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y135_SLICE_X4Y135_AO6),
.Q(CLBLL_L_X4Y135_SLICE_X4Y135_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y135_SLICE_X4Y135_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y135_SLICE_X4Y135_BO6),
.Q(CLBLL_L_X4Y135_SLICE_X4Y135_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y135_SLICE_X4Y135_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y135_SLICE_X4Y135_CO6),
.Q(CLBLL_L_X4Y135_SLICE_X4Y135_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfc0c0cff77ff77)
  ) CLBLL_L_X4Y135_SLICE_X4Y135_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X5Y137_SLICE_X6Y137_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLL_L_X4Y135_SLICE_X4Y135_A5Q),
.I4(CLBLM_R_X5Y138_SLICE_X7Y138_CQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y135_SLICE_X4Y135_DO5),
.O6(CLBLL_L_X4Y135_SLICE_X4Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffcffccf0f00000)
  ) CLBLL_L_X4Y135_SLICE_X4Y135_CLUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y135_SLICE_X4Y135_CQ),
.I2(CLBLM_R_X3Y135_SLICE_X3Y135_AQ),
.I3(CLBLM_R_X7Y135_SLICE_X9Y135_A5Q),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y144_SLICE_X9Y144_BO6),
.O5(CLBLL_L_X4Y135_SLICE_X4Y135_CO5),
.O6(CLBLL_L_X4Y135_SLICE_X4Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffececa0a0a0a0)
  ) CLBLL_L_X4Y135_SLICE_X4Y135_BLUT (
.I0(CLBLL_L_X4Y135_SLICE_X5Y135_DQ),
.I1(CLBLL_L_X4Y135_SLICE_X4Y135_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(CLBLM_L_X10Y134_SLICE_X13Y134_BQ),
.I5(CLBLM_R_X7Y144_SLICE_X9Y144_BO6),
.O5(CLBLL_L_X4Y135_SLICE_X4Y135_BO5),
.O6(CLBLL_L_X4Y135_SLICE_X4Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffcfcfcff000000)
  ) CLBLL_L_X4Y135_SLICE_X4Y135_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y137_SLICE_X9Y137_BQ),
.I2(CLBLL_L_X4Y135_SLICE_X4Y135_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X12Y133_SLICE_X16Y133_C5Q),
.I5(CLBLM_R_X7Y144_SLICE_X9Y144_BO6),
.O5(CLBLL_L_X4Y135_SLICE_X4Y135_AO5),
.O6(CLBLL_L_X4Y135_SLICE_X4Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y135_SLICE_X5Y135_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y135_SLICE_X5Y135_CO5),
.Q(CLBLL_L_X4Y135_SLICE_X5Y135_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y135_SLICE_X5Y135_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y135_SLICE_X5Y135_DO5),
.Q(CLBLL_L_X4Y135_SLICE_X5Y135_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y135_SLICE_X5Y135_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y135_SLICE_X5Y135_AO6),
.Q(CLBLL_L_X4Y135_SLICE_X5Y135_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y135_SLICE_X5Y135_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y135_SLICE_X5Y135_BO6),
.Q(CLBLL_L_X4Y135_SLICE_X5Y135_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y135_SLICE_X5Y135_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y135_SLICE_X5Y135_CO6),
.Q(CLBLL_L_X4Y135_SLICE_X5Y135_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y135_SLICE_X5Y135_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y135_SLICE_X5Y135_DO6),
.Q(CLBLL_L_X4Y135_SLICE_X5Y135_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hafa0afa0cfc0cfc0)
  ) CLBLL_L_X4Y135_SLICE_X5Y135_DLUT (
.I0(CLBLM_R_X7Y135_SLICE_X8Y135_AQ),
.I1(CLBLM_R_X7Y136_SLICE_X8Y136_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y101_IOB_X1Y102_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y135_SLICE_X5Y135_DO5),
.O6(CLBLL_L_X4Y135_SLICE_X5Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcccfccca0a0afaf)
  ) CLBLL_L_X4Y135_SLICE_X5Y135_CLUT (
.I0(CLBLM_R_X7Y137_SLICE_X9Y137_BQ),
.I1(CLBLM_L_X8Y134_SLICE_X10Y134_DO6),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLL_L_X4Y135_SLICE_X4Y135_CQ),
.I4(CLBLM_R_X5Y132_SLICE_X6Y132_AO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y135_SLICE_X5Y135_CO5),
.O6(CLBLL_L_X4Y135_SLICE_X5Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cf03cf03cc00)
  ) CLBLL_L_X4Y135_SLICE_X5Y135_BLUT (
.I0(1'b1),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLL_L_X4Y135_SLICE_X5Y135_D5Q),
.I4(CLBLM_R_X7Y137_SLICE_X9Y137_BQ),
.I5(CLBLM_R_X7Y135_SLICE_X9Y135_DO6),
.O5(CLBLL_L_X4Y135_SLICE_X5Y135_BO5),
.O6(CLBLL_L_X4Y135_SLICE_X5Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000ffa800a8)
  ) CLBLL_L_X4Y135_SLICE_X5Y135_ALUT (
.I0(CLBLM_L_X8Y138_SLICE_X10Y138_AQ),
.I1(CLBLM_L_X8Y134_SLICE_X11Y134_DQ),
.I2(CLBLL_L_X4Y135_SLICE_X5Y135_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLL_L_X4Y135_SLICE_X4Y135_AQ),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLL_L_X4Y135_SLICE_X5Y135_AO5),
.O6(CLBLL_L_X4Y135_SLICE_X5Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y136_SLICE_X4Y136_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y136_SLICE_X4Y136_DO5),
.Q(CLBLL_L_X4Y136_SLICE_X4Y136_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y136_SLICE_X4Y136_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y136_SLICE_X4Y136_AO6),
.Q(CLBLL_L_X4Y136_SLICE_X4Y136_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y136_SLICE_X4Y136_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y136_SLICE_X4Y136_BO6),
.Q(CLBLL_L_X4Y136_SLICE_X4Y136_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y136_SLICE_X4Y136_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y136_SLICE_X4Y136_CO6),
.Q(CLBLL_L_X4Y136_SLICE_X4Y136_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y136_SLICE_X4Y136_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y136_SLICE_X4Y136_DO6),
.Q(CLBLL_L_X4Y136_SLICE_X4Y136_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hc5c0c5c0ff0ff000)
  ) CLBLL_L_X4Y136_SLICE_X4Y136_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X5Y141_SLICE_X6Y141_A5Q),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y135_SLICE_X9Y135_A5Q),
.I4(CLBLL_L_X4Y136_SLICE_X4Y136_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y136_SLICE_X4Y136_DO5),
.O6(CLBLL_L_X4Y136_SLICE_X4Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0cccc00cc)
  ) CLBLL_L_X4Y136_SLICE_X4Y136_CLUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y136_SLICE_X4Y136_CQ),
.I2(CLBLL_L_X4Y137_SLICE_X4Y137_DQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_L_X8Y138_SLICE_X10Y138_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLL_L_X4Y136_SLICE_X4Y136_CO5),
.O6(CLBLL_L_X4Y136_SLICE_X4Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafaf0f0eaeac0c0)
  ) CLBLL_L_X4Y136_SLICE_X4Y136_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLL_L_X4Y136_SLICE_X4Y136_BQ),
.I2(CLBLM_R_X7Y144_SLICE_X9Y144_BO6),
.I3(1'b1),
.I4(CLBLM_R_X7Y132_SLICE_X8Y132_CQ),
.I5(CLBLL_L_X4Y136_SLICE_X4Y136_DQ),
.O5(CLBLL_L_X4Y136_SLICE_X4Y136_BO5),
.O6(CLBLL_L_X4Y136_SLICE_X4Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cca05f5f5f5f)
  ) CLBLL_L_X4Y136_SLICE_X4Y136_ALUT (
.I0(CLBLL_L_X4Y137_SLICE_X4Y137_CQ),
.I1(CLBLL_L_X4Y136_SLICE_X4Y136_BQ),
.I2(CLBLM_L_X12Y135_SLICE_X17Y135_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y136_SLICE_X4Y136_AO5),
.O6(CLBLL_L_X4Y136_SLICE_X4Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y136_SLICE_X5Y136_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y137_SLICE_X5Y137_AO6),
.Q(CLBLL_L_X4Y136_SLICE_X5Y136_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y136_SLICE_X5Y136_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y136_SLICE_X5Y136_AO6),
.Q(CLBLL_L_X4Y136_SLICE_X5Y136_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y136_SLICE_X5Y136_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y136_SLICE_X5Y136_BO6),
.Q(CLBLL_L_X4Y136_SLICE_X5Y136_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y136_SLICE_X5Y136_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y136_SLICE_X5Y136_CO6),
.Q(CLBLL_L_X4Y136_SLICE_X5Y136_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaf0f088008800)
  ) CLBLL_L_X4Y136_SLICE_X5Y136_DLUT (
.I0(CLBLM_R_X5Y136_SLICE_X7Y136_AQ),
.I1(CLBLM_R_X5Y137_SLICE_X6Y137_CQ),
.I2(RIOB33_X105Y127_IOB_X1Y127_I),
.I3(CLBLM_R_X5Y135_SLICE_X7Y135_DO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y136_SLICE_X5Y136_DO5),
.O6(CLBLL_L_X4Y136_SLICE_X5Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0eca0eca0eca0ec)
  ) CLBLL_L_X4Y136_SLICE_X5Y136_CLUT (
.I0(CLBLL_L_X4Y135_SLICE_X5Y135_AQ),
.I1(CLBLL_L_X4Y136_SLICE_X5Y136_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y133_SLICE_X8Y133_DO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y136_SLICE_X5Y136_CO5),
.O6(CLBLL_L_X4Y136_SLICE_X5Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0f5e4f5e4f5e4)
  ) CLBLL_L_X4Y136_SLICE_X5Y136_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLL_L_X4Y136_SLICE_X5Y136_BQ),
.I2(CLBLL_L_X4Y133_SLICE_X4Y133_AQ),
.I3(CLBLM_R_X7Y139_SLICE_X8Y139_AQ),
.I4(CLBLM_L_X12Y135_SLICE_X17Y135_AQ),
.I5(CLBLL_L_X4Y137_SLICE_X4Y137_CQ),
.O5(CLBLL_L_X4Y136_SLICE_X5Y136_BO5),
.O6(CLBLL_L_X4Y136_SLICE_X5Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccf0aaccccaaaa)
  ) CLBLL_L_X4Y136_SLICE_X5Y136_ALUT (
.I0(CLBLM_R_X11Y138_SLICE_X14Y138_BQ),
.I1(CLBLM_R_X5Y135_SLICE_X6Y135_CQ),
.I2(CLBLL_L_X4Y136_SLICE_X5Y136_AQ),
.I3(CLBLM_L_X12Y135_SLICE_X17Y135_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLL_L_X4Y137_SLICE_X4Y137_CQ),
.O5(CLBLL_L_X4Y136_SLICE_X5Y136_AO5),
.O6(CLBLL_L_X4Y136_SLICE_X5Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y137_SLICE_X4Y137_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y137_SLICE_X4Y137_AO5),
.Q(CLBLL_L_X4Y137_SLICE_X4Y137_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y137_SLICE_X4Y137_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y137_SLICE_X4Y137_DO5),
.Q(CLBLL_L_X4Y137_SLICE_X4Y137_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y137_SLICE_X4Y137_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y137_SLICE_X4Y137_AO6),
.Q(CLBLL_L_X4Y137_SLICE_X4Y137_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y137_SLICE_X4Y137_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y137_SLICE_X4Y137_BO6),
.Q(CLBLL_L_X4Y137_SLICE_X4Y137_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y137_SLICE_X4Y137_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y137_SLICE_X4Y137_CO6),
.Q(CLBLL_L_X4Y137_SLICE_X4Y137_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y137_SLICE_X4Y137_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y137_SLICE_X4Y137_DO6),
.Q(CLBLL_L_X4Y137_SLICE_X4Y137_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ff00ccccaaaa)
  ) CLBLL_L_X4Y137_SLICE_X4Y137_DLUT (
.I0(CLBLM_R_X5Y140_SLICE_X6Y140_AO6),
.I1(CLBLM_L_X10Y134_SLICE_X12Y134_CQ),
.I2(CLBLL_L_X4Y136_SLICE_X4Y136_AQ),
.I3(CLBLL_L_X4Y142_SLICE_X4Y142_BO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y137_SLICE_X4Y137_DO5),
.O6(CLBLL_L_X4Y137_SLICE_X4Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff005500000055)
  ) CLBLL_L_X4Y137_SLICE_X4Y137_CLUT (
.I0(CLBLL_L_X4Y136_SLICE_X4Y136_D5Q),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_L_X12Y135_SLICE_X17Y135_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLL_L_X4Y138_SLICE_X5Y138_AQ),
.O5(CLBLL_L_X4Y137_SLICE_X4Y137_CO5),
.O6(CLBLL_L_X4Y137_SLICE_X4Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hbabaeaea3030c0c0)
  ) CLBLL_L_X4Y137_SLICE_X4Y137_BLUT (
.I0(CLBLM_R_X5Y139_SLICE_X7Y139_AQ),
.I1(CLBLL_L_X4Y137_SLICE_X4Y137_BQ),
.I2(CLBLM_R_X7Y135_SLICE_X8Y135_DO5),
.I3(1'b1),
.I4(CLBLL_L_X4Y136_SLICE_X5Y136_DO5),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLL_L_X4Y137_SLICE_X4Y137_BO5),
.O6(CLBLL_L_X4Y137_SLICE_X4Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hafa0afa0cacacaca)
  ) CLBLL_L_X4Y137_SLICE_X4Y137_ALUT (
.I0(CLBLM_R_X7Y135_SLICE_X8Y135_BQ),
.I1(CLBLL_L_X4Y134_SLICE_X4Y134_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLL_L_X4Y139_SLICE_X4Y139_BO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y137_SLICE_X4Y137_AO5),
.O6(CLBLL_L_X4Y137_SLICE_X4Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y137_SLICE_X5Y137_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y137_SLICE_X5Y137_BO6),
.Q(CLBLL_L_X4Y137_SLICE_X5Y137_BQ),
.R(CLBLM_R_X7Y144_SLICE_X9Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000033313331)
  ) CLBLL_L_X4Y137_SLICE_X5Y137_DLUT (
.I0(CLBLM_R_X5Y140_SLICE_X6Y140_AO6),
.I1(CLBLL_L_X4Y138_SLICE_X5Y138_B5Q),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_L_X10Y134_SLICE_X12Y134_CQ),
.I4(1'b1),
.I5(CLBLL_L_X4Y134_SLICE_X4Y134_AQ),
.O5(CLBLL_L_X4Y137_SLICE_X5Y137_DO5),
.O6(CLBLL_L_X4Y137_SLICE_X5Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3100000020000000)
  ) CLBLL_L_X4Y137_SLICE_X5Y137_CLUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(CLBLL_L_X4Y144_SLICE_X4Y144_AO6),
.I2(CLBLM_L_X8Y136_SLICE_X10Y136_AQ),
.I3(RIOB33_X105Y133_IOB_X1Y134_I),
.I4(RIOB33_X105Y133_IOB_X1Y133_I),
.I5(CLBLL_L_X4Y136_SLICE_X5Y136_BQ),
.O5(CLBLL_L_X4Y137_SLICE_X5Y137_CO5),
.O6(CLBLL_L_X4Y137_SLICE_X5Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0ffffcccc)
  ) CLBLL_L_X4Y137_SLICE_X5Y137_BLUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y137_SLICE_X5Y137_BQ),
.I2(CLBLM_R_X3Y136_SLICE_X2Y136_AQ),
.I3(1'b1),
.I4(CLBLM_R_X7Y138_SLICE_X9Y138_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLL_L_X4Y137_SLICE_X5Y137_BO5),
.O6(CLBLL_L_X4Y137_SLICE_X5Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd11dc100f0f0000)
  ) CLBLL_L_X4Y137_SLICE_X5Y137_ALUT (
.I0(CLBLM_L_X8Y137_SLICE_X10Y137_CO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X8Y138_SLICE_X10Y138_AQ),
.I3(CLBLM_R_X3Y136_SLICE_X3Y136_BQ),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y137_SLICE_X5Y137_AO5),
.O6(CLBLL_L_X4Y137_SLICE_X5Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y138_SLICE_X4Y138_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y138_SLICE_X4Y138_AO6),
.Q(CLBLL_L_X4Y138_SLICE_X4Y138_AQ),
.R(CLBLM_R_X7Y144_SLICE_X9Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y138_SLICE_X4Y138_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y138_SLICE_X4Y138_BO6),
.Q(CLBLL_L_X4Y138_SLICE_X4Y138_BQ),
.R(CLBLM_R_X7Y144_SLICE_X9Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00aa00aaf0faf0fa)
  ) CLBLL_L_X4Y138_SLICE_X4Y138_DLUT (
.I0(CLBLL_L_X4Y136_SLICE_X5Y136_AQ),
.I1(1'b1),
.I2(CLBLM_L_X10Y138_SLICE_X13Y138_BQ),
.I3(CLBLL_L_X4Y143_SLICE_X5Y143_AO5),
.I4(1'b1),
.I5(CLBLM_R_X7Y142_SLICE_X9Y142_CO6),
.O5(CLBLL_L_X4Y138_SLICE_X4Y138_DO5),
.O6(CLBLL_L_X4Y138_SLICE_X4Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h4040500000000000)
  ) CLBLL_L_X4Y138_SLICE_X4Y138_CLUT (
.I0(CLBLL_L_X4Y144_SLICE_X4Y144_AO6),
.I1(CLBLL_L_X4Y139_SLICE_X4Y139_AQ),
.I2(RIOB33_X105Y133_IOB_X1Y133_I),
.I3(CLBLM_R_X7Y136_SLICE_X8Y136_BQ),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(RIOB33_X105Y133_IOB_X1Y134_I),
.O5(CLBLL_L_X4Y138_SLICE_X4Y138_CO5),
.O6(CLBLL_L_X4Y138_SLICE_X4Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5f5f5e4e4e4e4)
  ) CLBLL_L_X4Y138_SLICE_X4Y138_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLL_L_X4Y138_SLICE_X4Y138_BQ),
.I2(CLBLL_L_X4Y138_SLICE_X5Y138_B5Q),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X5Y139_SLICE_X7Y139_BQ),
.O5(CLBLL_L_X4Y138_SLICE_X4Y138_BO5),
.O6(CLBLL_L_X4Y138_SLICE_X4Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff3333fcfc3030)
  ) CLBLL_L_X4Y138_SLICE_X4Y138_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLL_L_X4Y138_SLICE_X4Y138_AQ),
.I3(1'b1),
.I4(CLBLL_L_X4Y139_SLICE_X4Y139_AQ),
.I5(CLBLM_L_X8Y136_SLICE_X11Y136_CQ),
.O5(CLBLL_L_X4Y138_SLICE_X4Y138_AO5),
.O6(CLBLL_L_X4Y138_SLICE_X4Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y138_SLICE_X5Y138_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y138_SLICE_X5Y138_AO5),
.Q(CLBLL_L_X4Y138_SLICE_X5Y138_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y138_SLICE_X5Y138_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y138_SLICE_X5Y138_CO6),
.Q(CLBLL_L_X4Y138_SLICE_X5Y138_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y138_SLICE_X5Y138_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y138_SLICE_X5Y138_AO6),
.Q(CLBLL_L_X4Y138_SLICE_X5Y138_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y138_SLICE_X5Y138_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y138_SLICE_X5Y138_BO6),
.Q(CLBLL_L_X4Y138_SLICE_X5Y138_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefeffffcc00ff00)
  ) CLBLL_L_X4Y138_SLICE_X5Y138_DLUT (
.I0(RIOB33_X105Y127_IOB_X1Y128_I),
.I1(RIOB33_X105Y129_IOB_X1Y129_I),
.I2(CLBLL_L_X4Y141_SLICE_X4Y141_DO6),
.I3(CLBLL_L_X4Y138_SLICE_X5Y138_AQ),
.I4(RIOB33_X105Y137_IOB_X1Y137_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y138_SLICE_X5Y138_DO5),
.O6(CLBLL_L_X4Y138_SLICE_X5Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h888888b8f000f000)
  ) CLBLL_L_X4Y138_SLICE_X5Y138_CLUT (
.I0(CLBLL_L_X4Y135_SLICE_X5Y135_BQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X8Y138_SLICE_X10Y138_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLL_L_X4Y137_SLICE_X5Y137_DO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y138_SLICE_X5Y138_CO5),
.O6(CLBLL_L_X4Y138_SLICE_X5Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f0ccf000f0cc)
  ) CLBLL_L_X4Y138_SLICE_X5Y138_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y139_SLICE_X7Y139_BQ),
.I2(CLBLL_L_X4Y136_SLICE_X5Y136_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y138_SLICE_X5Y138_BO5),
.O6(CLBLL_L_X4Y138_SLICE_X5Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfc3030eeaaeeaa)
  ) CLBLL_L_X4Y138_SLICE_X5Y138_ALUT (
.I0(CLBLM_R_X5Y137_SLICE_X6Y137_DO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X5Y142_SLICE_X6Y142_CO6),
.I3(CLBLL_L_X4Y138_SLICE_X4Y138_BQ),
.I4(CLBLM_R_X7Y141_SLICE_X8Y141_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y138_SLICE_X5Y138_AO5),
.O6(CLBLL_L_X4Y138_SLICE_X5Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y139_SLICE_X4Y139_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y139_SLICE_X4Y139_AO6),
.Q(CLBLL_L_X4Y139_SLICE_X4Y139_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h000b000b00080008)
  ) CLBLL_L_X4Y139_SLICE_X4Y139_DLUT (
.I0(CLBLL_L_X4Y135_SLICE_X4Y135_CQ),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(CLBLM_R_X3Y143_SLICE_X2Y143_AO5),
.I3(CLBLL_L_X2Y141_SLICE_X1Y141_AO5),
.I4(1'b1),
.I5(CLBLM_R_X7Y136_SLICE_X8Y136_CQ),
.O5(CLBLL_L_X4Y139_SLICE_X4Y139_DO5),
.O6(CLBLL_L_X4Y139_SLICE_X4Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffeeffcccceeee)
  ) CLBLL_L_X4Y139_SLICE_X4Y139_CLUT (
.I0(CLBLM_L_X8Y137_SLICE_X11Y137_AQ),
.I1(CLBLL_L_X4Y139_SLICE_X5Y139_CO6),
.I2(1'b1),
.I3(CLBLL_L_X4Y143_SLICE_X5Y143_AO6),
.I4(CLBLM_R_X3Y142_SLICE_X2Y142_AO6),
.I5(CLBLL_L_X4Y139_SLICE_X5Y139_BQ),
.O5(CLBLL_L_X4Y139_SLICE_X4Y139_CO5),
.O6(CLBLL_L_X4Y139_SLICE_X4Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLL_L_X4Y139_SLICE_X4Y139_BLUT (
.I0(CLBLL_L_X4Y138_SLICE_X4Y138_DO6),
.I1(CLBLM_R_X5Y139_SLICE_X7Y139_DO6),
.I2(CLBLM_R_X5Y140_SLICE_X6Y140_CO6),
.I3(CLBLM_R_X3Y142_SLICE_X2Y142_CO6),
.I4(CLBLM_R_X5Y140_SLICE_X6Y140_BO6),
.I5(CLBLL_L_X4Y139_SLICE_X4Y139_CO6),
.O5(CLBLL_L_X4Y139_SLICE_X4Y139_BO5),
.O6(CLBLL_L_X4Y139_SLICE_X4Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff50d8000050d8)
  ) CLBLL_L_X4Y139_SLICE_X4Y139_ALUT (
.I0(CLBLL_L_X4Y138_SLICE_X5Y138_CO5),
.I1(CLBLM_R_X5Y140_SLICE_X6Y140_AO6),
.I2(CLBLL_L_X4Y139_SLICE_X4Y139_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X10Y142_SLICE_X12Y142_CQ),
.O5(CLBLL_L_X4Y139_SLICE_X4Y139_AO5),
.O6(CLBLL_L_X4Y139_SLICE_X4Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y139_SLICE_X5Y139_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y139_SLICE_X5Y139_AO6),
.Q(CLBLL_L_X4Y139_SLICE_X5Y139_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y139_SLICE_X5Y139_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y139_SLICE_X5Y139_BO6),
.Q(CLBLL_L_X4Y139_SLICE_X5Y139_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000e200e2)
  ) CLBLL_L_X4Y139_SLICE_X5Y139_DLUT (
.I0(CLBLM_R_X5Y138_SLICE_X7Y138_BQ),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(CLBLM_R_X5Y134_SLICE_X6Y134_A5Q),
.I3(CLBLL_L_X2Y141_SLICE_X1Y141_AO5),
.I4(1'b1),
.I5(CLBLL_L_X4Y143_SLICE_X5Y143_BO6),
.O5(CLBLL_L_X4Y139_SLICE_X5Y139_DO5),
.O6(CLBLL_L_X4Y139_SLICE_X5Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h000c00000000000a)
  ) CLBLL_L_X4Y139_SLICE_X5Y139_CLUT (
.I0(CLBLM_R_X7Y135_SLICE_X9Y135_AQ),
.I1(CLBLL_L_X4Y138_SLICE_X5Y138_A5Q),
.I2(CLBLL_L_X4Y143_SLICE_X5Y143_BO5),
.I3(CLBLL_L_X2Y141_SLICE_X1Y141_AO5),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(RIOB33_X105Y135_IOB_X1Y136_I),
.O5(CLBLL_L_X4Y139_SLICE_X5Y139_CO5),
.O6(CLBLL_L_X4Y139_SLICE_X5Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f40504fffc0f0c)
  ) CLBLL_L_X4Y139_SLICE_X5Y139_BLUT (
.I0(CLBLM_L_X10Y139_SLICE_X13Y139_B5Q),
.I1(CLBLL_L_X4Y139_SLICE_X5Y139_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X11Y138_SLICE_X14Y138_BQ),
.I4(CLBLM_R_X7Y139_SLICE_X8Y139_AQ),
.I5(CLBLM_L_X12Y134_SLICE_X17Y134_AO6),
.O5(CLBLL_L_X4Y139_SLICE_X5Y139_BO5),
.O6(CLBLL_L_X4Y139_SLICE_X5Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hd8ddd8ddd888d888)
  ) CLBLL_L_X4Y139_SLICE_X5Y139_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLL_L_X4Y139_SLICE_X5Y139_BQ),
.I2(CLBLL_L_X4Y139_SLICE_X5Y139_AQ),
.I3(CLBLM_L_X8Y143_SLICE_X10Y143_DO5),
.I4(1'b1),
.I5(CLBLM_R_X7Y134_SLICE_X9Y134_AQ),
.O5(CLBLL_L_X4Y139_SLICE_X5Y139_AO5),
.O6(CLBLL_L_X4Y139_SLICE_X5Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff44ffffff4444)
  ) CLBLL_L_X4Y140_SLICE_X4Y140_DLUT (
.I0(CLBLL_L_X4Y143_SLICE_X5Y143_AO6),
.I1(CLBLM_R_X5Y139_SLICE_X6Y139_BQ),
.I2(1'b1),
.I3(CLBLM_R_X3Y142_SLICE_X2Y142_AO5),
.I4(CLBLL_L_X4Y139_SLICE_X4Y139_DO6),
.I5(CLBLL_L_X4Y135_SLICE_X4Y135_BQ),
.O5(CLBLL_L_X4Y140_SLICE_X4Y140_DO5),
.O6(CLBLL_L_X4Y140_SLICE_X4Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcdcc0500ffff0500)
  ) CLBLL_L_X4Y140_SLICE_X4Y140_CLUT (
.I0(CLBLL_L_X2Y140_SLICE_X1Y140_AO6),
.I1(RIOB33_X105Y129_IOB_X1Y129_I),
.I2(CLBLM_R_X3Y143_SLICE_X2Y143_AO6),
.I3(CLBLM_L_X8Y139_SLICE_X10Y139_DQ),
.I4(CLBLM_L_X8Y140_SLICE_X10Y140_AQ),
.I5(RIOB33_X105Y137_IOB_X1Y137_I),
.O5(CLBLL_L_X4Y140_SLICE_X4Y140_CO5),
.O6(CLBLL_L_X4Y140_SLICE_X4Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0404000004045500)
  ) CLBLL_L_X4Y140_SLICE_X4Y140_BLUT (
.I0(CLBLL_L_X4Y143_SLICE_X5Y143_BO5),
.I1(CLBLM_R_X5Y139_SLICE_X6Y139_BQ),
.I2(CLBLL_L_X2Y140_SLICE_X1Y140_AO6),
.I3(CLBLL_L_X4Y135_SLICE_X4Y135_BQ),
.I4(RIOB33_X105Y135_IOB_X1Y136_I),
.I5(CLBLM_R_X3Y141_SLICE_X3Y141_AO5),
.O5(CLBLL_L_X4Y140_SLICE_X4Y140_BO5),
.O6(CLBLL_L_X4Y140_SLICE_X4Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffeefffffffe)
  ) CLBLL_L_X4Y140_SLICE_X4Y140_ALUT (
.I0(CLBLL_L_X4Y139_SLICE_X4Y139_DO6),
.I1(CLBLL_L_X4Y140_SLICE_X5Y140_DO6),
.I2(LIOB33_X0Y65_IOB_X0Y66_I),
.I3(CLBLL_L_X4Y140_SLICE_X4Y140_BO6),
.I4(CLBLL_L_X4Y140_SLICE_X4Y140_CO6),
.I5(CLBLM_R_X3Y141_SLICE_X2Y141_AO6),
.O5(CLBLL_L_X4Y140_SLICE_X4Y140_AO5),
.O6(CLBLL_L_X4Y140_SLICE_X4Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000c0c00000a0a)
  ) CLBLL_L_X4Y140_SLICE_X5Y140_DLUT (
.I0(CLBLL_L_X4Y139_SLICE_X5Y139_AQ),
.I1(RIOB33_X105Y111_IOB_X1Y111_I),
.I2(CLBLM_R_X3Y143_SLICE_X3Y143_AO5),
.I3(1'b1),
.I4(CLBLL_L_X4Y143_SLICE_X5Y143_BO5),
.I5(RIOB33_X105Y135_IOB_X1Y136_I),
.O5(CLBLL_L_X4Y140_SLICE_X5Y140_DO5),
.O6(CLBLL_L_X4Y140_SLICE_X5Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00005d5d00000c0c)
  ) CLBLL_L_X4Y140_SLICE_X5Y140_CLUT (
.I0(CLBLL_L_X2Y140_SLICE_X1Y140_AO6),
.I1(CLBLM_R_X5Y138_SLICE_X7Y138_AQ),
.I2(CLBLM_R_X3Y143_SLICE_X3Y143_AO5),
.I3(1'b1),
.I4(CLBLM_R_X3Y143_SLICE_X2Y143_AO5),
.I5(CLBLL_L_X4Y135_SLICE_X4Y135_AQ),
.O5(CLBLL_L_X4Y140_SLICE_X5Y140_CO5),
.O6(CLBLL_L_X4Y140_SLICE_X5Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff0c0caeae)
  ) CLBLL_L_X4Y140_SLICE_X5Y140_BLUT (
.I0(RIOB33_X105Y109_IOB_X1Y110_I),
.I1(CLBLM_R_X5Y136_SLICE_X7Y136_CQ),
.I2(CLBLL_L_X4Y143_SLICE_X5Y143_AO6),
.I3(1'b1),
.I4(CLBLM_R_X5Y143_SLICE_X6Y143_BO6),
.I5(CLBLL_L_X4Y140_SLICE_X5Y140_CO6),
.O5(CLBLL_L_X4Y140_SLICE_X5Y140_BO5),
.O6(CLBLL_L_X4Y140_SLICE_X5Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000040000000)
  ) CLBLL_L_X4Y140_SLICE_X5Y140_ALUT (
.I0(RIOB33_X105Y131_IOB_X1Y132_I),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(CLBLM_R_X3Y138_SLICE_X3Y138_AQ),
.I3(RIOB33_X105Y133_IOB_X1Y134_I),
.I4(RIOB33_X105Y133_IOB_X1Y133_I),
.I5(CLBLM_R_X3Y143_SLICE_X2Y143_AO6),
.O5(CLBLL_L_X4Y140_SLICE_X5Y140_AO5),
.O6(CLBLL_L_X4Y140_SLICE_X5Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffa)
  ) CLBLL_L_X4Y141_SLICE_X4Y141_DLUT (
.I0(CLBLL_L_X4Y140_SLICE_X5Y140_DO6),
.I1(1'b1),
.I2(CLBLM_R_X7Y141_SLICE_X9Y141_DO6),
.I3(CLBLL_L_X4Y141_SLICE_X4Y141_CO6),
.I4(CLBLM_R_X3Y142_SLICE_X3Y142_DO6),
.I5(CLBLL_L_X4Y140_SLICE_X4Y140_DO6),
.O5(CLBLL_L_X4Y141_SLICE_X4Y141_DO5),
.O6(CLBLL_L_X4Y141_SLICE_X4Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcf0fcc00efafeeaa)
  ) CLBLL_L_X4Y141_SLICE_X4Y141_CLUT (
.I0(LIOB33_X0Y65_IOB_X0Y66_I),
.I1(CLBLM_R_X3Y139_SLICE_X2Y139_AO5),
.I2(CLBLL_L_X4Y143_SLICE_X4Y143_AO5),
.I3(CLBLM_L_X8Y140_SLICE_X10Y140_AQ),
.I4(CLBLM_L_X8Y139_SLICE_X10Y139_DQ),
.I5(CLBLM_R_X3Y141_SLICE_X2Y141_AO6),
.O5(CLBLL_L_X4Y141_SLICE_X4Y141_CO5),
.O6(CLBLL_L_X4Y141_SLICE_X4Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffafefffffaaee)
  ) CLBLL_L_X4Y141_SLICE_X4Y141_BLUT (
.I0(CLBLL_L_X4Y143_SLICE_X4Y143_DO6),
.I1(LIOB33_X0Y67_IOB_X0Y67_I),
.I2(CLBLL_L_X4Y143_SLICE_X5Y143_AO6),
.I3(CLBLM_R_X3Y141_SLICE_X2Y141_AO6),
.I4(CLBLL_L_X4Y141_SLICE_X4Y141_AO6),
.I5(CLBLM_L_X8Y139_SLICE_X10Y139_CQ),
.O5(CLBLL_L_X4Y141_SLICE_X4Y141_BO5),
.O6(CLBLL_L_X4Y141_SLICE_X4Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0030003011110000)
  ) CLBLL_L_X4Y141_SLICE_X4Y141_ALUT (
.I0(CLBLM_R_X3Y143_SLICE_X3Y143_AO6),
.I1(CLBLL_L_X4Y143_SLICE_X5Y143_BO5),
.I2(RIOB33_X105Y111_IOB_X1Y112_I),
.I3(CLBLM_R_X3Y143_SLICE_X3Y143_AO5),
.I4(CLBLM_R_X7Y137_SLICE_X8Y137_AQ),
.I5(RIOB33_X105Y135_IOB_X1Y136_I),
.O5(CLBLL_L_X4Y141_SLICE_X4Y141_AO5),
.O6(CLBLL_L_X4Y141_SLICE_X4Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffcfffe)
  ) CLBLL_L_X4Y141_SLICE_X5Y141_DLUT (
.I0(CLBLM_R_X5Y141_SLICE_X6Y141_BQ),
.I1(CLBLL_L_X4Y139_SLICE_X5Y139_DO6),
.I2(CLBLL_L_X4Y140_SLICE_X5Y140_AO6),
.I3(CLBLL_L_X4Y141_SLICE_X5Y141_CO6),
.I4(CLBLM_R_X3Y142_SLICE_X2Y142_AO6),
.I5(CLBLM_R_X5Y141_SLICE_X7Y141_CO6),
.O5(CLBLL_L_X4Y141_SLICE_X5Y141_DO5),
.O6(CLBLL_L_X4Y141_SLICE_X5Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h000002ce00000202)
  ) CLBLL_L_X4Y141_SLICE_X5Y141_CLUT (
.I0(CLBLL_L_X4Y138_SLICE_X4Y138_AQ),
.I1(RIOB33_X105Y135_IOB_X1Y136_I),
.I2(CLBLL_L_X2Y140_SLICE_X1Y140_AO6),
.I3(CLBLM_R_X3Y143_SLICE_X3Y143_AO5),
.I4(CLBLL_L_X4Y143_SLICE_X5Y143_BO5),
.I5(RIOB33_X105Y105_IOB_X1Y106_I),
.O5(CLBLL_L_X4Y141_SLICE_X5Y141_CO5),
.O6(CLBLL_L_X4Y141_SLICE_X5Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f2f0f20022f0f2)
  ) CLBLL_L_X4Y141_SLICE_X5Y141_BLUT (
.I0(LIOB33_X0Y67_IOB_X0Y68_I),
.I1(CLBLM_R_X3Y143_SLICE_X3Y143_AO5),
.I2(CLBLL_L_X4Y138_SLICE_X5Y138_AQ),
.I3(CLBLM_R_X3Y143_SLICE_X2Y143_AO6),
.I4(RIOB33_X105Y137_IOB_X1Y137_I),
.I5(RIOB33_X105Y129_IOB_X1Y129_I),
.O5(CLBLL_L_X4Y141_SLICE_X5Y141_BO5),
.O6(CLBLL_L_X4Y141_SLICE_X5Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h73ff50ff73735050)
  ) CLBLL_L_X4Y141_SLICE_X5Y141_ALUT (
.I0(CLBLM_R_X5Y143_SLICE_X6Y143_AO6),
.I1(CLBLM_R_X5Y143_SLICE_X6Y143_BO6),
.I2(CLBLM_R_X7Y137_SLICE_X8Y137_AQ),
.I3(CLBLL_L_X4Y143_SLICE_X5Y143_AO6),
.I4(RIOB33_X105Y111_IOB_X1Y112_I),
.I5(CLBLM_L_X8Y139_SLICE_X10Y139_CQ),
.O5(CLBLL_L_X4Y141_SLICE_X5Y141_AO5),
.O6(CLBLL_L_X4Y141_SLICE_X5Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000bb00bb)
  ) CLBLL_L_X4Y142_SLICE_X4Y142_DLUT (
.I0(CLBLM_R_X3Y142_SLICE_X3Y142_BO6),
.I1(CLBLM_R_X5Y143_SLICE_X6Y143_BO5),
.I2(1'b1),
.I3(CLBLL_L_X4Y143_SLICE_X4Y143_CO6),
.I4(1'b1),
.I5(CLBLL_L_X4Y141_SLICE_X5Y141_AO6),
.O5(CLBLL_L_X4Y142_SLICE_X4Y142_DO5),
.O6(CLBLL_L_X4Y142_SLICE_X4Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff2f222f222f22)
  ) CLBLL_L_X4Y142_SLICE_X4Y142_CLUT (
.I0(CLBLM_R_X7Y141_SLICE_X9Y141_BQ),
.I1(CLBLM_R_X5Y143_SLICE_X6Y143_BO5),
.I2(CLBLM_R_X3Y142_SLICE_X2Y142_AO6),
.I3(CLBLL_L_X4Y137_SLICE_X5Y137_BQ),
.I4(CLBLL_L_X4Y137_SLICE_X4Y137_DQ),
.I5(CLBLM_R_X3Y139_SLICE_X2Y139_AO5),
.O5(CLBLL_L_X4Y142_SLICE_X4Y142_CO5),
.O6(CLBLL_L_X4Y142_SLICE_X4Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffffce)
  ) CLBLL_L_X4Y142_SLICE_X4Y142_BLUT (
.I0(CLBLM_R_X5Y143_SLICE_X6Y143_BO5),
.I1(CLBLL_L_X4Y143_SLICE_X4Y143_CO6),
.I2(CLBLM_R_X3Y142_SLICE_X3Y142_BO6),
.I3(CLBLL_L_X4Y142_SLICE_X5Y142_CO6),
.I4(CLBLL_L_X4Y141_SLICE_X5Y141_AO6),
.I5(CLBLL_L_X4Y142_SLICE_X4Y142_CO6),
.O5(CLBLL_L_X4Y142_SLICE_X4Y142_BO5),
.O6(CLBLL_L_X4Y142_SLICE_X4Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f5f0f030753030)
  ) CLBLL_L_X4Y142_SLICE_X4Y142_ALUT (
.I0(CLBLM_R_X3Y143_SLICE_X3Y143_AO6),
.I1(RIOB33_X105Y137_IOB_X1Y137_I),
.I2(CLBLL_L_X4Y137_SLICE_X4Y137_DQ),
.I3(CLBLL_L_X4Y143_SLICE_X5Y143_BO6),
.I4(CLBLM_R_X7Y141_SLICE_X9Y141_BQ),
.I5(RIOB33_X105Y129_IOB_X1Y129_I),
.O5(CLBLL_L_X4Y142_SLICE_X4Y142_AO5),
.O6(CLBLL_L_X4Y142_SLICE_X4Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLL_L_X4Y142_SLICE_X5Y142_DLUT (
.I0(CLBLM_R_X3Y142_SLICE_X2Y142_CO6),
.I1(CLBLL_L_X4Y141_SLICE_X5Y141_DO6),
.I2(CLBLL_L_X4Y143_SLICE_X5Y143_CO6),
.I3(CLBLM_R_X3Y141_SLICE_X2Y141_DO6),
.I4(CLBLM_R_X7Y142_SLICE_X8Y142_BO6),
.I5(CLBLM_R_X5Y143_SLICE_X7Y143_BO6),
.O5(CLBLL_L_X4Y142_SLICE_X5Y142_DO5),
.O6(CLBLL_L_X4Y142_SLICE_X5Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0ace0aceffff0ace)
  ) CLBLL_L_X4Y142_SLICE_X5Y142_CLUT (
.I0(CLBLM_L_X8Y142_SLICE_X11Y142_AQ),
.I1(CLBLM_R_X7Y140_SLICE_X9Y140_AQ),
.I2(CLBLL_L_X4Y143_SLICE_X5Y143_AO5),
.I3(CLBLM_R_X5Y143_SLICE_X6Y143_AO5),
.I4(CLBLM_L_X8Y142_SLICE_X10Y142_AQ),
.I5(CLBLM_R_X3Y142_SLICE_X3Y142_AO6),
.O5(CLBLL_L_X4Y142_SLICE_X5Y142_CO5),
.O6(CLBLL_L_X4Y142_SLICE_X5Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000b08000000000)
  ) CLBLL_L_X4Y142_SLICE_X5Y142_BLUT (
.I0(CLBLM_L_X8Y142_SLICE_X10Y142_AQ),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(RIOB33_X105Y133_IOB_X1Y134_I),
.I3(CLBLM_L_X8Y142_SLICE_X11Y142_AQ),
.I4(CLBLL_L_X4Y144_SLICE_X4Y144_AO6),
.I5(RIOB33_X105Y133_IOB_X1Y133_I),
.O5(CLBLL_L_X4Y142_SLICE_X5Y142_BO5),
.O6(CLBLL_L_X4Y142_SLICE_X5Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff4fff4fffffff4)
  ) CLBLL_L_X4Y142_SLICE_X5Y142_ALUT (
.I0(CLBLM_R_X3Y142_SLICE_X2Y142_AO6),
.I1(CLBLL_L_X4Y137_SLICE_X5Y137_BQ),
.I2(CLBLL_L_X4Y142_SLICE_X4Y142_AO6),
.I3(CLBLL_L_X4Y142_SLICE_X5Y142_BO6),
.I4(CLBLM_R_X7Y140_SLICE_X9Y140_AQ),
.I5(CLBLM_R_X5Y143_SLICE_X6Y143_AO5),
.O5(CLBLL_L_X4Y142_SLICE_X5Y142_AO5),
.O6(CLBLL_L_X4Y142_SLICE_X5Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000030303300)
  ) CLBLL_L_X4Y143_SLICE_X4Y143_DLUT (
.I0(1'b1),
.I1(CLBLL_L_X2Y141_SLICE_X1Y141_AO5),
.I2(CLBLM_L_X8Y143_SLICE_X10Y143_CQ),
.I3(CLBLM_R_X3Y137_SLICE_X3Y137_CQ),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(CLBLM_R_X3Y143_SLICE_X2Y143_AO6),
.O5(CLBLL_L_X4Y143_SLICE_X4Y143_DO5),
.O6(CLBLL_L_X4Y143_SLICE_X4Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h50dcffff50dc50dc)
  ) CLBLL_L_X4Y143_SLICE_X4Y143_CLUT (
.I0(CLBLL_L_X4Y143_SLICE_X4Y143_AO6),
.I1(CLBLM_R_X3Y137_SLICE_X3Y137_CQ),
.I2(CLBLM_L_X8Y143_SLICE_X10Y143_CQ),
.I3(CLBLL_L_X4Y143_SLICE_X4Y143_AO5),
.I4(CLBLM_R_X3Y141_SLICE_X2Y141_AO6),
.I5(LIOB33_X0Y67_IOB_X0Y67_I),
.O5(CLBLL_L_X4Y143_SLICE_X4Y143_CO5),
.O6(CLBLL_L_X4Y143_SLICE_X4Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffeeffffffefff)
  ) CLBLL_L_X4Y143_SLICE_X4Y143_BLUT (
.I0(CLBLM_R_X3Y143_SLICE_X2Y143_AO5),
.I1(RIOB33_X105Y133_IOB_X1Y134_I),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(RIOB33_X105Y131_IOB_X1Y132_I),
.I4(RIOB33_X105Y133_IOB_X1Y133_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y143_SLICE_X4Y143_BO5),
.O6(CLBLL_L_X4Y143_SLICE_X4Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffdfffffffef)
  ) CLBLL_L_X4Y143_SLICE_X4Y143_ALUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(RIOB33_X105Y133_IOB_X1Y133_I),
.I2(RIOB33_X105Y133_IOB_X1Y134_I),
.I3(CLBLM_R_X3Y143_SLICE_X2Y143_AO6),
.I4(RIOB33_X105Y131_IOB_X1Y132_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y143_SLICE_X4Y143_AO5),
.O6(CLBLL_L_X4Y143_SLICE_X4Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000020000000)
  ) CLBLL_L_X4Y143_SLICE_X5Y143_DLUT (
.I0(RIOB33_X105Y133_IOB_X1Y134_I),
.I1(RIOB33_X105Y131_IOB_X1Y132_I),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(CLBLL_L_X4Y136_SLICE_X5Y136_CQ),
.I4(RIOB33_X105Y133_IOB_X1Y133_I),
.I5(CLBLM_R_X3Y143_SLICE_X2Y143_AO6),
.O5(CLBLL_L_X4Y143_SLICE_X5Y143_DO5),
.O6(CLBLL_L_X4Y143_SLICE_X5Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0a0f0a00cc00cc00)
  ) CLBLL_L_X4Y143_SLICE_X5Y143_CLUT (
.I0(CLBLM_L_X10Y141_SLICE_X12Y141_AQ),
.I1(RIOB33_X105Y131_IOB_X1Y132_I),
.I2(CLBLL_L_X4Y143_SLICE_X4Y143_BO6),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(CLBLM_R_X11Y141_SLICE_X15Y141_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y143_SLICE_X5Y143_CO5),
.O6(CLBLL_L_X4Y143_SLICE_X5Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffff7fffffff3)
  ) CLBLL_L_X4Y143_SLICE_X5Y143_BLUT (
.I0(RIOB33_X105Y135_IOB_X1Y136_I),
.I1(RIOB33_X105Y137_IOB_X1Y137_I),
.I2(RIOB33_X105Y129_IOB_X1Y130_I),
.I3(RIOB33_X105Y135_IOB_X1Y135_I),
.I4(RIOB33_X105Y129_IOB_X1Y129_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y143_SLICE_X5Y143_BO5),
.O6(CLBLL_L_X4Y143_SLICE_X5Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffeffffffbfffff)
  ) CLBLL_L_X4Y143_SLICE_X5Y143_ALUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(RIOB33_X105Y131_IOB_X1Y132_I),
.I2(RIOB33_X105Y133_IOB_X1Y133_I),
.I3(CLBLL_L_X4Y143_SLICE_X5Y143_BO6),
.I4(RIOB33_X105Y133_IOB_X1Y134_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y143_SLICE_X5Y143_AO5),
.O6(CLBLL_L_X4Y143_SLICE_X5Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y144_SLICE_X4Y144_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y144_SLICE_X4Y144_DO5),
.O6(CLBLL_L_X4Y144_SLICE_X4Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y144_SLICE_X4Y144_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y144_SLICE_X4Y144_CO5),
.O6(CLBLL_L_X4Y144_SLICE_X4Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y144_SLICE_X4Y144_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y144_SLICE_X4Y144_BO5),
.O6(CLBLL_L_X4Y144_SLICE_X4Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffff7ffffffff)
  ) CLBLL_L_X4Y144_SLICE_X4Y144_ALUT (
.I0(RIOB33_X105Y137_IOB_X1Y137_I),
.I1(RIOB33_X105Y131_IOB_X1Y132_I),
.I2(RIOB33_X105Y129_IOB_X1Y130_I),
.I3(RIOB33_X105Y135_IOB_X1Y135_I),
.I4(RIOB33_X105Y129_IOB_X1Y129_I),
.I5(RIOB33_X105Y135_IOB_X1Y136_I),
.O5(CLBLL_L_X4Y144_SLICE_X4Y144_AO5),
.O6(CLBLL_L_X4Y144_SLICE_X4Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y144_SLICE_X5Y144_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y144_SLICE_X5Y144_DO5),
.O6(CLBLL_L_X4Y144_SLICE_X5Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y144_SLICE_X5Y144_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y144_SLICE_X5Y144_CO5),
.O6(CLBLL_L_X4Y144_SLICE_X5Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y144_SLICE_X5Y144_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y144_SLICE_X5Y144_BO5),
.O6(CLBLL_L_X4Y144_SLICE_X5Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y144_SLICE_X5Y144_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y144_SLICE_X5Y144_AO5),
.O6(CLBLL_L_X4Y144_SLICE_X5Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y126_SLICE_X78Y126_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y126_SLICE_X78Y126_DO5),
.O6(CLBLL_L_X52Y126_SLICE_X78Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y126_SLICE_X78Y126_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y126_SLICE_X78Y126_CO5),
.O6(CLBLL_L_X52Y126_SLICE_X78Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y126_SLICE_X78Y126_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y126_SLICE_X78Y126_BO5),
.O6(CLBLL_L_X52Y126_SLICE_X78Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00ff00ff00ff)
  ) CLBLL_L_X52Y126_SLICE_X78Y126_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(RIOB33_X105Y123_IOB_X1Y124_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y126_SLICE_X78Y126_AO5),
.O6(CLBLL_L_X52Y126_SLICE_X78Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y126_SLICE_X79Y126_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y126_SLICE_X79Y126_DO5),
.O6(CLBLL_L_X52Y126_SLICE_X79Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y126_SLICE_X79Y126_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y126_SLICE_X79Y126_CO5),
.O6(CLBLL_L_X52Y126_SLICE_X79Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y126_SLICE_X79Y126_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y126_SLICE_X79Y126_BO5),
.O6(CLBLL_L_X52Y126_SLICE_X79Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y126_SLICE_X79Y126_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y126_SLICE_X79Y126_AO5),
.O6(CLBLL_L_X52Y126_SLICE_X79Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y131_SLICE_X10Y131_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y131_SLICE_X10Y131_BO6),
.Q(CLBLM_L_X8Y131_SLICE_X10Y131_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y131_SLICE_X10Y131_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y131_SLICE_X10Y131_AO6),
.Q(CLBLM_L_X8Y131_SLICE_X10Y131_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y131_SLICE_X10Y131_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y131_SLICE_X10Y131_DO5),
.O6(CLBLM_L_X8Y131_SLICE_X10Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5faf5faff5faf5fa)
  ) CLBLM_L_X8Y131_SLICE_X10Y131_CLUT (
.I0(CLBLM_L_X10Y131_SLICE_X13Y131_AQ),
.I1(1'b1),
.I2(CLBLM_L_X10Y137_SLICE_X12Y137_BQ),
.I3(CLBLM_L_X8Y135_SLICE_X11Y135_AQ),
.I4(1'b1),
.I5(CLBLL_L_X4Y132_SLICE_X5Y132_AQ),
.O5(CLBLM_L_X8Y131_SLICE_X10Y131_CO5),
.O6(CLBLM_L_X8Y131_SLICE_X10Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcf03ce0200005555)
  ) CLBLM_L_X8Y131_SLICE_X10Y131_BLUT (
.I0(CLBLM_L_X8Y131_SLICE_X11Y131_BQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X5Y132_SLICE_X7Y132_DO6),
.I3(CLBLM_L_X8Y135_SLICE_X11Y135_BQ),
.I4(CLBLM_L_X8Y131_SLICE_X10Y131_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X8Y131_SLICE_X10Y131_BO5),
.O6(CLBLM_L_X8Y131_SLICE_X10Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc55cc55cc50cc50)
  ) CLBLM_L_X8Y131_SLICE_X10Y131_ALUT (
.I0(CLBLM_R_X5Y133_SLICE_X7Y133_DO6),
.I1(CLBLM_L_X10Y137_SLICE_X12Y137_BQ),
.I2(CLBLM_L_X8Y131_SLICE_X10Y131_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLL_L_X4Y132_SLICE_X5Y132_AQ),
.O5(CLBLM_L_X8Y131_SLICE_X10Y131_AO5),
.O6(CLBLM_L_X8Y131_SLICE_X10Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y131_SLICE_X11Y131_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y131_SLICE_X11Y131_AO6),
.Q(CLBLM_L_X8Y131_SLICE_X11Y131_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y131_SLICE_X11Y131_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y131_SLICE_X11Y131_BO6),
.Q(CLBLM_L_X8Y131_SLICE_X11Y131_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h2100002121000021)
  ) CLBLM_L_X8Y131_SLICE_X11Y131_DLUT (
.I0(CLBLM_L_X8Y132_SLICE_X10Y132_AQ),
.I1(CLBLM_L_X8Y131_SLICE_X10Y131_CO6),
.I2(CLBLM_L_X10Y137_SLICE_X12Y137_B5Q),
.I3(CLBLM_L_X8Y133_SLICE_X10Y133_CQ),
.I4(CLBLM_R_X11Y146_SLICE_X14Y146_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y131_SLICE_X11Y131_DO5),
.O6(CLBLM_L_X8Y131_SLICE_X11Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000001)
  ) CLBLM_L_X8Y131_SLICE_X11Y131_CLUT (
.I0(CLBLM_L_X8Y132_SLICE_X11Y132_AQ),
.I1(CLBLM_L_X8Y132_SLICE_X10Y132_AQ),
.I2(CLBLM_L_X8Y131_SLICE_X10Y131_AQ),
.I3(CLBLM_L_X8Y133_SLICE_X10Y133_CQ),
.I4(CLBLM_L_X8Y131_SLICE_X11Y131_AQ),
.I5(CLBLM_L_X10Y131_SLICE_X13Y131_AQ),
.O5(CLBLM_L_X8Y131_SLICE_X11Y131_CO5),
.O6(CLBLM_L_X8Y131_SLICE_X11Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00ff55ee44)
  ) CLBLM_L_X8Y131_SLICE_X11Y131_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y131_SLICE_X11Y131_BQ),
.I2(1'b1),
.I3(CLBLM_R_X7Y134_SLICE_X8Y134_BQ),
.I4(CLBLM_R_X11Y132_SLICE_X15Y132_CO6),
.I5(CLBLM_R_X5Y133_SLICE_X7Y133_DO6),
.O5(CLBLM_L_X8Y131_SLICE_X11Y131_BO5),
.O6(CLBLM_L_X8Y131_SLICE_X11Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88bb88bb88bb8888)
  ) CLBLM_L_X8Y131_SLICE_X11Y131_ALUT (
.I0(CLBLM_R_X7Y132_SLICE_X9Y132_DQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(1'b1),
.I3(CLBLM_R_X5Y133_SLICE_X7Y133_DO6),
.I4(CLBLM_L_X8Y132_SLICE_X11Y132_AQ),
.I5(CLBLM_L_X8Y131_SLICE_X11Y131_AQ),
.O5(CLBLM_L_X8Y131_SLICE_X11Y131_AO5),
.O6(CLBLM_L_X8Y131_SLICE_X11Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y132_SLICE_X10Y132_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y132_SLICE_X10Y132_AO6),
.Q(CLBLM_L_X8Y132_SLICE_X10Y132_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y132_SLICE_X10Y132_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y132_SLICE_X10Y132_BO6),
.Q(CLBLM_L_X8Y132_SLICE_X10Y132_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaaa66aaaa)
  ) CLBLM_L_X8Y132_SLICE_X10Y132_DLUT (
.I0(CLBLM_R_X11Y133_SLICE_X15Y133_BQ),
.I1(CLBLM_L_X10Y130_SLICE_X12Y130_AQ),
.I2(1'b1),
.I3(CLBLM_L_X10Y131_SLICE_X12Y131_BQ),
.I4(CLBLL_L_X4Y135_SLICE_X5Y135_CQ),
.I5(CLBLM_R_X11Y131_SLICE_X15Y131_BQ),
.O5(CLBLM_L_X8Y132_SLICE_X10Y132_DO5),
.O6(CLBLM_L_X8Y132_SLICE_X10Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ddd0dddfdddf)
  ) CLBLM_L_X8Y132_SLICE_X10Y132_CLUT (
.I0(CLBLM_L_X8Y132_SLICE_X10Y132_DO6),
.I1(CLBLM_R_X5Y133_SLICE_X7Y133_AO6),
.I2(CLBLM_R_X7Y133_SLICE_X9Y133_DO6),
.I3(CLBLM_R_X5Y136_SLICE_X7Y136_DO6),
.I4(CLBLM_R_X5Y133_SLICE_X7Y133_CO6),
.I5(CLBLM_R_X7Y134_SLICE_X8Y134_C5Q),
.O5(CLBLM_L_X8Y132_SLICE_X10Y132_CO5),
.O6(CLBLM_L_X8Y132_SLICE_X10Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000aaaafc00)
  ) CLBLM_L_X8Y132_SLICE_X10Y132_BLUT (
.I0(CLBLM_L_X10Y137_SLICE_X12Y137_AQ),
.I1(CLBLM_L_X8Y132_SLICE_X10Y132_BQ),
.I2(CLBLM_L_X12Y132_SLICE_X17Y132_AQ),
.I3(CLBLM_L_X8Y138_SLICE_X10Y138_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_L_X8Y132_SLICE_X10Y132_BO5),
.O6(CLBLM_L_X8Y132_SLICE_X10Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00ff33cc00fc30)
  ) CLBLM_L_X8Y132_SLICE_X10Y132_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X8Y132_SLICE_X10Y132_AQ),
.I3(CLBLM_L_X8Y140_SLICE_X10Y140_BQ),
.I4(CLBLM_R_X5Y134_SLICE_X7Y134_DO6),
.I5(CLBLM_L_X10Y132_SLICE_X12Y132_BO6),
.O5(CLBLM_L_X8Y132_SLICE_X10Y132_AO5),
.O6(CLBLM_L_X8Y132_SLICE_X10Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y132_SLICE_X11Y132_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y132_SLICE_X11Y132_AO6),
.Q(CLBLM_L_X8Y132_SLICE_X11Y132_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y132_SLICE_X11Y132_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y132_SLICE_X11Y132_BO6),
.Q(CLBLM_L_X8Y132_SLICE_X11Y132_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y132_SLICE_X11Y132_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y132_SLICE_X11Y132_CO6),
.Q(CLBLM_L_X8Y132_SLICE_X11Y132_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffffbb)
  ) CLBLM_L_X8Y132_SLICE_X11Y132_DLUT (
.I0(CLBLL_L_X4Y132_SLICE_X5Y132_AQ),
.I1(CLBLM_L_X8Y131_SLICE_X11Y131_CO6),
.I2(1'b1),
.I3(CLBLM_L_X8Y133_SLICE_X10Y133_BQ),
.I4(CLBLM_R_X11Y132_SLICE_X15Y132_DO6),
.I5(CLBLM_L_X10Y133_SLICE_X12Y133_AQ),
.O5(CLBLM_L_X8Y132_SLICE_X11Y132_DO5),
.O6(CLBLM_L_X8Y132_SLICE_X11Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000000a800a8)
  ) CLBLM_L_X8Y132_SLICE_X11Y132_CLUT (
.I0(CLBLM_L_X8Y138_SLICE_X10Y138_AQ),
.I1(CLBLM_L_X8Y132_SLICE_X11Y132_CQ),
.I2(CLBLM_L_X8Y133_SLICE_X11Y133_CQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLL_L_X4Y136_SLICE_X4Y136_DQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y132_SLICE_X11Y132_CO5),
.O6(CLBLM_L_X8Y132_SLICE_X11Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa0afa0afa0afc0c)
  ) CLBLM_L_X8Y132_SLICE_X11Y132_BLUT (
.I0(CLBLM_L_X8Y132_SLICE_X11Y132_CQ),
.I1(CLBLM_L_X8Y132_SLICE_X11Y132_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y133_SLICE_X12Y133_AQ),
.I4(CLBLM_L_X8Y138_SLICE_X10Y138_AQ),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_L_X8Y132_SLICE_X11Y132_BO5),
.O6(CLBLM_L_X8Y132_SLICE_X11Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa33aa33aa30aa30)
  ) CLBLM_L_X8Y132_SLICE_X11Y132_ALUT (
.I0(CLBLM_L_X8Y132_SLICE_X11Y132_CQ),
.I1(CLBLM_R_X5Y133_SLICE_X7Y133_DO6),
.I2(CLBLM_L_X8Y132_SLICE_X11Y132_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLM_L_X8Y133_SLICE_X10Y133_BQ),
.O5(CLBLM_L_X8Y132_SLICE_X11Y132_AO5),
.O6(CLBLM_L_X8Y132_SLICE_X11Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y133_SLICE_X10Y133_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y133_SLICE_X10Y133_AO6),
.Q(CLBLM_L_X8Y133_SLICE_X10Y133_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y133_SLICE_X10Y133_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y133_SLICE_X10Y133_BO6),
.Q(CLBLM_L_X8Y133_SLICE_X10Y133_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y133_SLICE_X10Y133_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y133_SLICE_X10Y133_CO6),
.Q(CLBLM_L_X8Y133_SLICE_X10Y133_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h1300131313001313)
  ) CLBLM_L_X8Y133_SLICE_X10Y133_DLUT (
.I0(CLBLM_R_X5Y132_SLICE_X7Y132_DO6),
.I1(CLBLM_L_X8Y133_SLICE_X10Y133_AQ),
.I2(CLBLM_R_X7Y134_SLICE_X8Y134_C5Q),
.I3(CLBLM_R_X5Y133_SLICE_X7Y133_DO6),
.I4(CLBLM_L_X8Y132_SLICE_X10Y132_DO6),
.I5(1'b1),
.O5(CLBLM_L_X8Y133_SLICE_X10Y133_DO5),
.O6(CLBLM_L_X8Y133_SLICE_X10Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5f4f405050404)
  ) CLBLM_L_X8Y133_SLICE_X10Y133_CLUT (
.I0(CLBLM_R_X5Y134_SLICE_X7Y134_DO6),
.I1(CLBLM_L_X8Y133_SLICE_X10Y133_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(CLBLM_L_X8Y132_SLICE_X10Y132_AQ),
.I5(CLBLM_L_X8Y133_SLICE_X10Y133_AQ),
.O5(CLBLM_L_X8Y133_SLICE_X10Y133_CO5),
.O6(CLBLM_L_X8Y133_SLICE_X10Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00aafcaafc)
  ) CLBLM_L_X8Y133_SLICE_X10Y133_BLUT (
.I0(CLBLM_R_X5Y137_SLICE_X7Y137_B5Q),
.I1(CLBLM_L_X8Y133_SLICE_X10Y133_BQ),
.I2(CLBLM_L_X8Y131_SLICE_X10Y131_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLM_R_X5Y133_SLICE_X7Y133_DO6),
.O5(CLBLM_L_X8Y133_SLICE_X10Y133_BO5),
.O6(CLBLM_L_X8Y133_SLICE_X10Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hddddccdd11110011)
  ) CLBLM_L_X8Y133_SLICE_X10Y133_ALUT (
.I0(CLBLM_L_X8Y133_SLICE_X10Y133_DO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(1'b1),
.I3(RIOB33_X105Y141_IOB_X1Y142_I),
.I4(CLBLM_R_X7Y131_SLICE_X9Y131_AQ),
.I5(CLBLM_L_X10Y139_SLICE_X13Y139_B5Q),
.O5(CLBLM_L_X8Y133_SLICE_X10Y133_AO5),
.O6(CLBLM_L_X8Y133_SLICE_X10Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y133_SLICE_X11Y133_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y133_SLICE_X11Y133_AO6),
.Q(CLBLM_L_X8Y133_SLICE_X11Y133_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y133_SLICE_X11Y133_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y133_SLICE_X11Y133_BO6),
.Q(CLBLM_L_X8Y133_SLICE_X11Y133_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y133_SLICE_X11Y133_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y133_SLICE_X11Y133_CO6),
.Q(CLBLM_L_X8Y133_SLICE_X11Y133_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h000001ab000054fe)
  ) CLBLM_L_X8Y133_SLICE_X11Y133_DLUT (
.I0(CLBLM_R_X5Y132_SLICE_X7Y132_DO6),
.I1(CLBLM_R_X11Y131_SLICE_X15Y131_BQ),
.I2(CLBLM_L_X10Y133_SLICE_X12Y133_DO6),
.I3(CLBLM_L_X10Y141_SLICE_X12Y141_CQ),
.I4(CLBLM_L_X8Y134_SLICE_X11Y134_DQ),
.I5(CLBLM_L_X8Y137_SLICE_X11Y137_BQ),
.O5(CLBLM_L_X8Y133_SLICE_X11Y133_DO5),
.O6(CLBLM_L_X8Y133_SLICE_X11Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f000fff0f00033)
  ) CLBLM_L_X8Y133_SLICE_X11Y133_CLUT (
.I0(1'b1),
.I1(RIOB33_X105Y141_IOB_X1Y142_I),
.I2(CLBLM_R_X7Y142_SLICE_X9Y142_BQ),
.I3(CLBLM_L_X10Y131_SLICE_X12Y131_DO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y131_SLICE_X9Y131_AQ),
.O5(CLBLM_L_X8Y133_SLICE_X11Y133_CO5),
.O6(CLBLM_L_X8Y133_SLICE_X11Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0f5a0f5a0)
  ) CLBLM_L_X8Y133_SLICE_X11Y133_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(1'b1),
.I2(CLBLM_R_X5Y132_SLICE_X7Y132_AQ),
.I3(CLBLM_R_X13Y137_SLICE_X18Y137_AQ),
.I4(1'b1),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X8Y133_SLICE_X11Y133_BO5),
.O6(CLBLM_L_X8Y133_SLICE_X11Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffa50ea40)
  ) CLBLM_L_X8Y133_SLICE_X11Y133_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y138_SLICE_X10Y138_AQ),
.I2(CLBLM_L_X8Y133_SLICE_X11Y133_AQ),
.I3(CLBLM_L_X10Y131_SLICE_X13Y131_BQ),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLM_L_X8Y134_SLICE_X10Y134_CO6),
.O5(CLBLM_L_X8Y133_SLICE_X11Y133_AO5),
.O6(CLBLM_L_X8Y133_SLICE_X11Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y134_SLICE_X10Y134_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y134_SLICE_X13Y134_CO6),
.Q(CLBLM_L_X8Y134_SLICE_X10Y134_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y134_SLICE_X10Y134_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y134_SLICE_X10Y134_AO6),
.Q(CLBLM_L_X8Y134_SLICE_X10Y134_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hefff500000000000)
  ) CLBLM_L_X8Y134_SLICE_X10Y134_DLUT (
.I0(CLBLM_R_X5Y132_SLICE_X7Y132_DO6),
.I1(CLBLM_L_X10Y131_SLICE_X12Y131_BQ),
.I2(CLBLM_L_X10Y130_SLICE_X12Y130_AQ),
.I3(CLBLM_R_X11Y131_SLICE_X15Y131_BQ),
.I4(CLBLL_L_X4Y135_SLICE_X5Y135_CQ),
.I5(CLBLM_L_X8Y134_SLICE_X10Y134_BO6),
.O5(CLBLM_L_X8Y134_SLICE_X10Y134_DO5),
.O6(CLBLM_L_X8Y134_SLICE_X10Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ee00ae00ea00aa)
  ) CLBLM_L_X8Y134_SLICE_X10Y134_CLUT (
.I0(CLBLM_L_X8Y137_SLICE_X11Y137_CO5),
.I1(CLBLL_L_X4Y139_SLICE_X4Y139_BO6),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLM_R_X7Y134_SLICE_X9Y134_DO6),
.I4(CLBLM_R_X11Y136_SLICE_X15Y136_BQ),
.I5(CLBLM_L_X8Y135_SLICE_X10Y135_AQ),
.O5(CLBLM_L_X8Y134_SLICE_X10Y134_CO5),
.O6(CLBLM_L_X8Y134_SLICE_X10Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h000f0000aa00aacc)
  ) CLBLM_L_X8Y134_SLICE_X10Y134_BLUT (
.I0(CLBLL_L_X4Y136_SLICE_X4Y136_CQ),
.I1(CLBLM_R_X7Y133_SLICE_X8Y133_BQ),
.I2(CLBLM_R_X11Y140_SLICE_X15Y140_CQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y134_SLICE_X10Y134_BO5),
.O6(CLBLM_L_X8Y134_SLICE_X10Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa33300000)
  ) CLBLM_L_X8Y134_SLICE_X10Y134_ALUT (
.I0(CLBLM_R_X11Y135_SLICE_X15Y135_AQ),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_L_X8Y134_SLICE_X10Y134_AQ),
.I3(CLBLM_L_X8Y133_SLICE_X10Y133_AQ),
.I4(CLBLM_L_X8Y138_SLICE_X10Y138_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y134_SLICE_X10Y134_AO5),
.O6(CLBLM_L_X8Y134_SLICE_X10Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y134_SLICE_X11Y134_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y134_SLICE_X11Y134_AO6),
.Q(CLBLM_L_X8Y134_SLICE_X11Y134_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y134_SLICE_X11Y134_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y134_SLICE_X11Y134_BO6),
.Q(CLBLM_L_X8Y134_SLICE_X11Y134_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y134_SLICE_X11Y134_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y134_SLICE_X11Y134_CO6),
.Q(CLBLM_L_X8Y134_SLICE_X11Y134_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y134_SLICE_X11Y134_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y134_SLICE_X11Y134_DO6),
.Q(CLBLM_L_X8Y134_SLICE_X11Y134_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f022223333)
  ) CLBLM_L_X8Y134_SLICE_X11Y134_DLUT (
.I0(CLBLM_R_X7Y131_SLICE_X9Y131_AQ),
.I1(CLBLM_L_X8Y133_SLICE_X11Y133_DO6),
.I2(CLBLM_L_X8Y140_SLICE_X11Y140_AQ),
.I3(1'b1),
.I4(RIOB33_X105Y141_IOB_X1Y142_I),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y134_SLICE_X11Y134_DO5),
.O6(CLBLM_L_X8Y134_SLICE_X11Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000fa0af808)
  ) CLBLM_L_X8Y134_SLICE_X11Y134_CLUT (
.I0(CLBLM_L_X8Y138_SLICE_X10Y138_AQ),
.I1(CLBLM_L_X8Y134_SLICE_X11Y134_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X5Y137_SLICE_X6Y137_BQ),
.I4(CLBLM_R_X11Y133_SLICE_X15Y133_DQ),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_L_X8Y134_SLICE_X11Y134_CO5),
.O6(CLBLM_L_X8Y134_SLICE_X11Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haf05af05ae04ae04)
  ) CLBLM_L_X8Y134_SLICE_X11Y134_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y134_SLICE_X11Y134_BQ),
.I2(CLBLM_R_X5Y134_SLICE_X7Y134_DO6),
.I3(CLBLM_R_X5Y136_SLICE_X6Y136_BQ),
.I4(1'b1),
.I5(CLBLM_L_X8Y133_SLICE_X10Y133_CQ),
.O5(CLBLM_L_X8Y134_SLICE_X11Y134_BO5),
.O6(CLBLM_L_X8Y134_SLICE_X11Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3c0f3c0f3c0e2e2)
  ) CLBLM_L_X8Y134_SLICE_X11Y134_ALUT (
.I0(CLBLM_L_X8Y134_SLICE_X11Y134_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X7Y132_SLICE_X9Y132_BQ),
.I3(CLBLM_R_X7Y132_SLICE_X9Y132_CQ),
.I4(CLBLM_L_X8Y138_SLICE_X10Y138_AQ),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_L_X8Y134_SLICE_X11Y134_AO5),
.O6(CLBLM_L_X8Y134_SLICE_X11Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y135_SLICE_X10Y135_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y135_SLICE_X13Y135_AO6),
.Q(CLBLM_L_X8Y135_SLICE_X10Y135_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y135_SLICE_X10Y135_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y135_SLICE_X10Y135_AO6),
.Q(CLBLM_L_X8Y135_SLICE_X10Y135_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y135_SLICE_X10Y135_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y135_SLICE_X10Y135_BO6),
.Q(CLBLM_L_X8Y135_SLICE_X10Y135_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000800000)
  ) CLBLM_L_X8Y135_SLICE_X10Y135_DLUT (
.I0(CLBLM_L_X8Y135_SLICE_X10Y135_CO5),
.I1(RIOB33_X105Y121_IOB_X1Y121_I),
.I2(CLBLM_L_X10Y137_SLICE_X12Y137_AQ),
.I3(CLBLM_R_X11Y132_SLICE_X15Y132_DO6),
.I4(CLBLM_L_X8Y135_SLICE_X11Y135_DO5),
.I5(CLBLM_R_X5Y135_SLICE_X6Y135_AQ),
.O5(CLBLM_L_X8Y135_SLICE_X10Y135_DO5),
.O6(CLBLM_L_X8Y135_SLICE_X10Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h505050500000f0c0)
  ) CLBLM_L_X8Y135_SLICE_X10Y135_CLUT (
.I0(CLBLM_R_X3Y140_SLICE_X2Y140_DO6),
.I1(CLBLM_R_X11Y135_SLICE_X15Y135_AQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_L_X8Y135_SLICE_X11Y135_CQ),
.I4(CLBLM_R_X11Y136_SLICE_X14Y136_DQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y135_SLICE_X10Y135_CO5),
.O6(CLBLM_L_X8Y135_SLICE_X10Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0ccf0ccf000f000)
  ) CLBLM_L_X8Y135_SLICE_X10Y135_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y135_SLICE_X10Y135_BQ),
.I2(CLBLM_L_X8Y135_SLICE_X10Y135_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X8Y135_SLICE_X10Y135_BO5),
.O6(CLBLM_L_X8Y135_SLICE_X10Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hddd8ddd8ddd88888)
  ) CLBLM_L_X8Y135_SLICE_X10Y135_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X11Y135_SLICE_X14Y135_BQ),
.I2(CLBLM_L_X8Y135_SLICE_X10Y135_AQ),
.I3(CLBLM_L_X10Y137_SLICE_X13Y137_CO6),
.I4(CLBLM_L_X8Y138_SLICE_X10Y138_AQ),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_L_X8Y135_SLICE_X10Y135_AO5),
.O6(CLBLM_L_X8Y135_SLICE_X10Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y135_SLICE_X11Y135_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y135_SLICE_X11Y135_AO5),
.Q(CLBLM_L_X8Y135_SLICE_X11Y135_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y135_SLICE_X11Y135_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y135_SLICE_X11Y135_BO5),
.Q(CLBLM_L_X8Y135_SLICE_X11Y135_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y135_SLICE_X11Y135_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y135_SLICE_X11Y135_AO6),
.Q(CLBLM_L_X8Y135_SLICE_X11Y135_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y135_SLICE_X11Y135_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y135_SLICE_X11Y135_BO6),
.Q(CLBLM_L_X8Y135_SLICE_X11Y135_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y135_SLICE_X11Y135_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y135_SLICE_X11Y135_CO6),
.Q(CLBLM_L_X8Y135_SLICE_X11Y135_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0a0c0800003333)
  ) CLBLM_L_X8Y135_SLICE_X11Y135_DLUT (
.I0(CLBLL_L_X4Y134_SLICE_X4Y134_AQ),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y134_SLICE_X12Y134_CQ),
.I4(CLBLM_L_X8Y138_SLICE_X10Y138_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y135_SLICE_X11Y135_DO5),
.O6(CLBLM_L_X8Y135_SLICE_X11Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccdd0011cccc0000)
  ) CLBLM_L_X8Y135_SLICE_X11Y135_CLUT (
.I0(CLBLM_L_X10Y136_SLICE_X13Y136_AO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(1'b1),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_L_X8Y135_SLICE_X11Y135_B5Q),
.I5(CLBLM_R_X13Y137_SLICE_X18Y137_AQ),
.O5(CLBLM_L_X8Y135_SLICE_X11Y135_CO5),
.O6(CLBLM_L_X8Y135_SLICE_X11Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0aaf0aaccaaccaa)
  ) CLBLM_L_X8Y135_SLICE_X11Y135_BLUT (
.I0(RIOB33_X105Y125_IOB_X1Y126_I),
.I1(CLBLM_L_X12Y142_SLICE_X16Y142_AQ),
.I2(CLBLM_R_X3Y136_SLICE_X3Y136_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y135_SLICE_X11Y135_BO5),
.O6(CLBLM_L_X8Y135_SLICE_X11Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafa5050ee44aa00)
  ) CLBLM_L_X8Y135_SLICE_X11Y135_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_L_X8Y135_SLICE_X10Y135_A5Q),
.I3(CLBLM_R_X11Y134_SLICE_X14Y134_AQ),
.I4(CLBLM_L_X8Y136_SLICE_X10Y136_CQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y135_SLICE_X11Y135_AO5),
.O6(CLBLM_L_X8Y135_SLICE_X11Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y136_SLICE_X10Y136_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y136_SLICE_X10Y136_AO6),
.Q(CLBLM_L_X8Y136_SLICE_X10Y136_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y136_SLICE_X10Y136_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y136_SLICE_X10Y136_BO6),
.Q(CLBLM_L_X8Y136_SLICE_X10Y136_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y136_SLICE_X10Y136_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y136_SLICE_X10Y136_CO6),
.Q(CLBLM_L_X8Y136_SLICE_X10Y136_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y136_SLICE_X10Y136_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y136_SLICE_X10Y136_DO6),
.Q(CLBLM_L_X8Y136_SLICE_X10Y136_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffccffccfff0ffa0)
  ) CLBLM_L_X8Y136_SLICE_X10Y136_DLUT (
.I0(CLBLM_L_X8Y138_SLICE_X10Y138_AQ),
.I1(CLBLM_R_X5Y137_SLICE_X7Y137_CQ),
.I2(CLBLM_L_X8Y136_SLICE_X10Y136_DQ),
.I3(CLBLM_R_X7Y134_SLICE_X9Y134_CO6),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y136_SLICE_X10Y136_DO5),
.O6(CLBLM_L_X8Y136_SLICE_X10Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff00000a0a0a0a)
  ) CLBLM_L_X8Y136_SLICE_X10Y136_CLUT (
.I0(CLBLM_L_X10Y135_SLICE_X13Y135_B5Q),
.I1(1'b1),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(1'b1),
.I4(CLBLM_L_X8Y139_SLICE_X10Y139_DQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y136_SLICE_X10Y136_CO5),
.O6(CLBLM_L_X8Y136_SLICE_X10Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffc8ff00ffc8)
  ) CLBLM_L_X8Y136_SLICE_X10Y136_BLUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_L_X8Y136_SLICE_X10Y136_BQ),
.I2(CLBLM_L_X8Y138_SLICE_X10Y138_AQ),
.I3(CLBLM_L_X10Y136_SLICE_X13Y136_BO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y132_SLICE_X9Y132_D5Q),
.O5(CLBLM_L_X8Y136_SLICE_X10Y136_BO5),
.O6(CLBLM_L_X8Y136_SLICE_X10Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff72fff0007200f0)
  ) CLBLM_L_X8Y136_SLICE_X10Y136_ALUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_L_X8Y135_SLICE_X10Y135_CO6),
.I2(CLBLM_L_X8Y136_SLICE_X10Y136_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y138_SLICE_X10Y138_AQ),
.I5(CLBLL_L_X4Y137_SLICE_X4Y137_CQ),
.O5(CLBLM_L_X8Y136_SLICE_X10Y136_AO5),
.O6(CLBLM_L_X8Y136_SLICE_X10Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y136_SLICE_X11Y136_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y136_SLICE_X11Y136_AO6),
.Q(CLBLM_L_X8Y136_SLICE_X11Y136_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y136_SLICE_X11Y136_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y136_SLICE_X11Y136_BO6),
.Q(CLBLM_L_X8Y136_SLICE_X11Y136_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y136_SLICE_X11Y136_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y136_SLICE_X11Y136_CO6),
.Q(CLBLM_L_X8Y136_SLICE_X11Y136_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'heeee0000000fffff)
  ) CLBLM_L_X8Y136_SLICE_X11Y136_DLUT (
.I0(CLBLM_L_X10Y135_SLICE_X13Y135_B5Q),
.I1(CLBLM_L_X10Y138_SLICE_X13Y138_CQ),
.I2(CLBLM_L_X8Y136_SLICE_X11Y136_BQ),
.I3(CLBLM_R_X5Y137_SLICE_X7Y137_CQ),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y136_SLICE_X11Y136_DO5),
.O6(CLBLM_L_X8Y136_SLICE_X11Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0000033cc)
  ) CLBLM_L_X8Y136_SLICE_X11Y136_CLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y137_SLICE_X11Y137_DO6),
.I2(CLBLM_L_X8Y134_SLICE_X11Y134_AQ),
.I3(CLBLM_L_X10Y137_SLICE_X13Y137_AQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y136_SLICE_X11Y136_CO5),
.O6(CLBLM_L_X8Y136_SLICE_X11Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55fa50ee44ea40)
  ) CLBLM_L_X8Y136_SLICE_X11Y136_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y136_SLICE_X11Y136_BQ),
.I2(CLBLM_L_X8Y138_SLICE_X10Y138_AQ),
.I3(CLBLM_R_X3Y137_SLICE_X3Y137_BQ),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLM_L_X10Y138_SLICE_X12Y138_CO6),
.O5(CLBLM_L_X8Y136_SLICE_X11Y136_BO5),
.O6(CLBLM_L_X8Y136_SLICE_X11Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff050005ff0a000a)
  ) CLBLM_L_X8Y136_SLICE_X11Y136_ALUT (
.I0(CLBLM_R_X7Y138_SLICE_X8Y138_CQ),
.I1(1'b1),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y132_SLICE_X11Y132_AQ),
.I5(CLBLM_L_X8Y138_SLICE_X11Y138_CO6),
.O5(CLBLM_L_X8Y136_SLICE_X11Y136_AO5),
.O6(CLBLM_L_X8Y136_SLICE_X11Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y137_SLICE_X10Y137_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y137_SLICE_X10Y137_AO6),
.Q(CLBLM_L_X8Y137_SLICE_X10Y137_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000008000)
  ) CLBLM_L_X8Y137_SLICE_X10Y137_DLUT (
.I0(CLBLM_R_X7Y137_SLICE_X8Y137_DO6),
.I1(CLBLM_L_X10Y136_SLICE_X12Y136_CO6),
.I2(CLBLM_L_X8Y135_SLICE_X10Y135_DO6),
.I3(CLBLM_R_X5Y135_SLICE_X7Y135_CO5),
.I4(CLBLM_L_X8Y137_SLICE_X10Y137_BO5),
.I5(CLBLM_L_X10Y145_SLICE_X12Y145_CO6),
.O5(CLBLM_L_X8Y137_SLICE_X10Y137_DO5),
.O6(CLBLM_L_X8Y137_SLICE_X10Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000100033332333)
  ) CLBLM_L_X8Y137_SLICE_X10Y137_CLUT (
.I0(CLBLM_L_X10Y139_SLICE_X13Y139_AQ),
.I1(CLBLL_L_X4Y136_SLICE_X5Y136_A5Q),
.I2(CLBLM_R_X5Y136_SLICE_X7Y136_BQ),
.I3(CLBLM_R_X7Y136_SLICE_X9Y136_CQ),
.I4(CLBLM_R_X11Y139_SLICE_X15Y139_CQ),
.I5(CLBLM_L_X8Y135_SLICE_X10Y135_BQ),
.O5(CLBLM_L_X8Y137_SLICE_X10Y137_CO5),
.O6(CLBLM_L_X8Y137_SLICE_X10Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00330033ffcfffcf)
  ) CLBLM_L_X8Y137_SLICE_X10Y137_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y136_SLICE_X9Y136_CQ),
.I2(CLBLM_L_X10Y139_SLICE_X13Y139_AQ),
.I3(CLBLM_R_X5Y136_SLICE_X7Y136_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y137_SLICE_X10Y137_BO5),
.O6(CLBLM_L_X8Y137_SLICE_X10Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffccff00fcccf000)
  ) CLBLM_L_X8Y137_SLICE_X10Y137_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y135_SLICE_X15Y135_BQ),
.I2(CLBLM_L_X8Y137_SLICE_X10Y137_AQ),
.I3(CLBLM_R_X7Y144_SLICE_X9Y144_BO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X10Y137_SLICE_X13Y137_AQ),
.O5(CLBLM_L_X8Y137_SLICE_X10Y137_AO5),
.O6(CLBLM_L_X8Y137_SLICE_X10Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y137_SLICE_X11Y137_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y137_SLICE_X11Y137_AO6),
.Q(CLBLM_L_X8Y137_SLICE_X11Y137_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y137_SLICE_X11Y137_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y137_SLICE_X11Y137_BO6),
.Q(CLBLM_L_X8Y137_SLICE_X11Y137_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff6ccc00006ccc)
  ) CLBLM_L_X8Y137_SLICE_X11Y137_DLUT (
.I0(CLBLM_L_X10Y139_SLICE_X13Y139_AQ),
.I1(CLBLM_R_X5Y137_SLICE_X7Y137_BQ),
.I2(CLBLM_R_X11Y139_SLICE_X15Y139_CQ),
.I3(CLBLM_L_X8Y137_SLICE_X10Y137_BO6),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(CLBLM_R_X7Y139_SLICE_X8Y139_BQ),
.O5(CLBLM_L_X8Y137_SLICE_X11Y137_DO5),
.O6(CLBLM_L_X8Y137_SLICE_X11Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'heeeeccfc00003333)
  ) CLBLM_L_X8Y137_SLICE_X11Y137_CLUT (
.I0(CLBLM_R_X7Y136_SLICE_X9Y136_BO5),
.I1(CLBLL_L_X4Y134_SLICE_X4Y134_AQ),
.I2(CLBLM_R_X5Y141_SLICE_X7Y141_DO6),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_L_X10Y134_SLICE_X12Y134_CQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y137_SLICE_X11Y137_CO5),
.O6(CLBLM_L_X8Y137_SLICE_X11Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0eff0e000e000e)
  ) CLBLM_L_X8Y137_SLICE_X11Y137_BLUT (
.I0(CLBLM_L_X10Y137_SLICE_X12Y137_CQ),
.I1(CLBLM_L_X8Y137_SLICE_X11Y137_BQ),
.I2(CLBLM_R_X5Y132_SLICE_X7Y132_DO6),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLM_R_X7Y137_SLICE_X9Y137_AQ),
.O5(CLBLM_L_X8Y137_SLICE_X11Y137_BO5),
.O6(CLBLM_L_X8Y137_SLICE_X11Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbb888b8bbb888b8)
  ) CLBLM_L_X8Y137_SLICE_X11Y137_ALUT (
.I0(CLBLM_L_X10Y137_SLICE_X12Y137_B5Q),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X8Y137_SLICE_X11Y137_AQ),
.I3(CLBLM_L_X8Y143_SLICE_X10Y143_DO5),
.I4(CLBLM_R_X11Y137_SLICE_X14Y137_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y137_SLICE_X11Y137_AO5),
.O6(CLBLM_L_X8Y137_SLICE_X11Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y138_SLICE_X10Y138_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y138_SLICE_X10Y138_DO5),
.Q(CLBLM_L_X8Y138_SLICE_X10Y138_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y138_SLICE_X10Y138_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y138_SLICE_X10Y138_AO6),
.Q(CLBLM_L_X8Y138_SLICE_X10Y138_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y138_SLICE_X10Y138_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y138_SLICE_X10Y138_BO6),
.Q(CLBLM_L_X8Y138_SLICE_X10Y138_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y138_SLICE_X10Y138_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y138_SLICE_X10Y138_CO6),
.Q(CLBLM_L_X8Y138_SLICE_X10Y138_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y138_SLICE_X10Y138_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y138_SLICE_X10Y138_DO6),
.Q(CLBLM_L_X8Y138_SLICE_X10Y138_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc0fcc0faa00aaf0)
  ) CLBLM_L_X8Y138_SLICE_X10Y138_DLUT (
.I0(CLBLM_L_X10Y135_SLICE_X13Y135_B5Q),
.I1(CLBLM_L_X8Y138_SLICE_X10Y138_CQ),
.I2(RIOB33_X105Y119_IOB_X1Y119_I),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y138_SLICE_X10Y138_D5Q),
.I5(1'b1),
.O5(CLBLM_L_X8Y138_SLICE_X10Y138_DO5),
.O6(CLBLM_L_X8Y138_SLICE_X10Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000000a500a5)
  ) CLBLM_L_X8Y138_SLICE_X10Y138_CLUT (
.I0(CLBLM_L_X8Y136_SLICE_X11Y136_AQ),
.I1(1'b1),
.I2(CLBLM_L_X8Y136_SLICE_X11Y136_DO5),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_L_X8Y142_SLICE_X10Y142_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y138_SLICE_X10Y138_CO5),
.O6(CLBLM_L_X8Y138_SLICE_X10Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000ff006c6c)
  ) CLBLM_L_X8Y138_SLICE_X10Y138_BLUT (
.I0(CLBLM_R_X7Y138_SLICE_X9Y138_CO6),
.I1(CLBLM_L_X8Y138_SLICE_X10Y138_BQ),
.I2(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I3(CLBLM_R_X7Y139_SLICE_X8Y139_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X11Y135_SLICE_X14Y135_AQ),
.O5(CLBLM_L_X8Y138_SLICE_X10Y138_BO5),
.O6(CLBLM_L_X8Y138_SLICE_X10Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00aa03aa00)
  ) CLBLM_L_X8Y138_SLICE_X10Y138_ALUT (
.I0(CLBLL_L_X4Y138_SLICE_X4Y138_AQ),
.I1(CLBLM_L_X8Y138_SLICE_X10Y138_DQ),
.I2(CLBLM_L_X8Y138_SLICE_X10Y138_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y119_IOB_X1Y119_I),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_L_X8Y138_SLICE_X10Y138_AO5),
.O6(CLBLM_L_X8Y138_SLICE_X10Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y138_SLICE_X11Y138_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y138_SLICE_X11Y138_AO6),
.Q(CLBLM_L_X8Y138_SLICE_X11Y138_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y138_SLICE_X11Y138_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y138_SLICE_X11Y138_BO6),
.Q(CLBLM_L_X8Y138_SLICE_X11Y138_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3cc33cc3c33cc33c)
  ) CLBLM_L_X8Y138_SLICE_X11Y138_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y142_SLICE_X12Y142_DQ),
.I2(CLBLM_L_X12Y139_SLICE_X16Y139_A5Q),
.I3(CLBLM_R_X7Y135_SLICE_X8Y135_CQ),
.I4(1'b1),
.I5(CLBLM_L_X8Y138_SLICE_X11Y138_AQ),
.O5(CLBLM_L_X8Y138_SLICE_X11Y138_DO5),
.O6(CLBLM_L_X8Y138_SLICE_X11Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc8888333f333f)
  ) CLBLM_L_X8Y138_SLICE_X11Y138_CLUT (
.I0(CLBLM_L_X8Y139_SLICE_X11Y139_AQ),
.I1(RIOB33_X105Y121_IOB_X1Y121_I),
.I2(CLBLM_L_X10Y137_SLICE_X12Y137_AQ),
.I3(CLBLM_R_X5Y140_SLICE_X7Y140_BQ),
.I4(CLBLM_L_X10Y135_SLICE_X12Y135_BQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y138_SLICE_X11Y138_CO5),
.O6(CLBLM_L_X8Y138_SLICE_X11Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf044f044f044f044)
  ) CLBLM_L_X8Y138_SLICE_X11Y138_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X8Y138_SLICE_X11Y138_BQ),
.I2(CLBLM_L_X8Y138_SLICE_X11Y138_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y138_SLICE_X11Y138_BO5),
.O6(CLBLM_L_X8Y138_SLICE_X11Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf044f088f044f088)
  ) CLBLM_L_X8Y138_SLICE_X11Y138_ALUT (
.I0(CLBLM_L_X8Y138_SLICE_X11Y138_DO6),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_L_X8Y139_SLICE_X11Y139_BQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y136_SLICE_X13Y136_CO6),
.I5(1'b1),
.O5(CLBLM_L_X8Y138_SLICE_X11Y138_AO5),
.O6(CLBLM_L_X8Y138_SLICE_X11Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y139_SLICE_X10Y139_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y139_SLICE_X10Y139_AO6),
.Q(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y139_SLICE_X10Y139_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y139_SLICE_X10Y139_BO6),
.Q(CLBLM_L_X8Y139_SLICE_X10Y139_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y139_SLICE_X10Y139_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y139_SLICE_X10Y139_CO6),
.Q(CLBLM_L_X8Y139_SLICE_X10Y139_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y139_SLICE_X10Y139_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y139_SLICE_X10Y139_DO6),
.Q(CLBLM_L_X8Y139_SLICE_X10Y139_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0055555050)
  ) CLBLM_L_X8Y139_SLICE_X10Y139_DLUT (
.I0(CLBLL_L_X4Y133_SLICE_X5Y133_BO6),
.I1(1'b1),
.I2(CLBLM_L_X8Y139_SLICE_X10Y139_DQ),
.I3(CLBLM_L_X12Y140_SLICE_X17Y140_BQ),
.I4(CLBLM_R_X5Y137_SLICE_X7Y137_B5Q),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y139_SLICE_X10Y139_DO5),
.O6(CLBLM_L_X8Y139_SLICE_X10Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0afafafa0acacac)
  ) CLBLM_L_X8Y139_SLICE_X10Y139_CLUT (
.I0(CLBLM_L_X8Y138_SLICE_X11Y138_BQ),
.I1(CLBLM_L_X8Y139_SLICE_X10Y139_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X12Y134_SLICE_X17Y134_AO6),
.I4(CLBLM_L_X10Y139_SLICE_X13Y139_B5Q),
.I5(CLBLM_R_X5Y139_SLICE_X7Y139_AQ),
.O5(CLBLM_L_X8Y139_SLICE_X10Y139_CO5),
.O6(CLBLM_L_X8Y139_SLICE_X10Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0030300303)
  ) CLBLM_L_X8Y139_SLICE_X10Y139_BLUT (
.I0(1'b1),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_L_X8Y139_SLICE_X11Y139_CO6),
.I3(CLBLM_R_X11Y141_SLICE_X15Y141_BQ),
.I4(CLBLL_L_X4Y135_SLICE_X5Y135_BQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y139_SLICE_X10Y139_BO5),
.O6(CLBLM_L_X8Y139_SLICE_X10Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa0faa0faa00)
  ) CLBLM_L_X8Y139_SLICE_X10Y139_ALUT (
.I0(CLBLM_L_X8Y139_SLICE_X10Y139_CQ),
.I1(1'b1),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X11Y136_SLICE_X14Y136_CO5),
.I5(CLBLM_R_X11Y139_SLICE_X15Y139_DQ),
.O5(CLBLM_L_X8Y139_SLICE_X10Y139_AO5),
.O6(CLBLM_L_X8Y139_SLICE_X10Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y139_SLICE_X11Y139_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y139_SLICE_X11Y139_AO6),
.Q(CLBLM_L_X8Y139_SLICE_X11Y139_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y139_SLICE_X11Y139_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y139_SLICE_X11Y139_BO6),
.Q(CLBLM_L_X8Y139_SLICE_X11Y139_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfc0000f8fc1100)
  ) CLBLM_L_X8Y139_SLICE_X11Y139_DLUT (
.I0(CLBLM_L_X10Y139_SLICE_X13Y139_AQ),
.I1(CLBLM_L_X8Y141_SLICE_X10Y141_CQ),
.I2(CLBLM_R_X7Y139_SLICE_X8Y139_A5Q),
.I3(CLBLM_R_X11Y139_SLICE_X15Y139_CQ),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(CLBLM_L_X10Y138_SLICE_X12Y138_DO6),
.O5(CLBLM_L_X8Y139_SLICE_X11Y139_DO5),
.O6(CLBLM_L_X8Y139_SLICE_X11Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h03ff03ff0bdd03ff)
  ) CLBLM_L_X8Y139_SLICE_X11Y139_CLUT (
.I0(CLBLM_L_X10Y139_SLICE_X13Y139_AQ),
.I1(CLBLM_L_X8Y144_SLICE_X11Y144_AQ),
.I2(CLBLM_R_X5Y140_SLICE_X7Y140_BQ),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(CLBLM_R_X11Y139_SLICE_X15Y139_CQ),
.I5(CLBLM_L_X10Y138_SLICE_X12Y138_DO6),
.O5(CLBLM_L_X8Y139_SLICE_X11Y139_CO5),
.O6(CLBLM_L_X8Y139_SLICE_X11Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8888bb888888bb88)
  ) CLBLM_L_X8Y139_SLICE_X11Y139_BLUT (
.I0(CLBLM_R_X7Y144_SLICE_X8Y144_BQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(1'b1),
.I3(CLBLM_L_X10Y135_SLICE_X12Y135_BQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y139_SLICE_X11Y139_BO5),
.O6(CLBLM_L_X8Y139_SLICE_X11Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hb8b8b888bbbbbb88)
  ) CLBLM_L_X8Y139_SLICE_X11Y139_ALUT (
.I0(CLBLM_L_X10Y142_SLICE_X12Y142_DQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X8Y139_SLICE_X11Y139_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_L_X8Y138_SLICE_X10Y138_AQ),
.I5(CLBLM_L_X8Y139_SLICE_X11Y139_CO6),
.O5(CLBLM_L_X8Y139_SLICE_X11Y139_AO5),
.O6(CLBLM_L_X8Y139_SLICE_X11Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y140_SLICE_X10Y140_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y140_SLICE_X10Y140_AO5),
.Q(CLBLM_L_X8Y140_SLICE_X10Y140_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y140_SLICE_X10Y140_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y140_SLICE_X10Y140_AO6),
.Q(CLBLM_L_X8Y140_SLICE_X10Y140_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y140_SLICE_X10Y140_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y140_SLICE_X10Y140_BO6),
.Q(CLBLM_L_X8Y140_SLICE_X10Y140_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y140_SLICE_X10Y140_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y140_SLICE_X10Y140_CO6),
.Q(CLBLM_L_X8Y140_SLICE_X10Y140_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y140_SLICE_X10Y140_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y140_SLICE_X10Y140_DO6),
.Q(CLBLM_L_X8Y140_SLICE_X10Y140_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0012121212)
  ) CLBLM_L_X8Y140_SLICE_X10Y140_DLUT (
.I0(CLBLM_R_X7Y138_SLICE_X8Y138_BQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_L_X8Y136_SLICE_X11Y136_DO6),
.I3(CLBLM_R_X7Y143_SLICE_X9Y143_CQ),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y140_SLICE_X10Y140_DO5),
.O6(CLBLM_L_X8Y140_SLICE_X10Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5e4e4a0a0e4e4)
  ) CLBLM_L_X8Y140_SLICE_X10Y140_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y140_SLICE_X10Y140_CQ),
.I2(CLBLM_R_X11Y140_SLICE_X14Y140_CQ),
.I3(1'b1),
.I4(CLBLM_L_X8Y143_SLICE_X10Y143_DO5),
.I5(CLBLM_L_X10Y142_SLICE_X12Y142_DQ),
.O5(CLBLM_L_X8Y140_SLICE_X10Y140_CO5),
.O6(CLBLM_L_X8Y140_SLICE_X10Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00cacacaca)
  ) CLBLM_L_X8Y140_SLICE_X10Y140_BLUT (
.I0(CLBLM_R_X11Y141_SLICE_X15Y141_DQ),
.I1(CLBLM_L_X8Y140_SLICE_X10Y140_BQ),
.I2(CLBLM_L_X8Y143_SLICE_X10Y143_DO6),
.I3(CLBLM_L_X8Y142_SLICE_X10Y142_BQ),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y140_SLICE_X10Y140_BO5),
.O6(CLBLM_L_X8Y140_SLICE_X10Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccaaccaaf0fff000)
  ) CLBLM_L_X8Y140_SLICE_X10Y140_ALUT (
.I0(CLBLL_L_X4Y141_SLICE_X4Y141_DO6),
.I1(CLBLM_L_X8Y132_SLICE_X11Y132_BQ),
.I2(CLBLM_L_X10Y143_SLICE_X12Y143_BQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X3Y140_SLICE_X2Y140_DO6),
.I5(1'b1),
.O5(CLBLM_L_X8Y140_SLICE_X10Y140_AO5),
.O6(CLBLM_L_X8Y140_SLICE_X10Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y140_SLICE_X11Y140_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y140_SLICE_X11Y140_AO5),
.Q(CLBLM_L_X8Y140_SLICE_X11Y140_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y140_SLICE_X11Y140_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y140_SLICE_X11Y140_AO6),
.Q(CLBLM_L_X8Y140_SLICE_X11Y140_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y140_SLICE_X11Y140_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y140_SLICE_X11Y140_BO6),
.Q(CLBLM_L_X8Y140_SLICE_X11Y140_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffdffffffffffff)
  ) CLBLM_L_X8Y140_SLICE_X11Y140_DLUT (
.I0(CLBLM_L_X8Y140_SLICE_X11Y140_CO5),
.I1(CLBLM_L_X8Y136_SLICE_X11Y136_CQ),
.I2(CLBLM_R_X7Y144_SLICE_X8Y144_CQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_L_X8Y141_SLICE_X10Y141_DQ),
.I5(CLBLM_L_X10Y142_SLICE_X12Y142_DQ),
.O5(CLBLM_L_X8Y140_SLICE_X11Y140_DO5),
.O6(CLBLM_L_X8Y140_SLICE_X11Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffefef30303030)
  ) CLBLM_L_X8Y140_SLICE_X11Y140_CLUT (
.I0(CLBLM_L_X10Y137_SLICE_X13Y137_BQ),
.I1(RIOB33_X105Y121_IOB_X1Y121_I),
.I2(CLBLM_R_X11Y136_SLICE_X14Y136_DQ),
.I3(1'b1),
.I4(CLBLM_R_X7Y144_SLICE_X8Y144_CQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y140_SLICE_X11Y140_CO5),
.O6(CLBLM_L_X8Y140_SLICE_X11Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff5fff4c005f004c)
  ) CLBLM_L_X8Y140_SLICE_X11Y140_BLUT (
.I0(CLBLM_L_X12Y134_SLICE_X17Y134_AO6),
.I1(CLBLM_L_X8Y140_SLICE_X11Y140_BQ),
.I2(CLBLM_L_X10Y139_SLICE_X13Y139_B5Q),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X11Y136_SLICE_X14Y136_AQ),
.I5(CLBLM_L_X8Y141_SLICE_X10Y141_CQ),
.O5(CLBLM_L_X8Y140_SLICE_X11Y140_BO5),
.O6(CLBLM_L_X8Y140_SLICE_X11Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hd1c0d1c0ff33cc00)
  ) CLBLM_L_X8Y140_SLICE_X11Y140_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X7Y138_SLICE_X8Y138_BQ),
.I3(CLBLM_L_X12Y140_SLICE_X16Y140_DQ),
.I4(CLBLM_R_X7Y134_SLICE_X8Y134_BQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y140_SLICE_X11Y140_AO5),
.O6(CLBLM_L_X8Y140_SLICE_X11Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y141_SLICE_X10Y141_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y141_SLICE_X10Y141_AO6),
.Q(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y141_SLICE_X10Y141_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y141_SLICE_X10Y141_BO6),
.Q(CLBLM_L_X8Y141_SLICE_X10Y141_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y141_SLICE_X10Y141_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y141_SLICE_X10Y141_CO6),
.Q(CLBLM_L_X8Y141_SLICE_X10Y141_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y141_SLICE_X10Y141_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y141_SLICE_X10Y141_DO6),
.Q(CLBLM_L_X8Y141_SLICE_X10Y141_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa00cc00cc)
  ) CLBLM_L_X8Y141_SLICE_X10Y141_DLUT (
.I0(CLBLM_R_X11Y141_SLICE_X15Y141_DQ),
.I1(CLBLM_L_X10Y142_SLICE_X12Y142_DQ),
.I2(1'b1),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y141_SLICE_X10Y141_DO5),
.O6(CLBLM_L_X8Y141_SLICE_X10Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000000cc00cc)
  ) CLBLM_L_X8Y141_SLICE_X10Y141_CLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y141_SLICE_X10Y141_CQ),
.I2(1'b1),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_L_X8Y142_SLICE_X10Y142_CQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y141_SLICE_X10Y141_CO5),
.O6(CLBLM_L_X8Y141_SLICE_X10Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000a8a8a8a8)
  ) CLBLM_L_X8Y141_SLICE_X10Y141_BLUT (
.I0(CLBLM_L_X8Y143_SLICE_X10Y143_DO6),
.I1(CLBLM_L_X8Y141_SLICE_X10Y141_BQ),
.I2(CLBLM_L_X10Y140_SLICE_X13Y140_BQ),
.I3(1'b1),
.I4(CLBLM_R_X5Y140_SLICE_X7Y140_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y141_SLICE_X10Y141_BO5),
.O6(CLBLM_L_X8Y141_SLICE_X10Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffccf0cca0)
  ) CLBLM_L_X8Y141_SLICE_X10Y141_ALUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_L_X8Y141_SLICE_X10Y141_BQ),
.I2(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y138_SLICE_X10Y138_AQ),
.I5(CLBLM_L_X8Y134_SLICE_X10Y134_CO6),
.O5(CLBLM_L_X8Y141_SLICE_X10Y141_AO5),
.O6(CLBLM_L_X8Y141_SLICE_X10Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y141_SLICE_X11Y141_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y141_SLICE_X11Y141_AO6),
.Q(CLBLM_L_X8Y141_SLICE_X11Y141_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y141_SLICE_X11Y141_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y141_SLICE_X11Y141_BO6),
.Q(CLBLM_L_X8Y141_SLICE_X11Y141_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y141_SLICE_X11Y141_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y141_SLICE_X11Y141_CO6),
.Q(CLBLM_L_X8Y141_SLICE_X11Y141_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccf0ccf000005f5f)
  ) CLBLM_L_X8Y141_SLICE_X11Y141_DLUT (
.I0(CLBLM_R_X5Y139_SLICE_X7Y139_AQ),
.I1(CLBLM_R_X11Y139_SLICE_X14Y139_AQ),
.I2(CLBLL_L_X4Y142_SLICE_X5Y142_DO6),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X11Y138_SLICE_X14Y138_DQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y141_SLICE_X11Y141_DO5),
.O6(CLBLM_L_X8Y141_SLICE_X11Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000d0c0d0c0)
  ) CLBLM_L_X8Y141_SLICE_X11Y141_CLUT (
.I0(RIOB33_X105Y121_IOB_X1Y121_I),
.I1(CLBLM_L_X8Y141_SLICE_X11Y141_CQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X11Y136_SLICE_X14Y136_DQ),
.I4(CLBLM_L_X8Y142_SLICE_X11Y142_DQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y141_SLICE_X11Y141_CO5),
.O6(CLBLM_L_X8Y141_SLICE_X11Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'he4f5e4a0f5f5a0a0)
  ) CLBLM_L_X8Y141_SLICE_X11Y141_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y141_SLICE_X11Y141_BQ),
.I2(CLBLM_R_X13Y141_SLICE_X19Y141_BQ),
.I3(CLBLM_L_X12Y135_SLICE_X17Y135_AQ),
.I4(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I5(CLBLL_L_X4Y137_SLICE_X4Y137_CQ),
.O5(CLBLM_L_X8Y141_SLICE_X11Y141_BO5),
.O6(CLBLM_L_X8Y141_SLICE_X11Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88dddd88ddd8ddd8)
  ) CLBLM_L_X8Y141_SLICE_X11Y141_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y141_SLICE_X11Y141_BQ),
.I2(CLBLM_L_X8Y141_SLICE_X11Y141_AQ),
.I3(CLBLM_L_X10Y141_SLICE_X13Y141_DO6),
.I4(CLBLM_R_X7Y138_SLICE_X8Y138_BQ),
.I5(CLBLM_L_X8Y143_SLICE_X10Y143_DO5),
.O5(CLBLM_L_X8Y141_SLICE_X11Y141_AO5),
.O6(CLBLM_L_X8Y141_SLICE_X11Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y142_SLICE_X10Y142_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y142_SLICE_X10Y142_DO5),
.Q(CLBLM_L_X8Y142_SLICE_X10Y142_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y142_SLICE_X10Y142_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y142_SLICE_X10Y142_AO6),
.Q(CLBLM_L_X8Y142_SLICE_X10Y142_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y142_SLICE_X10Y142_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y142_SLICE_X10Y142_BO6),
.Q(CLBLM_L_X8Y142_SLICE_X10Y142_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y142_SLICE_X10Y142_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y142_SLICE_X10Y142_CO6),
.Q(CLBLM_L_X8Y142_SLICE_X10Y142_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y142_SLICE_X10Y142_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y142_SLICE_X10Y142_DO6),
.Q(CLBLM_L_X8Y142_SLICE_X10Y142_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3c0f3c0eeeeaaaa)
  ) CLBLM_L_X8Y142_SLICE_X10Y142_DLUT (
.I0(CLBLM_L_X8Y143_SLICE_X11Y143_AO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X7Y140_SLICE_X9Y140_BQ),
.I3(CLBLM_R_X7Y140_SLICE_X8Y140_DO6),
.I4(CLBLM_R_X5Y141_SLICE_X7Y141_BQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y142_SLICE_X10Y142_DO5),
.O6(CLBLM_L_X8Y142_SLICE_X10Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfecefece32023202)
  ) CLBLM_L_X8Y142_SLICE_X10Y142_CLUT (
.I0(CLBLM_L_X8Y142_SLICE_X10Y142_CQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X8Y143_SLICE_X10Y143_DO5),
.I3(CLBLM_L_X8Y139_SLICE_X10Y139_BQ),
.I4(1'b1),
.I5(CLBLM_L_X8Y142_SLICE_X10Y142_D5Q),
.O5(CLBLM_L_X8Y142_SLICE_X10Y142_CO5),
.O6(CLBLM_L_X8Y142_SLICE_X10Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc5500cccc5505)
  ) CLBLM_L_X8Y142_SLICE_X10Y142_BLUT (
.I0(CLBLM_R_X11Y144_SLICE_X14Y144_AQ),
.I1(CLBLL_L_X4Y135_SLICE_X4Y135_A5Q),
.I2(CLBLM_L_X10Y142_SLICE_X12Y142_CQ),
.I3(CLBLM_L_X8Y142_SLICE_X10Y142_D5Q),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.O5(CLBLM_L_X8Y142_SLICE_X10Y142_BO5),
.O6(CLBLM_L_X8Y142_SLICE_X10Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8888ddd8ddd8ddd8)
  ) CLBLM_L_X8Y142_SLICE_X10Y142_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X11Y142_SLICE_X14Y142_AQ),
.I2(CLBLM_L_X8Y142_SLICE_X10Y142_AQ),
.I3(CLBLM_R_X7Y140_SLICE_X9Y140_BQ),
.I4(CLBLM_L_X12Y135_SLICE_X17Y135_AQ),
.I5(CLBLL_L_X4Y137_SLICE_X4Y137_CQ),
.O5(CLBLM_L_X8Y142_SLICE_X10Y142_AO5),
.O6(CLBLM_L_X8Y142_SLICE_X10Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y142_SLICE_X11Y142_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y142_SLICE_X11Y142_AO6),
.Q(CLBLM_L_X8Y142_SLICE_X11Y142_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y142_SLICE_X11Y142_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y142_SLICE_X11Y142_BO6),
.Q(CLBLM_L_X8Y142_SLICE_X11Y142_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y142_SLICE_X11Y142_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y142_SLICE_X11Y142_CO6),
.Q(CLBLM_L_X8Y142_SLICE_X11Y142_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y142_SLICE_X11Y142_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y142_SLICE_X11Y142_DO6),
.Q(CLBLM_L_X8Y142_SLICE_X11Y142_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaffffaaaa0300)
  ) CLBLM_L_X8Y142_SLICE_X11Y142_DLUT (
.I0(CLBLM_L_X10Y134_SLICE_X12Y134_AQ),
.I1(CLBLM_R_X7Y141_SLICE_X8Y141_CO6),
.I2(CLBLM_R_X7Y139_SLICE_X9Y139_CO6),
.I3(CLBLM_L_X10Y145_SLICE_X13Y145_BO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y143_SLICE_X11Y143_BO6),
.O5(CLBLM_L_X8Y142_SLICE_X11Y142_DO5),
.O6(CLBLM_L_X8Y142_SLICE_X11Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0f000fff000000)
  ) CLBLM_L_X8Y142_SLICE_X11Y142_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_L_X10Y144_SLICE_X12Y144_AO5),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X12Y140_SLICE_X17Y140_CQ),
.I5(CLBLM_R_X7Y142_SLICE_X9Y142_AQ),
.O5(CLBLM_L_X8Y142_SLICE_X11Y142_CO5),
.O6(CLBLM_L_X8Y142_SLICE_X11Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbfb0b0bfefe0e0e)
  ) CLBLM_L_X8Y142_SLICE_X11Y142_BLUT (
.I0(CLBLM_L_X10Y145_SLICE_X13Y145_BO6),
.I1(CLBLM_L_X8Y142_SLICE_X11Y142_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(CLBLM_R_X7Y133_SLICE_X8Y133_BQ),
.I5(CLBLM_L_X8Y143_SLICE_X11Y143_CO6),
.O5(CLBLM_L_X8Y142_SLICE_X11Y142_BO5),
.O6(CLBLM_L_X8Y142_SLICE_X11Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8888ddd8ddd8ddd8)
  ) CLBLM_L_X8Y142_SLICE_X11Y142_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X11Y141_SLICE_X15Y141_CQ),
.I2(CLBLM_L_X8Y142_SLICE_X11Y142_AQ),
.I3(CLBLM_R_X5Y139_SLICE_X7Y139_AQ),
.I4(CLBLM_L_X12Y135_SLICE_X17Y135_AQ),
.I5(CLBLL_L_X4Y137_SLICE_X4Y137_CQ),
.O5(CLBLM_L_X8Y142_SLICE_X11Y142_AO5),
.O6(CLBLM_L_X8Y142_SLICE_X11Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y143_SLICE_X10Y143_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y143_SLICE_X10Y143_AO6),
.Q(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y143_SLICE_X10Y143_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y143_SLICE_X10Y143_BO6),
.Q(CLBLM_L_X8Y143_SLICE_X10Y143_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y143_SLICE_X10Y143_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y143_SLICE_X10Y143_CO6),
.Q(CLBLM_L_X8Y143_SLICE_X10Y143_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaa2a2aaaaaa22)
  ) CLBLM_L_X8Y143_SLICE_X10Y143_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X11Y136_SLICE_X14Y136_DQ),
.I2(CLBLM_R_X11Y141_SLICE_X15Y141_AQ),
.I3(CLBLM_R_X7Y144_SLICE_X8Y144_CQ),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y143_SLICE_X10Y143_DO5),
.O6(CLBLM_L_X8Y143_SLICE_X10Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff550055ff440044)
  ) CLBLM_L_X8Y143_SLICE_X10Y143_CLUT (
.I0(CLBLL_L_X4Y133_SLICE_X5Y133_BO6),
.I1(CLBLM_L_X8Y143_SLICE_X10Y143_CQ),
.I2(1'b1),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X11Y143_SLICE_X14Y143_AQ),
.I5(CLBLL_L_X4Y137_SLICE_X4Y137_A5Q),
.O5(CLBLM_L_X8Y143_SLICE_X10Y143_CO5),
.O6(CLBLM_L_X8Y143_SLICE_X10Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hacafacafaca0aca0)
  ) CLBLM_L_X8Y143_SLICE_X10Y143_BLUT (
.I0(CLBLM_L_X8Y140_SLICE_X10Y140_DQ),
.I1(CLBLM_L_X8Y143_SLICE_X10Y143_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y143_SLICE_X10Y143_DO5),
.I4(1'b1),
.I5(CLBLM_L_X8Y141_SLICE_X10Y141_DQ),
.O5(CLBLM_L_X8Y143_SLICE_X10Y143_BO5),
.O6(CLBLM_L_X8Y143_SLICE_X10Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbaa1100baba1010)
  ) CLBLM_L_X8Y143_SLICE_X10Y143_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y121_IOB_X1Y121_I),
.I2(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.I3(CLBLM_L_X10Y142_SLICE_X12Y142_CQ),
.I4(CLBLM_R_X3Y137_SLICE_X2Y137_AQ),
.I5(CLBLM_R_X11Y143_SLICE_X14Y143_DO6),
.O5(CLBLM_L_X8Y143_SLICE_X10Y143_AO5),
.O6(CLBLM_L_X8Y143_SLICE_X10Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y143_SLICE_X11Y143_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y143_SLICE_X11Y143_DO5),
.O6(CLBLM_L_X8Y143_SLICE_X11Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0300030003000300)
  ) CLBLM_L_X8Y143_SLICE_X11Y143_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y144_SLICE_X8Y144_BQ),
.I2(CLBLM_R_X7Y144_SLICE_X8Y144_AQ),
.I3(CLBLM_R_X7Y143_SLICE_X9Y143_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y143_SLICE_X11Y143_CO5),
.O6(CLBLM_L_X8Y143_SLICE_X11Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6666646466666460)
  ) CLBLM_L_X8Y143_SLICE_X11Y143_BLUT (
.I0(CLBLM_L_X8Y144_SLICE_X11Y144_BO5),
.I1(CLBLM_L_X8Y142_SLICE_X11Y142_DQ),
.I2(CLBLM_L_X10Y142_SLICE_X12Y142_CQ),
.I3(CLBLM_L_X8Y142_SLICE_X10Y142_D5Q),
.I4(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.I5(CLBLM_R_X11Y144_SLICE_X14Y144_AQ),
.O5(CLBLM_L_X8Y143_SLICE_X11Y143_BO5),
.O6(CLBLM_L_X8Y143_SLICE_X11Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h55aadf0000000000)
  ) CLBLM_L_X8Y143_SLICE_X11Y143_ALUT (
.I0(CLBLM_L_X8Y144_SLICE_X11Y144_BO5),
.I1(CLBLM_R_X11Y143_SLICE_X14Y143_DO6),
.I2(CLBLM_R_X11Y144_SLICE_X14Y144_AQ),
.I3(CLBLM_L_X8Y142_SLICE_X10Y142_D5Q),
.I4(CLBLM_L_X10Y141_SLICE_X12Y141_C5Q),
.I5(CLBLM_R_X7Y143_SLICE_X8Y143_BO5),
.O5(CLBLM_L_X8Y143_SLICE_X11Y143_AO5),
.O6(CLBLM_L_X8Y143_SLICE_X11Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y144_SLICE_X10Y144_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y144_SLICE_X10Y144_DO5),
.O6(CLBLM_L_X8Y144_SLICE_X10Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y144_SLICE_X10Y144_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y144_SLICE_X10Y144_CO5),
.O6(CLBLM_L_X8Y144_SLICE_X10Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y144_SLICE_X10Y144_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y144_SLICE_X10Y144_BO5),
.O6(CLBLM_L_X8Y144_SLICE_X10Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y144_SLICE_X10Y144_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y144_SLICE_X10Y144_AO5),
.O6(CLBLM_L_X8Y144_SLICE_X10Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y144_SLICE_X11Y144_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y144_SLICE_X11Y144_AO6),
.Q(CLBLM_L_X8Y144_SLICE_X11Y144_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y144_SLICE_X11Y144_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y144_SLICE_X11Y144_DO5),
.O6(CLBLM_L_X8Y144_SLICE_X11Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000020)
  ) CLBLM_L_X8Y144_SLICE_X11Y144_CLUT (
.I0(CLBLM_R_X7Y143_SLICE_X9Y143_BQ),
.I1(CLBLM_R_X7Y144_SLICE_X8Y144_AQ),
.I2(CLBLM_L_X10Y141_SLICE_X12Y141_C5Q),
.I3(CLBLM_R_X7Y144_SLICE_X8Y144_BQ),
.I4(CLBLM_L_X8Y142_SLICE_X10Y142_D5Q),
.I5(CLBLM_L_X8Y142_SLICE_X11Y142_BQ),
.O5(CLBLM_L_X8Y144_SLICE_X11Y144_CO5),
.O6(CLBLM_L_X8Y144_SLICE_X11Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333332300000050)
  ) CLBLM_L_X8Y144_SLICE_X11Y144_BLUT (
.I0(CLBLM_R_X7Y144_SLICE_X8Y144_BQ),
.I1(CLBLM_L_X10Y145_SLICE_X13Y145_BO6),
.I2(CLBLM_R_X7Y143_SLICE_X9Y143_BQ),
.I3(CLBLM_R_X7Y144_SLICE_X8Y144_AQ),
.I4(CLBLM_L_X8Y142_SLICE_X11Y142_BQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y144_SLICE_X11Y144_BO5),
.O6(CLBLM_L_X8Y144_SLICE_X11Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0a000aff0a000a)
  ) CLBLM_L_X8Y144_SLICE_X11Y144_ALUT (
.I0(CLBLM_L_X8Y144_SLICE_X11Y144_AQ),
.I1(1'b1),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y143_SLICE_X9Y143_BQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y144_SLICE_X11Y144_AO5),
.O6(CLBLM_L_X8Y144_SLICE_X11Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y130_SLICE_X12Y130_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y130_SLICE_X12Y130_AO6),
.Q(CLBLM_L_X10Y130_SLICE_X12Y130_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y130_SLICE_X12Y130_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y130_SLICE_X12Y130_DO5),
.O6(CLBLM_L_X10Y130_SLICE_X12Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y130_SLICE_X12Y130_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y130_SLICE_X12Y130_CO5),
.O6(CLBLM_L_X10Y130_SLICE_X12Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00002000ffff8000)
  ) CLBLM_L_X10Y130_SLICE_X12Y130_BLUT (
.I0(CLBLL_L_X4Y135_SLICE_X5Y135_CQ),
.I1(CLBLM_L_X10Y131_SLICE_X12Y131_BQ),
.I2(CLBLM_L_X10Y130_SLICE_X12Y130_AQ),
.I3(CLBLM_R_X11Y131_SLICE_X15Y131_BQ),
.I4(CLBLM_R_X5Y132_SLICE_X7Y132_DO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y130_SLICE_X12Y130_BO5),
.O6(CLBLM_L_X10Y130_SLICE_X12Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00cca5cc00)
  ) CLBLM_L_X10Y130_SLICE_X12Y130_ALUT (
.I0(CLBLM_L_X10Y130_SLICE_X12Y130_BO5),
.I1(CLBLM_L_X12Y132_SLICE_X17Y132_AQ),
.I2(CLBLM_L_X10Y130_SLICE_X12Y130_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X11Y140_SLICE_X15Y140_CQ),
.O5(CLBLM_L_X10Y130_SLICE_X12Y130_AO5),
.O6(CLBLM_L_X10Y130_SLICE_X12Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y130_SLICE_X13Y130_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y130_SLICE_X13Y130_DO5),
.O6(CLBLM_L_X10Y130_SLICE_X13Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y130_SLICE_X13Y130_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y130_SLICE_X13Y130_CO5),
.O6(CLBLM_L_X10Y130_SLICE_X13Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y130_SLICE_X13Y130_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y130_SLICE_X13Y130_BO5),
.O6(CLBLM_L_X10Y130_SLICE_X13Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0b43333ffff)
  ) CLBLM_L_X10Y130_SLICE_X13Y130_ALUT (
.I0(CLBLL_L_X4Y135_SLICE_X5Y135_CQ),
.I1(CLBLM_R_X11Y131_SLICE_X15Y131_BQ),
.I2(CLBLM_L_X8Y131_SLICE_X11Y131_BQ),
.I3(CLBLM_L_X10Y131_SLICE_X12Y131_BQ),
.I4(CLBLM_L_X10Y130_SLICE_X12Y130_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y130_SLICE_X13Y130_AO5),
.O6(CLBLM_L_X10Y130_SLICE_X13Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y131_SLICE_X12Y131_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y131_SLICE_X12Y131_BO6),
.Q(CLBLM_L_X10Y131_SLICE_X12Y131_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000035353a35)
  ) CLBLM_L_X10Y131_SLICE_X12Y131_DLUT (
.I0(CLBLM_L_X10Y133_SLICE_X13Y133_AQ),
.I1(CLBLM_L_X8Y135_SLICE_X11Y135_AQ),
.I2(CLBLM_R_X5Y132_SLICE_X7Y132_DO6),
.I3(CLBLM_L_X10Y131_SLICE_X12Y131_CO6),
.I4(CLBLM_L_X10Y131_SLICE_X12Y131_AO5),
.I5(CLBLM_L_X8Y133_SLICE_X11Y133_CQ),
.O5(CLBLM_L_X10Y131_SLICE_X12Y131_DO5),
.O6(CLBLM_L_X10Y131_SLICE_X12Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h30303030fd02ff00)
  ) CLBLM_L_X10Y131_SLICE_X12Y131_CLUT (
.I0(CLBLM_L_X10Y130_SLICE_X12Y130_AQ),
.I1(CLBLL_L_X4Y135_SLICE_X5Y135_CQ),
.I2(CLBLM_L_X10Y131_SLICE_X12Y131_BQ),
.I3(CLBLM_L_X8Y131_SLICE_X10Y131_A5Q),
.I4(CLBLM_R_X11Y131_SLICE_X15Y131_BQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y131_SLICE_X12Y131_CO5),
.O6(CLBLM_L_X10Y131_SLICE_X12Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0faf0f8000a0008)
  ) CLBLM_L_X10Y131_SLICE_X12Y131_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X10Y131_SLICE_X12Y131_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X11Y140_SLICE_X15Y140_CQ),
.I4(CLBLM_L_X10Y130_SLICE_X12Y130_BO6),
.I5(CLBLM_L_X8Y131_SLICE_X10Y131_A5Q),
.O5(CLBLM_L_X10Y131_SLICE_X12Y131_BO5),
.O6(CLBLM_L_X10Y131_SLICE_X12Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0b4f0f0aaaaffff)
  ) CLBLM_L_X10Y131_SLICE_X12Y131_ALUT (
.I0(CLBLM_R_X11Y131_SLICE_X15Y131_BQ),
.I1(CLBLM_L_X10Y131_SLICE_X12Y131_BQ),
.I2(CLBLM_L_X10Y133_SLICE_X13Y133_AQ),
.I3(CLBLL_L_X4Y135_SLICE_X5Y135_CQ),
.I4(CLBLM_L_X10Y130_SLICE_X12Y130_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y131_SLICE_X12Y131_AO5),
.O6(CLBLM_L_X10Y131_SLICE_X12Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y131_SLICE_X13Y131_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y131_SLICE_X13Y131_AO6),
.Q(CLBLM_L_X10Y131_SLICE_X13Y131_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y131_SLICE_X13Y131_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y131_SLICE_X13Y131_BO6),
.Q(CLBLM_L_X10Y131_SLICE_X13Y131_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y131_SLICE_X13Y131_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y131_SLICE_X13Y131_CO6),
.Q(CLBLM_L_X10Y131_SLICE_X13Y131_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfe0202fefd0101fd)
  ) CLBLM_L_X10Y131_SLICE_X13Y131_DLUT (
.I0(CLBLM_R_X11Y131_SLICE_X14Y131_AO6),
.I1(CLBLM_R_X3Y139_SLICE_X3Y139_BO6),
.I2(CLBLM_R_X5Y133_SLICE_X7Y133_CO6),
.I3(CLBLM_L_X8Y135_SLICE_X11Y135_AQ),
.I4(CLBLM_L_X12Y136_SLICE_X16Y136_B5Q),
.I5(CLBLM_L_X10Y131_SLICE_X12Y131_AO6),
.O5(CLBLM_L_X10Y131_SLICE_X13Y131_DO5),
.O6(CLBLM_L_X10Y131_SLICE_X13Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f000ff00aa)
  ) CLBLM_L_X10Y131_SLICE_X13Y131_CLUT (
.I0(CLBLM_L_X10Y133_SLICE_X13Y133_AQ),
.I1(1'b1),
.I2(CLBLM_L_X8Y131_SLICE_X11Y131_AQ),
.I3(CLBLM_R_X5Y132_SLICE_X7Y132_DO6),
.I4(CLBLM_L_X10Y131_SLICE_X13Y131_CQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y131_SLICE_X13Y131_CO5),
.O6(CLBLM_L_X10Y131_SLICE_X13Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f0eef000f0ee)
  ) CLBLM_L_X10Y131_SLICE_X13Y131_BLUT (
.I0(CLBLM_L_X10Y131_SLICE_X13Y131_CQ),
.I1(CLBLM_L_X10Y131_SLICE_X13Y131_BQ),
.I2(CLBLM_L_X10Y131_SLICE_X13Y131_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X5Y132_SLICE_X7Y132_DO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y131_SLICE_X13Y131_BO5),
.O6(CLBLM_L_X10Y131_SLICE_X13Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd11dd11dc10dc10)
  ) CLBLM_L_X10Y131_SLICE_X13Y131_ALUT (
.I0(CLBLM_R_X5Y133_SLICE_X7Y133_DO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y131_SLICE_X13Y131_AQ),
.I3(CLBLM_R_X11Y132_SLICE_X14Y132_AQ),
.I4(1'b1),
.I5(CLBLM_R_X11Y133_SLICE_X15Y133_CQ),
.O5(CLBLM_L_X10Y131_SLICE_X13Y131_AO5),
.O6(CLBLM_L_X10Y131_SLICE_X13Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h77bb77bbddeeddee)
  ) CLBLM_L_X10Y132_SLICE_X12Y132_DLUT (
.I0(CLBLM_L_X10Y133_SLICE_X12Y133_AQ),
.I1(CLBLM_L_X10Y134_SLICE_X12Y134_AQ),
.I2(1'b1),
.I3(CLBLM_R_X7Y134_SLICE_X8Y134_C5Q),
.I4(1'b1),
.I5(CLBLM_R_X13Y137_SLICE_X18Y137_A5Q),
.O5(CLBLM_L_X10Y132_SLICE_X12Y132_DO5),
.O6(CLBLM_L_X10Y132_SLICE_X12Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h11dd10df11dd10df)
  ) CLBLM_L_X10Y132_SLICE_X12Y132_CLUT (
.I0(CLBLM_L_X10Y131_SLICE_X12Y131_CO5),
.I1(CLBLM_R_X5Y133_SLICE_X7Y133_CO6),
.I2(CLBLM_R_X5Y136_SLICE_X7Y136_DO6),
.I3(CLBLM_R_X11Y146_SLICE_X14Y146_AQ),
.I4(CLBLM_R_X7Y133_SLICE_X9Y133_DO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y132_SLICE_X12Y132_CO5),
.O6(CLBLM_L_X10Y132_SLICE_X12Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5a5f5a5fcccccccc)
  ) CLBLM_L_X10Y132_SLICE_X12Y132_BLUT (
.I0(CLBLM_L_X10Y133_SLICE_X12Y133_CQ),
.I1(CLBLM_L_X12Y136_SLICE_X16Y136_CQ),
.I2(CLBLM_L_X10Y133_SLICE_X12Y133_BQ),
.I3(CLBLM_L_X8Y132_SLICE_X11Y132_DO6),
.I4(1'b1),
.I5(CLBLM_R_X5Y132_SLICE_X7Y132_BO5),
.O5(CLBLM_L_X10Y132_SLICE_X12Y132_BO5),
.O6(CLBLM_L_X10Y132_SLICE_X12Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0802000004010000)
  ) CLBLM_L_X10Y132_SLICE_X12Y132_ALUT (
.I0(CLBLM_L_X8Y134_SLICE_X11Y134_BQ),
.I1(CLBLM_L_X12Y136_SLICE_X16Y136_CQ),
.I2(CLBLM_L_X10Y132_SLICE_X13Y132_DO6),
.I3(CLBLM_L_X10Y132_SLICE_X12Y132_BO6),
.I4(CLBLM_L_X8Y131_SLICE_X11Y131_DO6),
.I5(CLBLM_L_X12Y136_SLICE_X16Y136_B5Q),
.O5(CLBLM_L_X10Y132_SLICE_X12Y132_AO5),
.O6(CLBLM_L_X10Y132_SLICE_X12Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf7fdfbfef7fdfbfe)
  ) CLBLM_L_X10Y132_SLICE_X13Y132_DLUT (
.I0(CLBLM_R_X11Y134_SLICE_X15Y134_CQ),
.I1(CLBLM_L_X10Y141_SLICE_X12Y141_CQ),
.I2(CLBLM_L_X10Y132_SLICE_X12Y132_DO6),
.I3(CLBLM_R_X11Y133_SLICE_X15Y133_CQ),
.I4(CLBLM_L_X10Y134_SLICE_X13Y134_B5Q),
.I5(1'b1),
.O5(CLBLM_L_X10Y132_SLICE_X13Y132_DO5),
.O6(CLBLM_L_X10Y132_SLICE_X13Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h4e4e4e0f1b1b1b0f)
  ) CLBLM_L_X10Y132_SLICE_X13Y132_CLUT (
.I0(CLBLM_R_X5Y133_SLICE_X7Y133_CO6),
.I1(CLBLM_L_X10Y137_SLICE_X12Y137_CQ),
.I2(CLBLM_L_X10Y134_SLICE_X13Y134_B5Q),
.I3(CLBLM_R_X5Y136_SLICE_X7Y136_DO6),
.I4(CLBLM_R_X7Y133_SLICE_X9Y133_DO6),
.I5(CLBLM_R_X11Y132_SLICE_X15Y132_AO6),
.O5(CLBLM_L_X10Y132_SLICE_X13Y132_CO5),
.O6(CLBLM_L_X10Y132_SLICE_X13Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaac3555555c3)
  ) CLBLM_L_X10Y132_SLICE_X13Y132_BLUT (
.I0(CLBLM_L_X10Y137_SLICE_X12Y137_B5Q),
.I1(CLBLM_L_X10Y133_SLICE_X12Y133_DO5),
.I2(CLBLM_L_X10Y130_SLICE_X13Y130_AO6),
.I3(CLBLM_R_X3Y139_SLICE_X3Y139_BO6),
.I4(CLBLM_R_X5Y133_SLICE_X7Y133_CO6),
.I5(CLBLM_L_X10Y141_SLICE_X12Y141_CQ),
.O5(CLBLM_L_X10Y132_SLICE_X13Y132_BO5),
.O6(CLBLM_L_X10Y132_SLICE_X13Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_L_X10Y132_SLICE_X13Y132_ALUT (
.I0(CLBLM_L_X10Y131_SLICE_X13Y131_DO6),
.I1(CLBLM_R_X11Y131_SLICE_X14Y131_CO6),
.I2(CLBLM_L_X10Y132_SLICE_X12Y132_CO6),
.I3(CLBLM_L_X10Y132_SLICE_X13Y132_BO6),
.I4(CLBLM_L_X8Y132_SLICE_X10Y132_CO6),
.I5(CLBLM_L_X10Y132_SLICE_X13Y132_CO6),
.O5(CLBLM_L_X10Y132_SLICE_X13Y132_AO5),
.O6(CLBLM_L_X10Y132_SLICE_X13Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y133_SLICE_X12Y133_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y133_SLICE_X12Y133_AO6),
.Q(CLBLM_L_X10Y133_SLICE_X12Y133_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y133_SLICE_X12Y133_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y133_SLICE_X12Y133_BO6),
.Q(CLBLM_L_X10Y133_SLICE_X12Y133_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y133_SLICE_X12Y133_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y133_SLICE_X12Y133_CO6),
.Q(CLBLM_L_X10Y133_SLICE_X12Y133_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffff0ffccccc9cc)
  ) CLBLM_L_X10Y133_SLICE_X12Y133_DLUT (
.I0(CLBLM_R_X11Y131_SLICE_X15Y131_BQ),
.I1(CLBLM_L_X8Y137_SLICE_X11Y137_BQ),
.I2(CLBLL_L_X4Y135_SLICE_X5Y135_CQ),
.I3(CLBLM_L_X10Y131_SLICE_X12Y131_BQ),
.I4(CLBLM_L_X10Y130_SLICE_X12Y130_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y133_SLICE_X12Y133_DO5),
.O6(CLBLM_L_X10Y133_SLICE_X12Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fef0fe000e000e)
  ) CLBLM_L_X10Y133_SLICE_X12Y133_CLUT (
.I0(CLBLM_L_X10Y133_SLICE_X12Y133_BQ),
.I1(CLBLM_L_X10Y133_SLICE_X12Y133_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X5Y132_SLICE_X7Y132_DO6),
.I4(1'b1),
.I5(CLBLM_R_X11Y133_SLICE_X15Y133_CQ),
.O5(CLBLM_L_X10Y133_SLICE_X12Y133_CO5),
.O6(CLBLM_L_X10Y133_SLICE_X12Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000fe0efe0e)
  ) CLBLM_L_X10Y133_SLICE_X12Y133_BLUT (
.I0(CLBLM_L_X8Y131_SLICE_X11Y131_AQ),
.I1(CLBLM_L_X10Y133_SLICE_X12Y133_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y134_SLICE_X12Y134_BQ),
.I4(1'b1),
.I5(CLBLM_R_X5Y133_SLICE_X7Y133_DO6),
.O5(CLBLM_L_X10Y133_SLICE_X12Y133_BO5),
.O6(CLBLM_L_X10Y133_SLICE_X12Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00ccfaccfa)
  ) CLBLM_L_X10Y133_SLICE_X12Y133_ALUT (
.I0(CLBLM_L_X8Y134_SLICE_X11Y134_BQ),
.I1(CLBLL_L_X4Y134_SLICE_X4Y134_AQ),
.I2(CLBLM_L_X10Y133_SLICE_X12Y133_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLM_R_X5Y133_SLICE_X7Y133_DO6),
.O5(CLBLM_L_X10Y133_SLICE_X12Y133_AO5),
.O6(CLBLM_L_X10Y133_SLICE_X12Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y133_SLICE_X13Y133_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y133_SLICE_X13Y133_AO6),
.Q(CLBLM_L_X10Y133_SLICE_X13Y133_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y133_SLICE_X13Y133_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y133_SLICE_X13Y133_BO6),
.Q(CLBLM_L_X10Y133_SLICE_X13Y133_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000f0f09090909)
  ) CLBLM_L_X10Y133_SLICE_X13Y133_DLUT (
.I0(CLBLM_L_X10Y137_SLICE_X12Y137_CQ),
.I1(CLBLM_R_X11Y132_SLICE_X15Y132_AO6),
.I2(CLBLM_L_X10Y133_SLICE_X13Y133_BQ),
.I3(1'b1),
.I4(CLBLM_L_X10Y134_SLICE_X13Y134_B5Q),
.I5(CLBLM_R_X5Y132_SLICE_X7Y132_DO6),
.O5(CLBLM_L_X10Y133_SLICE_X13Y133_DO5),
.O6(CLBLM_L_X10Y133_SLICE_X13Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000001)
  ) CLBLM_L_X10Y133_SLICE_X13Y133_CLUT (
.I0(CLBLM_L_X10Y131_SLICE_X13Y131_BQ),
.I1(CLBLM_L_X10Y137_SLICE_X12Y137_CQ),
.I2(CLBLM_L_X10Y131_SLICE_X13Y131_CQ),
.I3(CLBLM_L_X8Y137_SLICE_X11Y137_BQ),
.I4(CLBLM_L_X10Y133_SLICE_X13Y133_AQ),
.I5(CLBLM_R_X11Y132_SLICE_X14Y132_AQ),
.O5(CLBLM_L_X10Y133_SLICE_X13Y133_CO5),
.O6(CLBLM_L_X10Y133_SLICE_X13Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hdcdddcdd10111011)
  ) CLBLM_L_X10Y133_SLICE_X13Y133_BLUT (
.I0(CLBLM_L_X10Y133_SLICE_X13Y133_DO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X7Y131_SLICE_X9Y131_AQ),
.I3(RIOB33_X105Y141_IOB_X1Y142_I),
.I4(1'b1),
.I5(CLBLM_L_X10Y134_SLICE_X13Y134_BQ),
.O5(CLBLM_L_X10Y133_SLICE_X13Y133_BO5),
.O6(CLBLM_L_X10Y133_SLICE_X13Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffccfc00330030)
  ) CLBLM_L_X10Y133_SLICE_X13Y133_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y133_SLICE_X13Y133_AQ),
.I3(CLBLM_R_X5Y132_SLICE_X7Y132_DO6),
.I4(CLBLM_L_X8Y137_SLICE_X11Y137_BQ),
.I5(CLBLM_L_X10Y134_SLICE_X13Y134_A5Q),
.O5(CLBLM_L_X10Y133_SLICE_X13Y133_AO5),
.O6(CLBLM_L_X10Y133_SLICE_X13Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y134_SLICE_X12Y134_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y134_SLICE_X12Y134_AO6),
.Q(CLBLM_L_X10Y134_SLICE_X12Y134_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y134_SLICE_X12Y134_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y134_SLICE_X12Y134_BO6),
.Q(CLBLM_L_X10Y134_SLICE_X12Y134_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y134_SLICE_X12Y134_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y134_SLICE_X12Y134_CO6),
.Q(CLBLM_L_X10Y134_SLICE_X12Y134_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y134_SLICE_X12Y134_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y134_SLICE_X12Y134_DO6),
.Q(CLBLM_L_X10Y134_SLICE_X12Y134_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0030303030)
  ) CLBLM_L_X10Y134_SLICE_X12Y134_DLUT (
.I0(1'b1),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_L_X10Y134_SLICE_X12Y134_DQ),
.I3(CLBLM_L_X10Y134_SLICE_X13Y134_B5Q),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y134_SLICE_X12Y134_DO5),
.O6(CLBLM_L_X10Y134_SLICE_X12Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f000440044)
  ) CLBLM_L_X10Y134_SLICE_X12Y134_CLUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_L_X10Y134_SLICE_X12Y134_CQ),
.I2(CLBLM_L_X10Y134_SLICE_X12Y134_DQ),
.I3(CLBLM_L_X8Y138_SLICE_X10Y138_AQ),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y134_SLICE_X12Y134_CO5),
.O6(CLBLM_L_X10Y134_SLICE_X12Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffddff8800dd0088)
  ) CLBLM_L_X10Y134_SLICE_X12Y134_BLUT (
.I0(CLBLM_L_X8Y143_SLICE_X10Y143_DO6),
.I1(CLBLM_L_X10Y134_SLICE_X12Y134_BQ),
.I2(1'b1),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y140_SLICE_X12Y140_A5Q),
.I5(CLBLM_R_X11Y134_SLICE_X14Y134_CQ),
.O5(CLBLM_L_X10Y134_SLICE_X12Y134_BO5),
.O6(CLBLM_L_X10Y134_SLICE_X12Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00ccffccf0)
  ) CLBLM_L_X10Y134_SLICE_X12Y134_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y140_SLICE_X12Y140_AQ),
.I2(CLBLM_L_X10Y134_SLICE_X12Y134_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y133_SLICE_X12Y133_AQ),
.I5(CLBLM_R_X5Y133_SLICE_X7Y133_DO6),
.O5(CLBLM_L_X10Y134_SLICE_X12Y134_AO5),
.O6(CLBLM_L_X10Y134_SLICE_X12Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y134_SLICE_X13Y134_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y140_SLICE_X13Y140_AO6),
.Q(CLBLM_L_X10Y134_SLICE_X13Y134_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y134_SLICE_X13Y134_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y134_SLICE_X13Y134_BO5),
.Q(CLBLM_L_X10Y134_SLICE_X13Y134_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y134_SLICE_X13Y134_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y134_SLICE_X13Y134_AO6),
.Q(CLBLM_L_X10Y134_SLICE_X13Y134_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y134_SLICE_X13Y134_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y134_SLICE_X13Y134_BO6),
.Q(CLBLM_L_X10Y134_SLICE_X13Y134_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffddffff)
  ) CLBLM_L_X10Y134_SLICE_X13Y134_DLUT (
.I0(CLBLL_L_X4Y139_SLICE_X4Y139_BO6),
.I1(CLBLM_R_X13Y138_SLICE_X18Y138_BO6),
.I2(1'b1),
.I3(CLBLL_L_X4Y142_SLICE_X5Y142_DO6),
.I4(CLBLM_L_X8Y135_SLICE_X10Y135_CO6),
.I5(CLBLM_R_X5Y136_SLICE_X7Y136_DO6),
.O5(CLBLM_L_X10Y134_SLICE_X13Y134_DO5),
.O6(CLBLM_L_X10Y134_SLICE_X13Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfe54aa00fcfc0000)
  ) CLBLM_L_X10Y134_SLICE_X13Y134_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y135_SLICE_X12Y135_AQ),
.I2(CLBLM_R_X5Y140_SLICE_X7Y140_BQ),
.I3(CLBLM_R_X11Y134_SLICE_X15Y134_BQ),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y134_SLICE_X13Y134_CO5),
.O6(CLBLM_L_X10Y134_SLICE_X13Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00aaaaf0f0cccc)
  ) CLBLM_L_X10Y134_SLICE_X13Y134_BLUT (
.I0(CLBLM_L_X10Y137_SLICE_X13Y137_DO6),
.I1(CLBLM_L_X10Y134_SLICE_X13Y134_A5Q),
.I2(CLBLM_L_X10Y133_SLICE_X13Y133_BQ),
.I3(CLBLM_L_X10Y137_SLICE_X13Y137_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y134_SLICE_X13Y134_BO5),
.O6(CLBLM_L_X10Y134_SLICE_X13Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfceefc30302230)
  ) CLBLM_L_X10Y134_SLICE_X13Y134_ALUT (
.I0(CLBLM_L_X10Y134_SLICE_X13Y134_DO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y134_SLICE_X13Y134_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_L_X8Y138_SLICE_X10Y138_AQ),
.I5(CLBLM_R_X11Y134_SLICE_X15Y134_CQ),
.O5(CLBLM_L_X10Y134_SLICE_X13Y134_AO5),
.O6(CLBLM_L_X10Y134_SLICE_X13Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y135_SLICE_X12Y135_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y135_SLICE_X12Y135_BO5),
.Q(CLBLM_L_X10Y135_SLICE_X12Y135_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y135_SLICE_X12Y135_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y135_SLICE_X12Y135_AO6),
.Q(CLBLM_L_X10Y135_SLICE_X12Y135_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y135_SLICE_X12Y135_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y135_SLICE_X12Y135_BO6),
.Q(CLBLM_L_X10Y135_SLICE_X12Y135_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000002020202)
  ) CLBLM_L_X10Y135_SLICE_X12Y135_DLUT (
.I0(CLBLM_R_X5Y134_SLICE_X6Y134_AQ),
.I1(CLBLM_R_X11Y135_SLICE_X14Y135_AQ),
.I2(RIOB33_X105Y117_IOB_X1Y118_I),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X8Y138_SLICE_X10Y138_AQ),
.O5(CLBLM_L_X10Y135_SLICE_X12Y135_DO5),
.O6(CLBLM_L_X10Y135_SLICE_X12Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0c0f0d000005050)
  ) CLBLM_L_X10Y135_SLICE_X12Y135_CLUT (
.I0(CLBLL_L_X4Y134_SLICE_X4Y134_AQ),
.I1(CLBLM_L_X10Y137_SLICE_X12Y137_AQ),
.I2(CLBLM_L_X8Y135_SLICE_X11Y135_DO6),
.I3(CLBLM_R_X5Y140_SLICE_X7Y140_BQ),
.I4(CLBLM_L_X8Y135_SLICE_X10Y135_CO6),
.I5(RIOB33_X105Y121_IOB_X1Y121_I),
.O5(CLBLM_L_X10Y135_SLICE_X12Y135_CO5),
.O6(CLBLM_L_X10Y135_SLICE_X12Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f000aaaaaacccc)
  ) CLBLM_L_X10Y135_SLICE_X12Y135_BLUT (
.I0(CLBLM_L_X12Y135_SLICE_X16Y135_DQ),
.I1(CLBLM_R_X11Y139_SLICE_X15Y139_A5Q),
.I2(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y135_SLICE_X12Y135_BO5),
.O6(CLBLM_L_X10Y135_SLICE_X12Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffcec3020)
  ) CLBLM_L_X10Y135_SLICE_X12Y135_ALUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y135_SLICE_X12Y135_AQ),
.I3(CLBLM_L_X8Y138_SLICE_X10Y138_AQ),
.I4(CLBLM_R_X7Y132_SLICE_X8Y132_AQ),
.I5(CLBLM_L_X10Y135_SLICE_X12Y135_CO6),
.O5(CLBLM_L_X10Y135_SLICE_X12Y135_AO5),
.O6(CLBLM_L_X10Y135_SLICE_X12Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y135_SLICE_X13Y135_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y135_SLICE_X13Y135_BO5),
.Q(CLBLM_L_X10Y135_SLICE_X13Y135_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y135_SLICE_X13Y135_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y135_SLICE_X13Y135_BO6),
.Q(CLBLM_L_X10Y135_SLICE_X13Y135_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffcfffffffc)
  ) CLBLM_L_X10Y135_SLICE_X13Y135_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y133_SLICE_X11Y133_BQ),
.I2(CLBLM_L_X12Y135_SLICE_X16Y135_DQ),
.I3(CLBLM_R_X11Y134_SLICE_X14Y134_DQ),
.I4(CLBLM_L_X10Y135_SLICE_X13Y135_B5Q),
.I5(1'b1),
.O5(CLBLM_L_X10Y135_SLICE_X13Y135_DO5),
.O6(CLBLM_L_X10Y135_SLICE_X13Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000fdfdfddd)
  ) CLBLM_L_X10Y135_SLICE_X13Y135_CLUT (
.I0(CLBLM_R_X11Y135_SLICE_X15Y135_CO5),
.I1(CLBLL_L_X4Y142_SLICE_X5Y142_DO6),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLM_L_X10Y138_SLICE_X13Y138_CQ),
.I4(CLBLM_L_X10Y135_SLICE_X13Y135_B5Q),
.I5(CLBLM_L_X8Y137_SLICE_X11Y137_CO5),
.O5(CLBLM_L_X10Y135_SLICE_X13Y135_CO5),
.O6(CLBLM_L_X10Y135_SLICE_X13Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5a0a0ba10ba10)
  ) CLBLM_L_X10Y135_SLICE_X13Y135_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X11Y134_SLICE_X14Y134_DQ),
.I3(CLBLM_R_X11Y138_SLICE_X14Y138_BQ),
.I4(RIOB33_X105Y103_IOB_X1Y103_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y135_SLICE_X13Y135_BO5),
.O6(CLBLM_L_X10Y135_SLICE_X13Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfecc3200fa00fa00)
  ) CLBLM_L_X10Y135_SLICE_X13Y135_ALUT (
.I0(CLBLM_L_X10Y135_SLICE_X13Y135_B5Q),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X11Y135_SLICE_X14Y135_DQ),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(CLBLM_L_X10Y133_SLICE_X13Y133_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y135_SLICE_X13Y135_AO5),
.O6(CLBLM_L_X10Y135_SLICE_X13Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y136_SLICE_X12Y136_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y136_SLICE_X14Y136_CO6),
.Q(CLBLM_L_X10Y136_SLICE_X12Y136_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y136_SLICE_X12Y136_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y136_SLICE_X12Y136_AO6),
.Q(CLBLM_L_X10Y136_SLICE_X12Y136_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y136_SLICE_X12Y136_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y136_SLICE_X12Y136_BO6),
.Q(CLBLM_L_X10Y136_SLICE_X12Y136_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd88dd88cd88cd88)
  ) CLBLM_L_X10Y136_SLICE_X12Y136_DLUT (
.I0(CLBLL_L_X4Y134_SLICE_X4Y134_AQ),
.I1(CLBLM_L_X8Y138_SLICE_X11Y138_CO6),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_L_X10Y134_SLICE_X12Y134_CQ),
.I4(1'b1),
.I5(CLBLL_L_X4Y142_SLICE_X4Y142_BO6),
.O5(CLBLM_L_X10Y136_SLICE_X12Y136_DO5),
.O6(CLBLM_L_X10Y136_SLICE_X12Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000001fffffffc)
  ) CLBLM_L_X10Y136_SLICE_X12Y136_CLUT (
.I0(CLBLM_L_X10Y134_SLICE_X13Y134_AQ),
.I1(CLBLL_L_X4Y136_SLICE_X4Y136_CQ),
.I2(CLBLM_R_X5Y138_SLICE_X6Y138_BQ),
.I3(CLBLM_R_X11Y136_SLICE_X14Y136_BQ),
.I4(CLBLM_L_X10Y136_SLICE_X12Y136_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y136_SLICE_X12Y136_CO5),
.O6(CLBLM_L_X10Y136_SLICE_X12Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f000ee0000)
  ) CLBLM_L_X10Y136_SLICE_X12Y136_BLUT (
.I0(CLBLM_L_X10Y136_SLICE_X12Y136_DO6),
.I1(CLBLM_L_X10Y136_SLICE_X12Y136_BQ),
.I2(CLBLM_L_X10Y136_SLICE_X12Y136_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_L_X8Y138_SLICE_X10Y138_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y136_SLICE_X12Y136_BO5),
.O6(CLBLM_L_X10Y136_SLICE_X12Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccf0cc50ccf0cc50)
  ) CLBLM_L_X10Y136_SLICE_X12Y136_ALUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_L_X10Y134_SLICE_X13Y134_AQ),
.I2(CLBLM_L_X10Y136_SLICE_X12Y136_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y138_SLICE_X10Y138_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y136_SLICE_X12Y136_AO5),
.O6(CLBLM_L_X10Y136_SLICE_X12Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000400000)
  ) CLBLM_L_X10Y136_SLICE_X13Y136_DLUT (
.I0(CLBLM_R_X13Y135_SLICE_X18Y135_BQ),
.I1(CLBLM_R_X7Y134_SLICE_X8Y134_DO6),
.I2(CLBLM_L_X8Y140_SLICE_X11Y140_AQ),
.I3(RIOB33_X105Y133_IOB_X1Y134_I),
.I4(CLBLM_L_X8Y143_SLICE_X10Y143_DO6),
.I5(CLBLM_L_X10Y136_SLICE_X12Y136_CO5),
.O5(CLBLM_L_X10Y136_SLICE_X13Y136_DO5),
.O6(CLBLM_L_X10Y136_SLICE_X13Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa88aa80aaaaaaa2)
  ) CLBLM_L_X10Y136_SLICE_X13Y136_CLUT (
.I0(RIOB33_X105Y121_IOB_X1Y121_I),
.I1(CLBLM_L_X10Y136_SLICE_X12Y136_CO5),
.I2(CLBLL_L_X4Y141_SLICE_X4Y141_DO6),
.I3(CLBLM_R_X13Y137_SLICE_X18Y137_AQ),
.I4(CLBLM_R_X13Y138_SLICE_X18Y138_BO6),
.I5(CLBLM_L_X10Y134_SLICE_X13Y134_AQ),
.O5(CLBLM_L_X10Y136_SLICE_X13Y136_CO5),
.O6(CLBLM_L_X10Y136_SLICE_X13Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h08cc0ccc00c000c0)
  ) CLBLM_L_X10Y136_SLICE_X13Y136_BLUT (
.I0(CLBLL_L_X4Y141_SLICE_X4Y141_DO6),
.I1(CLBLM_L_X12Y135_SLICE_X17Y135_BO5),
.I2(CLBLL_L_X4Y134_SLICE_X4Y134_AQ),
.I3(CLBLM_L_X8Y136_SLICE_X11Y136_DO5),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_L_X10Y134_SLICE_X12Y134_CQ),
.O5(CLBLM_L_X10Y136_SLICE_X13Y136_BO5),
.O6(CLBLM_L_X10Y136_SLICE_X13Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_L_X10Y136_SLICE_X13Y136_ALUT (
.I0(CLBLM_R_X7Y139_SLICE_X8Y139_A5Q),
.I1(CLBLM_R_X11Y137_SLICE_X15Y137_BO6),
.I2(CLBLM_L_X10Y135_SLICE_X13Y135_DO6),
.I3(CLBLM_R_X11Y136_SLICE_X15Y136_BQ),
.I4(CLBLM_L_X10Y141_SLICE_X13Y141_BQ),
.I5(CLBLM_R_X7Y139_SLICE_X9Y139_A5Q),
.O5(CLBLM_L_X10Y136_SLICE_X13Y136_AO5),
.O6(CLBLM_L_X10Y136_SLICE_X13Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y137_SLICE_X12Y137_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y137_SLICE_X12Y137_BO5),
.Q(CLBLM_L_X10Y137_SLICE_X12Y137_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y137_SLICE_X12Y137_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y137_SLICE_X12Y137_AO6),
.Q(CLBLM_L_X10Y137_SLICE_X12Y137_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y137_SLICE_X12Y137_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y137_SLICE_X12Y137_BO6),
.Q(CLBLM_L_X10Y137_SLICE_X12Y137_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y137_SLICE_X12Y137_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y137_SLICE_X12Y137_CO6),
.Q(CLBLM_L_X10Y137_SLICE_X12Y137_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffafffa)
  ) CLBLM_L_X10Y137_SLICE_X12Y137_DLUT (
.I0(CLBLM_R_X7Y132_SLICE_X8Y132_BQ),
.I1(1'b1),
.I2(CLBLM_R_X11Y138_SLICE_X15Y138_B5Q),
.I3(CLBLM_R_X11Y133_SLICE_X14Y133_CQ),
.I4(1'b1),
.I5(CLBLM_L_X8Y135_SLICE_X10Y135_BQ),
.O5(CLBLM_L_X10Y137_SLICE_X12Y137_DO5),
.O6(CLBLM_L_X10Y137_SLICE_X12Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf055f044f055f044)
  ) CLBLM_L_X10Y137_SLICE_X12Y137_CLUT (
.I0(CLBLM_R_X5Y132_SLICE_X7Y132_DO6),
.I1(CLBLM_L_X10Y137_SLICE_X12Y137_CQ),
.I2(CLBLM_L_X8Y140_SLICE_X11Y140_BQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X11Y133_SLICE_X15Y133_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y137_SLICE_X12Y137_CO5),
.O6(CLBLM_L_X10Y137_SLICE_X12Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fff000ccaaccaa)
  ) CLBLM_L_X10Y137_SLICE_X12Y137_BLUT (
.I0(CLBLM_L_X10Y136_SLICE_X12Y136_A5Q),
.I1(CLBLL_L_X4Y137_SLICE_X5Y137_BQ),
.I2(CLBLM_L_X10Y143_SLICE_X12Y143_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X12Y136_SLICE_X17Y136_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X10Y137_SLICE_X12Y137_BO5),
.O6(CLBLM_L_X10Y137_SLICE_X12Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00fafac8c8)
  ) CLBLM_L_X10Y137_SLICE_X12Y137_ALUT (
.I0(CLBLM_L_X8Y137_SLICE_X11Y137_DO6),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_L_X10Y137_SLICE_X12Y137_AQ),
.I3(CLBLM_R_X11Y142_SLICE_X15Y142_BQ),
.I4(CLBLM_L_X8Y138_SLICE_X10Y138_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y137_SLICE_X12Y137_AO5),
.O6(CLBLM_L_X10Y137_SLICE_X12Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y137_SLICE_X13Y137_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y137_SLICE_X13Y137_AO6),
.Q(CLBLM_L_X10Y137_SLICE_X13Y137_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y137_SLICE_X13Y137_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y137_SLICE_X13Y137_BO6),
.Q(CLBLM_L_X10Y137_SLICE_X13Y137_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h1221122184488448)
  ) CLBLM_L_X10Y137_SLICE_X13Y137_DLUT (
.I0(CLBLM_R_X11Y137_SLICE_X14Y137_AQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_L_X10Y137_SLICE_X13Y137_BQ),
.I3(CLBLL_L_X4Y138_SLICE_X5Y138_BQ),
.I4(1'b1),
.I5(CLBLM_L_X10Y134_SLICE_X13Y134_BQ),
.O5(CLBLM_L_X10Y137_SLICE_X13Y137_DO5),
.O6(CLBLM_L_X10Y137_SLICE_X13Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfb00ae00ff00aa00)
  ) CLBLM_L_X10Y137_SLICE_X13Y137_CLUT (
.I0(CLBLM_L_X10Y141_SLICE_X13Y141_BQ),
.I1(CLBLM_L_X10Y139_SLICE_X13Y139_AQ),
.I2(CLBLM_R_X11Y139_SLICE_X15Y139_CQ),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(CLBLM_R_X11Y138_SLICE_X15Y138_B5Q),
.I5(CLBLM_L_X8Y137_SLICE_X10Y137_BO6),
.O5(CLBLM_L_X10Y137_SLICE_X13Y137_CO5),
.O6(CLBLM_L_X10Y137_SLICE_X13Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haabbbbaa00111100)
  ) CLBLM_L_X10Y137_SLICE_X13Y137_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(1'b1),
.I3(CLBLM_R_X11Y137_SLICE_X14Y137_CO6),
.I4(CLBLM_R_X11Y137_SLICE_X14Y137_AQ),
.I5(CLBLM_L_X8Y135_SLICE_X11Y135_A5Q),
.O5(CLBLM_L_X10Y137_SLICE_X13Y137_BO5),
.O6(CLBLM_L_X10Y137_SLICE_X13Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaf0005aafa0050)
  ) CLBLM_L_X10Y137_SLICE_X13Y137_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(1'b1),
.I2(CLBLM_L_X8Y139_SLICE_X10Y139_BQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_L_X12Y137_SLICE_X16Y137_AQ),
.I5(CLBLM_L_X10Y138_SLICE_X12Y138_CO6),
.O5(CLBLM_L_X10Y137_SLICE_X13Y137_AO5),
.O6(CLBLM_L_X10Y137_SLICE_X13Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y138_SLICE_X12Y138_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y137_SLICE_X14Y137_BO6),
.Q(CLBLM_L_X10Y138_SLICE_X12Y138_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y138_SLICE_X12Y138_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y138_SLICE_X12Y138_AO6),
.Q(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hafafafafafafafaf)
  ) CLBLM_L_X10Y138_SLICE_X12Y138_DLUT (
.I0(CLBLM_R_X7Y136_SLICE_X9Y136_CQ),
.I1(1'b1),
.I2(CLBLM_R_X5Y136_SLICE_X7Y136_BQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y138_SLICE_X12Y138_DO5),
.O6(CLBLM_L_X10Y138_SLICE_X12Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0d0f000f202)
  ) CLBLM_L_X10Y138_SLICE_X12Y138_CLUT (
.I0(CLBLM_L_X10Y139_SLICE_X13Y139_AQ),
.I1(CLBLM_R_X11Y139_SLICE_X15Y139_CQ),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLM_R_X11Y136_SLICE_X15Y136_BQ),
.I4(CLBLM_L_X10Y138_SLICE_X12Y138_DO6),
.I5(CLBLM_L_X8Y138_SLICE_X11Y138_BQ),
.O5(CLBLM_L_X10Y138_SLICE_X12Y138_CO5),
.O6(CLBLM_L_X10Y138_SLICE_X12Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff02fdfffff3f3)
  ) CLBLM_L_X10Y138_SLICE_X12Y138_BLUT (
.I0(CLBLM_R_X5Y136_SLICE_X7Y136_BQ),
.I1(CLBLM_R_X7Y136_SLICE_X9Y136_CQ),
.I2(CLBLM_L_X10Y139_SLICE_X13Y139_AQ),
.I3(CLBLM_L_X10Y139_SLICE_X13Y139_BQ),
.I4(CLBLM_R_X11Y139_SLICE_X15Y139_CQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y138_SLICE_X12Y138_BO5),
.O6(CLBLM_L_X10Y138_SLICE_X12Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc05055050)
  ) CLBLM_L_X10Y138_SLICE_X12Y138_ALUT (
.I0(CLBLM_R_X11Y135_SLICE_X14Y135_AQ),
.I1(CLBLM_R_X11Y133_SLICE_X14Y133_BQ),
.I2(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I3(1'b1),
.I4(CLBLM_R_X7Y138_SLICE_X9Y138_CO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y138_SLICE_X12Y138_AO5),
.O6(CLBLM_L_X10Y138_SLICE_X12Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y138_SLICE_X13Y138_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y138_SLICE_X13Y138_AO6),
.Q(CLBLM_L_X10Y138_SLICE_X13Y138_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y138_SLICE_X13Y138_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y138_SLICE_X13Y138_BO6),
.Q(CLBLM_L_X10Y138_SLICE_X13Y138_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y138_SLICE_X13Y138_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y138_SLICE_X13Y138_CO6),
.Q(CLBLM_L_X10Y138_SLICE_X13Y138_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff33df13cc00ec20)
  ) CLBLM_L_X10Y138_SLICE_X13Y138_DLUT (
.I0(CLBLM_R_X7Y136_SLICE_X9Y136_CQ),
.I1(RIOB33_X105Y121_IOB_X1Y121_I),
.I2(CLBLM_R_X11Y139_SLICE_X14Y139_DO6),
.I3(CLBLM_L_X10Y135_SLICE_X12Y135_BQ),
.I4(CLBLM_R_X5Y136_SLICE_X7Y136_BQ),
.I5(CLBLM_L_X10Y139_SLICE_X12Y139_BQ),
.O5(CLBLM_L_X10Y138_SLICE_X13Y138_DO5),
.O6(CLBLM_L_X10Y138_SLICE_X13Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00fafac8c8)
  ) CLBLM_L_X10Y138_SLICE_X13Y138_CLUT (
.I0(CLBLM_L_X8Y138_SLICE_X10Y138_AQ),
.I1(CLBLM_L_X10Y138_SLICE_X13Y138_CQ),
.I2(RIOB33_X105Y117_IOB_X1Y118_I),
.I3(CLBLM_R_X13Y136_SLICE_X18Y136_BQ),
.I4(CLBLM_L_X10Y138_SLICE_X13Y138_DO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y138_SLICE_X13Y138_CO5),
.O6(CLBLM_L_X10Y138_SLICE_X13Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00eeee0000)
  ) CLBLM_L_X10Y138_SLICE_X13Y138_BLUT (
.I0(CLBLM_R_X11Y140_SLICE_X15Y140_DQ),
.I1(CLBLM_L_X10Y138_SLICE_X13Y138_BQ),
.I2(1'b1),
.I3(CLBLM_R_X7Y136_SLICE_X9Y136_CQ),
.I4(CLBLM_L_X8Y143_SLICE_X10Y143_DO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y138_SLICE_X13Y138_BO5),
.O6(CLBLM_L_X10Y138_SLICE_X13Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffc4c8c4c8c4c8)
  ) CLBLM_L_X10Y138_SLICE_X13Y138_ALUT (
.I0(CLBLM_L_X10Y139_SLICE_X13Y139_DO6),
.I1(CLBLM_L_X12Y135_SLICE_X17Y135_BO5),
.I2(CLBLM_L_X10Y138_SLICE_X13Y138_AQ),
.I3(CLBLM_L_X10Y136_SLICE_X13Y136_CO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X10Y140_SLICE_X13Y140_BQ),
.O5(CLBLM_L_X10Y138_SLICE_X13Y138_AO5),
.O6(CLBLM_L_X10Y138_SLICE_X13Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y139_SLICE_X12Y139_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y139_SLICE_X12Y139_AO6),
.Q(CLBLM_L_X10Y139_SLICE_X12Y139_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y139_SLICE_X12Y139_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y139_SLICE_X12Y139_BO6),
.Q(CLBLM_L_X10Y139_SLICE_X12Y139_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333333333333332)
  ) CLBLM_L_X10Y139_SLICE_X12Y139_DLUT (
.I0(CLBLM_L_X10Y140_SLICE_X12Y140_BQ),
.I1(CLBLM_R_X13Y141_SLICE_X19Y141_BQ),
.I2(CLBLM_L_X10Y137_SLICE_X12Y137_DO6),
.I3(CLBLM_L_X10Y139_SLICE_X12Y139_CO6),
.I4(CLBLM_L_X8Y141_SLICE_X10Y141_CQ),
.I5(CLBLM_L_X10Y139_SLICE_X13Y139_BQ),
.O5(CLBLM_L_X10Y139_SLICE_X12Y139_DO5),
.O6(CLBLM_L_X10Y139_SLICE_X12Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_L_X10Y139_SLICE_X12Y139_CLUT (
.I0(CLBLM_R_X11Y139_SLICE_X14Y139_BQ),
.I1(CLBLM_R_X5Y137_SLICE_X7Y137_BQ),
.I2(CLBLM_L_X10Y139_SLICE_X12Y139_BQ),
.I3(CLBLM_L_X8Y138_SLICE_X11Y138_BQ),
.I4(CLBLM_L_X10Y134_SLICE_X12Y134_DQ),
.I5(CLBLM_L_X8Y144_SLICE_X11Y144_AQ),
.O5(CLBLM_L_X10Y139_SLICE_X12Y139_CO5),
.O6(CLBLM_L_X10Y139_SLICE_X12Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0cff0c000c000c)
  ) CLBLM_L_X10Y139_SLICE_X12Y139_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y139_SLICE_X12Y139_BQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLM_L_X8Y136_SLICE_X11Y136_CQ),
.O5(CLBLM_L_X10Y139_SLICE_X12Y139_BO5),
.O6(CLBLM_L_X10Y139_SLICE_X12Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccfffaffff)
  ) CLBLM_L_X10Y139_SLICE_X12Y139_ALUT (
.I0(RIOB33_X105Y135_IOB_X1Y135_I),
.I1(CLBLM_L_X10Y140_SLICE_X12Y140_BQ),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(CLBLM_R_X13Y139_SLICE_X18Y139_BO6),
.I4(RIOB33_X105Y135_IOB_X1Y136_I),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y139_SLICE_X12Y139_AO5),
.O6(CLBLM_L_X10Y139_SLICE_X12Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y139_SLICE_X13Y139_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y139_SLICE_X13Y139_BO5),
.Q(CLBLM_L_X10Y139_SLICE_X13Y139_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y139_SLICE_X13Y139_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y139_SLICE_X13Y139_AO6),
.Q(CLBLM_L_X10Y139_SLICE_X13Y139_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y139_SLICE_X13Y139_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y139_SLICE_X13Y139_BO6),
.Q(CLBLM_L_X10Y139_SLICE_X13Y139_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y139_SLICE_X13Y139_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y139_SLICE_X13Y139_CO6),
.Q(CLBLM_L_X10Y139_SLICE_X13Y139_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h56fca9039a3065cf)
  ) CLBLM_L_X10Y139_SLICE_X13Y139_DLUT (
.I0(CLBLM_L_X8Y137_SLICE_X10Y137_BO6),
.I1(CLBLM_L_X10Y140_SLICE_X13Y140_CQ),
.I2(CLBLM_L_X10Y139_SLICE_X12Y139_DO6),
.I3(CLBLM_R_X11Y139_SLICE_X14Y139_DO6),
.I4(CLBLM_L_X12Y135_SLICE_X17Y135_AQ),
.I5(CLBLM_R_X13Y141_SLICE_X19Y141_BQ),
.O5(CLBLM_L_X10Y139_SLICE_X13Y139_DO5),
.O6(CLBLM_L_X10Y139_SLICE_X13Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f000fff0f00033)
  ) CLBLM_L_X10Y139_SLICE_X13Y139_CLUT (
.I0(1'b1),
.I1(RIOB33_X105Y141_IOB_X1Y142_I),
.I2(CLBLM_L_X8Y142_SLICE_X11Y142_AQ),
.I3(CLBLM_R_X11Y135_SLICE_X15Y135_DO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y131_SLICE_X9Y131_AQ),
.O5(CLBLM_L_X10Y139_SLICE_X13Y139_CO5),
.O6(CLBLM_L_X10Y139_SLICE_X13Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f000ccccccaaaa)
  ) CLBLM_L_X10Y139_SLICE_X13Y139_BLUT (
.I0(CLBLM_R_X7Y136_SLICE_X8Y136_AQ),
.I1(CLBLM_L_X10Y139_SLICE_X13Y139_BQ),
.I2(CLBLM_R_X11Y144_SLICE_X15Y144_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y139_SLICE_X13Y139_BO5),
.O6(CLBLM_L_X10Y139_SLICE_X13Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0030300000)
  ) CLBLM_L_X10Y139_SLICE_X13Y139_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y139_SLICE_X9Y139_AQ),
.I2(CLBLM_L_X10Y139_SLICE_X13Y139_AQ),
.I3(CLBLM_L_X10Y139_SLICE_X12Y139_BQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y139_SLICE_X13Y139_AO5),
.O6(CLBLM_L_X10Y139_SLICE_X13Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y140_SLICE_X12Y140_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y141_SLICE_X12Y141_BO6),
.Q(CLBLM_L_X10Y140_SLICE_X12Y140_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y140_SLICE_X12Y140_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y140_SLICE_X12Y140_AO6),
.Q(CLBLM_L_X10Y140_SLICE_X12Y140_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y140_SLICE_X12Y140_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y140_SLICE_X12Y140_BO6),
.Q(CLBLM_L_X10Y140_SLICE_X12Y140_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y140_SLICE_X12Y140_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y140_SLICE_X12Y140_CO6),
.Q(CLBLM_L_X10Y140_SLICE_X12Y140_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffffdf)
  ) CLBLM_L_X10Y140_SLICE_X12Y140_DLUT (
.I0(CLBLM_L_X10Y140_SLICE_X12Y140_A5Q),
.I1(CLBLM_R_X11Y140_SLICE_X14Y140_DO6),
.I2(CLBLM_R_X11Y141_SLICE_X15Y141_DQ),
.I3(CLBLM_R_X11Y140_SLICE_X15Y140_BQ),
.I4(CLBLM_L_X10Y140_SLICE_X12Y140_BO5),
.I5(CLBLM_L_X10Y140_SLICE_X13Y140_BQ),
.O5(CLBLM_L_X10Y140_SLICE_X12Y140_DO5),
.O6(CLBLM_L_X10Y140_SLICE_X12Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaafcfcfc00)
  ) CLBLM_L_X10Y140_SLICE_X12Y140_CLUT (
.I0(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I1(CLBLM_L_X10Y140_SLICE_X12Y140_CQ),
.I2(CLBLM_L_X10Y136_SLICE_X12Y136_DO6),
.I3(CLBLM_L_X8Y138_SLICE_X10Y138_AQ),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y140_SLICE_X12Y140_CO5),
.O6(CLBLM_L_X10Y140_SLICE_X12Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf088f088ffaaffff)
  ) CLBLM_L_X10Y140_SLICE_X12Y140_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X10Y140_SLICE_X12Y140_BQ),
.I2(CLBLM_L_X10Y140_SLICE_X12Y140_CQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y140_SLICE_X11Y140_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y140_SLICE_X12Y140_BO5),
.O6(CLBLM_L_X10Y140_SLICE_X12Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffc8ffc800c800c8)
  ) CLBLM_L_X10Y140_SLICE_X12Y140_ALUT (
.I0(CLBLM_L_X12Y140_SLICE_X16Y140_DQ),
.I1(CLBLM_L_X8Y143_SLICE_X10Y143_DO6),
.I2(CLBLM_L_X10Y140_SLICE_X12Y140_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLM_L_X10Y141_SLICE_X12Y141_CQ),
.O5(CLBLM_L_X10Y140_SLICE_X12Y140_AO5),
.O6(CLBLM_L_X10Y140_SLICE_X12Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y140_SLICE_X13Y140_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y140_SLICE_X13Y140_CO5),
.Q(CLBLM_L_X10Y140_SLICE_X13Y140_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y140_SLICE_X13Y140_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y140_SLICE_X13Y140_BO6),
.Q(CLBLM_L_X10Y140_SLICE_X13Y140_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y140_SLICE_X13Y140_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y140_SLICE_X13Y140_CO6),
.Q(CLBLM_L_X10Y140_SLICE_X13Y140_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y140_SLICE_X13Y140_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y140_SLICE_X13Y140_DO6),
.Q(CLBLM_L_X10Y140_SLICE_X13Y140_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc05055050)
  ) CLBLM_L_X10Y140_SLICE_X13Y140_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X7Y133_SLICE_X9Y133_CQ),
.I2(CLBLM_R_X11Y141_SLICE_X15Y141_DQ),
.I3(1'b1),
.I4(CLBLM_L_X10Y134_SLICE_X13Y134_CO5),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y140_SLICE_X13Y140_DO5),
.O6(CLBLM_L_X10Y140_SLICE_X13Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa0caa0cccffcc00)
  ) CLBLM_L_X10Y140_SLICE_X13Y140_CLUT (
.I0(CLBLM_R_X11Y140_SLICE_X15Y140_DQ),
.I1(CLBLM_L_X10Y140_SLICE_X13Y140_CQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X5Y141_SLICE_X7Y141_DO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y140_SLICE_X13Y140_CO5),
.O6(CLBLM_L_X10Y140_SLICE_X13Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0d1d1c0c0e2e2)
  ) CLBLM_L_X10Y140_SLICE_X13Y140_BLUT (
.I0(CLBLM_L_X12Y138_SLICE_X16Y138_DQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X5Y138_SLICE_X6Y138_BQ),
.I3(1'b1),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_L_X10Y140_SLICE_X13Y140_AO5),
.O5(CLBLM_L_X10Y140_SLICE_X13Y140_BO5),
.O6(CLBLM_L_X10Y140_SLICE_X13Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0eef000eeee0000)
  ) CLBLM_L_X10Y140_SLICE_X13Y140_ALUT (
.I0(CLBLM_L_X10Y135_SLICE_X12Y135_BQ),
.I1(CLBLM_L_X10Y140_SLICE_X12Y140_CQ),
.I2(CLBLM_R_X3Y138_SLICE_X3Y138_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y140_SLICE_X13Y140_AO5),
.O6(CLBLM_L_X10Y140_SLICE_X13Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y141_SLICE_X12Y141_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y141_SLICE_X12Y141_CO5),
.Q(CLBLM_L_X10Y141_SLICE_X12Y141_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y141_SLICE_X12Y141_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y141_SLICE_X12Y141_AO6),
.Q(CLBLM_L_X10Y141_SLICE_X12Y141_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y141_SLICE_X12Y141_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y141_SLICE_X12Y141_CO6),
.Q(CLBLM_L_X10Y141_SLICE_X12Y141_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0004000000000000)
  ) CLBLM_L_X10Y141_SLICE_X12Y141_DLUT (
.I0(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I1(CLBLM_L_X12Y144_SLICE_X17Y144_AQ),
.I2(CLBLM_R_X11Y141_SLICE_X15Y141_AQ),
.I3(CLBLM_R_X11Y139_SLICE_X15Y139_DQ),
.I4(CLBLM_L_X10Y141_SLICE_X12Y141_BO5),
.I5(CLBLM_L_X8Y140_SLICE_X11Y140_CO5),
.O5(CLBLM_L_X10Y141_SLICE_X12Y141_DO5),
.O6(CLBLM_L_X10Y141_SLICE_X12Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd88dd88faf0faf0)
  ) CLBLM_L_X10Y141_SLICE_X12Y141_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X11Y135_SLICE_X14Y135_AQ),
.I2(CLBLM_L_X10Y145_SLICE_X13Y145_CO6),
.I3(CLBLM_L_X10Y138_SLICE_X12Y138_A5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y141_SLICE_X12Y141_CO5),
.O6(CLBLM_L_X10Y141_SLICE_X12Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hae04ae0400003333)
  ) CLBLM_L_X10Y141_SLICE_X12Y141_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X11Y141_SLICE_X14Y141_AQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X7Y135_SLICE_X9Y135_AQ),
.I4(CLBLM_L_X12Y140_SLICE_X16Y140_DQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y141_SLICE_X12Y141_BO5),
.O6(CLBLM_L_X10Y141_SLICE_X12Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffc000c0ffeaaaea)
  ) CLBLM_L_X10Y141_SLICE_X12Y141_ALUT (
.I0(CLBLM_L_X10Y141_SLICE_X12Y141_DO6),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_L_X10Y141_SLICE_X12Y141_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y131_SLICE_X10Y131_AQ),
.I5(CLBLM_L_X10Y140_SLICE_X12Y140_DO6),
.O5(CLBLM_L_X10Y141_SLICE_X12Y141_AO5),
.O6(CLBLM_L_X10Y141_SLICE_X12Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y141_SLICE_X13Y141_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y141_SLICE_X13Y141_AO5),
.Q(CLBLM_L_X10Y141_SLICE_X13Y141_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y141_SLICE_X13Y141_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y141_SLICE_X13Y141_AO6),
.Q(CLBLM_L_X10Y141_SLICE_X13Y141_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y141_SLICE_X13Y141_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y141_SLICE_X13Y141_BO6),
.Q(CLBLM_L_X10Y141_SLICE_X13Y141_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y141_SLICE_X13Y141_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y141_SLICE_X13Y141_CO6),
.Q(CLBLM_L_X10Y141_SLICE_X13Y141_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000080000000000)
  ) CLBLM_L_X10Y141_SLICE_X13Y141_DLUT (
.I0(CLBLM_R_X7Y140_SLICE_X8Y140_DO6),
.I1(CLBLM_L_X12Y141_SLICE_X17Y141_BO6),
.I2(CLBLM_R_X13Y137_SLICE_X18Y137_DO6),
.I3(CLBLM_R_X11Y143_SLICE_X14Y143_BO6),
.I4(CLBLL_L_X4Y141_SLICE_X4Y141_DO6),
.I5(CLBLM_L_X10Y136_SLICE_X13Y136_DO6),
.O5(CLBLM_L_X10Y141_SLICE_X13Y141_DO5),
.O6(CLBLM_L_X10Y141_SLICE_X13Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa0fff0ccc)
  ) CLBLM_L_X10Y141_SLICE_X13Y141_CLUT (
.I0(CLBLM_L_X12Y136_SLICE_X16Y136_DQ),
.I1(CLBLM_L_X10Y141_SLICE_X13Y141_CQ),
.I2(CLBLM_L_X10Y139_SLICE_X13Y139_B5Q),
.I3(CLBLM_L_X12Y134_SLICE_X17Y134_AO6),
.I4(CLBLM_L_X8Y138_SLICE_X10Y138_BQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y141_SLICE_X13Y141_CO5),
.O6(CLBLM_L_X10Y141_SLICE_X13Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfccc3000fccc3000)
  ) CLBLM_L_X10Y141_SLICE_X13Y141_BLUT (
.I0(1'b1),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_L_X12Y136_SLICE_X16Y136_AQ),
.I4(CLBLM_L_X10Y141_SLICE_X12Y141_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y141_SLICE_X13Y141_BO5),
.O6(CLBLM_L_X10Y141_SLICE_X13Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fff000aaffaa00)
  ) CLBLM_L_X10Y141_SLICE_X13Y141_ALUT (
.I0(CLBLM_R_X11Y142_SLICE_X15Y142_CQ),
.I1(1'b1),
.I2(CLBLL_L_X4Y134_SLICE_X5Y134_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y143_IOB_X1Y144_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y141_SLICE_X13Y141_AO5),
.O6(CLBLM_L_X10Y141_SLICE_X13Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y142_SLICE_X12Y142_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y142_SLICE_X12Y142_AO6),
.Q(CLBLM_L_X10Y142_SLICE_X12Y142_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y142_SLICE_X12Y142_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y142_SLICE_X12Y142_BO6),
.Q(CLBLM_L_X10Y142_SLICE_X12Y142_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y142_SLICE_X12Y142_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y142_SLICE_X12Y142_CO6),
.Q(CLBLM_L_X10Y142_SLICE_X12Y142_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y142_SLICE_X12Y142_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y142_SLICE_X12Y142_DO6),
.Q(CLBLM_L_X10Y142_SLICE_X12Y142_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hafaaafaa05000500)
  ) CLBLM_L_X10Y142_SLICE_X12Y142_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(1'b1),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X7Y135_SLICE_X8Y135_CQ),
.I4(1'b1),
.I5(CLBLM_L_X10Y142_SLICE_X13Y142_BQ),
.O5(CLBLM_L_X10Y142_SLICE_X12Y142_DO5),
.O6(CLBLM_L_X10Y142_SLICE_X12Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hbb11aa00fe54aa00)
  ) CLBLM_L_X10Y142_SLICE_X12Y142_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y142_SLICE_X12Y142_CQ),
.I2(CLBLM_L_X10Y145_SLICE_X13Y145_BO6),
.I3(CLBLM_L_X8Y133_SLICE_X10Y133_BQ),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(CLBLM_R_X11Y143_SLICE_X14Y143_BO6),
.O5(CLBLM_L_X10Y142_SLICE_X12Y142_CO5),
.O6(CLBLM_L_X10Y142_SLICE_X12Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf4fff4f0040f0400)
  ) CLBLM_L_X10Y142_SLICE_X12Y142_BLUT (
.I0(CLBLM_L_X10Y145_SLICE_X13Y145_BO6),
.I1(CLBLM_L_X10Y142_SLICE_X12Y142_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y144_SLICE_X11Y144_CO6),
.I4(CLBLM_L_X10Y142_SLICE_X13Y142_AQ),
.I5(CLBLM_L_X8Y140_SLICE_X11Y140_A5Q),
.O5(CLBLM_L_X10Y142_SLICE_X12Y142_BO5),
.O6(CLBLM_L_X10Y142_SLICE_X12Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff734000007340)
  ) CLBLM_L_X10Y142_SLICE_X12Y142_ALUT (
.I0(CLBLM_L_X10Y145_SLICE_X13Y145_BO6),
.I1(CLBLM_L_X8Y144_SLICE_X11Y144_CO6),
.I2(CLBLM_L_X10Y142_SLICE_X12Y142_AQ),
.I3(CLBLM_L_X10Y143_SLICE_X12Y143_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLL_L_X4Y136_SLICE_X5Y136_CQ),
.O5(CLBLM_L_X10Y142_SLICE_X12Y142_AO5),
.O6(CLBLM_L_X10Y142_SLICE_X12Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y142_SLICE_X13Y142_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y142_SLICE_X13Y142_AO6),
.Q(CLBLM_L_X10Y142_SLICE_X13Y142_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y142_SLICE_X13Y142_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y142_SLICE_X13Y142_BO6),
.Q(CLBLM_L_X10Y142_SLICE_X13Y142_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y142_SLICE_X13Y142_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y142_SLICE_X13Y142_CO6),
.Q(CLBLM_L_X10Y142_SLICE_X13Y142_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hc3c3c9c3c3c3c9c3)
  ) CLBLM_L_X10Y142_SLICE_X13Y142_DLUT (
.I0(CLBLM_L_X10Y142_SLICE_X13Y142_BQ),
.I1(CLBLM_L_X10Y142_SLICE_X13Y142_CQ),
.I2(CLBLM_L_X10Y144_SLICE_X13Y144_DO6),
.I3(CLBLM_L_X10Y144_SLICE_X13Y144_CO6),
.I4(CLBLM_L_X10Y145_SLICE_X12Y145_CO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y142_SLICE_X13Y142_DO5),
.O6(CLBLM_L_X10Y142_SLICE_X13Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00dddddd00dd00dd)
  ) CLBLM_L_X10Y142_SLICE_X13Y142_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y138_SLICE_X10Y138_BQ),
.I2(1'b1),
.I3(CLBLM_R_X11Y144_SLICE_X14Y144_DO6),
.I4(CLBLM_L_X10Y142_SLICE_X13Y142_DO6),
.I5(CLBLM_L_X10Y144_SLICE_X12Y144_AO6),
.O5(CLBLM_L_X10Y142_SLICE_X13Y142_CO5),
.O6(CLBLM_L_X10Y142_SLICE_X13Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf4fff4f0040f0400)
  ) CLBLM_L_X10Y142_SLICE_X13Y142_BLUT (
.I0(CLBLM_L_X10Y145_SLICE_X13Y145_BO6),
.I1(CLBLM_L_X10Y142_SLICE_X13Y142_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y144_SLICE_X11Y144_CO6),
.I4(CLBLM_L_X10Y142_SLICE_X12Y142_AQ),
.I5(CLBLM_L_X10Y133_SLICE_X12Y133_CQ),
.O5(CLBLM_L_X10Y142_SLICE_X13Y142_BO5),
.O6(CLBLM_L_X10Y142_SLICE_X13Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaee0044faee5044)
  ) CLBLM_L_X10Y142_SLICE_X13Y142_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y142_SLICE_X13Y142_BQ),
.I2(CLBLM_L_X10Y142_SLICE_X13Y142_AQ),
.I3(CLBLM_L_X8Y144_SLICE_X11Y144_CO6),
.I4(CLBLM_L_X10Y135_SLICE_X12Y135_AQ),
.I5(CLBLM_L_X10Y145_SLICE_X13Y145_BO6),
.O5(CLBLM_L_X10Y142_SLICE_X13Y142_AO5),
.O6(CLBLM_L_X10Y142_SLICE_X13Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y143_SLICE_X12Y143_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y143_SLICE_X12Y143_AO6),
.Q(CLBLM_L_X10Y143_SLICE_X12Y143_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y143_SLICE_X12Y143_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y143_SLICE_X12Y143_BO6),
.Q(CLBLM_L_X10Y143_SLICE_X12Y143_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y143_SLICE_X12Y143_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y143_SLICE_X12Y143_CO6),
.Q(CLBLM_L_X10Y143_SLICE_X12Y143_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hc3c3c9c3c3c3c3c9)
  ) CLBLM_L_X10Y143_SLICE_X12Y143_DLUT (
.I0(CLBLM_L_X10Y143_SLICE_X12Y143_BQ),
.I1(CLBLM_L_X10Y143_SLICE_X12Y143_AQ),
.I2(CLBLM_L_X10Y144_SLICE_X13Y144_DO6),
.I3(CLBLM_L_X10Y145_SLICE_X12Y145_BO6),
.I4(CLBLM_L_X10Y145_SLICE_X12Y145_CO6),
.I5(CLBLM_R_X11Y144_SLICE_X15Y144_BQ),
.O5(CLBLM_L_X10Y143_SLICE_X12Y143_DO5),
.O6(CLBLM_L_X10Y143_SLICE_X12Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8282ffff008200ff)
  ) CLBLM_L_X10Y143_SLICE_X12Y143_CLUT (
.I0(CLBLM_L_X10Y144_SLICE_X12Y144_AO6),
.I1(CLBLM_L_X10Y143_SLICE_X12Y143_CQ),
.I2(CLBLM_L_X10Y143_SLICE_X13Y143_BO6),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X11Y144_SLICE_X14Y144_DO6),
.I5(CLBLM_L_X10Y145_SLICE_X12Y145_AQ),
.O5(CLBLM_L_X10Y143_SLICE_X12Y143_CO5),
.O6(CLBLM_L_X10Y143_SLICE_X12Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa00f0aaaaccf0)
  ) CLBLM_L_X10Y143_SLICE_X12Y143_BLUT (
.I0(CLBLL_L_X4Y137_SLICE_X4Y137_BQ),
.I1(CLBLM_L_X10Y143_SLICE_X12Y143_BQ),
.I2(CLBLM_L_X10Y145_SLICE_X13Y145_AQ),
.I3(CLBLM_L_X8Y144_SLICE_X11Y144_CO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X10Y145_SLICE_X13Y145_BO6),
.O5(CLBLM_L_X10Y143_SLICE_X12Y143_BO5),
.O6(CLBLM_L_X10Y143_SLICE_X12Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h50ff000050ff50ff)
  ) CLBLM_L_X10Y143_SLICE_X12Y143_ALUT (
.I0(CLBLM_L_X10Y143_SLICE_X12Y143_DO6),
.I1(1'b1),
.I2(CLBLM_L_X10Y144_SLICE_X12Y144_AO6),
.I3(CLBLM_R_X11Y144_SLICE_X14Y144_DO6),
.I4(CLBLM_R_X5Y134_SLICE_X6Y134_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y143_SLICE_X12Y143_AO5),
.O6(CLBLM_L_X10Y143_SLICE_X12Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y143_SLICE_X13Y143_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y77_IOB_X0Y77_I),
.D(CLBLM_L_X10Y133_SLICE_X12Y133_BQ),
.Q(CLBLM_L_X10Y143_SLICE_X13Y143_AQ),
.R(CLBLM_L_X12Y144_SLICE_X16Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y143_SLICE_X13Y143_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y77_IOB_X0Y77_I),
.D(CLBLM_R_X7Y135_SLICE_X8Y135_CQ),
.Q(CLBLM_L_X10Y143_SLICE_X13Y143_BQ),
.R(CLBLM_L_X12Y144_SLICE_X16Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h2222222222222222)
  ) CLBLM_L_X10Y143_SLICE_X13Y143_DLUT (
.I0(CLBLM_L_X10Y143_SLICE_X13Y143_AO6),
.I1(CLBLM_L_X10Y142_SLICE_X13Y142_CQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y143_SLICE_X13Y143_DO5),
.O6(CLBLM_L_X10Y143_SLICE_X13Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc39cc39cc39cc33)
  ) CLBLM_L_X10Y143_SLICE_X13Y143_CLUT (
.I0(CLBLM_L_X10Y142_SLICE_X13Y142_AQ),
.I1(CLBLM_R_X11Y142_SLICE_X15Y142_CQ),
.I2(CLBLM_L_X10Y145_SLICE_X12Y145_CO6),
.I3(CLBLM_L_X10Y144_SLICE_X13Y144_DO6),
.I4(CLBLM_L_X10Y143_SLICE_X13Y143_DO6),
.I5(CLBLM_R_X11Y143_SLICE_X14Y143_CO5),
.O5(CLBLM_L_X10Y143_SLICE_X13Y143_CO5),
.O6(CLBLM_L_X10Y143_SLICE_X13Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000ff1fffdf)
  ) CLBLM_L_X10Y143_SLICE_X13Y143_BLUT (
.I0(CLBLM_L_X10Y143_SLICE_X13Y143_DO6),
.I1(CLBLM_R_X11Y142_SLICE_X15Y142_CQ),
.I2(CLBLM_L_X10Y142_SLICE_X12Y142_BQ),
.I3(CLBLM_L_X10Y145_SLICE_X12Y145_CO6),
.I4(CLBLM_R_X11Y143_SLICE_X14Y143_CO5),
.I5(CLBLM_L_X10Y144_SLICE_X13Y144_DO6),
.O5(CLBLM_L_X10Y143_SLICE_X13Y143_BO5),
.O6(CLBLM_L_X10Y143_SLICE_X13Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000300020)
  ) CLBLM_L_X10Y143_SLICE_X13Y143_ALUT (
.I0(CLBLM_R_X11Y144_SLICE_X14Y144_AQ),
.I1(CLBLM_R_X11Y144_SLICE_X15Y144_BQ),
.I2(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.I3(CLBLM_L_X10Y144_SLICE_X13Y144_AQ),
.I4(CLBLM_L_X10Y142_SLICE_X12Y142_CQ),
.I5(CLBLM_L_X10Y143_SLICE_X12Y143_AQ),
.O5(CLBLM_L_X10Y143_SLICE_X13Y143_AO5),
.O6(CLBLM_L_X10Y143_SLICE_X13Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y144_SLICE_X12Y144_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y144_SLICE_X14Y144_BO6),
.Q(CLBLM_L_X10Y144_SLICE_X12Y144_AQ),
.R(CLBLM_R_X7Y144_SLICE_X9Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y144_SLICE_X12Y144_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y144_SLICE_X12Y144_DO5),
.O6(CLBLM_L_X10Y144_SLICE_X12Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha5a52d78a5f02d78)
  ) CLBLM_L_X10Y144_SLICE_X12Y144_CLUT (
.I0(CLBLM_L_X8Y142_SLICE_X11Y142_DQ),
.I1(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.I2(CLBLM_L_X8Y135_SLICE_X10Y135_CO6),
.I3(CLBLM_L_X8Y142_SLICE_X10Y142_D5Q),
.I4(CLBLM_R_X11Y144_SLICE_X14Y144_AQ),
.I5(CLBLM_L_X10Y142_SLICE_X12Y142_CQ),
.O5(CLBLM_L_X10Y144_SLICE_X12Y144_CO5),
.O6(CLBLM_L_X10Y144_SLICE_X12Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ffff2300ffff)
  ) CLBLM_L_X10Y144_SLICE_X12Y144_BLUT (
.I0(CLBLM_L_X10Y145_SLICE_X12Y145_BO5),
.I1(CLBLM_L_X10Y144_SLICE_X12Y144_CO6),
.I2(CLBLM_L_X10Y141_SLICE_X12Y141_C5Q),
.I3(CLBLM_R_X7Y142_SLICE_X9Y142_AQ),
.I4(CLBLM_R_X11Y143_SLICE_X14Y143_AQ),
.I5(CLBLM_L_X10Y144_SLICE_X12Y144_AO5),
.O5(CLBLM_L_X10Y144_SLICE_X12Y144_BO5),
.O6(CLBLM_L_X10Y144_SLICE_X12Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0e0000aabb)
  ) CLBLM_L_X10Y144_SLICE_X12Y144_ALUT (
.I0(CLBLM_L_X8Y142_SLICE_X10Y142_D5Q),
.I1(CLBLM_L_X10Y142_SLICE_X12Y142_CQ),
.I2(CLBLM_R_X11Y143_SLICE_X14Y143_DO6),
.I3(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.I4(CLBLM_R_X11Y144_SLICE_X14Y144_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y144_SLICE_X12Y144_AO5),
.O6(CLBLM_L_X10Y144_SLICE_X12Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y144_SLICE_X13Y144_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y144_SLICE_X13Y144_AO6),
.Q(CLBLM_L_X10Y144_SLICE_X13Y144_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0fffff0e0fffff)
  ) CLBLM_L_X10Y144_SLICE_X13Y144_DLUT (
.I0(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.I1(CLBLM_L_X8Y142_SLICE_X10Y142_D5Q),
.I2(CLBLM_L_X10Y141_SLICE_X12Y141_C5Q),
.I3(CLBLM_R_X11Y144_SLICE_X14Y144_AQ),
.I4(CLBLM_L_X8Y144_SLICE_X11Y144_BO5),
.I5(CLBLM_L_X10Y142_SLICE_X12Y142_CQ),
.O5(CLBLM_L_X10Y144_SLICE_X13Y144_DO5),
.O6(CLBLM_L_X10Y144_SLICE_X13Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0808101008881000)
  ) CLBLM_L_X10Y144_SLICE_X13Y144_CLUT (
.I0(CLBLM_R_X11Y144_SLICE_X15Y144_BQ),
.I1(CLBLM_L_X10Y143_SLICE_X12Y143_AQ),
.I2(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.I3(CLBLM_R_X11Y144_SLICE_X14Y144_AQ),
.I4(CLBLM_L_X10Y144_SLICE_X13Y144_AQ),
.I5(CLBLM_L_X10Y142_SLICE_X12Y142_CQ),
.O5(CLBLM_L_X10Y144_SLICE_X13Y144_CO5),
.O6(CLBLM_L_X10Y144_SLICE_X13Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5515555555555545)
  ) CLBLM_L_X10Y144_SLICE_X13Y144_BLUT (
.I0(CLBLM_L_X10Y144_SLICE_X13Y144_DO6),
.I1(CLBLM_L_X10Y143_SLICE_X12Y143_AQ),
.I2(CLBLM_L_X10Y142_SLICE_X12Y142_AQ),
.I3(CLBLM_L_X10Y145_SLICE_X12Y145_CO6),
.I4(CLBLM_R_X11Y144_SLICE_X15Y144_BQ),
.I5(CLBLM_L_X10Y145_SLICE_X12Y145_BO6),
.O5(CLBLM_L_X10Y144_SLICE_X13Y144_BO5),
.O6(CLBLM_L_X10Y144_SLICE_X13Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0502010ffff3333)
  ) CLBLM_L_X10Y144_SLICE_X13Y144_ALUT (
.I0(CLBLM_L_X10Y144_SLICE_X13Y144_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y144_SLICE_X12Y144_AO6),
.I3(CLBLM_L_X10Y144_SLICE_X13Y144_BO6),
.I4(CLBLM_L_X8Y144_SLICE_X11Y144_AQ),
.I5(CLBLM_R_X11Y144_SLICE_X14Y144_DO6),
.O5(CLBLM_L_X10Y144_SLICE_X13Y144_AO5),
.O6(CLBLM_L_X10Y144_SLICE_X13Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y145_SLICE_X12Y145_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y145_SLICE_X12Y145_AO6),
.Q(CLBLM_L_X10Y145_SLICE_X12Y145_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y145_SLICE_X12Y145_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y145_SLICE_X12Y145_DO5),
.O6(CLBLM_L_X10Y145_SLICE_X12Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0055ffff005fffff)
  ) CLBLM_L_X10Y145_SLICE_X12Y145_CLUT (
.I0(CLBLM_L_X8Y142_SLICE_X11Y142_DQ),
.I1(1'b1),
.I2(CLBLM_L_X10Y142_SLICE_X12Y142_CQ),
.I3(CLBLM_L_X10Y145_SLICE_X12Y145_AO5),
.I4(CLBLM_L_X8Y144_SLICE_X11Y144_BO5),
.I5(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.O5(CLBLM_L_X10Y145_SLICE_X12Y145_CO5),
.O6(CLBLM_L_X10Y145_SLICE_X12Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0303ffffffffffcc)
  ) CLBLM_L_X10Y145_SLICE_X12Y145_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y142_SLICE_X12Y142_CQ),
.I2(CLBLM_R_X11Y144_SLICE_X14Y144_AQ),
.I3(CLBLM_L_X8Y142_SLICE_X10Y142_D5Q),
.I4(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y145_SLICE_X12Y145_BO5),
.O6(CLBLM_L_X10Y145_SLICE_X12Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafa505033000000)
  ) CLBLM_L_X10Y145_SLICE_X12Y145_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y141_SLICE_X12Y141_C5Q),
.I2(CLBLM_L_X12Y143_SLICE_X16Y143_BQ),
.I3(CLBLM_L_X8Y142_SLICE_X10Y142_D5Q),
.I4(CLBLM_R_X11Y144_SLICE_X14Y144_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y145_SLICE_X12Y145_AO5),
.O6(CLBLM_L_X10Y145_SLICE_X12Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y145_SLICE_X13Y145_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y145_SLICE_X13Y145_AO6),
.Q(CLBLM_L_X10Y145_SLICE_X13Y145_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y145_SLICE_X13Y145_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y145_SLICE_X13Y145_DO5),
.O6(CLBLM_L_X10Y145_SLICE_X13Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000bf00bc)
  ) CLBLM_L_X10Y145_SLICE_X13Y145_CLUT (
.I0(CLBLM_L_X8Y144_SLICE_X11Y144_CO6),
.I1(CLBLM_L_X10Y141_SLICE_X12Y141_C5Q),
.I2(CLBLM_R_X11Y142_SLICE_X15Y142_AQ),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(CLBLM_L_X10Y145_SLICE_X13Y145_BO5),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y145_SLICE_X13Y145_CO5),
.O6(CLBLM_L_X10Y145_SLICE_X13Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000300000020)
  ) CLBLM_L_X10Y145_SLICE_X13Y145_BLUT (
.I0(CLBLM_L_X8Y144_SLICE_X11Y144_BO5),
.I1(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.I2(CLBLM_R_X11Y144_SLICE_X14Y144_AQ),
.I3(CLBLM_L_X8Y142_SLICE_X10Y142_D5Q),
.I4(CLBLM_L_X10Y142_SLICE_X12Y142_CQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y145_SLICE_X13Y145_BO5),
.O6(CLBLM_L_X10Y145_SLICE_X13Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffff320000ff32)
  ) CLBLM_L_X10Y145_SLICE_X13Y145_ALUT (
.I0(CLBLM_R_X11Y142_SLICE_X15Y142_AQ),
.I1(CLBLM_L_X8Y144_SLICE_X11Y144_CO6),
.I2(CLBLM_L_X10Y145_SLICE_X13Y145_AQ),
.I3(CLBLM_L_X10Y145_SLICE_X13Y145_BO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y144_SLICE_X8Y144_CQ),
.O5(CLBLM_L_X10Y145_SLICE_X13Y145_AO5),
.O6(CLBLM_L_X10Y145_SLICE_X13Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y146_SLICE_X12Y146_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y146_SLICE_X12Y146_DO5),
.O6(CLBLM_L_X10Y146_SLICE_X12Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y146_SLICE_X12Y146_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y146_SLICE_X12Y146_CO5),
.O6(CLBLM_L_X10Y146_SLICE_X12Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y146_SLICE_X12Y146_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y146_SLICE_X12Y146_BO5),
.O6(CLBLM_L_X10Y146_SLICE_X12Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc30fc30ff00ffff)
  ) CLBLM_L_X10Y146_SLICE_X12Y146_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X5Y136_SLICE_X7Y136_DO5),
.I3(CLBLM_L_X10Y143_SLICE_X13Y143_BQ),
.I4(RIOB33_X105Y143_IOB_X1Y143_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y146_SLICE_X12Y146_AO5),
.O6(CLBLM_L_X10Y146_SLICE_X12Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y146_SLICE_X13Y146_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y146_SLICE_X13Y146_DO5),
.O6(CLBLM_L_X10Y146_SLICE_X13Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y146_SLICE_X13Y146_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y146_SLICE_X13Y146_CO5),
.O6(CLBLM_L_X10Y146_SLICE_X13Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y146_SLICE_X13Y146_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y146_SLICE_X13Y146_BO5),
.O6(CLBLM_L_X10Y146_SLICE_X13Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y146_SLICE_X13Y146_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y146_SLICE_X13Y146_AO5),
.O6(CLBLM_L_X10Y146_SLICE_X13Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y132_SLICE_X16Y132_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y132_SLICE_X16Y132_AO6),
.Q(CLBLM_L_X12Y132_SLICE_X16Y132_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y132_SLICE_X16Y132_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y132_SLICE_X16Y132_BO6),
.Q(CLBLM_L_X12Y132_SLICE_X16Y132_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y132_SLICE_X16Y132_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y132_SLICE_X16Y132_CO6),
.Q(CLBLM_L_X12Y132_SLICE_X16Y132_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00003333)
  ) CLBLM_L_X12Y132_SLICE_X16Y132_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X12Y136_SLICE_X16Y136_CQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X11Y132_SLICE_X15Y132_AO5),
.I5(CLBLM_R_X5Y134_SLICE_X7Y134_DO6),
.O5(CLBLM_L_X12Y132_SLICE_X16Y132_DO5),
.O6(CLBLM_L_X12Y132_SLICE_X16Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff550055ff050005)
  ) CLBLM_L_X12Y132_SLICE_X16Y132_CLUT (
.I0(CLBLM_R_X11Y132_SLICE_X15Y132_BO6),
.I1(1'b1),
.I2(RIOB33_X105Y141_IOB_X1Y142_I),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X12Y136_SLICE_X17Y136_DQ),
.I5(CLBLM_R_X7Y131_SLICE_X9Y131_AQ),
.O5(CLBLM_L_X12Y132_SLICE_X16Y132_CO5),
.O6(CLBLM_L_X12Y132_SLICE_X16Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haafe0054aafe0054)
  ) CLBLM_L_X12Y132_SLICE_X16Y132_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X12Y132_SLICE_X16Y132_BQ),
.I2(CLBLM_R_X11Y133_SLICE_X14Y133_AQ),
.I3(CLBLM_R_X5Y134_SLICE_X7Y134_DO6),
.I4(CLBLM_R_X11Y138_SLICE_X14Y138_CQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y132_SLICE_X16Y132_BO5),
.O6(CLBLM_L_X12Y132_SLICE_X16Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heeececeeaaa0a0aa)
  ) CLBLM_L_X12Y132_SLICE_X16Y132_ALUT (
.I0(CLBLM_L_X12Y144_SLICE_X16Y144_AO6),
.I1(CLBLM_L_X12Y136_SLICE_X16Y136_CQ),
.I2(CLBLM_L_X12Y132_SLICE_X16Y132_AQ),
.I3(CLBLM_L_X12Y132_SLICE_X16Y132_DO6),
.I4(CLBLM_L_X10Y132_SLICE_X13Y132_AO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X12Y132_SLICE_X16Y132_AO5),
.O6(CLBLM_L_X12Y132_SLICE_X16Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y132_SLICE_X17Y132_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y132_SLICE_X17Y132_AO6),
.Q(CLBLM_L_X12Y132_SLICE_X17Y132_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y132_SLICE_X17Y132_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y132_SLICE_X17Y132_DO5),
.O6(CLBLM_L_X12Y132_SLICE_X17Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y132_SLICE_X17Y132_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y132_SLICE_X17Y132_CO5),
.O6(CLBLM_L_X12Y132_SLICE_X17Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfcfdfdf0f0f0f0)
  ) CLBLM_L_X12Y132_SLICE_X17Y132_BLUT (
.I0(CLBLM_L_X12Y136_SLICE_X16Y136_CQ),
.I1(CLBLM_R_X5Y132_SLICE_X7Y132_DO6),
.I2(CLBLM_L_X12Y132_SLICE_X17Y132_AQ),
.I3(1'b1),
.I4(CLBLM_R_X11Y132_SLICE_X15Y132_AO5),
.I5(CLBLM_L_X12Y133_SLICE_X16Y133_DO5),
.O5(CLBLM_L_X12Y132_SLICE_X17Y132_BO5),
.O6(CLBLM_L_X12Y132_SLICE_X17Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heeccaa00eeceaa0a)
  ) CLBLM_L_X12Y132_SLICE_X17Y132_ALUT (
.I0(CLBLM_L_X12Y144_SLICE_X16Y144_AO6),
.I1(CLBLM_L_X12Y141_SLICE_X17Y141_AQ),
.I2(CLBLM_L_X10Y132_SLICE_X13Y132_AO6),
.I3(CLBLM_L_X12Y132_SLICE_X17Y132_BO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X12Y133_SLICE_X16Y133_DO5),
.O5(CLBLM_L_X12Y132_SLICE_X17Y132_AO5),
.O6(CLBLM_L_X12Y132_SLICE_X17Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y133_SLICE_X16Y133_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y133_SLICE_X16Y133_CO5),
.Q(CLBLM_L_X12Y133_SLICE_X16Y133_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y133_SLICE_X16Y133_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y133_SLICE_X16Y133_AO6),
.Q(CLBLM_L_X12Y133_SLICE_X16Y133_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y133_SLICE_X16Y133_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y133_SLICE_X16Y133_BO6),
.Q(CLBLM_L_X12Y133_SLICE_X16Y133_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y133_SLICE_X16Y133_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y133_SLICE_X16Y133_CO6),
.Q(CLBLM_L_X12Y133_SLICE_X16Y133_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h99959995000f000f)
  ) CLBLM_L_X12Y133_SLICE_X16Y133_DLUT (
.I0(CLBLM_R_X7Y132_SLICE_X9Y132_BQ),
.I1(CLBLM_L_X12Y137_SLICE_X16Y137_AQ),
.I2(CLBLM_R_X13Y138_SLICE_X18Y138_BO6),
.I3(CLBLL_L_X4Y142_SLICE_X4Y142_BO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y133_SLICE_X16Y133_DO5),
.O6(CLBLM_L_X12Y133_SLICE_X16Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcfc0c0afa0afa0)
  ) CLBLM_L_X12Y133_SLICE_X16Y133_CLUT (
.I0(CLBLM_R_X11Y131_SLICE_X14Y131_BQ),
.I1(CLBLM_L_X12Y133_SLICE_X16Y133_AQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X11Y136_SLICE_X15Y136_B5Q),
.I4(RIOB33_X105Y103_IOB_X1Y104_I),
.I5(1'b1),
.O5(CLBLM_L_X12Y133_SLICE_X16Y133_CO5),
.O6(CLBLM_L_X12Y133_SLICE_X16Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcaff0a00ca000a)
  ) CLBLM_L_X12Y133_SLICE_X16Y133_BLUT (
.I0(CLBLM_R_X13Y133_SLICE_X18Y133_AQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_L_X10Y135_SLICE_X12Y135_DO6),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X12Y133_SLICE_X16Y133_BQ),
.I5(CLBLM_L_X8Y133_SLICE_X11Y133_CQ),
.O5(CLBLM_L_X12Y133_SLICE_X16Y133_BO5),
.O6(CLBLM_L_X12Y133_SLICE_X16Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffb3800000b380)
  ) CLBLM_L_X12Y133_SLICE_X16Y133_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X10Y135_SLICE_X12Y135_DO6),
.I2(CLBLM_L_X12Y133_SLICE_X16Y133_AQ),
.I3(CLBLM_L_X12Y133_SLICE_X17Y133_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X11Y140_SLICE_X14Y140_BQ),
.O5(CLBLM_L_X12Y133_SLICE_X16Y133_AO5),
.O6(CLBLM_L_X12Y133_SLICE_X16Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y133_SLICE_X17Y133_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y133_SLICE_X17Y133_AO6),
.Q(CLBLM_L_X12Y133_SLICE_X17Y133_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y133_SLICE_X17Y133_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y133_SLICE_X17Y133_BO6),
.Q(CLBLM_L_X12Y133_SLICE_X17Y133_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y133_SLICE_X17Y133_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y133_SLICE_X17Y133_DO5),
.O6(CLBLM_L_X12Y133_SLICE_X17Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y133_SLICE_X17Y133_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y133_SLICE_X17Y133_CO5),
.O6(CLBLM_L_X12Y133_SLICE_X17Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc0cfa0af000fa0a)
  ) CLBLM_L_X12Y133_SLICE_X17Y133_BLUT (
.I0(CLBLM_R_X11Y134_SLICE_X14Y134_AQ),
.I1(CLBLM_L_X12Y133_SLICE_X17Y133_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X13Y134_SLICE_X19Y134_DQ),
.I4(CLBLM_L_X10Y135_SLICE_X12Y135_DO6),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X12Y133_SLICE_X17Y133_BO5),
.O6(CLBLM_L_X12Y133_SLICE_X17Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hd888ddddd8888888)
  ) CLBLM_L_X12Y133_SLICE_X17Y133_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X13Y137_SLICE_X18Y137_AQ),
.I2(CLBLM_L_X12Y133_SLICE_X17Y133_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_L_X10Y135_SLICE_X12Y135_DO6),
.I5(CLBLM_R_X13Y135_SLICE_X18Y135_BQ),
.O5(CLBLM_L_X12Y133_SLICE_X17Y133_AO5),
.O6(CLBLM_L_X12Y133_SLICE_X17Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y134_SLICE_X16Y134_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y77_IOB_X0Y77_I),
.D(CLBLM_L_X12Y133_SLICE_X16Y133_CQ),
.Q(CLBLM_L_X12Y134_SLICE_X16Y134_AQ),
.R(CLBLM_L_X12Y144_SLICE_X16Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5aff5affff5aff5a)
  ) CLBLM_L_X12Y134_SLICE_X16Y134_DLUT (
.I0(CLBLM_R_X13Y133_SLICE_X18Y133_AQ),
.I1(1'b1),
.I2(CLBLM_R_X13Y134_SLICE_X19Y134_CQ),
.I3(CLBLM_R_X13Y134_SLICE_X19Y134_AQ),
.I4(1'b1),
.I5(CLBLM_R_X11Y135_SLICE_X14Y135_BQ),
.O5(CLBLM_L_X12Y134_SLICE_X16Y134_DO5),
.O6(CLBLM_L_X12Y134_SLICE_X16Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5aa55aa5a55aa55a)
  ) CLBLM_L_X12Y134_SLICE_X16Y134_CLUT (
.I0(CLBLM_R_X7Y132_SLICE_X9Y132_BQ),
.I1(1'b1),
.I2(CLBLM_R_X13Y134_SLICE_X19Y134_CQ),
.I3(CLBLM_R_X11Y134_SLICE_X15Y134_BQ),
.I4(1'b1),
.I5(CLBLM_R_X11Y135_SLICE_X14Y135_BQ),
.O5(CLBLM_L_X12Y134_SLICE_X16Y134_CO5),
.O6(CLBLM_L_X12Y134_SLICE_X16Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hbfefbfeffbfefbfe)
  ) CLBLM_L_X12Y134_SLICE_X16Y134_BLUT (
.I0(CLBLM_L_X12Y134_SLICE_X16Y134_DO6),
.I1(CLBLM_R_X11Y134_SLICE_X14Y134_CQ),
.I2(CLBLM_L_X12Y135_SLICE_X16Y135_AQ),
.I3(CLBLM_R_X13Y134_SLICE_X19Y134_DQ),
.I4(1'b1),
.I5(CLBLM_L_X12Y135_SLICE_X16Y135_CQ),
.O5(CLBLM_L_X12Y134_SLICE_X16Y134_BO5),
.O6(CLBLM_L_X12Y134_SLICE_X16Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h4141141414144141)
  ) CLBLM_L_X12Y134_SLICE_X16Y134_ALUT (
.I0(CLBLM_L_X12Y135_SLICE_X17Y135_CQ),
.I1(CLBLM_R_X11Y134_SLICE_X15Y134_DO6),
.I2(CLBLM_L_X12Y135_SLICE_X16Y135_AQ),
.I3(1'b1),
.I4(CLBLM_R_X13Y134_SLICE_X19Y134_DQ),
.I5(CLBLM_L_X12Y134_SLICE_X16Y134_CO6),
.O5(CLBLM_L_X12Y134_SLICE_X16Y134_AO5),
.O6(CLBLM_L_X12Y134_SLICE_X16Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y134_SLICE_X17Y134_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y134_SLICE_X18Y134_AO6),
.Q(CLBLM_L_X12Y134_SLICE_X17Y134_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h33ffccffff33ffcc)
  ) CLBLM_L_X12Y134_SLICE_X17Y134_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X12Y139_SLICE_X17Y139_CQ),
.I2(1'b1),
.I3(CLBLM_R_X11Y134_SLICE_X15Y134_BQ),
.I4(CLBLM_R_X7Y133_SLICE_X9Y133_AQ),
.I5(CLBLM_L_X12Y135_SLICE_X16Y135_BQ),
.O5(CLBLM_L_X12Y134_SLICE_X17Y134_DO5),
.O6(CLBLM_L_X12Y134_SLICE_X17Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffff3c3c)
  ) CLBLM_L_X12Y134_SLICE_X17Y134_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y134_SLICE_X14Y134_BQ),
.I2(CLBLM_L_X8Y134_SLICE_X11Y134_AQ),
.I3(1'b1),
.I4(CLBLM_L_X12Y135_SLICE_X17Y135_DO6),
.I5(CLBLM_L_X12Y134_SLICE_X17Y134_DO6),
.O5(CLBLM_L_X12Y134_SLICE_X17Y134_CO5),
.O6(CLBLM_L_X12Y134_SLICE_X17Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000001)
  ) CLBLM_L_X12Y134_SLICE_X17Y134_BLUT (
.I0(CLBLM_R_X13Y134_SLICE_X19Y134_AQ),
.I1(CLBLM_R_X11Y134_SLICE_X14Y134_CQ),
.I2(CLBLM_L_X12Y133_SLICE_X16Y133_AQ),
.I3(CLBLM_L_X12Y135_SLICE_X16Y135_BQ),
.I4(CLBLM_R_X13Y135_SLICE_X18Y135_AQ),
.I5(CLBLM_L_X12Y133_SLICE_X17Y133_BQ),
.O5(CLBLM_L_X12Y134_SLICE_X17Y134_BO5),
.O6(CLBLM_L_X12Y134_SLICE_X17Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000d000e000)
  ) CLBLM_L_X12Y134_SLICE_X17Y134_ALUT (
.I0(CLBLM_R_X13Y134_SLICE_X18Y134_DO6),
.I1(CLBLM_L_X12Y134_SLICE_X16Y134_BO6),
.I2(CLBLM_L_X12Y138_SLICE_X17Y138_BO5),
.I3(CLBLM_L_X10Y135_SLICE_X12Y135_DO6),
.I4(CLBLM_L_X12Y133_SLICE_X16Y133_DO6),
.I5(CLBLM_L_X12Y134_SLICE_X17Y134_CO6),
.O5(CLBLM_L_X12Y134_SLICE_X17Y134_AO5),
.O6(CLBLM_L_X12Y134_SLICE_X17Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y135_SLICE_X16Y135_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y135_SLICE_X16Y135_AO6),
.Q(CLBLM_L_X12Y135_SLICE_X16Y135_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y135_SLICE_X16Y135_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y135_SLICE_X16Y135_BO6),
.Q(CLBLM_L_X12Y135_SLICE_X16Y135_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y135_SLICE_X16Y135_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y135_SLICE_X16Y135_CO6),
.Q(CLBLM_L_X12Y135_SLICE_X16Y135_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y135_SLICE_X16Y135_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y135_SLICE_X16Y135_DO6),
.Q(CLBLM_L_X12Y135_SLICE_X16Y135_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc55005500)
  ) CLBLM_L_X12Y135_SLICE_X16Y135_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X12Y135_SLICE_X16Y135_AQ),
.I2(1'b1),
.I3(CLBLM_L_X8Y135_SLICE_X11Y135_A5Q),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X12Y135_SLICE_X16Y135_DO5),
.O6(CLBLM_L_X12Y135_SLICE_X16Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0dd885500)
  ) CLBLM_L_X12Y135_SLICE_X16Y135_CLUT (
.I0(CLBLM_L_X10Y135_SLICE_X12Y135_DO6),
.I1(CLBLM_L_X12Y135_SLICE_X16Y135_CQ),
.I2(CLBLM_R_X11Y140_SLICE_X15Y140_CQ),
.I3(CLBLM_L_X12Y139_SLICE_X17Y139_CQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X12Y135_SLICE_X16Y135_CO5),
.O6(CLBLM_L_X12Y135_SLICE_X16Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffc0ffaa00c000aa)
  ) CLBLM_L_X12Y135_SLICE_X16Y135_BLUT (
.I0(CLBLM_R_X13Y136_SLICE_X18Y136_AQ),
.I1(CLBLM_L_X12Y135_SLICE_X16Y135_BQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y135_SLICE_X12Y135_DO6),
.I5(CLBLM_L_X8Y136_SLICE_X10Y136_AQ),
.O5(CLBLM_L_X12Y135_SLICE_X16Y135_BO5),
.O6(CLBLM_L_X12Y135_SLICE_X16Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffeccdc33320010)
  ) CLBLM_L_X12Y135_SLICE_X16Y135_ALUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X12Y135_SLICE_X16Y135_AQ),
.I3(CLBLM_L_X8Y138_SLICE_X10Y138_AQ),
.I4(CLBLL_L_X4Y135_SLICE_X5Y135_AQ),
.I5(CLBLM_L_X12Y142_SLICE_X16Y142_CQ),
.O5(CLBLM_L_X12Y135_SLICE_X16Y135_AO5),
.O6(CLBLM_L_X12Y135_SLICE_X16Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y135_SLICE_X17Y135_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y135_SLICE_X17Y135_BO6),
.Q(CLBLM_L_X12Y135_SLICE_X17Y135_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y135_SLICE_X17Y135_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y135_SLICE_X17Y135_AO6),
.Q(CLBLM_L_X12Y135_SLICE_X17Y135_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y135_SLICE_X17Y135_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y135_SLICE_X17Y135_CO6),
.Q(CLBLM_L_X12Y135_SLICE_X17Y135_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5f5ff5f5afaffafa)
  ) CLBLM_L_X12Y135_SLICE_X17Y135_DLUT (
.I0(CLBLM_L_X12Y133_SLICE_X16Y133_BQ),
.I1(1'b1),
.I2(CLBLM_R_X13Y136_SLICE_X18Y136_AQ),
.I3(1'b1),
.I4(CLBLM_L_X8Y132_SLICE_X11Y132_BQ),
.I5(CLBLM_R_X11Y139_SLICE_X14Y139_AQ),
.O5(CLBLM_L_X12Y135_SLICE_X17Y135_DO5),
.O6(CLBLM_L_X12Y135_SLICE_X17Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ddddff00d0d0)
  ) CLBLM_L_X12Y135_SLICE_X17Y135_CLUT (
.I0(CLBLM_L_X12Y134_SLICE_X16Y134_AO6),
.I1(CLBLM_L_X12Y133_SLICE_X16Y133_DO5),
.I2(RIOB33_X105Y117_IOB_X1Y118_I),
.I3(CLBLM_L_X12Y137_SLICE_X17Y137_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y138_SLICE_X10Y138_AQ),
.O5(CLBLM_L_X12Y135_SLICE_X17Y135_CO5),
.O6(CLBLM_L_X12Y135_SLICE_X17Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f04400ee00ee)
  ) CLBLM_L_X12Y135_SLICE_X17Y135_BLUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_L_X8Y138_SLICE_X10Y138_AQ),
.I2(CLBLM_L_X12Y135_SLICE_X17Y135_CQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X11Y135_SLICE_X15Y135_CO6),
.I5(1'b1),
.O5(CLBLM_L_X12Y135_SLICE_X17Y135_BO5),
.O6(CLBLM_L_X12Y135_SLICE_X17Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc30fc30dc10dc10)
  ) CLBLM_L_X12Y135_SLICE_X17Y135_ALUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X12Y135_SLICE_X17Y135_AQ),
.I3(CLBLM_L_X12Y135_SLICE_X16Y135_BQ),
.I4(1'b1),
.I5(CLBLM_L_X8Y138_SLICE_X10Y138_AQ),
.O5(CLBLM_L_X12Y135_SLICE_X17Y135_AO5),
.O6(CLBLM_L_X12Y135_SLICE_X17Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y136_SLICE_X16Y136_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y136_SLICE_X16Y136_BO5),
.Q(CLBLM_L_X12Y136_SLICE_X16Y136_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y136_SLICE_X16Y136_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y136_SLICE_X16Y136_CO5),
.Q(CLBLM_L_X12Y136_SLICE_X16Y136_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y136_SLICE_X16Y136_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y136_SLICE_X16Y136_AO6),
.Q(CLBLM_L_X12Y136_SLICE_X16Y136_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y136_SLICE_X16Y136_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y136_SLICE_X16Y136_BO6),
.Q(CLBLM_L_X12Y136_SLICE_X16Y136_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y136_SLICE_X16Y136_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y136_SLICE_X16Y136_CO6),
.Q(CLBLM_L_X12Y136_SLICE_X16Y136_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y136_SLICE_X16Y136_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y136_SLICE_X16Y136_DO6),
.Q(CLBLM_L_X12Y136_SLICE_X16Y136_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hdddcdddc11101110)
  ) CLBLM_L_X12Y136_SLICE_X16Y136_DLUT (
.I0(CLBLM_R_X5Y132_SLICE_X7Y132_DO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X12Y136_SLICE_X16Y136_DQ),
.I3(CLBLM_L_X12Y132_SLICE_X16Y132_BQ),
.I4(1'b1),
.I5(CLBLM_L_X12Y138_SLICE_X17Y138_BQ),
.O5(CLBLM_L_X12Y136_SLICE_X16Y136_DO5),
.O6(CLBLM_L_X12Y136_SLICE_X16Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0ccf0ccaaffaa00)
  ) CLBLM_L_X12Y136_SLICE_X16Y136_CLUT (
.I0(CLBLM_L_X12Y132_SLICE_X16Y132_AQ),
.I1(CLBLM_L_X12Y138_SLICE_X17Y138_A5Q),
.I2(CLBLM_L_X10Y130_SLICE_X12Y130_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X13Y140_SLICE_X18Y140_CQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y136_SLICE_X16Y136_CO5),
.O6(CLBLM_L_X12Y136_SLICE_X16Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcfc0c0afa0afa0)
  ) CLBLM_L_X12Y136_SLICE_X16Y136_BLUT (
.I0(CLBLM_R_X7Y136_SLICE_X8Y136_CQ),
.I1(CLBLM_L_X12Y132_SLICE_X16Y132_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X12Y138_SLICE_X17Y138_BQ),
.I4(RIOB33_X105Y103_IOB_X1Y104_I),
.I5(1'b1),
.O5(CLBLM_L_X12Y136_SLICE_X16Y136_BO5),
.O6(CLBLM_L_X12Y136_SLICE_X16Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf044f044f044f044)
  ) CLBLM_L_X12Y136_SLICE_X16Y136_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X7Y139_SLICE_X8Y139_BQ),
.I2(CLBLM_R_X13Y135_SLICE_X18Y135_BQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y136_SLICE_X16Y136_AO5),
.O6(CLBLM_L_X12Y136_SLICE_X16Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y136_SLICE_X17Y136_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y136_SLICE_X17Y136_BO6),
.Q(CLBLM_L_X12Y136_SLICE_X17Y136_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y136_SLICE_X17Y136_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y136_SLICE_X17Y136_AO6),
.Q(CLBLM_L_X12Y136_SLICE_X17Y136_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y136_SLICE_X17Y136_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y136_SLICE_X17Y136_CO6),
.Q(CLBLM_L_X12Y136_SLICE_X17Y136_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y136_SLICE_X17Y136_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y136_SLICE_X17Y136_DO6),
.Q(CLBLM_L_X12Y136_SLICE_X17Y136_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffccccfffff0a0)
  ) CLBLM_L_X12Y136_SLICE_X17Y136_DLUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_R_X11Y136_SLICE_X15Y136_B5Q),
.I2(CLBLM_L_X12Y136_SLICE_X17Y136_DQ),
.I3(CLBLM_L_X8Y138_SLICE_X10Y138_AQ),
.I4(CLBLM_R_X11Y136_SLICE_X15Y136_CO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X12Y136_SLICE_X17Y136_DO5),
.O6(CLBLM_L_X12Y136_SLICE_X17Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffeeeaffff4440)
  ) CLBLM_L_X12Y136_SLICE_X17Y136_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X12Y136_SLICE_X17Y136_CQ),
.I2(RIOB33_X105Y117_IOB_X1Y118_I),
.I3(CLBLM_L_X8Y138_SLICE_X10Y138_AQ),
.I4(CLBLM_R_X11Y136_SLICE_X15Y136_CO6),
.I5(CLBLM_R_X13Y143_SLICE_X18Y143_BQ),
.O5(CLBLM_L_X12Y136_SLICE_X17Y136_CO5),
.O6(CLBLM_L_X12Y136_SLICE_X17Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'heeec2220aaa0aaa0)
  ) CLBLM_L_X12Y136_SLICE_X17Y136_BLUT (
.I0(RIOB33_X105Y121_IOB_X1Y121_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X12Y137_SLICE_X17Y137_CQ),
.I3(CLBLM_R_X11Y136_SLICE_X15Y136_AQ),
.I4(CLBLM_R_X3Y136_SLICE_X3Y136_CQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y136_SLICE_X17Y136_BO5),
.O6(CLBLM_L_X12Y136_SLICE_X17Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaaffa000aa00a0)
  ) CLBLM_L_X12Y136_SLICE_X17Y136_ALUT (
.I0(CLBLM_L_X8Y143_SLICE_X10Y143_DO6),
.I1(1'b1),
.I2(CLBLM_L_X12Y136_SLICE_X17Y136_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X11Y138_SLICE_X14Y138_CQ),
.I5(CLBLM_R_X13Y137_SLICE_X19Y137_CQ),
.O5(CLBLM_L_X12Y136_SLICE_X17Y136_AO5),
.O6(CLBLM_L_X12Y136_SLICE_X17Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y137_SLICE_X16Y137_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y137_SLICE_X16Y137_BO6),
.Q(CLBLM_L_X12Y137_SLICE_X16Y137_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y137_SLICE_X16Y137_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y137_SLICE_X16Y137_AO6),
.Q(CLBLM_L_X12Y137_SLICE_X16Y137_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y137_SLICE_X16Y137_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y137_SLICE_X16Y137_CO6),
.Q(CLBLM_L_X12Y137_SLICE_X16Y137_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y137_SLICE_X16Y137_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y137_SLICE_X16Y137_DO6),
.Q(CLBLM_L_X12Y137_SLICE_X16Y137_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaafff0ffaaffc0)
  ) CLBLM_L_X12Y137_SLICE_X16Y137_DLUT (
.I0(CLBLL_L_X4Y136_SLICE_X4Y136_D5Q),
.I1(CLBLM_L_X8Y138_SLICE_X10Y138_AQ),
.I2(CLBLM_L_X12Y137_SLICE_X16Y137_DQ),
.I3(CLBLM_R_X11Y137_SLICE_X14Y137_DO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_L_X12Y137_SLICE_X16Y137_DO5),
.O6(CLBLM_L_X12Y137_SLICE_X16Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f000cc0088)
  ) CLBLM_L_X12Y137_SLICE_X16Y137_CLUT (
.I0(CLBLM_L_X12Y132_SLICE_X16Y132_AQ),
.I1(CLBLM_L_X8Y138_SLICE_X10Y138_AQ),
.I2(CLBLM_L_X12Y137_SLICE_X16Y137_DQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_L_X12Y137_SLICE_X16Y137_CQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X12Y137_SLICE_X16Y137_CO5),
.O6(CLBLM_L_X12Y137_SLICE_X16Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hef23fe320000f0f0)
  ) CLBLM_L_X12Y137_SLICE_X16Y137_BLUT (
.I0(CLBLM_R_X13Y143_SLICE_X18Y143_AO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X11Y139_SLICE_X15Y139_BQ),
.I3(CLBLM_L_X8Y135_SLICE_X10Y135_BQ),
.I4(CLBLM_L_X12Y137_SLICE_X16Y137_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X12Y137_SLICE_X16Y137_BO5),
.O6(CLBLM_L_X12Y137_SLICE_X16Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffa00faffc800c8)
  ) CLBLM_L_X12Y137_SLICE_X16Y137_ALUT (
.I0(CLBLM_L_X12Y137_SLICE_X16Y137_CQ),
.I1(CLBLM_L_X8Y138_SLICE_X10Y138_AQ),
.I2(CLBLM_L_X12Y137_SLICE_X16Y137_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X11Y139_SLICE_X14Y139_B5Q),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_L_X12Y137_SLICE_X16Y137_AO5),
.O6(CLBLM_L_X12Y137_SLICE_X16Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y137_SLICE_X17Y137_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y137_SLICE_X17Y137_BO6),
.Q(CLBLM_L_X12Y137_SLICE_X17Y137_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y137_SLICE_X17Y137_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y137_SLICE_X17Y137_AO6),
.Q(CLBLM_L_X12Y137_SLICE_X17Y137_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y137_SLICE_X17Y137_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y137_SLICE_X17Y137_CO6),
.Q(CLBLM_L_X12Y137_SLICE_X17Y137_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc33cc33cc3ccc3c)
  ) CLBLM_L_X12Y137_SLICE_X17Y137_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X13Y136_SLICE_X18Y136_CQ),
.I2(CLBLM_R_X13Y137_SLICE_X18Y137_AQ),
.I3(CLBLM_L_X12Y139_SLICE_X16Y139_CQ),
.I4(1'b1),
.I5(CLBLM_L_X10Y136_SLICE_X13Y136_AO6),
.O5(CLBLM_L_X12Y137_SLICE_X17Y137_DO5),
.O6(CLBLM_L_X12Y137_SLICE_X17Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0ffccaa88)
  ) CLBLM_L_X12Y137_SLICE_X17Y137_CLUT (
.I0(CLBLM_L_X8Y138_SLICE_X10Y138_AQ),
.I1(CLBLM_L_X12Y137_SLICE_X17Y137_CQ),
.I2(CLBLM_R_X11Y139_SLICE_X15Y139_CQ),
.I3(CLBLM_L_X8Y137_SLICE_X11Y137_CO6),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X12Y137_SLICE_X17Y137_CO5),
.O6(CLBLM_L_X12Y137_SLICE_X17Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'he2e2e2c0555555ff)
  ) CLBLM_L_X12Y137_SLICE_X17Y137_BLUT (
.I0(RIOB33_X105Y121_IOB_X1Y121_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X12Y135_SLICE_X16Y135_CQ),
.I3(CLBLM_R_X5Y137_SLICE_X7Y137_CQ),
.I4(CLBLM_R_X13Y137_SLICE_X19Y137_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y137_SLICE_X17Y137_BO5),
.O6(CLBLM_L_X12Y137_SLICE_X17Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00ccaacca0)
  ) CLBLM_L_X12Y137_SLICE_X17Y137_ALUT (
.I0(CLBLM_L_X8Y138_SLICE_X10Y138_AQ),
.I1(CLBLM_R_X11Y136_SLICE_X15Y136_AQ),
.I2(CLBLM_L_X12Y137_SLICE_X17Y137_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y136_SLICE_X8Y136_DO6),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_L_X12Y137_SLICE_X17Y137_AO5),
.O6(CLBLM_L_X12Y137_SLICE_X17Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y138_SLICE_X16Y138_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y138_SLICE_X16Y138_AO6),
.Q(CLBLM_L_X12Y138_SLICE_X16Y138_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y138_SLICE_X16Y138_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y138_SLICE_X16Y138_BO6),
.Q(CLBLM_L_X12Y138_SLICE_X16Y138_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y138_SLICE_X16Y138_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y138_SLICE_X16Y138_CO6),
.Q(CLBLM_L_X12Y138_SLICE_X16Y138_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y138_SLICE_X16Y138_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y138_SLICE_X16Y138_DO6),
.Q(CLBLM_L_X12Y138_SLICE_X16Y138_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc05500550)
  ) CLBLM_L_X12Y138_SLICE_X16Y138_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X12Y137_SLICE_X17Y137_A5Q),
.I2(CLBLM_R_X11Y138_SLICE_X14Y138_CQ),
.I3(CLBLM_R_X11Y137_SLICE_X14Y137_BO5),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X12Y138_SLICE_X16Y138_DO5),
.O6(CLBLM_L_X12Y138_SLICE_X16Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf1f00100f4f00400)
  ) CLBLM_L_X12Y138_SLICE_X16Y138_CLUT (
.I0(CLBLM_L_X10Y145_SLICE_X12Y145_AQ),
.I1(CLBLM_L_X12Y138_SLICE_X17Y138_CO6),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_L_X12Y139_SLICE_X16Y139_A5Q),
.I5(CLBLM_L_X12Y138_SLICE_X16Y138_CQ),
.O5(CLBLM_L_X12Y138_SLICE_X16Y138_CO5),
.O6(CLBLM_L_X12Y138_SLICE_X16Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f0eef000f000)
  ) CLBLM_L_X12Y138_SLICE_X16Y138_BLUT (
.I0(CLBLM_L_X12Y138_SLICE_X16Y138_BQ),
.I1(CLBLM_L_X12Y138_SLICE_X17Y138_BO6),
.I2(CLBLM_L_X12Y137_SLICE_X16Y137_CQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y145_SLICE_X12Y145_AQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X12Y138_SLICE_X16Y138_BO5),
.O6(CLBLM_L_X12Y138_SLICE_X16Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffd3331ffff3333)
  ) CLBLM_L_X12Y138_SLICE_X16Y138_ALUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(RIOB33_X105Y135_IOB_X1Y136_I),
.I3(CLBLM_R_X13Y139_SLICE_X18Y139_BO6),
.I4(CLBLM_L_X12Y138_SLICE_X17Y138_A5Q),
.I5(RIOB33_X105Y135_IOB_X1Y135_I),
.O5(CLBLM_L_X12Y138_SLICE_X16Y138_AO5),
.O6(CLBLM_L_X12Y138_SLICE_X16Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y138_SLICE_X17Y138_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y139_SLICE_X16Y139_BO6),
.Q(CLBLM_L_X12Y138_SLICE_X17Y138_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y138_SLICE_X17Y138_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y138_SLICE_X17Y138_AO6),
.Q(CLBLM_L_X12Y138_SLICE_X17Y138_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y138_SLICE_X17Y138_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y140_SLICE_X15Y140_AO6),
.Q(CLBLM_L_X12Y138_SLICE_X17Y138_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000fafa0000ffcc)
  ) CLBLM_L_X12Y138_SLICE_X17Y138_DLUT (
.I0(CLBLM_L_X10Y136_SLICE_X12Y136_BQ),
.I1(CLBLM_L_X12Y137_SLICE_X17Y137_AQ),
.I2(CLBLM_L_X12Y137_SLICE_X16Y137_DQ),
.I3(CLBLM_L_X12Y136_SLICE_X17Y136_DQ),
.I4(CLBLM_R_X11Y138_SLICE_X14Y138_DQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y138_SLICE_X17Y138_DO5),
.O6(CLBLM_L_X12Y138_SLICE_X17Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0222000002222222)
  ) CLBLM_L_X12Y138_SLICE_X17Y138_CLUT (
.I0(CLBLM_R_X13Y138_SLICE_X18Y138_AQ),
.I1(CLBLM_L_X10Y135_SLICE_X12Y135_DO6),
.I2(CLBLM_L_X12Y138_SLICE_X16Y138_BQ),
.I3(CLBLM_L_X12Y138_SLICE_X16Y138_CQ),
.I4(CLBLM_L_X12Y138_SLICE_X17Y138_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y138_SLICE_X17Y138_CO5),
.O6(CLBLM_L_X12Y138_SLICE_X17Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00400000c0000000)
  ) CLBLM_L_X12Y138_SLICE_X17Y138_BLUT (
.I0(CLBLM_L_X10Y135_SLICE_X12Y135_DO6),
.I1(CLBLM_R_X13Y138_SLICE_X18Y138_AQ),
.I2(CLBLM_L_X12Y138_SLICE_X17Y138_AQ),
.I3(CLBLM_L_X12Y138_SLICE_X16Y138_BQ),
.I4(CLBLM_L_X12Y138_SLICE_X16Y138_CQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y138_SLICE_X17Y138_BO5),
.O6(CLBLM_L_X12Y138_SLICE_X17Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0004040808)
  ) CLBLM_L_X12Y138_SLICE_X17Y138_ALUT (
.I0(CLBLM_L_X12Y138_SLICE_X17Y138_AQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_L_X10Y145_SLICE_X12Y145_AQ),
.I3(CLBLM_L_X10Y139_SLICE_X13Y139_AQ),
.I4(CLBLM_L_X12Y138_SLICE_X17Y138_CO5),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X12Y138_SLICE_X17Y138_AO5),
.O6(CLBLM_L_X12Y138_SLICE_X17Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y139_SLICE_X16Y139_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y139_SLICE_X17Y139_BO6),
.Q(CLBLM_L_X12Y139_SLICE_X16Y139_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y139_SLICE_X16Y139_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y139_SLICE_X16Y139_AO6),
.Q(CLBLM_L_X12Y139_SLICE_X16Y139_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y139_SLICE_X16Y139_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y139_SLICE_X16Y139_CO6),
.Q(CLBLM_L_X12Y139_SLICE_X16Y139_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc30ec20f0f0a0a0)
  ) CLBLM_L_X12Y139_SLICE_X16Y139_DLUT (
.I0(CLBLM_L_X8Y136_SLICE_X10Y136_DQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLM_L_X12Y139_SLICE_X17Y139_CQ),
.I4(CLBLM_R_X7Y139_SLICE_X8Y139_BQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y139_SLICE_X16Y139_DO5),
.O6(CLBLM_L_X12Y139_SLICE_X16Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0055550000)
  ) CLBLM_L_X12Y139_SLICE_X16Y139_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_L_X12Y140_SLICE_X17Y140_AQ),
.I4(CLBLM_R_X7Y139_SLICE_X8Y139_A5Q),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X12Y139_SLICE_X16Y139_CO5),
.O6(CLBLM_L_X12Y139_SLICE_X16Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0ccf088cccc8888)
  ) CLBLM_L_X12Y139_SLICE_X16Y139_BLUT (
.I0(CLBLM_R_X7Y139_SLICE_X8Y139_A5Q),
.I1(RIOB33_X105Y121_IOB_X1Y121_I),
.I2(CLBLM_L_X12Y139_SLICE_X16Y139_CQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X11Y137_SLICE_X15Y137_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y139_SLICE_X16Y139_BO5),
.O6(CLBLM_L_X12Y139_SLICE_X16Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffccffccffcc00)
  ) CLBLM_L_X12Y139_SLICE_X16Y139_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X12Y134_SLICE_X17Y134_AQ),
.I2(1'b1),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X11Y139_SLICE_X15Y139_BQ),
.I5(CLBLM_R_X13Y141_SLICE_X18Y141_AO6),
.O5(CLBLM_L_X12Y139_SLICE_X16Y139_AO5),
.O6(CLBLM_L_X12Y139_SLICE_X16Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y139_SLICE_X17Y139_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y139_SLICE_X17Y139_AO6),
.Q(CLBLM_L_X12Y139_SLICE_X17Y139_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y139_SLICE_X17Y139_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y139_SLICE_X17Y139_CO6),
.Q(CLBLM_L_X12Y139_SLICE_X17Y139_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555505055445544)
  ) CLBLM_L_X12Y139_SLICE_X17Y139_DLUT (
.I0(CLBLM_R_X11Y138_SLICE_X14Y138_DQ),
.I1(CLBLM_L_X12Y135_SLICE_X17Y135_A5Q),
.I2(CLBLL_L_X4Y138_SLICE_X5Y138_B5Q),
.I3(CLBLM_L_X8Y136_SLICE_X10Y136_BQ),
.I4(CLBLM_L_X12Y139_SLICE_X17Y139_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y139_SLICE_X17Y139_DO5),
.O6(CLBLM_L_X12Y139_SLICE_X17Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaac0c0aaaaff00)
  ) CLBLM_L_X12Y139_SLICE_X17Y139_CLUT (
.I0(CLBLM_L_X10Y144_SLICE_X13Y144_AQ),
.I1(CLBLM_L_X12Y139_SLICE_X17Y139_CQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_L_X12Y133_SLICE_X16Y133_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X10Y135_SLICE_X12Y135_DO6),
.O5(CLBLM_L_X12Y139_SLICE_X17Y139_CO5),
.O6(CLBLM_L_X12Y139_SLICE_X17Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hce02ce0200003030)
  ) CLBLM_L_X12Y139_SLICE_X17Y139_BLUT (
.I0(CLBLM_L_X8Y141_SLICE_X10Y141_DQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_L_X12Y140_SLICE_X16Y140_CQ),
.I4(CLBLM_L_X10Y145_SLICE_X12Y145_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y139_SLICE_X17Y139_BO5),
.O6(CLBLM_L_X12Y139_SLICE_X17Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffd8d8d888)
  ) CLBLM_L_X12Y139_SLICE_X17Y139_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X13Y139_SLICE_X18Y139_AQ),
.I2(CLBLM_L_X12Y139_SLICE_X17Y139_AQ),
.I3(CLBLM_L_X8Y138_SLICE_X10Y138_AQ),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLM_L_X10Y135_SLICE_X12Y135_CO6),
.O5(CLBLM_L_X12Y139_SLICE_X17Y139_AO5),
.O6(CLBLM_L_X12Y139_SLICE_X17Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y140_SLICE_X16Y140_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y140_SLICE_X16Y140_AO6),
.Q(CLBLM_L_X12Y140_SLICE_X16Y140_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y140_SLICE_X16Y140_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y140_SLICE_X16Y140_BO6),
.Q(CLBLM_L_X12Y140_SLICE_X16Y140_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y140_SLICE_X16Y140_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y140_SLICE_X16Y140_CO6),
.Q(CLBLM_L_X12Y140_SLICE_X16Y140_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y140_SLICE_X16Y140_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y140_SLICE_X16Y140_DO6),
.Q(CLBLM_L_X12Y140_SLICE_X16Y140_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000005500550)
  ) CLBLM_L_X12Y140_SLICE_X16Y140_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(1'b1),
.I2(CLBLM_L_X12Y139_SLICE_X16Y139_BO5),
.I3(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I4(CLBLM_L_X12Y139_SLICE_X16Y139_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X12Y140_SLICE_X16Y140_DO5),
.O6(CLBLM_L_X12Y140_SLICE_X16Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa0000f0f0)
  ) CLBLM_L_X12Y140_SLICE_X16Y140_CLUT (
.I0(CLBLM_L_X8Y140_SLICE_X10Y140_AQ),
.I1(1'b1),
.I2(CLBLM_L_X12Y141_SLICE_X16Y141_BQ),
.I3(1'b1),
.I4(CLBLM_R_X13Y141_SLICE_X18Y141_AO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X12Y140_SLICE_X16Y140_CO5),
.O6(CLBLM_L_X12Y140_SLICE_X16Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000c0cff00aaaa)
  ) CLBLM_L_X12Y140_SLICE_X16Y140_BLUT (
.I0(CLBLM_L_X12Y143_SLICE_X16Y143_CQ),
.I1(CLBLM_L_X12Y140_SLICE_X16Y140_BQ),
.I2(CLBLM_R_X13Y143_SLICE_X18Y143_AO6),
.I3(CLBLM_R_X5Y138_SLICE_X7Y138_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X12Y143_SLICE_X17Y143_CO5),
.O5(CLBLM_L_X12Y140_SLICE_X16Y140_BO5),
.O6(CLBLM_L_X12Y140_SLICE_X16Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffa800a8ffa800a8)
  ) CLBLM_L_X12Y140_SLICE_X16Y140_ALUT (
.I0(CLBLM_L_X8Y143_SLICE_X10Y143_DO6),
.I1(CLBLM_L_X12Y138_SLICE_X16Y138_DQ),
.I2(CLBLM_L_X12Y140_SLICE_X16Y140_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X13Y135_SLICE_X18Y135_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y140_SLICE_X16Y140_AO5),
.O6(CLBLM_L_X12Y140_SLICE_X16Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y140_SLICE_X17Y140_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y140_SLICE_X17Y140_AO6),
.Q(CLBLM_L_X12Y140_SLICE_X17Y140_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y140_SLICE_X17Y140_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y140_SLICE_X17Y140_BO6),
.Q(CLBLM_L_X12Y140_SLICE_X17Y140_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y140_SLICE_X17Y140_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y140_SLICE_X17Y140_CO6),
.Q(CLBLM_L_X12Y140_SLICE_X17Y140_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcc3033cfcc3033)
  ) CLBLM_L_X12Y140_SLICE_X17Y140_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X13Y144_SLICE_X18Y144_CO6),
.I2(CLBLM_R_X13Y141_SLICE_X18Y141_BO5),
.I3(CLBLM_L_X12Y140_SLICE_X17Y140_BQ),
.I4(CLBLM_L_X12Y140_SLICE_X17Y140_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y140_SLICE_X17Y140_DO5),
.O6(CLBLM_L_X12Y140_SLICE_X17Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f04444ff00)
  ) CLBLM_L_X12Y140_SLICE_X17Y140_CLUT (
.I0(CLBLM_R_X13Y143_SLICE_X18Y143_AO6),
.I1(CLBLM_L_X12Y140_SLICE_X17Y140_CQ),
.I2(CLBLM_L_X12Y136_SLICE_X16Y136_AQ),
.I3(CLBLM_L_X12Y140_SLICE_X17Y140_BQ),
.I4(CLBLM_L_X12Y143_SLICE_X17Y143_CO5),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X12Y140_SLICE_X17Y140_CO5),
.O6(CLBLM_L_X12Y140_SLICE_X17Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcff3033fcfe3032)
  ) CLBLM_L_X12Y140_SLICE_X17Y140_BLUT (
.I0(CLBLM_L_X12Y142_SLICE_X16Y142_CQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X13Y143_SLICE_X18Y143_AO6),
.I3(CLBLM_L_X12Y143_SLICE_X17Y143_CO5),
.I4(CLBLM_L_X8Y141_SLICE_X11Y141_CQ),
.I5(CLBLM_L_X12Y140_SLICE_X17Y140_BQ),
.O5(CLBLM_L_X12Y140_SLICE_X17Y140_BO5),
.O6(CLBLM_L_X12Y140_SLICE_X17Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ccff4455ccff)
  ) CLBLM_L_X12Y140_SLICE_X17Y140_ALUT (
.I0(CLBLM_L_X12Y140_SLICE_X17Y140_DO6),
.I1(CLBLM_L_X8Y134_SLICE_X11Y134_BQ),
.I2(1'b1),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X12Y143_SLICE_X17Y143_DO6),
.I5(CLBLM_R_X13Y141_SLICE_X18Y141_AO5),
.O5(CLBLM_L_X12Y140_SLICE_X17Y140_AO5),
.O6(CLBLM_L_X12Y140_SLICE_X17Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y141_SLICE_X16Y141_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y141_SLICE_X16Y141_AO6),
.Q(CLBLM_L_X12Y141_SLICE_X16Y141_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y141_SLICE_X16Y141_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y141_SLICE_X16Y141_BO6),
.Q(CLBLM_L_X12Y141_SLICE_X16Y141_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0d0f0d0ff2f0f2f0)
  ) CLBLM_L_X12Y141_SLICE_X16Y141_DLUT (
.I0(CLBLM_R_X11Y140_SLICE_X14Y140_AQ),
.I1(CLBLM_R_X13Y141_SLICE_X18Y141_BO5),
.I2(CLBLM_R_X13Y144_SLICE_X18Y144_CO6),
.I3(CLBLM_L_X12Y141_SLICE_X16Y141_CO6),
.I4(1'b1),
.I5(CLBLM_L_X12Y141_SLICE_X16Y141_AQ),
.O5(CLBLM_L_X12Y141_SLICE_X16Y141_DO5),
.O6(CLBLM_L_X12Y141_SLICE_X16Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00034002c000c000)
  ) CLBLM_L_X12Y141_SLICE_X16Y141_CLUT (
.I0(CLBLM_R_X13Y144_SLICE_X18Y144_AQ),
.I1(CLBLM_L_X12Y140_SLICE_X17Y140_AQ),
.I2(CLBLM_L_X12Y142_SLICE_X17Y142_AQ),
.I3(CLBLM_L_X12Y142_SLICE_X16Y142_AQ),
.I4(CLBLM_R_X13Y140_SLICE_X18Y140_BQ),
.I5(CLBLM_L_X12Y142_SLICE_X16Y142_BQ),
.O5(CLBLM_L_X12Y141_SLICE_X16Y141_CO5),
.O6(CLBLM_L_X12Y141_SLICE_X16Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff0ff0000f000e0)
  ) CLBLM_L_X12Y141_SLICE_X16Y141_BLUT (
.I0(CLBLM_R_X13Y140_SLICE_X18Y140_BQ),
.I1(CLBLM_L_X12Y142_SLICE_X16Y142_BQ),
.I2(CLBLM_L_X12Y139_SLICE_X16Y139_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X13Y144_SLICE_X18Y144_AQ),
.I5(CLBLM_L_X12Y143_SLICE_X17Y143_BQ),
.O5(CLBLM_L_X12Y141_SLICE_X16Y141_BO5),
.O6(CLBLM_L_X12Y141_SLICE_X16Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h33bb33bb030b030b)
  ) CLBLM_L_X12Y141_SLICE_X16Y141_ALUT (
.I0(CLBLM_L_X12Y141_SLICE_X16Y141_DO6),
.I1(CLBLM_L_X12Y143_SLICE_X17Y143_DO6),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X13Y141_SLICE_X18Y141_AO5),
.I4(1'b1),
.I5(CLBLM_L_X8Y141_SLICE_X10Y141_DQ),
.O5(CLBLM_L_X12Y141_SLICE_X16Y141_AO5),
.O6(CLBLM_L_X12Y141_SLICE_X16Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y141_SLICE_X17Y141_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y141_SLICE_X17Y141_AO6),
.Q(CLBLM_L_X12Y141_SLICE_X17Y141_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h44574455ffffffff)
  ) CLBLM_L_X12Y141_SLICE_X17Y141_DLUT (
.I0(CLBLM_R_X13Y144_SLICE_X18Y144_AQ),
.I1(CLBLM_L_X12Y143_SLICE_X17Y143_BQ),
.I2(CLBLM_R_X13Y140_SLICE_X18Y140_BQ),
.I3(CLBLM_L_X12Y142_SLICE_X16Y142_BQ),
.I4(CLBLM_R_X13Y140_SLICE_X19Y140_AQ),
.I5(CLBLM_L_X12Y140_SLICE_X16Y140_CQ),
.O5(CLBLM_L_X12Y141_SLICE_X17Y141_DO5),
.O6(CLBLM_L_X12Y141_SLICE_X17Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hddddcccc5dd548c0)
  ) CLBLM_L_X12Y141_SLICE_X17Y141_CLUT (
.I0(CLBLM_L_X12Y143_SLICE_X17Y143_AQ),
.I1(CLBLM_R_X13Y140_SLICE_X18Y140_CQ),
.I2(CLBLM_R_X13Y141_SLICE_X18Y141_CO6),
.I3(CLBLM_L_X12Y136_SLICE_X17Y136_A5Q),
.I4(CLBLM_L_X12Y141_SLICE_X17Y141_BO5),
.I5(CLBLM_L_X12Y141_SLICE_X17Y141_DO6),
.O5(CLBLM_L_X12Y141_SLICE_X17Y141_CO5),
.O6(CLBLM_L_X12Y141_SLICE_X17Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h1111115500003300)
  ) CLBLM_L_X12Y141_SLICE_X17Y141_BLUT (
.I0(CLBLM_L_X12Y142_SLICE_X17Y142_AQ),
.I1(CLBLM_L_X12Y142_SLICE_X16Y142_BQ),
.I2(1'b1),
.I3(CLBLM_R_X13Y140_SLICE_X18Y140_BQ),
.I4(CLBLM_R_X13Y144_SLICE_X18Y144_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y141_SLICE_X17Y141_BO5),
.O6(CLBLM_L_X12Y141_SLICE_X17Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0f3f3c0c0c0d1)
  ) CLBLM_L_X12Y141_SLICE_X17Y141_ALUT (
.I0(CLBLM_R_X13Y140_SLICE_X18Y140_BQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X13Y140_SLICE_X19Y140_AQ),
.I3(CLBLM_L_X12Y142_SLICE_X16Y142_BQ),
.I4(CLBLM_R_X13Y144_SLICE_X18Y144_AQ),
.I5(CLBLM_L_X12Y143_SLICE_X17Y143_BQ),
.O5(CLBLM_L_X12Y141_SLICE_X17Y141_AO5),
.O6(CLBLM_L_X12Y141_SLICE_X17Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y142_SLICE_X16Y142_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y139_SLICE_X16Y139_DO6),
.Q(CLBLM_L_X12Y142_SLICE_X16Y142_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y142_SLICE_X16Y142_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y142_SLICE_X16Y142_AO6),
.Q(CLBLM_L_X12Y142_SLICE_X16Y142_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y142_SLICE_X16Y142_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y142_SLICE_X16Y142_BO6),
.Q(CLBLM_L_X12Y142_SLICE_X16Y142_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y142_SLICE_X16Y142_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y142_SLICE_X16Y142_CO6),
.Q(CLBLM_L_X12Y142_SLICE_X16Y142_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000fdefffff)
  ) CLBLM_L_X12Y142_SLICE_X16Y142_DLUT (
.I0(CLBLM_L_X12Y142_SLICE_X17Y142_AQ),
.I1(CLBLM_R_X13Y141_SLICE_X18Y141_BO5),
.I2(CLBLM_R_X13Y141_SLICE_X18Y141_CO5),
.I3(CLBLM_L_X12Y140_SLICE_X17Y140_AQ),
.I4(CLBLM_R_X11Y140_SLICE_X14Y140_BQ),
.I5(CLBLM_R_X13Y144_SLICE_X18Y144_CO6),
.O5(CLBLM_L_X12Y142_SLICE_X16Y142_DO5),
.O6(CLBLM_L_X12Y142_SLICE_X16Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0afa0a0acafaca0)
  ) CLBLM_L_X12Y142_SLICE_X16Y142_CLUT (
.I0(CLBLM_L_X10Y142_SLICE_X12Y142_AQ),
.I1(CLBLM_L_X12Y142_SLICE_X16Y142_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X12Y143_SLICE_X17Y143_CO5),
.I4(CLBLM_L_X12Y140_SLICE_X16Y140_BQ),
.I5(CLBLM_R_X13Y143_SLICE_X18Y143_AO6),
.O5(CLBLM_L_X12Y142_SLICE_X16Y142_CO5),
.O6(CLBLM_L_X12Y142_SLICE_X16Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hafaeaaae05040004)
  ) CLBLM_L_X12Y142_SLICE_X16Y142_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X12Y142_SLICE_X16Y142_BQ),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLM_R_X13Y141_SLICE_X19Y141_CO6),
.I4(CLBLM_R_X13Y140_SLICE_X18Y140_BQ),
.I5(CLBLM_R_X5Y135_SLICE_X7Y135_A5Q),
.O5(CLBLM_L_X12Y142_SLICE_X16Y142_BO5),
.O6(CLBLM_L_X12Y142_SLICE_X16Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00cc00ff84cca5ff)
  ) CLBLM_L_X12Y142_SLICE_X16Y142_ALUT (
.I0(CLBLM_L_X12Y142_SLICE_X16Y142_DO6),
.I1(CLBLM_R_X11Y144_SLICE_X15Y144_BQ),
.I2(CLBLM_L_X12Y142_SLICE_X16Y142_AQ),
.I3(CLBLM_L_X12Y143_SLICE_X17Y143_DO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X13Y141_SLICE_X18Y141_AO5),
.O5(CLBLM_L_X12Y142_SLICE_X16Y142_AO5),
.O6(CLBLM_L_X12Y142_SLICE_X16Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y142_SLICE_X17Y142_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y142_SLICE_X17Y142_AO6),
.Q(CLBLM_L_X12Y142_SLICE_X17Y142_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y142_SLICE_X17Y142_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y142_SLICE_X17Y142_BO6),
.Q(CLBLM_L_X12Y142_SLICE_X17Y142_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0ff0d2f078)
  ) CLBLM_L_X12Y142_SLICE_X17Y142_DLUT (
.I0(CLBLM_L_X12Y140_SLICE_X17Y140_CQ),
.I1(CLBLM_L_X12Y140_SLICE_X17Y140_AQ),
.I2(CLBLM_L_X12Y142_SLICE_X17Y142_AQ),
.I3(CLBLM_R_X13Y141_SLICE_X18Y141_BO5),
.I4(CLBLM_R_X13Y141_SLICE_X18Y141_CO5),
.I5(CLBLM_R_X13Y144_SLICE_X18Y144_CO6),
.O5(CLBLM_L_X12Y142_SLICE_X17Y142_DO5),
.O6(CLBLM_L_X12Y142_SLICE_X17Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h040000000c000c00)
  ) CLBLM_L_X12Y142_SLICE_X17Y142_CLUT (
.I0(CLBLM_L_X12Y143_SLICE_X17Y143_AQ),
.I1(CLBLM_R_X13Y144_SLICE_X18Y144_AQ),
.I2(CLBLM_R_X13Y140_SLICE_X19Y140_AQ),
.I3(CLBLM_L_X12Y143_SLICE_X17Y143_BQ),
.I4(CLBLM_R_X13Y141_SLICE_X19Y141_CO6),
.I5(1'b1),
.O5(CLBLM_L_X12Y142_SLICE_X17Y142_CO5),
.O6(CLBLM_L_X12Y142_SLICE_X17Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h55055505dd0d7707)
  ) CLBLM_L_X12Y142_SLICE_X17Y142_BLUT (
.I0(CLBLM_L_X12Y143_SLICE_X17Y143_DO6),
.I1(CLBLM_L_X12Y142_SLICE_X17Y142_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y141_SLICE_X13Y141_BQ),
.I4(CLBLM_R_X13Y142_SLICE_X18Y142_BO6),
.I5(CLBLM_R_X13Y141_SLICE_X18Y141_AO5),
.O5(CLBLM_L_X12Y142_SLICE_X17Y142_BO5),
.O6(CLBLM_L_X12Y142_SLICE_X17Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h51515151f351f351)
  ) CLBLM_L_X12Y142_SLICE_X17Y142_ALUT (
.I0(CLBLM_L_X12Y143_SLICE_X17Y143_DO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X11Y141_SLICE_X15Y141_AQ),
.I3(CLBLM_L_X12Y142_SLICE_X17Y142_DO6),
.I4(1'b1),
.I5(CLBLM_R_X13Y141_SLICE_X18Y141_AO5),
.O5(CLBLM_L_X12Y142_SLICE_X17Y142_AO5),
.O6(CLBLM_L_X12Y142_SLICE_X17Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y143_SLICE_X16Y143_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y143_SLICE_X16Y143_AO6),
.Q(CLBLM_L_X12Y143_SLICE_X16Y143_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y143_SLICE_X16Y143_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y143_SLICE_X16Y143_BO6),
.Q(CLBLM_L_X12Y143_SLICE_X16Y143_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y143_SLICE_X16Y143_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y143_SLICE_X16Y143_CO6),
.Q(CLBLM_L_X12Y143_SLICE_X16Y143_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y143_SLICE_X16Y143_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y143_SLICE_X16Y143_DO5),
.O6(CLBLM_L_X12Y143_SLICE_X16Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff4f4000004f40)
  ) CLBLM_L_X12Y143_SLICE_X16Y143_CLUT (
.I0(CLBLM_R_X13Y143_SLICE_X18Y143_AO6),
.I1(CLBLM_L_X12Y143_SLICE_X16Y143_CQ),
.I2(CLBLM_L_X12Y143_SLICE_X17Y143_CO5),
.I3(CLBLM_R_X11Y142_SLICE_X14Y142_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y139_SLICE_X10Y139_BQ),
.O5(CLBLM_L_X12Y143_SLICE_X16Y143_CO5),
.O6(CLBLM_L_X12Y143_SLICE_X16Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffd00fdffff00ff)
  ) CLBLM_L_X12Y143_SLICE_X16Y143_BLUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(RIOB33_X105Y135_IOB_X1Y135_I),
.I2(CLBLM_R_X13Y139_SLICE_X18Y139_BO6),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X12Y141_SLICE_X16Y141_BQ),
.I5(RIOB33_X105Y135_IOB_X1Y136_I),
.O5(CLBLM_L_X12Y143_SLICE_X16Y143_BO5),
.O6(CLBLM_L_X12Y143_SLICE_X16Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffeff33333233)
  ) CLBLM_L_X12Y143_SLICE_X16Y143_ALUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X13Y139_SLICE_X18Y139_BO6),
.I3(RIOB33_X105Y135_IOB_X1Y135_I),
.I4(RIOB33_X105Y135_IOB_X1Y136_I),
.I5(CLBLM_L_X12Y142_SLICE_X16Y142_A5Q),
.O5(CLBLM_L_X12Y143_SLICE_X16Y143_AO5),
.O6(CLBLM_L_X12Y143_SLICE_X16Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y143_SLICE_X17Y143_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y143_SLICE_X17Y143_AO6),
.Q(CLBLM_L_X12Y143_SLICE_X17Y143_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y143_SLICE_X17Y143_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y143_SLICE_X17Y143_BO6),
.Q(CLBLM_L_X12Y143_SLICE_X17Y143_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00ff0075007d)
  ) CLBLM_L_X12Y143_SLICE_X17Y143_DLUT (
.I0(CLBLM_R_X13Y141_SLICE_X19Y141_CO5),
.I1(CLBLM_R_X13Y140_SLICE_X18Y140_BQ),
.I2(CLBLM_L_X12Y142_SLICE_X16Y142_BQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X13Y144_SLICE_X18Y144_AQ),
.I5(CLBLM_R_X13Y144_SLICE_X18Y144_BO6),
.O5(CLBLM_L_X12Y143_SLICE_X17Y143_DO5),
.O6(CLBLM_L_X12Y143_SLICE_X17Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h2f3f3f3f00c000c0)
  ) CLBLM_L_X12Y143_SLICE_X17Y143_CLUT (
.I0(CLBLM_R_X13Y141_SLICE_X19Y141_CO5),
.I1(CLBLM_R_X13Y140_SLICE_X19Y140_AQ),
.I2(CLBLM_R_X13Y137_SLICE_X18Y137_CO5),
.I3(CLBLM_L_X12Y143_SLICE_X17Y143_BQ),
.I4(CLBLM_R_X13Y144_SLICE_X18Y144_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y143_SLICE_X17Y143_CO5),
.O6(CLBLM_L_X12Y143_SLICE_X17Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa03aa0caa03aa03)
  ) CLBLM_L_X12Y143_SLICE_X17Y143_BLUT (
.I0(CLBLM_R_X7Y141_SLICE_X9Y141_BQ),
.I1(CLBLM_L_X12Y143_SLICE_X17Y143_BQ),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X12Y142_SLICE_X17Y142_CO6),
.I5(CLBLM_L_X12Y143_SLICE_X17Y143_CO6),
.O5(CLBLM_L_X12Y143_SLICE_X17Y143_BO5),
.O6(CLBLM_L_X12Y143_SLICE_X17Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffa5550ffba5510)
  ) CLBLM_L_X12Y143_SLICE_X17Y143_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X13Y144_SLICE_X18Y144_BO6),
.I2(CLBLM_L_X12Y143_SLICE_X17Y143_AQ),
.I3(CLBLM_L_X12Y142_SLICE_X17Y142_CO6),
.I4(CLBLM_L_X8Y137_SLICE_X11Y137_AQ),
.I5(CLBLM_R_X13Y141_SLICE_X18Y141_AO5),
.O5(CLBLM_L_X12Y143_SLICE_X17Y143_AO5),
.O6(CLBLM_L_X12Y143_SLICE_X17Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y144_SLICE_X16Y144_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y77_IOB_X0Y77_I),
.D(CLBLM_L_X10Y141_SLICE_X12Y141_C5Q),
.Q(CLBLM_L_X12Y144_SLICE_X16Y144_AQ),
.R(CLBLM_L_X12Y144_SLICE_X16Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y144_SLICE_X16Y144_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y144_SLICE_X16Y144_DO5),
.O6(CLBLM_L_X12Y144_SLICE_X16Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y144_SLICE_X16Y144_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y144_SLICE_X16Y144_CO5),
.O6(CLBLM_L_X12Y144_SLICE_X16Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y144_SLICE_X16Y144_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y144_SLICE_X16Y144_BO5),
.O6(CLBLM_L_X12Y144_SLICE_X16Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00ff000f000f)
  ) CLBLM_L_X12Y144_SLICE_X16Y144_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(RIOB33_X105Y141_IOB_X1Y142_I),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLM_R_X7Y131_SLICE_X9Y131_AQ),
.O5(CLBLM_L_X12Y144_SLICE_X16Y144_AO5),
.O6(CLBLM_L_X12Y144_SLICE_X16Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y144_SLICE_X17Y144_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y144_SLICE_X17Y144_AO6),
.Q(CLBLM_L_X12Y144_SLICE_X17Y144_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y144_SLICE_X17Y144_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y144_SLICE_X17Y144_DO5),
.O6(CLBLM_L_X12Y144_SLICE_X17Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y144_SLICE_X17Y144_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y144_SLICE_X17Y144_CO5),
.O6(CLBLM_L_X12Y144_SLICE_X17Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y144_SLICE_X17Y144_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y144_SLICE_X17Y144_BO5),
.O6(CLBLM_L_X12Y144_SLICE_X17Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf055f000f3f3f3f3)
  ) CLBLM_L_X12Y144_SLICE_X17Y144_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(RIOB33_X105Y143_IOB_X1Y143_I),
.I2(CLBLM_R_X13Y143_SLICE_X18Y143_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y140_SLICE_X11Y140_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y144_SLICE_X17Y144_AO5),
.O6(CLBLM_L_X12Y144_SLICE_X17Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y146_SLICE_X16Y146_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y146_SLICE_X16Y146_DO5),
.O6(CLBLM_L_X12Y146_SLICE_X16Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y146_SLICE_X16Y146_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y146_SLICE_X16Y146_CO5),
.O6(CLBLM_L_X12Y146_SLICE_X16Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y146_SLICE_X16Y146_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y146_SLICE_X16Y146_BO5),
.O6(CLBLM_L_X12Y146_SLICE_X16Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff00fffcfc3030)
  ) CLBLM_L_X12Y146_SLICE_X16Y146_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X12Y142_SLICE_X16Y142_A5Q),
.I3(RIOB33_X105Y143_IOB_X1Y143_I),
.I4(CLBLM_L_X12Y144_SLICE_X16Y144_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y146_SLICE_X16Y146_AO5),
.O6(CLBLM_L_X12Y146_SLICE_X16Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y146_SLICE_X17Y146_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y146_SLICE_X17Y146_DO5),
.O6(CLBLM_L_X12Y146_SLICE_X17Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y146_SLICE_X17Y146_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y146_SLICE_X17Y146_CO5),
.O6(CLBLM_L_X12Y146_SLICE_X17Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y146_SLICE_X17Y146_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y146_SLICE_X17Y146_BO5),
.O6(CLBLM_L_X12Y146_SLICE_X17Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y146_SLICE_X17Y146_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y146_SLICE_X17Y146_AO5),
.O6(CLBLM_L_X12Y146_SLICE_X17Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y133_SLICE_X2Y133_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y133_SLICE_X2Y133_DO5),
.O6(CLBLM_R_X3Y133_SLICE_X2Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffb3b3b3ffa0a0a0)
  ) CLBLM_R_X3Y133_SLICE_X2Y133_CLUT (
.I0(CLBLL_L_X4Y142_SLICE_X5Y142_DO6),
.I1(CLBLL_L_X4Y135_SLICE_X4Y135_DO5),
.I2(LIOB33_X0Y51_IOB_X0Y51_I),
.I3(LIOB33_X0Y53_IOB_X0Y53_I),
.I4(CLBLM_R_X5Y141_SLICE_X7Y141_DO6),
.I5(CLBLM_R_X5Y140_SLICE_X6Y140_AO6),
.O5(CLBLM_R_X3Y133_SLICE_X2Y133_CO5),
.O6(CLBLM_R_X3Y133_SLICE_X2Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ec00ff00a000)
  ) CLBLM_R_X3Y133_SLICE_X2Y133_BLUT (
.I0(CLBLL_L_X4Y135_SLICE_X5Y135_C5Q),
.I1(CLBLL_L_X4Y133_SLICE_X4Y133_BO5),
.I2(CLBLL_L_X4Y139_SLICE_X4Y139_BO6),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X3Y133_SLICE_X2Y133_CO6),
.I5(CLBLM_R_X3Y140_SLICE_X2Y140_DO6),
.O5(CLBLM_R_X3Y133_SLICE_X2Y133_BO5),
.O6(CLBLM_R_X3Y133_SLICE_X2Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffcfffffffaff)
  ) CLBLM_R_X3Y133_SLICE_X2Y133_ALUT (
.I0(CLBLM_R_X5Y141_SLICE_X7Y141_DO6),
.I1(CLBLL_L_X4Y142_SLICE_X5Y142_DO6),
.I2(RIOB33_X105Y129_IOB_X1Y129_I),
.I3(RIOB33_X105Y137_IOB_X1Y137_I),
.I4(RIOB33_X105Y127_IOB_X1Y128_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y133_SLICE_X2Y133_AO5),
.O6(CLBLM_R_X3Y133_SLICE_X2Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y133_SLICE_X3Y133_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y133_SLICE_X3Y133_AO6),
.Q(CLBLM_R_X3Y133_SLICE_X3Y133_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y133_SLICE_X3Y133_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y133_SLICE_X3Y133_DO5),
.O6(CLBLM_R_X3Y133_SLICE_X3Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y133_SLICE_X3Y133_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y133_SLICE_X3Y133_CO5),
.O6(CLBLM_R_X3Y133_SLICE_X3Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y133_SLICE_X3Y133_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y133_SLICE_X3Y133_BO5),
.O6(CLBLM_R_X3Y133_SLICE_X3Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'habba0110aaaa0000)
  ) CLBLM_R_X3Y133_SLICE_X3Y133_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLL_L_X4Y134_SLICE_X4Y134_BQ),
.I2(CLBLM_R_X3Y133_SLICE_X3Y133_AQ),
.I3(CLBLM_R_X3Y137_SLICE_X3Y137_AQ),
.I4(CLBLL_L_X4Y132_SLICE_X5Y132_AQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X3Y133_SLICE_X3Y133_AO5),
.O6(CLBLM_R_X3Y133_SLICE_X3Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y135_SLICE_X2Y135_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y135_SLICE_X2Y135_DO5),
.O6(CLBLM_R_X3Y135_SLICE_X2Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y135_SLICE_X2Y135_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y135_SLICE_X2Y135_CO5),
.O6(CLBLM_R_X3Y135_SLICE_X2Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y135_SLICE_X2Y135_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y135_SLICE_X2Y135_BO5),
.O6(CLBLM_R_X3Y135_SLICE_X2Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y135_SLICE_X2Y135_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y135_SLICE_X2Y135_AO5),
.O6(CLBLM_R_X3Y135_SLICE_X2Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y135_SLICE_X3Y135_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y135_SLICE_X3Y135_AO6),
.Q(CLBLM_R_X3Y135_SLICE_X3Y135_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y135_SLICE_X3Y135_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y135_SLICE_X3Y135_BO6),
.Q(CLBLM_R_X3Y135_SLICE_X3Y135_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y135_SLICE_X3Y135_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y135_SLICE_X3Y135_DO5),
.O6(CLBLM_R_X3Y135_SLICE_X3Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8888000088880000)
  ) CLBLM_R_X3Y135_SLICE_X3Y135_CLUT (
.I0(CLBLM_R_X3Y137_SLICE_X3Y137_AQ),
.I1(CLBLM_R_X3Y136_SLICE_X3Y136_AQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X3Y133_SLICE_X3Y133_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y135_SLICE_X3Y135_CO5),
.O6(CLBLM_R_X3Y135_SLICE_X3Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0dddd8888)
  ) CLBLM_R_X3Y135_SLICE_X3Y135_BLUT (
.I0(CLBLL_L_X4Y133_SLICE_X5Y133_BO6),
.I1(CLBLM_R_X3Y135_SLICE_X3Y135_BQ),
.I2(CLBLM_R_X3Y133_SLICE_X3Y133_AQ),
.I3(1'b1),
.I4(CLBLM_R_X5Y135_SLICE_X6Y135_D5Q),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X3Y135_SLICE_X3Y135_BO5),
.O6(CLBLM_R_X3Y135_SLICE_X3Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0002022020)
  ) CLBLM_R_X3Y135_SLICE_X3Y135_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLL_L_X4Y134_SLICE_X4Y134_BQ),
.I2(CLBLM_R_X3Y135_SLICE_X3Y135_AQ),
.I3(CLBLM_R_X7Y142_SLICE_X9Y142_AQ),
.I4(CLBLM_R_X3Y135_SLICE_X3Y135_CO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X3Y135_SLICE_X3Y135_AO5),
.O6(CLBLM_R_X3Y135_SLICE_X3Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y136_SLICE_X2Y136_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y136_SLICE_X2Y136_AO6),
.Q(CLBLM_R_X3Y136_SLICE_X2Y136_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y136_SLICE_X2Y136_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y136_SLICE_X2Y136_DO5),
.O6(CLBLM_R_X3Y136_SLICE_X2Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_R_X3Y136_SLICE_X2Y136_CLUT (
.I0(CLBLM_R_X3Y136_SLICE_X3Y136_AQ),
.I1(CLBLM_R_X3Y135_SLICE_X3Y135_AQ),
.I2(CLBLM_R_X3Y137_SLICE_X2Y137_BQ),
.I3(CLBLM_R_X3Y133_SLICE_X3Y133_AQ),
.I4(CLBLM_R_X3Y136_SLICE_X3Y136_DQ),
.I5(CLBLM_R_X3Y137_SLICE_X3Y137_AQ),
.O5(CLBLM_R_X3Y136_SLICE_X2Y136_CO5),
.O6(CLBLM_R_X3Y136_SLICE_X2Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h80000000c0000000)
  ) CLBLM_R_X3Y136_SLICE_X2Y136_BLUT (
.I0(CLBLM_R_X3Y137_SLICE_X2Y137_BQ),
.I1(CLBLM_R_X3Y135_SLICE_X3Y135_AQ),
.I2(CLBLM_R_X3Y137_SLICE_X3Y137_AQ),
.I3(CLBLM_R_X3Y133_SLICE_X3Y133_AQ),
.I4(CLBLM_R_X3Y136_SLICE_X3Y136_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y136_SLICE_X2Y136_BO5),
.O6(CLBLM_R_X3Y136_SLICE_X2Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000012001200)
  ) CLBLM_R_X3Y136_SLICE_X2Y136_ALUT (
.I0(CLBLM_R_X3Y137_SLICE_X3Y137_BO5),
.I1(CLBLL_L_X4Y134_SLICE_X4Y134_BQ),
.I2(CLBLM_R_X3Y136_SLICE_X2Y136_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLL_L_X4Y135_SLICE_X5Y135_C5Q),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X3Y136_SLICE_X2Y136_AO5),
.O6(CLBLM_R_X3Y136_SLICE_X2Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y136_SLICE_X3Y136_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y136_SLICE_X3Y136_AO6),
.Q(CLBLM_R_X3Y136_SLICE_X3Y136_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y136_SLICE_X3Y136_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y136_SLICE_X3Y136_BO6),
.Q(CLBLM_R_X3Y136_SLICE_X3Y136_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y136_SLICE_X3Y136_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y136_SLICE_X3Y136_CO6),
.Q(CLBLM_R_X3Y136_SLICE_X3Y136_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y136_SLICE_X3Y136_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y136_SLICE_X3Y136_DO6),
.Q(CLBLM_R_X3Y136_SLICE_X3Y136_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc05cc00cc50cc00)
  ) CLBLM_R_X3Y136_SLICE_X3Y136_DLUT (
.I0(CLBLL_L_X4Y134_SLICE_X4Y134_BQ),
.I1(CLBLM_L_X8Y135_SLICE_X10Y135_A5Q),
.I2(CLBLM_R_X3Y136_SLICE_X2Y136_BO6),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X3Y136_SLICE_X3Y136_DQ),
.O5(CLBLM_R_X3Y136_SLICE_X3Y136_DO5),
.O6(CLBLM_R_X3Y136_SLICE_X3Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hdf13ff33ec20cc00)
  ) CLBLM_R_X3Y136_SLICE_X3Y136_CLUT (
.I0(CLBLM_R_X3Y136_SLICE_X2Y136_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X3Y136_SLICE_X3Y136_BQ),
.I3(CLBLM_R_X7Y137_SLICE_X8Y137_CQ),
.I4(CLBLM_R_X3Y137_SLICE_X3Y137_BO5),
.I5(CLBLL_L_X4Y134_SLICE_X4Y134_BQ),
.O5(CLBLM_R_X3Y136_SLICE_X3Y136_CO5),
.O6(CLBLM_R_X3Y136_SLICE_X3Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf666fcccf000f000)
  ) CLBLM_R_X3Y136_SLICE_X3Y136_BLUT (
.I0(CLBLM_R_X3Y137_SLICE_X3Y137_BO5),
.I1(CLBLM_R_X3Y136_SLICE_X3Y136_BQ),
.I2(CLBLM_R_X5Y135_SLICE_X6Y135_D5Q),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X3Y136_SLICE_X2Y136_AQ),
.I5(CLBLM_R_X3Y137_SLICE_X3Y137_AO5),
.O5(CLBLM_R_X3Y136_SLICE_X3Y136_BO5),
.O6(CLBLM_R_X3Y136_SLICE_X3Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbe3cfaf0aa00aa00)
  ) CLBLM_R_X3Y136_SLICE_X3Y136_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X3Y133_SLICE_X3Y133_AQ),
.I2(CLBLM_R_X3Y136_SLICE_X3Y136_AQ),
.I3(CLBLM_R_X3Y139_SLICE_X3Y139_AQ),
.I4(CLBLM_R_X3Y137_SLICE_X3Y137_AQ),
.I5(CLBLM_R_X3Y137_SLICE_X3Y137_AO5),
.O5(CLBLM_R_X3Y136_SLICE_X3Y136_AO5),
.O6(CLBLM_R_X3Y136_SLICE_X3Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y137_SLICE_X2Y137_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y137_SLICE_X2Y137_AO6),
.Q(CLBLM_R_X3Y137_SLICE_X2Y137_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y137_SLICE_X2Y137_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y137_SLICE_X2Y137_BO6),
.Q(CLBLM_R_X3Y137_SLICE_X2Y137_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y137_SLICE_X2Y137_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y137_SLICE_X2Y137_DO5),
.O6(CLBLM_R_X3Y137_SLICE_X2Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y137_SLICE_X2Y137_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y137_SLICE_X2Y137_CO5),
.O6(CLBLM_R_X3Y137_SLICE_X2Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc005acccc0000)
  ) CLBLM_R_X3Y137_SLICE_X2Y137_BLUT (
.I0(CLBLM_R_X3Y136_SLICE_X2Y136_BO5),
.I1(CLBLM_R_X7Y138_SLICE_X8Y138_AQ),
.I2(CLBLM_R_X3Y137_SLICE_X2Y137_BQ),
.I3(CLBLL_L_X4Y134_SLICE_X4Y134_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X3Y137_SLICE_X2Y137_BO5),
.O6(CLBLM_R_X3Y137_SLICE_X2Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h888b888888b88888)
  ) CLBLM_R_X3Y137_SLICE_X2Y137_ALUT (
.I0(CLBLM_L_X10Y143_SLICE_X12Y143_CQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X3Y137_SLICE_X2Y137_AQ),
.I3(CLBLL_L_X4Y134_SLICE_X4Y134_BQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X3Y136_SLICE_X2Y136_CO6),
.O5(CLBLM_R_X3Y137_SLICE_X2Y137_AO5),
.O6(CLBLM_R_X3Y137_SLICE_X2Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y137_SLICE_X3Y137_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y137_SLICE_X3Y137_AO6),
.Q(CLBLM_R_X3Y137_SLICE_X3Y137_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y137_SLICE_X3Y137_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y137_SLICE_X3Y137_BO6),
.Q(CLBLM_R_X3Y137_SLICE_X3Y137_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y137_SLICE_X3Y137_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y137_SLICE_X3Y137_CO6),
.Q(CLBLM_R_X3Y137_SLICE_X3Y137_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6969969696696996)
  ) CLBLM_R_X3Y137_SLICE_X3Y137_DLUT (
.I0(CLBLL_L_X4Y142_SLICE_X5Y142_DO6),
.I1(CLBLM_R_X5Y142_SLICE_X6Y142_CO6),
.I2(CLBLL_L_X4Y141_SLICE_X4Y141_DO6),
.I3(CLBLM_R_X3Y139_SLICE_X2Y139_AO5),
.I4(CLBLL_L_X4Y142_SLICE_X4Y142_BO6),
.I5(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.O5(CLBLM_R_X3Y137_SLICE_X3Y137_DO5),
.O6(CLBLM_R_X3Y137_SLICE_X3Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haafeaafe00540054)
  ) CLBLM_R_X3Y137_SLICE_X3Y137_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X3Y137_SLICE_X3Y137_CQ),
.I2(CLBLM_R_X3Y137_SLICE_X3Y137_BQ),
.I3(CLBLL_L_X4Y133_SLICE_X5Y133_BO6),
.I4(1'b1),
.I5(CLBLM_L_X8Y140_SLICE_X10Y140_A5Q),
.O5(CLBLM_R_X3Y137_SLICE_X3Y137_CO5),
.O6(CLBLM_R_X3Y137_SLICE_X3Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccaaccaac0c00000)
  ) CLBLM_R_X3Y137_SLICE_X3Y137_BLUT (
.I0(CLBLL_L_X4Y137_SLICE_X4Y137_BQ),
.I1(CLBLM_R_X3Y136_SLICE_X3Y136_DQ),
.I2(CLBLM_R_X3Y136_SLICE_X2Y136_BO6),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X3Y137_SLICE_X2Y137_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y137_SLICE_X3Y137_BO5),
.O6(CLBLM_R_X3Y137_SLICE_X3Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h888d888800550000)
  ) CLBLM_R_X3Y137_SLICE_X3Y137_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y142_SLICE_X11Y142_BQ),
.I2(CLBLM_R_X3Y137_SLICE_X3Y137_AQ),
.I3(CLBLL_L_X4Y134_SLICE_X4Y134_BQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y137_SLICE_X3Y137_AO5),
.O6(CLBLM_R_X3Y137_SLICE_X3Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y138_SLICE_X2Y138_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y138_SLICE_X2Y138_DO5),
.O6(CLBLM_R_X3Y138_SLICE_X2Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y138_SLICE_X2Y138_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y138_SLICE_X2Y138_CO5),
.O6(CLBLM_R_X3Y138_SLICE_X2Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000000000a00c)
  ) CLBLM_R_X3Y138_SLICE_X2Y138_BLUT (
.I0(LIOB33_X0Y57_IOB_X0Y57_I),
.I1(CLBLM_R_X3Y135_SLICE_X3Y135_BQ),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(RIOB33_X105Y131_IOB_X1Y132_I),
.I4(CLBLM_R_X3Y138_SLICE_X2Y138_AO6),
.I5(CLBLM_R_X3Y143_SLICE_X2Y143_AO6),
.O5(CLBLM_R_X3Y138_SLICE_X2Y138_BO5),
.O6(CLBLM_R_X3Y138_SLICE_X2Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0fff0ff0fff0ff)
  ) CLBLM_R_X3Y138_SLICE_X2Y138_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(RIOB33_X105Y133_IOB_X1Y134_I),
.I3(RIOB33_X105Y133_IOB_X1Y133_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y138_SLICE_X2Y138_AO5),
.O6(CLBLM_R_X3Y138_SLICE_X2Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y138_SLICE_X3Y138_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y138_SLICE_X3Y138_AO6),
.Q(CLBLM_R_X3Y138_SLICE_X3Y138_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y138_SLICE_X3Y138_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y138_SLICE_X3Y138_DO5),
.O6(CLBLM_R_X3Y138_SLICE_X3Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y138_SLICE_X3Y138_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y138_SLICE_X3Y138_CO5),
.O6(CLBLM_R_X3Y138_SLICE_X3Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y138_SLICE_X3Y138_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y138_SLICE_X3Y138_BO5),
.O6(CLBLM_R_X3Y138_SLICE_X3Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccfc00f0ccfc00f0)
  ) CLBLM_R_X3Y138_SLICE_X3Y138_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X3Y138_SLICE_X3Y138_AQ),
.I3(CLBLM_R_X7Y133_SLICE_X8Y133_DO6),
.I4(CLBLL_L_X4Y137_SLICE_X4Y137_D5Q),
.I5(1'b1),
.O5(CLBLM_R_X3Y138_SLICE_X3Y138_AO5),
.O6(CLBLM_R_X3Y138_SLICE_X3Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000002f2f2222)
  ) CLBLM_R_X3Y139_SLICE_X2Y139_DLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X3Y143_SLICE_X3Y143_AO5),
.I2(CLBLM_R_X3Y143_SLICE_X3Y143_AO6),
.I3(1'b1),
.I4(CLBLL_L_X4Y133_SLICE_X5Y133_AQ),
.I5(CLBLM_R_X3Y143_SLICE_X2Y143_AO6),
.O5(CLBLM_R_X3Y139_SLICE_X2Y139_DO5),
.O6(CLBLM_R_X3Y139_SLICE_X2Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffefffffffee)
  ) CLBLM_R_X3Y139_SLICE_X2Y139_CLUT (
.I0(CLBLM_R_X3Y138_SLICE_X2Y138_BO6),
.I1(CLBLM_R_X3Y139_SLICE_X3Y139_CO6),
.I2(CLBLM_R_X3Y142_SLICE_X2Y142_AO6),
.I3(CLBLL_L_X4Y138_SLICE_X4Y138_CO6),
.I4(CLBLM_R_X3Y139_SLICE_X2Y139_DO6),
.I5(CLBLM_R_X5Y138_SLICE_X6Y138_AQ),
.O5(CLBLM_R_X3Y139_SLICE_X2Y139_CO5),
.O6(CLBLM_R_X3Y139_SLICE_X2Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0705ffff0300)
  ) CLBLM_R_X3Y139_SLICE_X2Y139_BLUT (
.I0(CLBLL_L_X2Y140_SLICE_X1Y140_AO6),
.I1(CLBLM_R_X3Y143_SLICE_X3Y143_AO5),
.I2(CLBLM_R_X3Y143_SLICE_X2Y143_AO6),
.I3(LIOB33_X0Y65_IOB_X0Y65_I),
.I4(CLBLM_R_X3Y139_SLICE_X2Y139_AO6),
.I5(CLBLM_R_X3Y139_SLICE_X3Y139_AQ),
.O5(CLBLM_R_X3Y139_SLICE_X2Y139_BO5),
.O6(CLBLM_R_X3Y139_SLICE_X2Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd00dd00dddddddd)
  ) CLBLM_R_X3Y139_SLICE_X2Y139_ALUT (
.I0(RIOB33_X105Y137_IOB_X1Y137_I),
.I1(RIOB33_X105Y129_IOB_X1Y129_I),
.I2(1'b1),
.I3(CLBLM_L_X8Y140_SLICE_X10Y140_A5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y139_SLICE_X2Y139_AO5),
.O6(CLBLM_R_X3Y139_SLICE_X2Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y139_SLICE_X3Y139_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y139_SLICE_X3Y139_AO6),
.Q(CLBLM_R_X3Y139_SLICE_X3Y139_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcfdfcf00005500)
  ) CLBLM_R_X3Y139_SLICE_X3Y139_DLUT (
.I0(CLBLM_R_X3Y143_SLICE_X2Y143_AO6),
.I1(RIOB33_X105Y129_IOB_X1Y129_I),
.I2(RIOB33_X105Y137_IOB_X1Y137_I),
.I3(CLBLM_R_X3Y139_SLICE_X3Y139_AQ),
.I4(CLBLL_L_X2Y140_SLICE_X1Y140_AO6),
.I5(CLBLM_L_X8Y140_SLICE_X10Y140_A5Q),
.O5(CLBLM_R_X3Y139_SLICE_X3Y139_DO5),
.O6(CLBLM_R_X3Y139_SLICE_X3Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0c0c0e2c0)
  ) CLBLM_R_X3Y139_SLICE_X3Y139_CLUT (
.I0(RIOB33_X105Y115_IOB_X1Y116_I),
.I1(CLBLM_R_X3Y139_SLICE_X2Y139_AO5),
.I2(CLBLL_L_X4Y137_SLICE_X4Y137_D5Q),
.I3(CLBLL_L_X2Y140_SLICE_X1Y140_AO5),
.I4(RIOB33_X105Y129_IOB_X1Y130_I),
.I5(RIOB33_X105Y135_IOB_X1Y135_I),
.O5(CLBLM_R_X3Y139_SLICE_X3Y139_CO5),
.O6(CLBLM_R_X3Y139_SLICE_X3Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000001)
  ) CLBLM_R_X3Y139_SLICE_X3Y139_BLUT (
.I0(CLBLM_R_X3Y141_SLICE_X3Y141_CO6),
.I1(CLBLM_R_X3Y140_SLICE_X3Y140_BO6),
.I2(CLBLM_R_X5Y140_SLICE_X6Y140_AO6),
.I3(CLBLL_L_X4Y139_SLICE_X4Y139_BO6),
.I4(CLBLL_L_X4Y142_SLICE_X5Y142_DO6),
.I5(CLBLM_R_X5Y141_SLICE_X7Y141_DO6),
.O5(CLBLM_R_X3Y139_SLICE_X3Y139_BO5),
.O6(CLBLM_R_X3Y139_SLICE_X3Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00ccffccf0)
  ) CLBLM_R_X3Y139_SLICE_X3Y139_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I2(CLBLM_R_X3Y139_SLICE_X3Y139_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X5Y136_SLICE_X6Y136_DQ),
.I5(CLBLL_L_X4Y133_SLICE_X5Y133_BO6),
.O5(CLBLM_R_X3Y139_SLICE_X3Y139_AO5),
.O6(CLBLM_R_X3Y139_SLICE_X3Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffc)
  ) CLBLM_R_X3Y140_SLICE_X2Y140_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y142_SLICE_X2Y142_DO6),
.I2(CLBLM_R_X3Y140_SLICE_X3Y140_DO6),
.I3(CLBLL_L_X4Y140_SLICE_X5Y140_BO6),
.I4(CLBLM_R_X5Y140_SLICE_X7Y140_DO6),
.I5(CLBLM_R_X3Y140_SLICE_X2Y140_BO6),
.O5(CLBLM_R_X3Y140_SLICE_X2Y140_DO5),
.O6(CLBLM_R_X3Y140_SLICE_X2Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000800000000)
  ) CLBLM_R_X3Y140_SLICE_X2Y140_CLUT (
.I0(RIOB33_X105Y131_IOB_X1Y132_I),
.I1(CLBLM_R_X5Y136_SLICE_X6Y136_AQ),
.I2(CLBLM_R_X3Y143_SLICE_X2Y143_AO5),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(RIOB33_X105Y133_IOB_X1Y134_I),
.I5(RIOB33_X105Y133_IOB_X1Y133_I),
.O5(CLBLM_R_X3Y140_SLICE_X2Y140_CO5),
.O6(CLBLM_R_X3Y140_SLICE_X2Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffff3bff0a)
  ) CLBLM_R_X3Y140_SLICE_X2Y140_BLUT (
.I0(LIOB33_X0Y65_IOB_X0Y65_I),
.I1(CLBLM_R_X5Y143_SLICE_X6Y143_AO6),
.I2(CLBLM_R_X3Y141_SLICE_X2Y141_AO6),
.I3(CLBLM_R_X3Y139_SLICE_X3Y139_DO6),
.I4(CLBLL_L_X4Y136_SLICE_X4Y136_BQ),
.I5(CLBLM_R_X3Y140_SLICE_X2Y140_CO6),
.O5(CLBLM_R_X3Y140_SLICE_X2Y140_BO5),
.O6(CLBLM_R_X3Y140_SLICE_X2Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h000050500000dc50)
  ) CLBLM_R_X3Y140_SLICE_X2Y140_ALUT (
.I0(CLBLM_R_X3Y143_SLICE_X3Y143_AO6),
.I1(CLBLM_R_X5Y136_SLICE_X6Y136_AQ),
.I2(CLBLL_L_X4Y136_SLICE_X4Y136_BQ),
.I3(CLBLL_L_X2Y141_SLICE_X1Y141_AO6),
.I4(CLBLM_R_X3Y143_SLICE_X2Y143_AO5),
.I5(RIOB33_X105Y131_IOB_X1Y131_I),
.O5(CLBLM_R_X3Y140_SLICE_X2Y140_AO5),
.O6(CLBLM_R_X3Y140_SLICE_X2Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h55f555f500f000f0)
  ) CLBLM_R_X3Y140_SLICE_X3Y140_DLUT (
.I0(CLBLL_L_X4Y143_SLICE_X4Y143_BO5),
.I1(1'b1),
.I2(CLBLM_L_X10Y134_SLICE_X12Y134_BQ),
.I3(CLBLM_R_X7Y142_SLICE_X9Y142_CO6),
.I4(1'b1),
.I5(CLBLM_R_X11Y140_SLICE_X15Y140_C5Q),
.O5(CLBLM_R_X3Y140_SLICE_X3Y140_DO5),
.O6(CLBLM_R_X3Y140_SLICE_X3Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h03ab00aa03030000)
  ) CLBLM_R_X3Y140_SLICE_X3Y140_CLUT (
.I0(CLBLL_L_X2Y140_SLICE_X1Y140_AO5),
.I1(CLBLM_R_X3Y143_SLICE_X2Y143_AO6),
.I2(CLBLM_R_X3Y143_SLICE_X3Y143_AO6),
.I3(CLBLL_L_X4Y143_SLICE_X5Y143_BO5),
.I4(CLBLL_L_X4Y134_SLICE_X5Y134_BQ),
.I5(RIOB33_X105Y117_IOB_X1Y117_I),
.O5(CLBLM_R_X3Y140_SLICE_X3Y140_CO5),
.O6(CLBLM_R_X3Y140_SLICE_X3Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_R_X3Y140_SLICE_X3Y140_BLUT (
.I0(CLBLM_R_X3Y141_SLICE_X3Y141_BO6),
.I1(CLBLM_R_X3Y142_SLICE_X2Y142_DO6),
.I2(CLBLM_R_X5Y142_SLICE_X6Y142_AO6),
.I3(CLBLM_R_X5Y140_SLICE_X7Y140_DO6),
.I4(CLBLM_R_X3Y140_SLICE_X3Y140_AO6),
.I5(CLBLL_L_X4Y140_SLICE_X5Y140_BO6),
.O5(CLBLM_R_X3Y140_SLICE_X3Y140_BO5),
.O6(CLBLM_R_X3Y140_SLICE_X3Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafffafafefffefe)
  ) CLBLM_R_X3Y140_SLICE_X3Y140_ALUT (
.I0(CLBLM_R_X3Y139_SLICE_X2Y139_BO6),
.I1(CLBLM_L_X10Y134_SLICE_X12Y134_BQ),
.I2(CLBLM_R_X3Y140_SLICE_X2Y140_AO6),
.I3(CLBLL_L_X4Y143_SLICE_X4Y143_BO5),
.I4(CLBLM_R_X11Y140_SLICE_X15Y140_C5Q),
.I5(CLBLM_R_X7Y142_SLICE_X9Y142_CO6),
.O5(CLBLM_R_X3Y140_SLICE_X3Y140_AO5),
.O6(CLBLM_R_X3Y140_SLICE_X3Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffdfcf5f0)
  ) CLBLM_R_X3Y141_SLICE_X2Y141_DLUT (
.I0(CLBLM_R_X3Y141_SLICE_X2Y141_AO6),
.I1(CLBLM_R_X5Y141_SLICE_X6Y141_A5Q),
.I2(CLBLL_L_X2Y141_SLICE_X1Y141_CO6),
.I3(LIOB33_X0Y59_IOB_X0Y59_I),
.I4(CLBLM_R_X3Y139_SLICE_X2Y139_AO5),
.I5(CLBLM_R_X3Y141_SLICE_X2Y141_BO6),
.O5(CLBLM_R_X3Y141_SLICE_X2Y141_DO5),
.O6(CLBLM_R_X3Y141_SLICE_X2Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00aa00a000ee00ee)
  ) CLBLM_R_X3Y141_SLICE_X2Y141_CLUT (
.I0(CLBLM_R_X3Y143_SLICE_X2Y143_AO6),
.I1(CLBLL_L_X2Y141_SLICE_X1Y141_BO6),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(CLBLM_R_X3Y139_SLICE_X2Y139_AO5),
.I4(CLBLM_R_X3Y143_SLICE_X2Y143_AO5),
.I5(CLBLL_L_X2Y141_SLICE_X1Y141_AO6),
.O5(CLBLM_R_X3Y141_SLICE_X2Y141_CO5),
.O6(CLBLM_R_X3Y141_SLICE_X2Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000020000000000)
  ) CLBLM_R_X3Y141_SLICE_X2Y141_BLUT (
.I0(RIOB33_X105Y135_IOB_X1Y136_I),
.I1(RIOB33_X105Y129_IOB_X1Y130_I),
.I2(CLBLM_R_X3Y139_SLICE_X2Y139_AO5),
.I3(CLBLL_L_X2Y141_SLICE_X1Y141_AO6),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(RIOB33_X105Y135_IOB_X1Y135_I),
.O5(CLBLM_R_X3Y141_SLICE_X2Y141_BO5),
.O6(CLBLM_R_X3Y141_SLICE_X2Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff7fffffdffffff)
  ) CLBLM_R_X3Y141_SLICE_X2Y141_ALUT (
.I0(RIOB33_X105Y133_IOB_X1Y133_I),
.I1(RIOB33_X105Y131_IOB_X1Y132_I),
.I2(CLBLM_R_X3Y143_SLICE_X2Y143_AO6),
.I3(RIOB33_X105Y133_IOB_X1Y134_I),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y141_SLICE_X2Y141_AO5),
.O6(CLBLM_R_X3Y141_SLICE_X2Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000080800000c08)
  ) CLBLM_R_X3Y141_SLICE_X3Y141_DLUT (
.I0(CLBLM_R_X3Y143_SLICE_X2Y143_AO6),
.I1(CLBLM_R_X3Y142_SLICE_X2Y142_AO5),
.I2(CLBLM_R_X3Y139_SLICE_X2Y139_AO5),
.I3(CLBLL_L_X2Y141_SLICE_X1Y141_BO6),
.I4(CLBLM_R_X3Y143_SLICE_X3Y143_BO6),
.I5(CLBLL_L_X2Y141_SLICE_X1Y141_AO6),
.O5(CLBLM_R_X3Y141_SLICE_X3Y141_DO5),
.O6(CLBLM_R_X3Y141_SLICE_X3Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffffef)
  ) CLBLM_R_X3Y141_SLICE_X3Y141_CLUT (
.I0(CLBLL_L_X4Y142_SLICE_X5Y142_AO6),
.I1(CLBLL_L_X4Y141_SLICE_X4Y141_BO6),
.I2(CLBLM_R_X3Y142_SLICE_X3Y142_CO6),
.I3(CLBLM_R_X3Y142_SLICE_X3Y142_DO6),
.I4(CLBLL_L_X4Y140_SLICE_X4Y140_AO6),
.I5(CLBLM_R_X7Y141_SLICE_X9Y141_DO6),
.O5(CLBLM_R_X3Y141_SLICE_X3Y141_CO5),
.O6(CLBLM_R_X3Y141_SLICE_X3Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000001000000000)
  ) CLBLM_R_X3Y141_SLICE_X3Y141_BLUT (
.I0(CLBLM_R_X3Y143_SLICE_X3Y143_BO6),
.I1(CLBLM_R_X3Y141_SLICE_X2Y141_BO6),
.I2(CLBLM_R_X3Y142_SLICE_X2Y142_AO5),
.I3(CLBLM_R_X3Y143_SLICE_X3Y143_CO6),
.I4(CLBLM_R_X3Y141_SLICE_X3Y141_AO6),
.I5(CLBLM_R_X5Y143_SLICE_X6Y143_BO5),
.O5(CLBLM_R_X3Y141_SLICE_X3Y141_BO5),
.O6(CLBLM_R_X3Y141_SLICE_X3Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h20002000ffffafff)
  ) CLBLM_R_X3Y141_SLICE_X3Y141_ALUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(CLBLL_L_X4Y143_SLICE_X5Y143_BO6),
.I2(RIOB33_X105Y133_IOB_X1Y133_I),
.I3(RIOB33_X105Y131_IOB_X1Y132_I),
.I4(RIOB33_X105Y133_IOB_X1Y134_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y141_SLICE_X3Y141_AO5),
.O6(CLBLM_R_X3Y141_SLICE_X3Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000800000000)
  ) CLBLM_R_X3Y142_SLICE_X2Y142_DLUT (
.I0(CLBLM_R_X3Y142_SLICE_X2Y142_AO5),
.I1(CLBLM_R_X3Y142_SLICE_X3Y142_AO5),
.I2(CLBLM_R_X3Y143_SLICE_X3Y143_BO6),
.I3(CLBLM_R_X3Y143_SLICE_X3Y143_CO6),
.I4(CLBLM_R_X3Y141_SLICE_X2Y141_BO6),
.I5(CLBLL_L_X4Y143_SLICE_X4Y143_BO6),
.O5(CLBLM_R_X3Y142_SLICE_X2Y142_DO5),
.O6(CLBLM_R_X3Y142_SLICE_X2Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000004000000)
  ) CLBLM_R_X3Y142_SLICE_X2Y142_CLUT (
.I0(CLBLM_R_X3Y141_SLICE_X2Y141_BO6),
.I1(CLBLM_R_X3Y142_SLICE_X3Y142_AO5),
.I2(CLBLM_R_X3Y143_SLICE_X3Y143_BO6),
.I3(CLBLM_R_X3Y141_SLICE_X2Y141_CO6),
.I4(CLBLL_L_X4Y143_SLICE_X4Y143_BO6),
.I5(CLBLM_R_X3Y142_SLICE_X2Y142_BO6),
.O5(CLBLM_R_X3Y142_SLICE_X2Y142_CO5),
.O6(CLBLM_R_X3Y142_SLICE_X2Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0100000000400000)
  ) CLBLM_R_X3Y142_SLICE_X2Y142_BLUT (
.I0(CLBLL_L_X4Y143_SLICE_X5Y143_BO5),
.I1(RIOB33_X105Y133_IOB_X1Y134_I),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(RIOB33_X105Y131_IOB_X1Y132_I),
.I4(RIOB33_X105Y135_IOB_X1Y136_I),
.I5(RIOB33_X105Y133_IOB_X1Y133_I),
.O5(CLBLM_R_X3Y142_SLICE_X2Y142_BO5),
.O6(CLBLM_R_X3Y142_SLICE_X2Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hefffffffffffefff)
  ) CLBLM_R_X3Y142_SLICE_X2Y142_ALUT (
.I0(CLBLM_R_X3Y143_SLICE_X2Y143_AO5),
.I1(RIOB33_X105Y133_IOB_X1Y134_I),
.I2(RIOB33_X105Y133_IOB_X1Y133_I),
.I3(RIOB33_X105Y131_IOB_X1Y132_I),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y142_SLICE_X2Y142_AO5),
.O6(CLBLM_R_X3Y142_SLICE_X2Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000030000000000)
  ) CLBLM_R_X3Y142_SLICE_X3Y142_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y143_SLICE_X3Y143_CO6),
.I2(CLBLM_R_X3Y141_SLICE_X2Y141_BO6),
.I3(CLBLM_R_X3Y142_SLICE_X3Y142_AO5),
.I4(CLBLM_R_X3Y143_SLICE_X3Y143_BO6),
.I5(CLBLM_R_X3Y142_SLICE_X2Y142_AO5),
.O5(CLBLM_R_X3Y142_SLICE_X3Y142_DO5),
.O6(CLBLM_R_X3Y142_SLICE_X3Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffcfffffffffff)
  ) CLBLM_R_X3Y142_SLICE_X3Y142_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y143_SLICE_X3Y143_CO6),
.I2(CLBLM_R_X5Y143_SLICE_X6Y143_BO5),
.I3(CLBLM_R_X3Y142_SLICE_X3Y142_AO5),
.I4(CLBLM_R_X3Y143_SLICE_X3Y143_BO6),
.I5(CLBLM_R_X3Y142_SLICE_X2Y142_AO5),
.O5(CLBLM_R_X3Y142_SLICE_X3Y142_CO5),
.O6(CLBLM_R_X3Y142_SLICE_X3Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffdffffff)
  ) CLBLM_R_X3Y142_SLICE_X3Y142_BLUT (
.I0(CLBLL_L_X4Y143_SLICE_X5Y143_AO5),
.I1(CLBLM_R_X3Y143_SLICE_X3Y143_BO6),
.I2(CLBLM_R_X3Y141_SLICE_X3Y141_AO6),
.I3(CLBLM_R_X3Y142_SLICE_X2Y142_AO5),
.I4(CLBLL_L_X4Y143_SLICE_X5Y143_AO6),
.I5(CLBLM_R_X3Y143_SLICE_X3Y143_CO6),
.O5(CLBLM_R_X3Y142_SLICE_X3Y142_BO5),
.O6(CLBLM_R_X3Y142_SLICE_X3Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff7fffffff3e7f)
  ) CLBLM_R_X3Y142_SLICE_X3Y142_ALUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(RIOB33_X105Y131_IOB_X1Y132_I),
.I2(RIOB33_X105Y133_IOB_X1Y133_I),
.I3(RIOB33_X105Y133_IOB_X1Y134_I),
.I4(CLBLL_L_X4Y143_SLICE_X5Y143_BO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y142_SLICE_X3Y142_AO5),
.O6(CLBLM_R_X3Y142_SLICE_X3Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y143_SLICE_X2Y143_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y143_SLICE_X2Y143_DO5),
.O6(CLBLM_R_X3Y143_SLICE_X2Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y143_SLICE_X2Y143_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y143_SLICE_X2Y143_CO5),
.O6(CLBLM_R_X3Y143_SLICE_X2Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000c0008080000)
  ) CLBLM_R_X3Y143_SLICE_X2Y143_BLUT (
.I0(LIOB33_X0Y57_IOB_X0Y58_I),
.I1(CLBLL_L_X4Y143_SLICE_X5Y143_CO5),
.I2(CLBLM_R_X3Y143_SLICE_X2Y143_AO6),
.I3(LIOB33_X0Y63_IOB_X0Y63_I),
.I4(RIOB33_X105Y133_IOB_X1Y134_I),
.I5(RIOB33_X105Y133_IOB_X1Y133_I),
.O5(CLBLM_R_X3Y143_SLICE_X2Y143_BO5),
.O6(CLBLM_R_X3Y143_SLICE_X2Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffefffffffffffef)
  ) CLBLM_R_X3Y143_SLICE_X2Y143_ALUT (
.I0(RIOB33_X105Y135_IOB_X1Y136_I),
.I1(RIOB33_X105Y129_IOB_X1Y130_I),
.I2(RIOB33_X105Y137_IOB_X1Y137_I),
.I3(RIOB33_X105Y129_IOB_X1Y129_I),
.I4(RIOB33_X105Y135_IOB_X1Y135_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y143_SLICE_X2Y143_AO5),
.O6(CLBLM_R_X3Y143_SLICE_X2Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf2f1f2f0f0f0f0f0)
  ) CLBLM_R_X3Y143_SLICE_X3Y143_DLUT (
.I0(RIOB33_X105Y131_IOB_X1Y132_I),
.I1(CLBLL_L_X4Y143_SLICE_X5Y143_BO6),
.I2(CLBLM_R_X3Y141_SLICE_X2Y141_BO6),
.I3(RIOB33_X105Y133_IOB_X1Y133_I),
.I4(RIOB33_X105Y133_IOB_X1Y134_I),
.I5(RIOB33_X105Y131_IOB_X1Y131_I),
.O5(CLBLM_R_X3Y143_SLICE_X3Y143_DO5),
.O6(CLBLM_R_X3Y143_SLICE_X3Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccdcdcccccdccccc)
  ) CLBLM_R_X3Y143_SLICE_X3Y143_CLUT (
.I0(CLBLM_R_X3Y143_SLICE_X2Y143_AO6),
.I1(CLBLM_R_X3Y139_SLICE_X2Y139_AO5),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(RIOB33_X105Y133_IOB_X1Y134_I),
.I4(RIOB33_X105Y133_IOB_X1Y133_I),
.I5(RIOB33_X105Y131_IOB_X1Y131_I),
.O5(CLBLM_R_X3Y143_SLICE_X3Y143_CO5),
.O6(CLBLM_R_X3Y143_SLICE_X3Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000d5d008800aa)
  ) CLBLM_R_X3Y143_SLICE_X3Y143_BLUT (
.I0(RIOB33_X105Y133_IOB_X1Y133_I),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(CLBLM_R_X3Y143_SLICE_X2Y143_AO6),
.I3(CLBLM_R_X3Y143_SLICE_X2Y143_AO5),
.I4(RIOB33_X105Y131_IOB_X1Y132_I),
.I5(RIOB33_X105Y133_IOB_X1Y134_I),
.O5(CLBLM_R_X3Y143_SLICE_X3Y143_BO5),
.O6(CLBLM_R_X3Y143_SLICE_X3Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffbfbff7f7ffff)
  ) CLBLM_R_X3Y143_SLICE_X3Y143_ALUT (
.I0(RIOB33_X105Y133_IOB_X1Y133_I),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(RIOB33_X105Y133_IOB_X1Y134_I),
.I3(1'b1),
.I4(RIOB33_X105Y131_IOB_X1Y132_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y143_SLICE_X3Y143_AO5),
.O6(CLBLM_R_X3Y143_SLICE_X3Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y132_SLICE_X6Y132_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y132_SLICE_X6Y132_DO5),
.O6(CLBLM_R_X5Y132_SLICE_X6Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y132_SLICE_X6Y132_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y132_SLICE_X6Y132_CO5),
.O6(CLBLM_R_X5Y132_SLICE_X6Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y132_SLICE_X6Y132_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y132_SLICE_X6Y132_BO5),
.O6(CLBLM_R_X5Y132_SLICE_X6Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff7fffffffffffff)
  ) CLBLM_R_X5Y132_SLICE_X6Y132_ALUT (
.I0(CLBLL_L_X4Y133_SLICE_X4Y133_AQ),
.I1(CLBLM_R_X5Y132_SLICE_X7Y132_DO6),
.I2(CLBLM_R_X7Y132_SLICE_X8Y132_AQ),
.I3(CLBLM_L_X10Y132_SLICE_X12Y132_AO6),
.I4(CLBLM_R_X5Y132_SLICE_X7Y132_AQ),
.I5(CLBLM_R_X7Y132_SLICE_X8Y132_CQ),
.O5(CLBLM_R_X5Y132_SLICE_X6Y132_AO5),
.O6(CLBLM_R_X5Y132_SLICE_X6Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y132_SLICE_X7Y132_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y132_SLICE_X7Y132_AO6),
.Q(CLBLM_R_X5Y132_SLICE_X7Y132_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccddccddccddccdd)
  ) CLBLM_R_X5Y132_SLICE_X7Y132_DLUT (
.I0(CLBLM_R_X5Y136_SLICE_X7Y136_DO6),
.I1(CLBLM_R_X5Y133_SLICE_X7Y133_CO6),
.I2(1'b1),
.I3(CLBLM_R_X7Y133_SLICE_X9Y133_DO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y132_SLICE_X7Y132_DO5),
.O6(CLBLM_R_X5Y132_SLICE_X7Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00002000ffffd5ff)
  ) CLBLM_R_X5Y132_SLICE_X7Y132_CLUT (
.I0(CLBLM_R_X7Y132_SLICE_X8Y132_AQ),
.I1(CLBLM_R_X5Y132_SLICE_X7Y132_AQ),
.I2(CLBLL_L_X4Y133_SLICE_X4Y133_AQ),
.I3(CLBLM_R_X7Y132_SLICE_X8Y132_CQ),
.I4(CLBLM_R_X5Y132_SLICE_X7Y132_DO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y132_SLICE_X7Y132_CO5),
.O6(CLBLM_R_X5Y132_SLICE_X7Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h1300ccffa0000000)
  ) CLBLM_R_X5Y132_SLICE_X7Y132_BLUT (
.I0(CLBLL_L_X4Y133_SLICE_X4Y133_AQ),
.I1(CLBLM_R_X5Y134_SLICE_X7Y134_DO6),
.I2(CLBLM_R_X5Y132_SLICE_X7Y132_AQ),
.I3(CLBLM_R_X7Y132_SLICE_X8Y132_CQ),
.I4(CLBLM_R_X7Y132_SLICE_X8Y132_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y132_SLICE_X7Y132_BO5),
.O6(CLBLM_R_X5Y132_SLICE_X7Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa3300aaaa3000)
  ) CLBLM_R_X5Y132_SLICE_X7Y132_ALUT (
.I0(CLBLM_R_X7Y133_SLICE_X8Y133_AQ),
.I1(CLBLM_R_X11Y138_SLICE_X15Y138_BQ),
.I2(CLBLM_R_X5Y132_SLICE_X7Y132_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X5Y132_SLICE_X7Y132_CO6),
.O5(CLBLM_R_X5Y132_SLICE_X7Y132_AO5),
.O6(CLBLM_R_X5Y132_SLICE_X7Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafafafafafafafa)
  ) CLBLM_R_X5Y133_SLICE_X6Y133_DLUT (
.I0(CLBLM_R_X5Y137_SLICE_X7Y137_C5Q),
.I1(1'b1),
.I2(CLBLM_R_X5Y135_SLICE_X6Y135_DQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y133_SLICE_X6Y133_DO5),
.O6(CLBLM_R_X5Y133_SLICE_X6Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcece0a0affceff0a)
  ) CLBLM_R_X5Y133_SLICE_X6Y133_CLUT (
.I0(CLBLL_L_X4Y141_SLICE_X4Y141_DO6),
.I1(CLBLM_R_X3Y136_SLICE_X3Y136_CQ),
.I2(CLBLM_L_X12Y135_SLICE_X17Y135_CQ),
.I3(CLBLM_R_X3Y140_SLICE_X2Y140_DO6),
.I4(CLBLM_R_X5Y142_SLICE_X6Y142_CO6),
.I5(CLBLM_R_X5Y134_SLICE_X6Y134_CO5),
.O5(CLBLM_R_X5Y133_SLICE_X6Y133_CO5),
.O6(CLBLM_R_X5Y133_SLICE_X6Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffb)
  ) CLBLM_R_X5Y133_SLICE_X6Y133_BLUT (
.I0(CLBLM_L_X8Y140_SLICE_X11Y140_A5Q),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X5Y137_SLICE_X7Y137_B5Q),
.I3(CLBLM_R_X5Y135_SLICE_X6Y135_D5Q),
.I4(CLBLM_R_X5Y133_SLICE_X6Y133_AO6),
.I5(CLBLL_L_X4Y137_SLICE_X4Y137_A5Q),
.O5(CLBLM_R_X5Y133_SLICE_X6Y133_BO5),
.O6(CLBLM_R_X5Y133_SLICE_X6Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffefefffffffe)
  ) CLBLM_R_X5Y133_SLICE_X6Y133_ALUT (
.I0(CLBLM_R_X5Y135_SLICE_X6Y135_DQ),
.I1(CLBLM_R_X5Y136_SLICE_X6Y136_DQ),
.I2(CLBLM_R_X5Y137_SLICE_X7Y137_C5Q),
.I3(CLBLM_R_X5Y135_SLICE_X6Y135_D5Q),
.I4(CLBLM_R_X3Y137_SLICE_X3Y137_BQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y133_SLICE_X6Y133_AO5),
.O6(CLBLM_R_X5Y133_SLICE_X6Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfcfcfcfdfdfdfd)
  ) CLBLM_R_X5Y133_SLICE_X7Y133_DLUT (
.I0(CLBLM_R_X5Y136_SLICE_X7Y136_DO6),
.I1(CLBLM_R_X5Y135_SLICE_X7Y135_A5Q),
.I2(CLBLM_R_X5Y133_SLICE_X6Y133_BO6),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X7Y133_SLICE_X9Y133_DO6),
.O5(CLBLM_R_X5Y133_SLICE_X7Y133_DO5),
.O6(CLBLM_R_X5Y133_SLICE_X7Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffeeffff)
  ) CLBLM_R_X5Y133_SLICE_X7Y133_CLUT (
.I0(CLBLM_R_X5Y137_SLICE_X7Y137_C5Q),
.I1(CLBLL_L_X4Y137_SLICE_X4Y137_A5Q),
.I2(1'b1),
.I3(CLBLM_R_X5Y135_SLICE_X7Y135_A5Q),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X5Y133_SLICE_X7Y133_BO6),
.O5(CLBLM_R_X5Y133_SLICE_X7Y133_CO5),
.O6(CLBLM_R_X5Y133_SLICE_X7Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_R_X5Y133_SLICE_X7Y133_BLUT (
.I0(CLBLM_R_X5Y137_SLICE_X7Y137_B5Q),
.I1(CLBLM_R_X5Y135_SLICE_X6Y135_DQ),
.I2(CLBLM_R_X3Y137_SLICE_X3Y137_BQ),
.I3(CLBLM_R_X5Y135_SLICE_X6Y135_D5Q),
.I4(CLBLM_R_X5Y136_SLICE_X6Y136_DQ),
.I5(CLBLM_L_X8Y140_SLICE_X11Y140_A5Q),
.O5(CLBLM_R_X5Y133_SLICE_X7Y133_BO5),
.O6(CLBLM_R_X5Y133_SLICE_X7Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_R_X5Y133_SLICE_X7Y133_ALUT (
.I0(CLBLM_R_X5Y135_SLICE_X7Y135_A5Q),
.I1(CLBLM_R_X5Y135_SLICE_X6Y135_D5Q),
.I2(CLBLM_R_X3Y137_SLICE_X3Y137_BQ),
.I3(CLBLM_R_X5Y136_SLICE_X6Y136_DQ),
.I4(CLBLM_R_X5Y133_SLICE_X6Y133_DO6),
.I5(CLBLM_R_X5Y134_SLICE_X7Y134_AO6),
.O5(CLBLM_R_X5Y133_SLICE_X7Y133_AO5),
.O6(CLBLM_R_X5Y133_SLICE_X7Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y134_SLICE_X6Y134_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y134_SLICE_X6Y134_BO6),
.Q(CLBLM_R_X5Y134_SLICE_X6Y134_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y134_SLICE_X6Y134_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y134_SLICE_X6Y134_AO6),
.Q(CLBLM_R_X5Y134_SLICE_X6Y134_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haeaaafaaffffffff)
  ) CLBLM_R_X5Y134_SLICE_X6Y134_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y134_SLICE_X8Y134_CQ),
.I2(CLBLM_L_X12Y134_SLICE_X17Y134_AQ),
.I3(CLBLM_L_X10Y145_SLICE_X12Y145_AQ),
.I4(CLBLM_R_X5Y136_SLICE_X6Y136_CQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X5Y134_SLICE_X6Y134_DO5),
.O6(CLBLM_R_X5Y134_SLICE_X6Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa08aaf7f7f7f7)
  ) CLBLM_R_X5Y134_SLICE_X6Y134_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X5Y136_SLICE_X6Y136_CQ),
.I2(CLBLM_R_X7Y134_SLICE_X8Y134_CQ),
.I3(CLBLM_L_X10Y145_SLICE_X12Y145_AQ),
.I4(CLBLM_L_X12Y134_SLICE_X17Y134_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y134_SLICE_X6Y134_CO5),
.O6(CLBLM_R_X5Y134_SLICE_X6Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcd05dc500f0fffff)
  ) CLBLM_R_X5Y134_SLICE_X6Y134_BLUT (
.I0(CLBLM_R_X5Y134_SLICE_X6Y134_DO6),
.I1(CLBLM_R_X5Y137_SLICE_X7Y137_C5Q),
.I2(CLBLM_L_X12Y134_SLICE_X17Y134_AO6),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X5Y134_SLICE_X6Y134_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X5Y134_SLICE_X6Y134_BO5),
.O6(CLBLM_R_X5Y134_SLICE_X6Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaafcfcaaaafcfc)
  ) CLBLM_R_X5Y134_SLICE_X6Y134_ALUT (
.I0(LIOB33_X0Y79_IOB_X0Y79_I),
.I1(CLBLM_L_X10Y145_SLICE_X12Y145_AQ),
.I2(CLBLM_R_X5Y134_SLICE_X6Y134_AQ),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y134_SLICE_X6Y134_AO5),
.O6(CLBLM_R_X5Y134_SLICE_X6Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y134_SLICE_X7Y134_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y134_SLICE_X7Y134_BO6),
.Q(CLBLM_R_X5Y134_SLICE_X7Y134_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y134_SLICE_X7Y134_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y134_SLICE_X7Y134_CO6),
.Q(CLBLM_R_X5Y134_SLICE_X7Y134_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffeffffffff)
  ) CLBLM_R_X5Y134_SLICE_X7Y134_DLUT (
.I0(CLBLM_L_X8Y140_SLICE_X11Y140_A5Q),
.I1(CLBLM_R_X3Y139_SLICE_X3Y139_BO6),
.I2(CLBLM_R_X5Y135_SLICE_X7Y135_A5Q),
.I3(CLBLM_R_X5Y134_SLICE_X7Y134_AO5),
.I4(CLBLM_R_X5Y133_SLICE_X6Y133_AO5),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X5Y134_SLICE_X7Y134_DO5),
.O6(CLBLM_R_X5Y134_SLICE_X7Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0ccf0ccf0aaf0aa)
  ) CLBLM_R_X5Y134_SLICE_X7Y134_CLUT (
.I0(CLBLM_R_X5Y137_SLICE_X7Y137_C5Q),
.I1(CLBLM_R_X5Y134_SLICE_X7Y134_CQ),
.I2(CLBLM_R_X7Y139_SLICE_X8Y139_A5Q),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLL_L_X4Y133_SLICE_X5Y133_BO6),
.O5(CLBLM_R_X5Y134_SLICE_X7Y134_CO5),
.O6(CLBLM_R_X5Y134_SLICE_X7Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf6f00600fcf00c00)
  ) CLBLM_R_X5Y134_SLICE_X7Y134_BLUT (
.I0(CLBLM_R_X5Y136_SLICE_X6Y136_BQ),
.I1(CLBLM_R_X5Y134_SLICE_X7Y134_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y135_SLICE_X8Y135_DO6),
.I4(CLBLM_L_X8Y135_SLICE_X11Y135_AQ),
.I5(CLBLM_R_X5Y135_SLICE_X7Y135_CO6),
.O5(CLBLM_R_X5Y134_SLICE_X7Y134_BO5),
.O6(CLBLM_R_X5Y134_SLICE_X7Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffeeffffffaaaa)
  ) CLBLM_R_X5Y134_SLICE_X7Y134_ALUT (
.I0(CLBLM_R_X5Y137_SLICE_X7Y137_B5Q),
.I1(CLBLM_L_X8Y140_SLICE_X11Y140_A5Q),
.I2(1'b1),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLL_L_X4Y137_SLICE_X4Y137_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X5Y134_SLICE_X7Y134_AO5),
.O6(CLBLM_R_X5Y134_SLICE_X7Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y135_SLICE_X6Y135_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y135_SLICE_X6Y135_DO5),
.Q(CLBLM_R_X5Y135_SLICE_X6Y135_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y135_SLICE_X6Y135_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y135_SLICE_X6Y135_AO6),
.Q(CLBLM_R_X5Y135_SLICE_X6Y135_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y135_SLICE_X6Y135_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y135_SLICE_X6Y135_BO6),
.Q(CLBLM_R_X5Y135_SLICE_X6Y135_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y135_SLICE_X6Y135_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y135_SLICE_X6Y135_CO6),
.Q(CLBLM_R_X5Y135_SLICE_X6Y135_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y135_SLICE_X6Y135_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y135_SLICE_X6Y135_DO6),
.Q(CLBLM_R_X5Y135_SLICE_X6Y135_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0aaaaff00cccc)
  ) CLBLM_R_X5Y135_SLICE_X6Y135_DLUT (
.I0(CLBLM_R_X5Y135_SLICE_X7Y135_AQ),
.I1(CLBLM_R_X5Y136_SLICE_X6Y136_BQ),
.I2(CLBLM_R_X5Y136_SLICE_X6Y136_D5Q),
.I3(CLBLM_R_X5Y139_SLICE_X6Y139_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y135_SLICE_X6Y135_DO5),
.O6(CLBLM_R_X5Y135_SLICE_X6Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5e4e4f5a0e4a0)
  ) CLBLM_R_X5Y135_SLICE_X6Y135_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y135_SLICE_X6Y135_CQ),
.I2(CLBLM_R_X5Y135_SLICE_X6Y135_AQ),
.I3(CLBLM_L_X8Y138_SLICE_X10Y138_AQ),
.I4(CLBLM_R_X7Y135_SLICE_X9Y135_DO6),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_R_X5Y135_SLICE_X6Y135_CO5),
.O6(CLBLM_R_X5Y135_SLICE_X6Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000c030c030)
  ) CLBLM_R_X5Y135_SLICE_X6Y135_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y135_SLICE_X6Y135_BQ),
.I2(CLBLM_R_X5Y134_SLICE_X6Y134_CO6),
.I3(CLBLM_R_X5Y134_SLICE_X6Y134_BO5),
.I4(CLBLM_R_X7Y132_SLICE_X8Y132_BQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X5Y135_SLICE_X6Y135_BO5),
.O6(CLBLM_R_X5Y135_SLICE_X6Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccca050a0a0)
  ) CLBLM_R_X5Y135_SLICE_X6Y135_ALUT (
.I0(CLBLM_R_X5Y135_SLICE_X6Y135_AQ),
.I1(CLBLM_L_X12Y136_SLICE_X17Y136_AQ),
.I2(CLBLM_R_X5Y134_SLICE_X6Y134_CO6),
.I3(CLBLM_R_X5Y134_SLICE_X6Y134_BO5),
.I4(CLBLM_R_X5Y135_SLICE_X6Y135_BQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X5Y135_SLICE_X6Y135_AO5),
.O6(CLBLM_R_X5Y135_SLICE_X6Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y135_SLICE_X7Y135_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y135_SLICE_X7Y135_BO6),
.Q(CLBLM_R_X5Y135_SLICE_X7Y135_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y135_SLICE_X7Y135_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y135_SLICE_X7Y135_AO6),
.Q(CLBLM_R_X5Y135_SLICE_X7Y135_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_R_X5Y135_SLICE_X7Y135_DLUT (
.I0(CLBLM_R_X5Y137_SLICE_X7Y137_AQ),
.I1(CLBLM_R_X7Y135_SLICE_X8Y135_BQ),
.I2(CLBLM_R_X5Y134_SLICE_X7Y134_BQ),
.I3(CLBLM_R_X5Y136_SLICE_X6Y136_BQ),
.I4(CLBLM_R_X5Y135_SLICE_X7Y135_AQ),
.I5(CLBLM_R_X7Y134_SLICE_X8Y134_BQ),
.O5(CLBLM_R_X5Y135_SLICE_X7Y135_DO5),
.O6(CLBLM_R_X5Y135_SLICE_X7Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h88000000115533ff)
  ) CLBLM_R_X5Y135_SLICE_X7Y135_CLUT (
.I0(CLBLM_R_X5Y137_SLICE_X7Y137_AQ),
.I1(CLBLM_R_X7Y135_SLICE_X8Y135_BQ),
.I2(1'b1),
.I3(CLBLM_R_X7Y134_SLICE_X8Y134_BQ),
.I4(CLBLM_R_X5Y135_SLICE_X7Y135_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y135_SLICE_X7Y135_CO5),
.O6(CLBLM_R_X5Y135_SLICE_X7Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hafafa0a0cc000000)
  ) CLBLM_R_X5Y135_SLICE_X7Y135_BLUT (
.I0(CLBLM_L_X8Y134_SLICE_X11Y134_DQ),
.I1(CLBLM_R_X7Y135_SLICE_X8Y135_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y134_SLICE_X8Y134_BQ),
.I4(CLBLM_R_X5Y137_SLICE_X7Y137_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y135_SLICE_X7Y135_BO5),
.O6(CLBLM_R_X5Y135_SLICE_X7Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff484800004848)
  ) CLBLM_R_X5Y135_SLICE_X7Y135_ALUT (
.I0(CLBLM_R_X5Y135_SLICE_X7Y135_BO5),
.I1(CLBLM_R_X7Y135_SLICE_X8Y135_DO6),
.I2(CLBLM_R_X5Y135_SLICE_X7Y135_AQ),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y139_SLICE_X9Y139_AQ),
.O5(CLBLM_R_X5Y135_SLICE_X7Y135_AO5),
.O6(CLBLM_R_X5Y135_SLICE_X7Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y136_SLICE_X6Y136_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y136_SLICE_X6Y136_DO5),
.Q(CLBLM_R_X5Y136_SLICE_X6Y136_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y136_SLICE_X6Y136_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y136_SLICE_X6Y136_AO6),
.Q(CLBLM_R_X5Y136_SLICE_X6Y136_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y136_SLICE_X6Y136_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y136_SLICE_X6Y136_BO6),
.Q(CLBLM_R_X5Y136_SLICE_X6Y136_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y136_SLICE_X6Y136_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y136_SLICE_X6Y136_CO6),
.Q(CLBLM_R_X5Y136_SLICE_X6Y136_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y136_SLICE_X6Y136_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y136_SLICE_X6Y136_DO6),
.Q(CLBLM_R_X5Y136_SLICE_X6Y136_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff33cc00b8b8b8b8)
  ) CLBLM_R_X5Y136_SLICE_X6Y136_DLUT (
.I0(CLBLL_L_X4Y136_SLICE_X5Y136_BQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(RIOB33_X105Y127_IOB_X1Y127_I),
.I3(CLBLM_L_X10Y138_SLICE_X13Y138_CQ),
.I4(CLBLM_R_X5Y137_SLICE_X6Y137_CQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y136_SLICE_X6Y136_DO5),
.O6(CLBLM_R_X5Y136_SLICE_X6Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f08800f0f00000)
  ) CLBLM_R_X5Y136_SLICE_X6Y136_CLUT (
.I0(CLBLM_R_X5Y135_SLICE_X6Y135_BQ),
.I1(CLBLM_R_X5Y135_SLICE_X6Y135_AQ),
.I2(CLBLM_R_X7Y139_SLICE_X9Y139_A5Q),
.I3(CLBLM_R_X5Y134_SLICE_X6Y134_A5Q),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLL_L_X4Y138_SLICE_X5Y138_A5Q),
.O5(CLBLM_R_X5Y136_SLICE_X6Y136_CO5),
.O6(CLBLM_R_X5Y136_SLICE_X6Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hbeaabeaa3c003c00)
  ) CLBLM_R_X5Y136_SLICE_X6Y136_BLUT (
.I0(CLBLM_R_X5Y141_SLICE_X6Y141_CQ),
.I1(CLBLM_R_X5Y136_SLICE_X6Y136_BQ),
.I2(CLBLM_R_X5Y135_SLICE_X7Y135_CO6),
.I3(CLBLM_R_X7Y135_SLICE_X8Y135_DO5),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X5Y136_SLICE_X6Y136_BO5),
.O6(CLBLM_R_X5Y136_SLICE_X6Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfaeefaee50445044)
  ) CLBLM_R_X5Y136_SLICE_X6Y136_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y138_SLICE_X6Y138_CQ),
.I2(CLBLM_R_X5Y136_SLICE_X6Y136_AQ),
.I3(CLBLM_L_X8Y143_SLICE_X10Y143_DO5),
.I4(1'b1),
.I5(CLBLL_L_X4Y135_SLICE_X5Y135_CQ),
.O5(CLBLM_R_X5Y136_SLICE_X6Y136_AO5),
.O6(CLBLM_R_X5Y136_SLICE_X6Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y136_SLICE_X7Y136_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y136_SLICE_X7Y136_AO6),
.Q(CLBLM_R_X5Y136_SLICE_X7Y136_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y136_SLICE_X7Y136_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y136_SLICE_X7Y136_BO6),
.Q(CLBLM_R_X5Y136_SLICE_X7Y136_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y136_SLICE_X7Y136_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y136_SLICE_X7Y136_CO6),
.Q(CLBLM_R_X5Y136_SLICE_X7Y136_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffaaaa69969669)
  ) CLBLM_R_X5Y136_SLICE_X7Y136_DLUT (
.I0(CLBLM_R_X5Y140_SLICE_X6Y140_AO6),
.I1(CLBLL_L_X4Y139_SLICE_X4Y139_BO6),
.I2(CLBLM_R_X3Y137_SLICE_X3Y137_DO6),
.I3(CLBLM_R_X3Y140_SLICE_X2Y140_DO6),
.I4(CLBLM_R_X5Y141_SLICE_X7Y141_DO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y136_SLICE_X7Y136_DO5),
.O6(CLBLM_R_X5Y136_SLICE_X7Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f000eef0f0eeee)
  ) CLBLM_R_X5Y136_SLICE_X7Y136_CLUT (
.I0(CLBLM_R_X7Y139_SLICE_X8Y139_AQ),
.I1(CLBLM_R_X5Y136_SLICE_X7Y136_CQ),
.I2(CLBLM_R_X7Y134_SLICE_X8Y134_CQ),
.I3(CLBLM_L_X10Y139_SLICE_X13Y139_B5Q),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X12Y134_SLICE_X17Y134_AO6),
.O5(CLBLM_R_X5Y136_SLICE_X7Y136_CO5),
.O6(CLBLM_R_X5Y136_SLICE_X7Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa00cc0000)
  ) CLBLM_R_X5Y136_SLICE_X7Y136_BLUT (
.I0(CLBLM_R_X3Y137_SLICE_X2Y137_BQ),
.I1(CLBLM_R_X5Y136_SLICE_X7Y136_BQ),
.I2(1'b1),
.I3(CLBLM_R_X7Y139_SLICE_X9Y139_AQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X5Y136_SLICE_X7Y136_BO5),
.O6(CLBLM_R_X5Y136_SLICE_X7Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbeaafaaa3c00f000)
  ) CLBLM_R_X5Y136_SLICE_X7Y136_ALUT (
.I0(CLBLM_R_X7Y138_SLICE_X8Y138_CQ),
.I1(CLBLM_R_X5Y135_SLICE_X7Y135_DO6),
.I2(CLBLM_R_X5Y136_SLICE_X7Y136_AQ),
.I3(CLBLM_R_X7Y135_SLICE_X8Y135_DO5),
.I4(CLBLM_R_X5Y137_SLICE_X6Y137_CQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X5Y136_SLICE_X7Y136_AO5),
.O6(CLBLM_R_X5Y136_SLICE_X7Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y137_SLICE_X6Y137_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y137_SLICE_X6Y137_AO6),
.Q(CLBLM_R_X5Y137_SLICE_X6Y137_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y137_SLICE_X6Y137_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y137_SLICE_X6Y137_BO6),
.Q(CLBLM_R_X5Y137_SLICE_X6Y137_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y137_SLICE_X6Y137_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y137_SLICE_X6Y137_CO6),
.Q(CLBLM_R_X5Y137_SLICE_X6Y137_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h1333333320000000)
  ) CLBLM_R_X5Y137_SLICE_X6Y137_DLUT (
.I0(CLBLM_R_X5Y135_SLICE_X6Y135_BQ),
.I1(CLBLM_R_X5Y134_SLICE_X6Y134_DO6),
.I2(CLBLM_R_X5Y135_SLICE_X6Y135_AQ),
.I3(CLBLM_R_X5Y134_SLICE_X6Y134_A5Q),
.I4(CLBLM_L_X12Y134_SLICE_X17Y134_AO6),
.I5(CLBLL_L_X4Y138_SLICE_X5Y138_A5Q),
.O5(CLBLM_R_X5Y137_SLICE_X6Y137_DO5),
.O6(CLBLM_R_X5Y137_SLICE_X6Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hbeaa3c00beaa3c00)
  ) CLBLM_R_X5Y137_SLICE_X6Y137_CLUT (
.I0(CLBLM_R_X7Y143_SLICE_X8Y143_AQ),
.I1(CLBLM_R_X5Y137_SLICE_X6Y137_CQ),
.I2(CLBLM_R_X5Y135_SLICE_X7Y135_DO6),
.I3(CLBLM_R_X7Y135_SLICE_X8Y135_DO5),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y137_SLICE_X6Y137_CO5),
.O6(CLBLM_R_X5Y137_SLICE_X6Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'heccc2000cccc0000)
  ) CLBLM_R_X5Y137_SLICE_X6Y137_BLUT (
.I0(CLBLM_R_X7Y143_SLICE_X8Y143_A5Q),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLL_L_X4Y136_SLICE_X5Y136_CQ),
.I3(CLBLM_R_X7Y133_SLICE_X8Y133_CQ),
.I4(CLBLM_L_X8Y134_SLICE_X10Y134_AQ),
.I5(CLBLM_R_X3Y138_SLICE_X3Y138_AQ),
.O5(CLBLM_R_X5Y137_SLICE_X6Y137_BO5),
.O6(CLBLM_R_X5Y137_SLICE_X6Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00f7f78080)
  ) CLBLM_R_X5Y137_SLICE_X6Y137_ALUT (
.I0(CLBLL_L_X4Y137_SLICE_X4Y137_CQ),
.I1(CLBLM_L_X12Y135_SLICE_X17Y135_AQ),
.I2(CLBLM_R_X5Y137_SLICE_X6Y137_AQ),
.I3(CLBLM_R_X5Y137_SLICE_X6Y137_CQ),
.I4(CLBLM_L_X8Y138_SLICE_X10Y138_BQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X5Y137_SLICE_X6Y137_AO5),
.O6(CLBLM_R_X5Y137_SLICE_X6Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y137_SLICE_X7Y137_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y137_SLICE_X7Y137_BO5),
.Q(CLBLM_R_X5Y137_SLICE_X7Y137_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y137_SLICE_X7Y137_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y137_SLICE_X7Y137_CO5),
.Q(CLBLM_R_X5Y137_SLICE_X7Y137_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y137_SLICE_X7Y137_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y137_SLICE_X7Y137_AO6),
.Q(CLBLM_R_X5Y137_SLICE_X7Y137_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y137_SLICE_X7Y137_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y137_SLICE_X7Y137_BO6),
.Q(CLBLM_R_X5Y137_SLICE_X7Y137_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y137_SLICE_X7Y137_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y137_SLICE_X7Y137_CO6),
.Q(CLBLM_R_X5Y137_SLICE_X7Y137_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff1f3fffff5fff)
  ) CLBLM_R_X5Y137_SLICE_X7Y137_DLUT (
.I0(CLBLM_R_X5Y136_SLICE_X7Y136_AQ),
.I1(CLBLM_R_X5Y134_SLICE_X7Y134_BQ),
.I2(CLBLL_L_X4Y137_SLICE_X4Y137_BQ),
.I3(CLBLM_R_X5Y137_SLICE_X6Y137_CQ),
.I4(CLBLM_R_X5Y135_SLICE_X7Y135_CO5),
.I5(CLBLM_R_X5Y136_SLICE_X6Y136_BQ),
.O5(CLBLM_R_X5Y137_SLICE_X7Y137_DO5),
.O6(CLBLM_R_X5Y137_SLICE_X7Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hbaba1010ff55aa00)
  ) CLBLM_R_X5Y137_SLICE_X7Y137_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_L_X8Y139_SLICE_X11Y139_BQ),
.I3(CLBLM_R_X5Y138_SLICE_X7Y138_BQ),
.I4(CLBLM_R_X5Y134_SLICE_X7Y134_BQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y137_SLICE_X7Y137_CO5),
.O6(CLBLM_R_X5Y137_SLICE_X7Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f04444ccccff00)
  ) CLBLM_R_X5Y137_SLICE_X7Y137_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X5Y137_SLICE_X7Y137_BQ),
.I2(CLBLM_R_X7Y142_SLICE_X8Y142_AQ),
.I3(CLBLM_R_X5Y136_SLICE_X7Y136_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y137_SLICE_X7Y137_BO5),
.O6(CLBLM_R_X5Y137_SLICE_X7Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdecc5a00fcccf000)
  ) CLBLM_R_X5Y137_SLICE_X7Y137_ALUT (
.I0(CLBLM_R_X7Y134_SLICE_X8Y134_BQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X5Y137_SLICE_X7Y137_AQ),
.I3(CLBLM_R_X7Y135_SLICE_X8Y135_DO5),
.I4(CLBLM_R_X5Y137_SLICE_X6Y137_AQ),
.I5(CLBLM_R_X7Y135_SLICE_X8Y135_BQ),
.O5(CLBLM_R_X5Y137_SLICE_X7Y137_AO5),
.O6(CLBLM_R_X5Y137_SLICE_X7Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y138_SLICE_X6Y138_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y138_SLICE_X6Y138_AO6),
.Q(CLBLM_R_X5Y138_SLICE_X6Y138_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y138_SLICE_X6Y138_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y138_SLICE_X6Y138_BO6),
.Q(CLBLM_R_X5Y138_SLICE_X6Y138_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y138_SLICE_X6Y138_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y138_SLICE_X6Y138_CO6),
.Q(CLBLM_R_X5Y138_SLICE_X6Y138_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5f5f55550f0f0000)
  ) CLBLM_R_X5Y138_SLICE_X6Y138_DLUT (
.I0(CLBLM_R_X7Y142_SLICE_X9Y142_CO6),
.I1(1'b1),
.I2(CLBLL_L_X4Y143_SLICE_X4Y143_BO5),
.I3(1'b1),
.I4(CLBLM_R_X7Y137_SLICE_X9Y137_AQ),
.I5(CLBLM_L_X12Y136_SLICE_X17Y136_AQ),
.O5(CLBLM_R_X5Y138_SLICE_X6Y138_DO5),
.O6(CLBLM_R_X5Y138_SLICE_X6Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5f0f005050000)
  ) CLBLM_R_X5Y138_SLICE_X6Y138_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(1'b1),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(CLBLM_L_X10Y134_SLICE_X13Y134_BQ),
.I5(CLBLM_R_X5Y138_SLICE_X6Y138_AQ),
.O5(CLBLM_R_X5Y138_SLICE_X6Y138_CO5),
.O6(CLBLM_R_X5Y138_SLICE_X6Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccf5f5cccc0000)
  ) CLBLM_R_X5Y138_SLICE_X6Y138_BLUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLL_L_X4Y138_SLICE_X5Y138_A5Q),
.I2(CLBLM_L_X8Y138_SLICE_X10Y138_AQ),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X5Y138_SLICE_X6Y138_BQ),
.O5(CLBLM_R_X5Y138_SLICE_X6Y138_BO5),
.O6(CLBLM_R_X5Y138_SLICE_X6Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffa500000fa50)
  ) CLBLM_R_X5Y138_SLICE_X6Y138_ALUT (
.I0(CLBLM_L_X8Y143_SLICE_X10Y143_DO5),
.I1(1'b1),
.I2(CLBLM_R_X5Y138_SLICE_X6Y138_AQ),
.I3(CLBLM_L_X10Y137_SLICE_X13Y137_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X11Y138_SLICE_X15Y138_CQ),
.O5(CLBLM_R_X5Y138_SLICE_X6Y138_AO5),
.O6(CLBLM_R_X5Y138_SLICE_X6Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y138_SLICE_X7Y138_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y138_SLICE_X7Y138_AO6),
.Q(CLBLM_R_X5Y138_SLICE_X7Y138_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y138_SLICE_X7Y138_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y138_SLICE_X7Y138_BO6),
.Q(CLBLM_R_X5Y138_SLICE_X7Y138_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y138_SLICE_X7Y138_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y138_SLICE_X7Y138_CO6),
.Q(CLBLM_R_X5Y138_SLICE_X7Y138_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ff00aaaaffaa)
  ) CLBLM_R_X5Y138_SLICE_X7Y138_DLUT (
.I0(CLBLM_R_X5Y137_SLICE_X6Y137_AQ),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X11Y134_SLICE_X15Y134_AQ),
.I4(CLBLM_R_X5Y143_SLICE_X6Y143_AO5),
.I5(CLBLL_L_X4Y143_SLICE_X5Y143_AO5),
.O5(CLBLM_R_X5Y138_SLICE_X7Y138_DO5),
.O6(CLBLM_R_X5Y138_SLICE_X7Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f05500f0f0cccc)
  ) CLBLM_R_X5Y138_SLICE_X7Y138_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X5Y138_SLICE_X7Y138_CQ),
.I2(CLBLM_L_X12Y138_SLICE_X16Y138_CQ),
.I3(CLBLL_L_X4Y142_SLICE_X5Y142_DO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLL_L_X4Y138_SLICE_X5Y138_CO5),
.O5(CLBLM_R_X5Y138_SLICE_X7Y138_CO5),
.O6(CLBLM_R_X5Y138_SLICE_X7Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdf8fff00d080f00)
  ) CLBLM_R_X5Y138_SLICE_X7Y138_BLUT (
.I0(CLBLM_L_X10Y139_SLICE_X13Y139_B5Q),
.I1(CLBLM_R_X5Y138_SLICE_X7Y138_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I4(CLBLM_L_X12Y134_SLICE_X17Y134_AO6),
.I5(CLBLM_R_X7Y143_SLICE_X8Y143_A5Q),
.O5(CLBLM_R_X5Y138_SLICE_X7Y138_BO5),
.O6(CLBLM_R_X5Y138_SLICE_X7Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffccccccffc0c0c0)
  ) CLBLM_R_X5Y138_SLICE_X7Y138_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y144_SLICE_X9Y144_BO6),
.I2(CLBLM_R_X5Y138_SLICE_X7Y138_AQ),
.I3(CLBLM_L_X8Y137_SLICE_X10Y137_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y134_SLICE_X8Y134_AQ),
.O5(CLBLM_R_X5Y138_SLICE_X7Y138_AO5),
.O6(CLBLM_R_X5Y138_SLICE_X7Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y139_SLICE_X6Y139_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y139_SLICE_X6Y139_AO6),
.Q(CLBLM_R_X5Y139_SLICE_X6Y139_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y139_SLICE_X6Y139_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y139_SLICE_X6Y139_BO6),
.Q(CLBLM_R_X5Y139_SLICE_X6Y139_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00ba30aaaababa)
  ) CLBLM_R_X5Y139_SLICE_X6Y139_DLUT (
.I0(CLBLL_L_X4Y137_SLICE_X4Y137_AQ),
.I1(CLBLM_R_X3Y143_SLICE_X2Y143_AO6),
.I2(CLBLM_R_X5Y134_SLICE_X7Y134_CQ),
.I3(RIOB33_X105Y129_IOB_X1Y129_I),
.I4(CLBLL_L_X2Y140_SLICE_X1Y140_AO6),
.I5(RIOB33_X105Y137_IOB_X1Y137_I),
.O5(CLBLM_R_X5Y139_SLICE_X6Y139_DO5),
.O6(CLBLM_R_X5Y139_SLICE_X6Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h000a00ce000a000a)
  ) CLBLM_R_X5Y139_SLICE_X6Y139_CLUT (
.I0(CLBLM_L_X8Y137_SLICE_X10Y137_AQ),
.I1(CLBLM_R_X7Y137_SLICE_X8Y137_BQ),
.I2(CLBLL_L_X2Y140_SLICE_X1Y140_AO6),
.I3(CLBLM_R_X3Y143_SLICE_X2Y143_AO5),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(CLBLL_L_X2Y141_SLICE_X1Y141_AO6),
.O5(CLBLM_R_X5Y139_SLICE_X6Y139_CO5),
.O6(CLBLM_R_X5Y139_SLICE_X6Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f000eef0f0eeee)
  ) CLBLM_R_X5Y139_SLICE_X6Y139_BLUT (
.I0(CLBLM_L_X8Y142_SLICE_X10Y142_DQ),
.I1(CLBLM_R_X5Y139_SLICE_X6Y139_BQ),
.I2(CLBLM_R_X7Y131_SLICE_X9Y131_AQ),
.I3(CLBLM_L_X12Y134_SLICE_X17Y134_AO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X10Y139_SLICE_X13Y139_B5Q),
.O5(CLBLM_R_X5Y139_SLICE_X6Y139_BO5),
.O6(CLBLM_R_X5Y139_SLICE_X6Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00f5f5ff00a0a0)
  ) CLBLM_R_X5Y139_SLICE_X6Y139_ALUT (
.I0(CLBLM_L_X8Y143_SLICE_X10Y143_DO6),
.I1(1'b1),
.I2(CLBLM_R_X5Y139_SLICE_X6Y139_AQ),
.I3(CLBLM_R_X5Y134_SLICE_X6Y134_A5Q),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.O5(CLBLM_R_X5Y139_SLICE_X6Y139_AO5),
.O6(CLBLM_R_X5Y139_SLICE_X6Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y139_SLICE_X7Y139_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y139_SLICE_X7Y139_AO6),
.Q(CLBLM_R_X5Y139_SLICE_X7Y139_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y139_SLICE_X7Y139_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y139_SLICE_X7Y139_BO6),
.Q(CLBLM_R_X5Y139_SLICE_X7Y139_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y139_SLICE_X7Y139_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y139_SLICE_X7Y139_CO6),
.Q(CLBLM_R_X5Y139_SLICE_X7Y139_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0ace0ace0ace0ace)
  ) CLBLM_R_X5Y139_SLICE_X7Y139_DLUT (
.I0(CLBLM_R_X5Y139_SLICE_X6Y139_AQ),
.I1(CLBLM_R_X5Y139_SLICE_X7Y139_CQ),
.I2(CLBLM_R_X5Y143_SLICE_X6Y143_AO5),
.I3(CLBLM_R_X3Y142_SLICE_X3Y142_AO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y139_SLICE_X7Y139_DO5),
.O6(CLBLM_R_X5Y139_SLICE_X7Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0afa0acacacac)
  ) CLBLM_R_X5Y139_SLICE_X7Y139_CLUT (
.I0(CLBLM_R_X7Y134_SLICE_X9Y134_AQ),
.I1(CLBLM_R_X5Y139_SLICE_X7Y139_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLL_L_X4Y139_SLICE_X4Y139_BO6),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLL_L_X4Y138_SLICE_X5Y138_CO5),
.O5(CLBLM_R_X5Y139_SLICE_X7Y139_CO5),
.O6(CLBLM_R_X5Y139_SLICE_X7Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0afafa0a0)
  ) CLBLM_R_X5Y139_SLICE_X7Y139_BLUT (
.I0(CLBLM_R_X5Y139_SLICE_X7Y139_CQ),
.I1(1'b1),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(CLBLM_L_X10Y137_SLICE_X13Y137_BQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X5Y139_SLICE_X7Y139_BO5),
.O6(CLBLM_R_X5Y139_SLICE_X7Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff050005ff500050)
  ) CLBLM_R_X5Y139_SLICE_X7Y139_ALUT (
.I0(CLBLM_R_X11Y135_SLICE_X14Y135_AQ),
.I1(1'b1),
.I2(CLBLM_R_X5Y139_SLICE_X7Y139_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X5Y139_SLICE_X6Y139_AQ),
.I5(CLBLM_R_X7Y139_SLICE_X8Y139_DO6),
.O5(CLBLM_R_X5Y139_SLICE_X7Y139_AO5),
.O6(CLBLM_R_X5Y139_SLICE_X7Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff2222ffffff22)
  ) CLBLM_R_X5Y140_SLICE_X6Y140_DLUT (
.I0(CLBLM_L_X8Y140_SLICE_X11Y140_BQ),
.I1(CLBLL_L_X4Y143_SLICE_X5Y143_AO6),
.I2(1'b1),
.I3(CLBLM_R_X7Y143_SLICE_X8Y143_A5Q),
.I4(CLBLM_R_X5Y141_SLICE_X6Y141_DO6),
.I5(CLBLM_R_X3Y141_SLICE_X2Y141_AO5),
.O5(CLBLM_R_X5Y140_SLICE_X6Y140_DO5),
.O6(CLBLM_R_X5Y140_SLICE_X6Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0c0caeaeff0cffae)
  ) CLBLM_R_X5Y140_SLICE_X6Y140_CLUT (
.I0(CLBLM_L_X8Y141_SLICE_X11Y141_AQ),
.I1(CLBLM_R_X7Y133_SLICE_X8Y133_CQ),
.I2(CLBLM_R_X3Y141_SLICE_X2Y141_AO5),
.I3(RIOB33_X105Y109_IOB_X1Y109_I),
.I4(CLBLM_R_X3Y142_SLICE_X2Y142_AO5),
.I5(CLBLM_R_X5Y143_SLICE_X6Y143_BO6),
.O5(CLBLM_R_X5Y140_SLICE_X6Y140_CO5),
.O6(CLBLM_R_X5Y140_SLICE_X6Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffcfffffffe)
  ) CLBLM_R_X5Y140_SLICE_X6Y140_BLUT (
.I0(CLBLM_R_X5Y141_SLICE_X6Y141_CQ),
.I1(CLBLM_R_X3Y143_SLICE_X2Y143_BO6),
.I2(CLBLM_R_X5Y139_SLICE_X6Y139_DO6),
.I3(CLBLM_R_X7Y141_SLICE_X9Y141_CO6),
.I4(CLBLM_R_X3Y140_SLICE_X3Y140_CO6),
.I5(CLBLM_R_X5Y143_SLICE_X6Y143_AO6),
.O5(CLBLM_R_X5Y140_SLICE_X6Y140_BO5),
.O6(CLBLM_R_X5Y140_SLICE_X6Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_R_X5Y140_SLICE_X6Y140_ALUT (
.I0(CLBLM_R_X5Y140_SLICE_X6Y140_DO6),
.I1(CLBLM_R_X5Y138_SLICE_X6Y138_DO6),
.I2(CLBLM_R_X5Y140_SLICE_X7Y140_CO6),
.I3(CLBLM_R_X3Y142_SLICE_X2Y142_CO6),
.I4(CLBLM_R_X3Y139_SLICE_X2Y139_CO6),
.I5(CLBLM_R_X7Y140_SLICE_X9Y140_DO6),
.O5(CLBLM_R_X5Y140_SLICE_X6Y140_AO5),
.O6(CLBLM_R_X5Y140_SLICE_X6Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y140_SLICE_X7Y140_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y140_SLICE_X7Y140_AO6),
.Q(CLBLM_R_X5Y140_SLICE_X7Y140_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y140_SLICE_X7Y140_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y140_SLICE_X7Y140_BO6),
.Q(CLBLM_R_X5Y140_SLICE_X7Y140_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcecececeffceffce)
  ) CLBLM_R_X5Y140_SLICE_X7Y140_DLUT (
.I0(CLBLM_R_X5Y141_SLICE_X7Y141_AQ),
.I1(CLBLL_L_X4Y137_SLICE_X5Y137_CO6),
.I2(CLBLM_R_X5Y143_SLICE_X6Y143_AO5),
.I3(CLBLM_L_X8Y142_SLICE_X10Y142_BQ),
.I4(1'b1),
.I5(CLBLM_R_X7Y142_SLICE_X9Y142_CO5),
.O5(CLBLM_R_X5Y140_SLICE_X7Y140_DO5),
.O6(CLBLM_R_X5Y140_SLICE_X7Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0aceffff0ace0ace)
  ) CLBLM_R_X5Y140_SLICE_X7Y140_CLUT (
.I0(CLBLM_R_X5Y135_SLICE_X6Y135_AQ),
.I1(CLBLM_L_X8Y140_SLICE_X10Y140_CQ),
.I2(CLBLM_R_X5Y143_SLICE_X6Y143_BO5),
.I3(CLBLM_R_X5Y143_SLICE_X6Y143_AO6),
.I4(CLBLM_R_X3Y142_SLICE_X2Y142_AO5),
.I5(CLBLM_L_X10Y144_SLICE_X12Y144_AQ),
.O5(CLBLM_R_X5Y140_SLICE_X7Y140_CO5),
.O6(CLBLM_R_X5Y140_SLICE_X7Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccf0f0cccc0000)
  ) CLBLM_R_X5Y140_SLICE_X7Y140_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y141_SLICE_X6Y141_AQ),
.I2(CLBLM_R_X11Y138_SLICE_X15Y138_CQ),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X5Y140_SLICE_X7Y140_BO5),
.O6(CLBLM_R_X5Y140_SLICE_X7Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaf0ffaaaaf000)
  ) CLBLM_R_X5Y140_SLICE_X7Y140_ALUT (
.I0(CLBLM_R_X5Y136_SLICE_X6Y136_AQ),
.I1(1'b1),
.I2(CLBLM_L_X8Y138_SLICE_X10Y138_CQ),
.I3(CLBLM_L_X8Y143_SLICE_X10Y143_DO5),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X5Y140_SLICE_X7Y140_AQ),
.O5(CLBLM_R_X5Y140_SLICE_X7Y140_AO5),
.O6(CLBLM_R_X5Y140_SLICE_X7Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y141_SLICE_X6Y141_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y141_SLICE_X11Y141_DO6),
.Q(CLBLM_R_X5Y141_SLICE_X6Y141_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y141_SLICE_X6Y141_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y141_SLICE_X6Y141_AO6),
.Q(CLBLM_R_X5Y141_SLICE_X6Y141_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y141_SLICE_X6Y141_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y141_SLICE_X6Y141_BO6),
.Q(CLBLM_R_X5Y141_SLICE_X6Y141_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y141_SLICE_X6Y141_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y141_SLICE_X6Y141_CO6),
.Q(CLBLM_R_X5Y141_SLICE_X6Y141_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000c0c05000500)
  ) CLBLM_R_X5Y141_SLICE_X6Y141_DLUT (
.I0(CLBLL_L_X2Y140_SLICE_X1Y140_AO6),
.I1(RIOB33_X105Y107_IOB_X1Y108_I),
.I2(CLBLL_L_X4Y143_SLICE_X5Y143_BO5),
.I3(CLBLM_L_X8Y142_SLICE_X10Y142_CQ),
.I4(CLBLM_R_X3Y143_SLICE_X3Y143_AO5),
.I5(RIOB33_X105Y135_IOB_X1Y136_I),
.O5(CLBLM_R_X5Y141_SLICE_X6Y141_DO5),
.O6(CLBLM_R_X5Y141_SLICE_X6Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0eef0eef044f044)
  ) CLBLM_R_X5Y141_SLICE_X6Y141_CLUT (
.I0(CLBLM_L_X8Y143_SLICE_X10Y143_DO5),
.I1(CLBLM_R_X5Y141_SLICE_X6Y141_CQ),
.I2(CLBLM_R_X5Y141_SLICE_X6Y141_BQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLM_R_X7Y135_SLICE_X8Y135_CQ),
.O5(CLBLM_R_X5Y141_SLICE_X6Y141_CO5),
.O6(CLBLM_R_X5Y141_SLICE_X6Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcff0c0ffcf00c00)
  ) CLBLM_R_X5Y141_SLICE_X6Y141_BLUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y138_SLICE_X5Y138_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y143_SLICE_X10Y143_DO5),
.I4(CLBLM_R_X5Y141_SLICE_X7Y141_AQ),
.I5(CLBLM_R_X5Y141_SLICE_X6Y141_BQ),
.O5(CLBLM_R_X5Y141_SLICE_X6Y141_BO5),
.O6(CLBLM_R_X5Y141_SLICE_X6Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000f780f780)
  ) CLBLM_R_X5Y141_SLICE_X6Y141_ALUT (
.I0(CLBLL_L_X4Y137_SLICE_X4Y137_CQ),
.I1(CLBLM_L_X12Y135_SLICE_X17Y135_AQ),
.I2(CLBLM_R_X5Y141_SLICE_X6Y141_AQ),
.I3(CLBLM_R_X7Y137_SLICE_X8Y137_CQ),
.I4(CLBLL_L_X4Y135_SLICE_X4Y135_BQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X5Y141_SLICE_X6Y141_AO5),
.O6(CLBLM_R_X5Y141_SLICE_X6Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y141_SLICE_X7Y141_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y141_SLICE_X7Y141_AO6),
.Q(CLBLM_R_X5Y141_SLICE_X7Y141_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y141_SLICE_X7Y141_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y141_SLICE_X7Y141_BO6),
.Q(CLBLM_R_X5Y141_SLICE_X7Y141_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_R_X5Y141_SLICE_X7Y141_DLUT (
.I0(CLBLM_R_X5Y143_SLICE_X7Y143_CO6),
.I1(CLBLM_R_X7Y142_SLICE_X8Y142_DO6),
.I2(CLBLM_R_X5Y143_SLICE_X6Y143_DO6),
.I3(CLBLL_L_X2Y141_SLICE_X1Y141_DO6),
.I4(CLBLM_R_X5Y138_SLICE_X7Y138_DO6),
.I5(CLBLM_R_X3Y142_SLICE_X2Y142_CO6),
.O5(CLBLM_R_X5Y141_SLICE_X7Y141_DO5),
.O6(CLBLM_R_X5Y141_SLICE_X7Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000ace000000cc)
  ) CLBLM_R_X5Y141_SLICE_X7Y141_CLUT (
.I0(CLBLM_R_X7Y135_SLICE_X9Y135_BQ),
.I1(CLBLM_R_X7Y140_SLICE_X9Y140_CQ),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(CLBLM_R_X3Y143_SLICE_X3Y143_AO6),
.I4(CLBLM_R_X3Y143_SLICE_X2Y143_AO5),
.I5(CLBLL_L_X2Y141_SLICE_X1Y141_AO6),
.O5(CLBLM_R_X5Y141_SLICE_X7Y141_CO5),
.O6(CLBLM_R_X5Y141_SLICE_X7Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefe0e0ef0f00000)
  ) CLBLM_R_X5Y141_SLICE_X7Y141_BLUT (
.I0(CLBLM_L_X8Y140_SLICE_X11Y140_A5Q),
.I1(CLBLM_R_X5Y141_SLICE_X7Y141_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(CLBLM_R_X7Y135_SLICE_X9Y135_BQ),
.I5(CLBLL_L_X4Y133_SLICE_X5Y133_BO6),
.O5(CLBLM_R_X5Y141_SLICE_X7Y141_BO5),
.O6(CLBLM_R_X5Y141_SLICE_X7Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000fa50fa50)
  ) CLBLM_R_X5Y141_SLICE_X7Y141_ALUT (
.I0(CLBLM_L_X8Y143_SLICE_X10Y143_DO6),
.I1(1'b1),
.I2(CLBLM_R_X5Y141_SLICE_X7Y141_AQ),
.I3(CLBLM_R_X11Y139_SLICE_X15Y139_DQ),
.I4(CLBLM_R_X5Y137_SLICE_X7Y137_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X5Y141_SLICE_X7Y141_AO5),
.O6(CLBLM_R_X5Y141_SLICE_X7Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccfcccfceefeeefe)
  ) CLBLM_R_X5Y142_SLICE_X6Y142_DLUT (
.I0(CLBLM_R_X5Y141_SLICE_X7Y141_BQ),
.I1(CLBLL_L_X4Y141_SLICE_X5Y141_BO6),
.I2(CLBLM_R_X5Y141_SLICE_X6Y141_AQ),
.I3(CLBLM_R_X3Y142_SLICE_X3Y142_AO6),
.I4(1'b1),
.I5(CLBLL_L_X4Y143_SLICE_X4Y143_AO6),
.O5(CLBLM_R_X5Y142_SLICE_X6Y142_DO5),
.O6(CLBLM_R_X5Y142_SLICE_X6Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffff5fdfffff0fc)
  ) CLBLM_R_X5Y142_SLICE_X6Y142_CLUT (
.I0(CLBLM_R_X5Y143_SLICE_X6Y143_AO5),
.I1(CLBLM_R_X3Y141_SLICE_X3Y141_DO6),
.I2(CLBLM_R_X5Y142_SLICE_X7Y142_DO6),
.I3(CLBLM_R_X3Y143_SLICE_X3Y143_DO6),
.I4(CLBLM_R_X5Y142_SLICE_X6Y142_DO6),
.I5(CLBLM_L_X8Y140_SLICE_X10Y140_BQ),
.O5(CLBLM_R_X5Y142_SLICE_X6Y142_CO5),
.O6(CLBLM_R_X5Y142_SLICE_X6Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f3f0f0f2f3f2f2)
  ) CLBLM_R_X5Y142_SLICE_X6Y142_BLUT (
.I0(LIOB33_X0Y67_IOB_X0Y68_I),
.I1(CLBLM_R_X3Y143_SLICE_X2Y143_AO6),
.I2(CLBLL_L_X4Y138_SLICE_X5Y138_DO5),
.I3(CLBLM_R_X3Y143_SLICE_X3Y143_AO6),
.I4(CLBLM_R_X5Y141_SLICE_X7Y141_BQ),
.I5(CLBLM_R_X3Y143_SLICE_X3Y143_AO5),
.O5(CLBLM_R_X5Y142_SLICE_X6Y142_BO5),
.O6(CLBLM_R_X5Y142_SLICE_X6Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffefffefffffffe)
  ) CLBLM_R_X5Y142_SLICE_X6Y142_ALUT (
.I0(CLBLM_R_X5Y142_SLICE_X7Y142_CO6),
.I1(CLBLM_R_X5Y142_SLICE_X7Y142_BO6),
.I2(CLBLM_R_X5Y142_SLICE_X7Y142_AO6),
.I3(CLBLM_R_X5Y142_SLICE_X6Y142_BO6),
.I4(CLBLM_R_X5Y141_SLICE_X6Y141_AQ),
.I5(CLBLM_R_X3Y142_SLICE_X3Y142_AO6),
.O5(CLBLM_R_X5Y142_SLICE_X6Y142_AO5),
.O6(CLBLM_R_X5Y142_SLICE_X6Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff33ffbbff00ffaa)
  ) CLBLM_R_X5Y142_SLICE_X7Y142_DLUT (
.I0(CLBLM_R_X7Y134_SLICE_X9Y134_BQ),
.I1(CLBLM_R_X5Y143_SLICE_X6Y143_AO6),
.I2(1'b1),
.I3(CLBLM_R_X5Y142_SLICE_X7Y142_CO6),
.I4(CLBLM_R_X5Y143_SLICE_X6Y143_BO5),
.I5(CLBLM_R_X7Y143_SLICE_X9Y143_CQ),
.O5(CLBLM_R_X5Y142_SLICE_X7Y142_DO5),
.O6(CLBLM_R_X5Y142_SLICE_X7Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000cc000000f0)
  ) CLBLM_R_X5Y142_SLICE_X7Y142_CLUT (
.I0(1'b1),
.I1(RIOB33_X105Y113_IOB_X1Y113_I),
.I2(CLBLM_R_X5Y140_SLICE_X7Y140_AQ),
.I3(CLBLM_R_X3Y143_SLICE_X3Y143_AO5),
.I4(CLBLL_L_X4Y143_SLICE_X5Y143_BO5),
.I5(RIOB33_X105Y135_IOB_X1Y136_I),
.O5(CLBLM_R_X5Y142_SLICE_X7Y142_CO5),
.O6(CLBLM_R_X5Y142_SLICE_X7Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000054540404)
  ) CLBLM_R_X5Y142_SLICE_X7Y142_BLUT (
.I0(CLBLL_L_X4Y143_SLICE_X5Y143_BO5),
.I1(CLBLM_R_X7Y143_SLICE_X9Y143_CQ),
.I2(RIOB33_X105Y135_IOB_X1Y136_I),
.I3(1'b1),
.I4(CLBLM_R_X7Y134_SLICE_X9Y134_BQ),
.I5(CLBLM_R_X3Y143_SLICE_X3Y143_AO6),
.O5(CLBLM_R_X5Y142_SLICE_X7Y142_BO5),
.O6(CLBLM_R_X5Y142_SLICE_X7Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000800)
  ) CLBLM_R_X5Y142_SLICE_X7Y142_ALUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(CLBLM_L_X8Y140_SLICE_X10Y140_BQ),
.I2(CLBLM_R_X3Y143_SLICE_X2Y143_AO5),
.I3(RIOB33_X105Y133_IOB_X1Y133_I),
.I4(RIOB33_X105Y133_IOB_X1Y134_I),
.I5(RIOB33_X105Y131_IOB_X1Y132_I),
.O5(CLBLM_R_X5Y142_SLICE_X7Y142_AO5),
.O6(CLBLM_R_X5Y142_SLICE_X7Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffcfffe)
  ) CLBLM_R_X5Y143_SLICE_X6Y143_DLUT (
.I0(CLBLM_R_X5Y135_SLICE_X6Y135_BQ),
.I1(CLBLM_R_X5Y139_SLICE_X6Y139_CO6),
.I2(CLBLM_R_X5Y143_SLICE_X7Y143_DO6),
.I3(CLBLM_R_X5Y143_SLICE_X6Y143_CO6),
.I4(CLBLM_R_X5Y143_SLICE_X6Y143_BO5),
.I5(CLBLL_L_X4Y143_SLICE_X5Y143_DO6),
.O5(CLBLM_R_X5Y143_SLICE_X6Y143_DO5),
.O6(CLBLM_R_X5Y143_SLICE_X6Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000030002020000)
  ) CLBLM_R_X5Y143_SLICE_X6Y143_CLUT (
.I0(CLBLM_L_X10Y141_SLICE_X13Y141_CQ),
.I1(CLBLL_L_X2Y141_SLICE_X1Y141_AO5),
.I2(CLBLL_L_X4Y143_SLICE_X5Y143_BO5),
.I3(CLBLM_L_X8Y143_SLICE_X10Y143_BQ),
.I4(RIOB33_X105Y135_IOB_X1Y136_I),
.I5(RIOB33_X105Y131_IOB_X1Y131_I),
.O5(CLBLM_R_X5Y143_SLICE_X6Y143_CO5),
.O6(CLBLM_R_X5Y143_SLICE_X6Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffff7fffffdffff)
  ) CLBLM_R_X5Y143_SLICE_X6Y143_BLUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(RIOB33_X105Y131_IOB_X1Y132_I),
.I2(CLBLL_L_X4Y143_SLICE_X5Y143_BO6),
.I3(RIOB33_X105Y133_IOB_X1Y133_I),
.I4(RIOB33_X105Y133_IOB_X1Y134_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y143_SLICE_X6Y143_BO5),
.O6(CLBLM_R_X5Y143_SLICE_X6Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffdfffffffffdff)
  ) CLBLM_R_X5Y143_SLICE_X6Y143_ALUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(RIOB33_X105Y131_IOB_X1Y132_I),
.I2(CLBLM_R_X3Y143_SLICE_X2Y143_AO5),
.I3(RIOB33_X105Y133_IOB_X1Y133_I),
.I4(RIOB33_X105Y133_IOB_X1Y134_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y143_SLICE_X6Y143_AO5),
.O6(CLBLM_R_X5Y143_SLICE_X6Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000af000000a0)
  ) CLBLM_R_X5Y143_SLICE_X7Y143_DLUT (
.I0(RIOB33_X105Y107_IOB_X1Y107_I),
.I1(1'b1),
.I2(RIOB33_X105Y135_IOB_X1Y136_I),
.I3(CLBLM_R_X3Y143_SLICE_X3Y143_AO5),
.I4(CLBLL_L_X4Y143_SLICE_X5Y143_BO5),
.I5(CLBLL_L_X4Y138_SLICE_X4Y138_BQ),
.O5(CLBLM_R_X5Y143_SLICE_X7Y143_DO5),
.O6(CLBLM_R_X5Y143_SLICE_X7Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h73507350ffff7350)
  ) CLBLM_R_X5Y143_SLICE_X7Y143_CLUT (
.I0(CLBLM_R_X5Y143_SLICE_X7Y143_AO6),
.I1(CLBLL_L_X4Y143_SLICE_X4Y143_AO6),
.I2(RIOB33_X105Y115_IOB_X1Y115_I),
.I3(CLBLL_L_X4Y134_SLICE_X5Y134_CQ),
.I4(CLBLM_R_X7Y143_SLICE_X8Y143_CQ),
.I5(CLBLL_L_X4Y143_SLICE_X4Y143_AO5),
.O5(CLBLM_R_X5Y143_SLICE_X7Y143_CO5),
.O6(CLBLM_R_X5Y143_SLICE_X7Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h22f2ffff22f222f2)
  ) CLBLM_R_X5Y143_SLICE_X7Y143_BLUT (
.I0(CLBLL_L_X4Y134_SLICE_X5Y134_AQ),
.I1(CLBLL_L_X4Y143_SLICE_X4Y143_AO6),
.I2(CLBLM_R_X7Y142_SLICE_X8Y142_AQ),
.I3(CLBLL_L_X4Y143_SLICE_X4Y143_AO5),
.I4(CLBLM_R_X5Y143_SLICE_X7Y143_AO6),
.I5(RIOB33_X105Y113_IOB_X1Y114_I),
.O5(CLBLM_R_X5Y143_SLICE_X7Y143_BO5),
.O6(CLBLM_R_X5Y143_SLICE_X7Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfeffffffffffffff)
  ) CLBLM_R_X5Y143_SLICE_X7Y143_ALUT (
.I0(CLBLL_L_X4Y143_SLICE_X5Y143_BO5),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(RIOB33_X105Y133_IOB_X1Y134_I),
.I3(RIOB33_X105Y131_IOB_X1Y132_I),
.I4(RIOB33_X105Y135_IOB_X1Y136_I),
.I5(RIOB33_X105Y133_IOB_X1Y133_I),
.O5(CLBLM_R_X5Y143_SLICE_X7Y143_AO5),
.O6(CLBLM_R_X5Y143_SLICE_X7Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y131_SLICE_X8Y131_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y131_SLICE_X8Y131_DO5),
.O6(CLBLM_R_X7Y131_SLICE_X8Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y131_SLICE_X8Y131_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y131_SLICE_X8Y131_CO5),
.O6(CLBLM_R_X7Y131_SLICE_X8Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y131_SLICE_X8Y131_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y131_SLICE_X8Y131_BO5),
.O6(CLBLM_R_X7Y131_SLICE_X8Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y131_SLICE_X8Y131_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y131_SLICE_X8Y131_AO5),
.O6(CLBLM_R_X7Y131_SLICE_X8Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y131_SLICE_X9Y131_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y131_SLICE_X9Y131_AO6),
.Q(CLBLM_R_X7Y131_SLICE_X9Y131_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y131_SLICE_X9Y131_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y131_SLICE_X9Y131_BO6),
.Q(CLBLM_R_X7Y131_SLICE_X9Y131_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y131_SLICE_X9Y131_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y131_SLICE_X9Y131_DO5),
.O6(CLBLM_R_X7Y131_SLICE_X9Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y131_SLICE_X9Y131_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y131_SLICE_X9Y131_CO5),
.O6(CLBLM_R_X7Y131_SLICE_X9Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0fefe00000e0e)
  ) CLBLM_R_X7Y131_SLICE_X9Y131_BLUT (
.I0(CLBLM_L_X8Y131_SLICE_X10Y131_A5Q),
.I1(CLBLM_R_X7Y131_SLICE_X9Y131_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(CLBLM_R_X5Y134_SLICE_X7Y134_DO6),
.I5(CLBLM_R_X5Y136_SLICE_X6Y136_CQ),
.O5(CLBLM_R_X7Y131_SLICE_X9Y131_BO5),
.O6(CLBLM_R_X7Y131_SLICE_X9Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdcc310055005500)
  ) CLBLM_R_X7Y131_SLICE_X9Y131_ALUT (
.I0(RIOB33_X105Y141_IOB_X1Y142_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X7Y131_SLICE_X9Y131_AQ),
.I3(CLBLM_R_X11Y139_SLICE_X15Y139_A5Q),
.I4(CLBLM_L_X8Y131_SLICE_X11Y131_BQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y131_SLICE_X9Y131_AO5),
.O6(CLBLM_R_X7Y131_SLICE_X9Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y132_SLICE_X8Y132_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y132_SLICE_X8Y132_AO6),
.Q(CLBLM_R_X7Y132_SLICE_X8Y132_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y132_SLICE_X8Y132_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y132_SLICE_X8Y132_BO6),
.Q(CLBLM_R_X7Y132_SLICE_X8Y132_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y132_SLICE_X8Y132_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y132_SLICE_X8Y132_CO6),
.Q(CLBLM_R_X7Y132_SLICE_X8Y132_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y132_SLICE_X8Y132_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y132_SLICE_X8Y132_DO5),
.O6(CLBLM_R_X7Y132_SLICE_X8Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaee00ccaafb00f3)
  ) CLBLM_R_X7Y132_SLICE_X8Y132_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y132_SLICE_X8Y132_CQ),
.I2(CLBLM_R_X5Y132_SLICE_X7Y132_BO5),
.I3(CLBLM_R_X7Y132_SLICE_X8Y132_AO5),
.I4(CLBLM_R_X7Y144_SLICE_X8Y144_AQ),
.I5(CLBLM_R_X5Y132_SLICE_X7Y132_DO6),
.O5(CLBLM_R_X7Y132_SLICE_X8Y132_CO5),
.O6(CLBLM_R_X7Y132_SLICE_X8Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f04444f0f04444)
  ) CLBLM_R_X7Y132_SLICE_X8Y132_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X7Y132_SLICE_X8Y132_BQ),
.I2(CLBLM_R_X7Y134_SLICE_X8Y134_C5Q),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y132_SLICE_X8Y132_BO5),
.O6(CLBLM_R_X7Y132_SLICE_X8Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00022ffffff55)
  ) CLBLM_R_X7Y132_SLICE_X8Y132_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X5Y132_SLICE_X7Y132_BO6),
.I2(CLBLM_L_X8Y133_SLICE_X11Y133_AQ),
.I3(CLBLM_R_X11Y138_SLICE_X15Y138_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y132_SLICE_X8Y132_AO5),
.O6(CLBLM_R_X7Y132_SLICE_X8Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y132_SLICE_X9Y132_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y132_SLICE_X9Y132_DO5),
.Q(CLBLM_R_X7Y132_SLICE_X9Y132_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y132_SLICE_X9Y132_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y132_SLICE_X9Y132_AO6),
.Q(CLBLM_R_X7Y132_SLICE_X9Y132_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y132_SLICE_X9Y132_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y132_SLICE_X9Y132_BO6),
.Q(CLBLM_R_X7Y132_SLICE_X9Y132_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y132_SLICE_X9Y132_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y132_SLICE_X9Y132_CO6),
.Q(CLBLM_R_X7Y132_SLICE_X9Y132_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y132_SLICE_X9Y132_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y132_SLICE_X9Y132_DO6),
.Q(CLBLM_R_X7Y132_SLICE_X9Y132_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd88dd88f5a0f5a0)
  ) CLBLM_R_X7Y132_SLICE_X9Y132_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y132_SLICE_X10Y132_BQ),
.I2(CLBLM_R_X7Y137_SLICE_X8Y137_BQ),
.I3(RIOB33_X105Y101_IOB_X1Y101_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y132_SLICE_X9Y132_DO5),
.O6(CLBLM_R_X7Y132_SLICE_X9Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000aaaaf0c0)
  ) CLBLM_R_X7Y132_SLICE_X9Y132_CLUT (
.I0(CLBLL_L_X4Y134_SLICE_X4Y134_B5Q),
.I1(CLBLM_R_X7Y132_SLICE_X9Y132_CQ),
.I2(CLBLM_L_X8Y138_SLICE_X10Y138_AQ),
.I3(CLBLM_L_X12Y132_SLICE_X16Y132_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_R_X7Y132_SLICE_X9Y132_CO5),
.O6(CLBLM_R_X7Y132_SLICE_X9Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hafafafa0acacaca0)
  ) CLBLM_R_X7Y132_SLICE_X9Y132_BLUT (
.I0(CLBLM_R_X5Y135_SLICE_X6Y135_DQ),
.I1(CLBLM_R_X7Y132_SLICE_X9Y132_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_L_X8Y138_SLICE_X10Y138_AQ),
.I5(CLBLM_L_X8Y132_SLICE_X10Y132_BQ),
.O5(CLBLM_R_X7Y132_SLICE_X9Y132_BO5),
.O6(CLBLM_R_X7Y132_SLICE_X9Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hacafa0a0acafafaf)
  ) CLBLM_R_X7Y132_SLICE_X9Y132_ALUT (
.I0(CLBLM_L_X12Y132_SLICE_X16Y132_CQ),
.I1(CLBLL_L_X4Y135_SLICE_X4Y135_A5Q),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X5Y137_SLICE_X6Y137_BQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(LIOB33_X0Y53_IOB_X0Y53_I),
.O5(CLBLM_R_X7Y132_SLICE_X9Y132_AO5),
.O6(CLBLM_R_X7Y132_SLICE_X9Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y133_SLICE_X8Y133_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y133_SLICE_X8Y133_AO6),
.Q(CLBLM_R_X7Y133_SLICE_X8Y133_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y133_SLICE_X8Y133_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y133_SLICE_X8Y133_BO6),
.Q(CLBLM_R_X7Y133_SLICE_X8Y133_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y133_SLICE_X8Y133_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y133_SLICE_X8Y133_CO6),
.Q(CLBLM_R_X7Y133_SLICE_X8Y133_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'habaaffffababffff)
  ) CLBLM_R_X7Y133_SLICE_X8Y133_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(LIOB33_X0Y53_IOB_X0Y53_I),
.I2(CLBLM_R_X7Y135_SLICE_X9Y135_B5Q),
.I3(CLBLL_L_X4Y135_SLICE_X4Y135_A5Q),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X5Y137_SLICE_X6Y137_BQ),
.O5(CLBLM_R_X7Y133_SLICE_X8Y133_DO5),
.O6(CLBLM_R_X7Y133_SLICE_X8Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0fcfc0000cccc)
  ) CLBLM_R_X7Y133_SLICE_X8Y133_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y133_SLICE_X8Y133_CQ),
.I2(CLBLM_R_X11Y131_SLICE_X15Y131_BQ),
.I3(1'b1),
.I4(CLBLM_R_X7Y133_SLICE_X8Y133_DO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X7Y133_SLICE_X8Y133_CO5),
.O6(CLBLM_R_X7Y133_SLICE_X8Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff030003ff300030)
  ) CLBLM_R_X7Y133_SLICE_X8Y133_BLUT (
.I0(1'b1),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X7Y135_SLICE_X8Y135_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y133_SLICE_X9Y133_AQ),
.I5(CLBLM_L_X8Y139_SLICE_X11Y139_DO6),
.O5(CLBLM_R_X7Y133_SLICE_X8Y133_BO5),
.O6(CLBLM_R_X7Y133_SLICE_X8Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00fefe1010)
  ) CLBLM_R_X7Y133_SLICE_X8Y133_ALUT (
.I0(CLBLM_L_X8Y138_SLICE_X10Y138_AQ),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_R_X7Y133_SLICE_X8Y133_AQ),
.I3(CLBLM_R_X7Y134_SLICE_X9Y134_BQ),
.I4(CLBLM_L_X8Y139_SLICE_X11Y139_DO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X7Y133_SLICE_X8Y133_AO5),
.O6(CLBLM_R_X7Y133_SLICE_X8Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y133_SLICE_X9Y133_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y133_SLICE_X9Y133_AO6),
.Q(CLBLM_R_X7Y133_SLICE_X9Y133_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y133_SLICE_X9Y133_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y133_SLICE_X9Y133_BO6),
.Q(CLBLM_R_X7Y133_SLICE_X9Y133_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y133_SLICE_X9Y133_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y133_SLICE_X9Y133_CO6),
.Q(CLBLM_R_X7Y133_SLICE_X9Y133_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_R_X7Y133_SLICE_X9Y133_DLUT (
.I0(CLBLL_L_X4Y141_SLICE_X4Y141_DO6),
.I1(CLBLM_R_X3Y140_SLICE_X2Y140_DO6),
.I2(CLBLL_L_X4Y142_SLICE_X4Y142_BO6),
.I3(CLBLL_L_X4Y142_SLICE_X5Y142_DO6),
.I4(CLBLM_R_X5Y142_SLICE_X6Y142_CO6),
.I5(CLBLL_L_X4Y139_SLICE_X4Y139_BO6),
.O5(CLBLM_R_X7Y133_SLICE_X9Y133_DO5),
.O6(CLBLM_R_X7Y133_SLICE_X9Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffff0f0fcf8fcf8)
  ) CLBLM_R_X7Y133_SLICE_X9Y133_CLUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_R_X7Y133_SLICE_X9Y133_CQ),
.I2(CLBLM_R_X7Y134_SLICE_X9Y134_CO6),
.I3(CLBLM_L_X8Y138_SLICE_X10Y138_AQ),
.I4(CLBLL_L_X4Y133_SLICE_X5Y133_A5Q),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X7Y133_SLICE_X9Y133_CO5),
.O6(CLBLM_R_X7Y133_SLICE_X9Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0afa0aca0a0a0a0)
  ) CLBLM_R_X7Y133_SLICE_X9Y133_BLUT (
.I0(CLBLL_L_X4Y137_SLICE_X4Y137_A5Q),
.I1(CLBLM_R_X7Y133_SLICE_X9Y133_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_L_X10Y133_SLICE_X13Y133_BQ),
.I5(CLBLM_L_X8Y138_SLICE_X10Y138_AQ),
.O5(CLBLM_R_X7Y133_SLICE_X9Y133_BO5),
.O6(CLBLM_R_X7Y133_SLICE_X9Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hee44ee44ee44fa50)
  ) CLBLM_R_X7Y133_SLICE_X9Y133_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y133_SLICE_X9Y133_BQ),
.I2(CLBLM_R_X7Y133_SLICE_X9Y133_AQ),
.I3(CLBLM_R_X5Y134_SLICE_X7Y134_CQ),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLM_L_X8Y138_SLICE_X10Y138_AQ),
.O5(CLBLM_R_X7Y133_SLICE_X9Y133_AO5),
.O6(CLBLM_R_X7Y133_SLICE_X9Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y134_SLICE_X8Y134_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y134_SLICE_X8Y134_CO5),
.Q(CLBLM_R_X7Y134_SLICE_X8Y134_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y134_SLICE_X8Y134_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y134_SLICE_X8Y134_AO6),
.Q(CLBLM_R_X7Y134_SLICE_X8Y134_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y134_SLICE_X8Y134_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y134_SLICE_X8Y134_BO6),
.Q(CLBLM_R_X7Y134_SLICE_X8Y134_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y134_SLICE_X8Y134_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y134_SLICE_X8Y134_CO6),
.Q(CLBLM_R_X7Y134_SLICE_X8Y134_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5040f0c0afaf0f0f)
  ) CLBLM_R_X7Y134_SLICE_X8Y134_DLUT (
.I0(CLBLM_R_X7Y133_SLICE_X8Y133_AQ),
.I1(CLBLM_L_X10Y134_SLICE_X12Y134_CQ),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLL_L_X4Y134_SLICE_X4Y134_AQ),
.I4(CLBLM_R_X7Y139_SLICE_X8Y139_BQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y134_SLICE_X8Y134_DO5),
.O6(CLBLM_R_X7Y134_SLICE_X8Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'he4e4e4e4fafa5050)
  ) CLBLM_R_X7Y134_SLICE_X8Y134_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y136_SLICE_X6Y136_CQ),
.I2(CLBLM_L_X8Y134_SLICE_X10Y134_A5Q),
.I3(1'b1),
.I4(CLBLM_R_X7Y137_SLICE_X8Y137_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y134_SLICE_X8Y134_CO5),
.O6(CLBLM_R_X7Y134_SLICE_X8Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3fcffff030c0f0f)
  ) CLBLM_R_X7Y134_SLICE_X8Y134_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y134_SLICE_X8Y134_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y135_SLICE_X8Y135_BQ),
.I4(CLBLM_R_X7Y135_SLICE_X8Y135_DO6),
.I5(CLBLM_R_X13Y134_SLICE_X19Y134_CQ),
.O5(CLBLM_R_X7Y134_SLICE_X8Y134_BO5),
.O6(CLBLM_R_X7Y134_SLICE_X8Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f30003f3f00300)
  ) CLBLM_R_X7Y134_SLICE_X8Y134_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y134_SLICE_X8Y134_DO5),
.I4(CLBLM_R_X7Y135_SLICE_X9Y135_B5Q),
.I5(CLBLM_R_X7Y134_SLICE_X9Y134_AQ),
.O5(CLBLM_R_X7Y134_SLICE_X8Y134_AO5),
.O6(CLBLM_R_X7Y134_SLICE_X8Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y134_SLICE_X9Y134_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y134_SLICE_X9Y134_AO6),
.Q(CLBLM_R_X7Y134_SLICE_X9Y134_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y134_SLICE_X9Y134_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y134_SLICE_X9Y134_BO6),
.Q(CLBLM_R_X7Y134_SLICE_X9Y134_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffefefffe)
  ) CLBLM_R_X7Y134_SLICE_X9Y134_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y138_SLICE_X10Y138_AQ),
.I2(RIOB33_X105Y117_IOB_X1Y118_I),
.I3(CLBLM_L_X10Y134_SLICE_X12Y134_CQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLL_L_X4Y134_SLICE_X4Y134_AQ),
.O5(CLBLM_R_X7Y134_SLICE_X9Y134_DO5),
.O6(CLBLM_R_X7Y134_SLICE_X9Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ffff00008f00)
  ) CLBLM_R_X7Y134_SLICE_X9Y134_CLUT (
.I0(CLBLM_R_X7Y133_SLICE_X8Y133_AQ),
.I1(CLBLM_R_X7Y139_SLICE_X8Y139_BQ),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLM_R_X5Y140_SLICE_X6Y140_AO6),
.I4(CLBLM_R_X7Y134_SLICE_X9Y134_DO6),
.I5(CLBLM_L_X8Y137_SLICE_X11Y137_CO5),
.O5(CLBLM_R_X7Y134_SLICE_X9Y134_CO5),
.O6(CLBLM_R_X7Y134_SLICE_X9Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ddfff0f08800)
  ) CLBLM_R_X7Y134_SLICE_X9Y134_BLUT (
.I0(CLBLM_L_X10Y139_SLICE_X13Y139_B5Q),
.I1(CLBLM_R_X7Y134_SLICE_X9Y134_BQ),
.I2(CLBLM_R_X13Y134_SLICE_X19Y134_AQ),
.I3(CLBLM_L_X12Y134_SLICE_X17Y134_AO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y137_SLICE_X8Y137_CQ),
.O5(CLBLM_R_X7Y134_SLICE_X9Y134_BO5),
.O6(CLBLM_R_X7Y134_SLICE_X9Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff11ff4400110044)
  ) CLBLM_R_X7Y134_SLICE_X9Y134_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X7Y135_SLICE_X9Y135_CO5),
.I2(1'b1),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y138_SLICE_X9Y138_AQ),
.I5(CLBLM_R_X7Y132_SLICE_X9Y132_CQ),
.O5(CLBLM_R_X7Y134_SLICE_X9Y134_AO5),
.O6(CLBLM_R_X7Y134_SLICE_X9Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y135_SLICE_X8Y135_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y135_SLICE_X8Y135_AO6),
.Q(CLBLM_R_X7Y135_SLICE_X8Y135_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y135_SLICE_X8Y135_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y135_SLICE_X8Y135_BO6),
.Q(CLBLM_R_X7Y135_SLICE_X8Y135_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y135_SLICE_X8Y135_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y135_SLICE_X8Y135_CO6),
.Q(CLBLM_R_X7Y135_SLICE_X8Y135_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hc000c00040004000)
  ) CLBLM_R_X7Y135_SLICE_X8Y135_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X11Y139_SLICE_X15Y139_A5Q),
.I2(CLBLM_L_X10Y135_SLICE_X12Y135_B5Q),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y135_SLICE_X8Y135_DO5),
.O6(CLBLM_R_X7Y135_SLICE_X8Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0f5a0a0a0f5a0a0)
  ) CLBLM_R_X7Y135_SLICE_X8Y135_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(1'b1),
.I2(CLBLM_L_X10Y135_SLICE_X12Y135_B5Q),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLL_L_X4Y136_SLICE_X4Y136_DQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y135_SLICE_X8Y135_CO5),
.O6(CLBLM_R_X7Y135_SLICE_X8Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf7ff070fffff0f0f)
  ) CLBLM_R_X7Y135_SLICE_X8Y135_BLUT (
.I0(CLBLM_L_X10Y135_SLICE_X12Y135_B5Q),
.I1(CLBLM_R_X7Y135_SLICE_X8Y135_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X11Y139_SLICE_X15Y139_A5Q),
.I4(CLBLM_R_X7Y136_SLICE_X8Y136_AQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X7Y135_SLICE_X8Y135_BO5),
.O6(CLBLM_R_X7Y135_SLICE_X8Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f30003f0fc000c)
  ) CLBLM_R_X7Y135_SLICE_X8Y135_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y137_SLICE_X13Y137_CO6),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X5Y135_SLICE_X7Y135_AQ),
.I5(CLBLM_L_X8Y136_SLICE_X11Y136_CQ),
.O5(CLBLM_R_X7Y135_SLICE_X8Y135_AO5),
.O6(CLBLM_R_X7Y135_SLICE_X8Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y135_SLICE_X9Y135_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y134_SLICE_X10Y134_BO5),
.Q(CLBLM_R_X7Y135_SLICE_X9Y135_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y135_SLICE_X9Y135_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y136_SLICE_X9Y136_BO6),
.Q(CLBLM_R_X7Y135_SLICE_X9Y135_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y135_SLICE_X9Y135_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y135_SLICE_X9Y135_AO6),
.Q(CLBLM_R_X7Y135_SLICE_X9Y135_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y135_SLICE_X9Y135_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y135_SLICE_X9Y135_BO6),
.Q(CLBLM_R_X7Y135_SLICE_X9Y135_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa0af909fa0af909)
  ) CLBLM_R_X7Y135_SLICE_X9Y135_DLUT (
.I0(CLBLM_R_X7Y132_SLICE_X8Y132_BQ),
.I1(CLBLM_L_X10Y138_SLICE_X12Y138_BO5),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLM_R_X5Y137_SLICE_X7Y137_CQ),
.I4(CLBLM_R_X5Y136_SLICE_X7Y136_BQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y135_SLICE_X9Y135_DO5),
.O6(CLBLM_R_X7Y135_SLICE_X9Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f000cacacaca)
  ) CLBLM_R_X7Y135_SLICE_X9Y135_CLUT (
.I0(CLBLM_L_X8Y135_SLICE_X10Y135_AQ),
.I1(CLBLM_R_X11Y136_SLICE_X15Y136_BQ),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLM_R_X5Y135_SLICE_X6Y135_CQ),
.I4(CLBLM_L_X8Y135_SLICE_X11Y135_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X7Y135_SLICE_X9Y135_CO5),
.O6(CLBLM_R_X7Y135_SLICE_X9Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0ff000fc0cfc0c)
  ) CLBLM_R_X7Y135_SLICE_X9Y135_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y135_SLICE_X9Y135_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y135_SLICE_X11Y135_CQ),
.I4(CLBLM_L_X8Y136_SLICE_X11Y136_AQ),
.I5(CLBLM_L_X8Y143_SLICE_X10Y143_DO5),
.O5(CLBLM_R_X7Y135_SLICE_X9Y135_BO5),
.O6(CLBLM_R_X7Y135_SLICE_X9Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccaaaaccccf0f0)
  ) CLBLM_R_X7Y135_SLICE_X9Y135_ALUT (
.I0(CLBLL_L_X4Y135_SLICE_X5Y135_BQ),
.I1(CLBLM_L_X8Y133_SLICE_X10Y133_CQ),
.I2(CLBLM_R_X7Y135_SLICE_X9Y135_AQ),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y143_SLICE_X10Y143_DO5),
.O5(CLBLM_R_X7Y135_SLICE_X9Y135_AO5),
.O6(CLBLM_R_X7Y135_SLICE_X9Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y136_SLICE_X8Y136_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y136_SLICE_X8Y136_AO6),
.Q(CLBLM_R_X7Y136_SLICE_X8Y136_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y136_SLICE_X8Y136_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y136_SLICE_X8Y136_BO6),
.Q(CLBLM_R_X7Y136_SLICE_X8Y136_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y136_SLICE_X8Y136_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y136_SLICE_X8Y136_CO6),
.Q(CLBLM_R_X7Y136_SLICE_X8Y136_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'heeaafebaeeaafeba)
  ) CLBLM_R_X7Y136_SLICE_X8Y136_DLUT (
.I0(CLBLL_L_X4Y134_SLICE_X4Y134_AQ),
.I1(CLBLM_L_X10Y134_SLICE_X12Y134_CQ),
.I2(CLBLM_R_X5Y142_SLICE_X6Y142_CO6),
.I3(CLBLM_R_X7Y135_SLICE_X9Y135_CO6),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y136_SLICE_X8Y136_DO5),
.O6(CLBLM_R_X7Y136_SLICE_X8Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfeeefeeef000f000)
  ) CLBLM_R_X7Y136_SLICE_X8Y136_CLUT (
.I0(CLBLM_L_X8Y138_SLICE_X11Y138_AQ),
.I1(CLBLM_R_X7Y136_SLICE_X8Y136_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X12Y136_SLICE_X16Y136_BQ),
.I4(1'b1),
.I5(CLBLM_R_X7Y144_SLICE_X9Y144_BO6),
.O5(CLBLM_R_X7Y136_SLICE_X8Y136_CO5),
.O6(CLBLM_R_X7Y136_SLICE_X8Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfd0df808ff0ff000)
  ) CLBLM_R_X7Y136_SLICE_X8Y136_BLUT (
.I0(CLBLL_L_X4Y137_SLICE_X4Y137_CQ),
.I1(CLBLM_R_X7Y136_SLICE_X8Y136_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y136_SLICE_X12Y136_A5Q),
.I4(CLBLM_R_X11Y136_SLICE_X14Y136_AQ),
.I5(CLBLM_L_X12Y135_SLICE_X17Y135_AQ),
.O5(CLBLM_R_X7Y136_SLICE_X8Y136_BO5),
.O6(CLBLM_R_X7Y136_SLICE_X8Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfc5cfc5c0c5cfc5)
  ) CLBLM_R_X7Y136_SLICE_X8Y136_ALUT (
.I0(CLBLM_L_X12Y134_SLICE_X17Y134_AQ),
.I1(CLBLM_R_X11Y146_SLICE_X14Y146_AQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X5Y136_SLICE_X6Y136_CQ),
.I5(CLBLM_R_X7Y134_SLICE_X8Y134_CQ),
.O5(CLBLM_R_X7Y136_SLICE_X8Y136_AO5),
.O6(CLBLM_R_X7Y136_SLICE_X8Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y136_SLICE_X9Y136_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y136_SLICE_X9Y136_AO6),
.Q(CLBLM_R_X7Y136_SLICE_X9Y136_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y136_SLICE_X9Y136_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y136_SLICE_X9Y136_CO6),
.Q(CLBLM_R_X7Y136_SLICE_X9Y136_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8800880000000000)
  ) CLBLM_R_X7Y136_SLICE_X9Y136_DLUT (
.I0(CLBLM_L_X8Y138_SLICE_X11Y138_AQ),
.I1(CLBLM_R_X7Y135_SLICE_X8Y135_AQ),
.I2(1'b1),
.I3(CLBLM_R_X7Y135_SLICE_X8Y135_CQ),
.I4(1'b1),
.I5(CLBLM_R_X7Y135_SLICE_X9Y135_A5Q),
.O5(CLBLM_R_X7Y136_SLICE_X9Y136_DO5),
.O6(CLBLM_R_X7Y136_SLICE_X9Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa0caa0caa00aa00)
  ) CLBLM_R_X7Y136_SLICE_X9Y136_CLUT (
.I0(CLBLM_R_X7Y138_SLICE_X9Y138_AQ),
.I1(CLBLM_R_X7Y136_SLICE_X9Y136_CQ),
.I2(CLBLM_R_X7Y139_SLICE_X9Y139_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X7Y136_SLICE_X9Y136_CO5),
.O6(CLBLM_R_X7Y136_SLICE_X9Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc30fc30aaaaaa00)
  ) CLBLM_R_X7Y136_SLICE_X9Y136_BLUT (
.I0(RIOB33_X105Y121_IOB_X1Y121_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X7Y132_SLICE_X9Y132_AQ),
.I3(CLBLL_L_X4Y136_SLICE_X5Y136_A5Q),
.I4(CLBLM_R_X11Y136_SLICE_X15Y136_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y136_SLICE_X9Y136_BO5),
.O6(CLBLM_R_X7Y136_SLICE_X9Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffca80000fca8)
  ) CLBLM_R_X7Y136_SLICE_X9Y136_ALUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_R_X7Y136_SLICE_X8Y136_DO6),
.I2(CLBLM_R_X7Y136_SLICE_X9Y136_AQ),
.I3(CLBLM_L_X8Y138_SLICE_X10Y138_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X5Y138_SLICE_X6Y138_CQ),
.O5(CLBLM_R_X7Y136_SLICE_X9Y136_AO5),
.O6(CLBLM_R_X7Y136_SLICE_X9Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y137_SLICE_X8Y137_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y137_SLICE_X8Y137_AO6),
.Q(CLBLM_R_X7Y137_SLICE_X8Y137_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y137_SLICE_X8Y137_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y137_SLICE_X8Y137_BO6),
.Q(CLBLM_R_X7Y137_SLICE_X8Y137_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y137_SLICE_X8Y137_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y137_SLICE_X8Y137_CO6),
.Q(CLBLM_R_X7Y137_SLICE_X8Y137_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha000a00000000000)
  ) CLBLM_R_X7Y137_SLICE_X8Y137_DLUT (
.I0(CLBLM_R_X3Y138_SLICE_X3Y138_AQ),
.I1(1'b1),
.I2(CLBLM_R_X7Y143_SLICE_X8Y143_A5Q),
.I3(CLBLL_L_X4Y136_SLICE_X5Y136_CQ),
.I4(1'b1),
.I5(CLBLM_R_X7Y133_SLICE_X8Y133_CQ),
.O5(CLBLM_R_X7Y137_SLICE_X8Y137_DO5),
.O6(CLBLM_R_X7Y137_SLICE_X8Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00aa3caacc)
  ) CLBLM_R_X7Y137_SLICE_X8Y137_CLUT (
.I0(CLBLM_L_X12Y136_SLICE_X16Y136_C5Q),
.I1(CLBLM_R_X7Y137_SLICE_X8Y137_CQ),
.I2(CLBLL_L_X4Y137_SLICE_X5Y137_AO5),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y140_SLICE_X9Y140_BQ),
.I5(CLBLM_R_X11Y135_SLICE_X14Y135_AQ),
.O5(CLBLM_R_X7Y137_SLICE_X8Y137_CO5),
.O6(CLBLM_R_X7Y137_SLICE_X8Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa0afa0afc0cfc0c)
  ) CLBLM_R_X7Y137_SLICE_X8Y137_BLUT (
.I0(CLBLM_R_X7Y138_SLICE_X8Y138_CQ),
.I1(CLBLM_R_X7Y137_SLICE_X8Y137_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y141_SLICE_X13Y141_A5Q),
.I4(1'b1),
.I5(CLBLM_L_X8Y143_SLICE_X10Y143_DO5),
.O5(CLBLM_R_X7Y137_SLICE_X8Y137_BO5),
.O6(CLBLM_R_X7Y137_SLICE_X8Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffcfff0cccc0000)
  ) CLBLM_R_X7Y137_SLICE_X8Y137_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y136_SLICE_X10Y136_BQ),
.I2(CLBLM_R_X7Y137_SLICE_X8Y137_AQ),
.I3(CLBLM_R_X7Y133_SLICE_X8Y133_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y144_SLICE_X9Y144_BO6),
.O5(CLBLM_R_X7Y137_SLICE_X8Y137_AO5),
.O6(CLBLM_R_X7Y137_SLICE_X8Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y137_SLICE_X9Y137_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y137_SLICE_X9Y137_AO6),
.Q(CLBLM_R_X7Y137_SLICE_X9Y137_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y137_SLICE_X9Y137_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y137_SLICE_X9Y137_BO6),
.Q(CLBLM_R_X7Y137_SLICE_X9Y137_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff5fffffff)
  ) CLBLM_R_X7Y137_SLICE_X9Y137_DLUT (
.I0(CLBLM_L_X10Y137_SLICE_X13Y137_AQ),
.I1(1'b1),
.I2(CLBLL_L_X4Y135_SLICE_X5Y135_BQ),
.I3(CLBLM_R_X7Y137_SLICE_X9Y137_BQ),
.I4(CLBLM_L_X8Y139_SLICE_X10Y139_BQ),
.I5(CLBLM_R_X7Y133_SLICE_X8Y133_BQ),
.O5(CLBLM_R_X7Y137_SLICE_X9Y137_DO5),
.O6(CLBLM_R_X7Y137_SLICE_X9Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000404)
  ) CLBLM_R_X7Y137_SLICE_X9Y137_CLUT (
.I0(CLBLL_L_X4Y136_SLICE_X4Y136_DQ),
.I1(CLBLM_R_X7Y136_SLICE_X9Y136_DO6),
.I2(CLBLM_L_X12Y139_SLICE_X16Y139_A5Q),
.I3(1'b1),
.I4(CLBLM_R_X7Y137_SLICE_X9Y137_DO6),
.I5(CLBLM_L_X8Y140_SLICE_X11Y140_DO6),
.O5(CLBLM_R_X7Y137_SLICE_X9Y137_CO5),
.O6(CLBLM_R_X7Y137_SLICE_X9Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cf03cf03cc00)
  ) CLBLM_R_X7Y137_SLICE_X9Y137_BLUT (
.I0(1'b1),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_L_X10Y137_SLICE_X13Y137_BQ),
.I4(CLBLM_L_X8Y138_SLICE_X11Y138_AQ),
.I5(CLBLM_L_X10Y138_SLICE_X13Y138_DO6),
.O5(CLBLM_R_X7Y137_SLICE_X9Y137_BO5),
.O6(CLBLM_R_X7Y137_SLICE_X9Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbbbbbbb8888b8b8)
  ) CLBLM_R_X7Y137_SLICE_X9Y137_ALUT (
.I0(CLBLM_L_X10Y139_SLICE_X12Y139_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X7Y137_SLICE_X9Y137_AQ),
.I3(1'b1),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X7Y137_SLICE_X9Y137_CO6),
.O5(CLBLM_R_X7Y137_SLICE_X9Y137_AO5),
.O6(CLBLM_R_X7Y137_SLICE_X9Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y138_SLICE_X8Y138_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y138_SLICE_X8Y138_AO6),
.Q(CLBLM_R_X7Y138_SLICE_X8Y138_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y138_SLICE_X8Y138_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y138_SLICE_X8Y138_BO6),
.Q(CLBLM_R_X7Y138_SLICE_X8Y138_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y138_SLICE_X8Y138_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y138_SLICE_X8Y138_CO6),
.Q(CLBLM_R_X7Y138_SLICE_X8Y138_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff7fffffff)
  ) CLBLM_R_X7Y138_SLICE_X8Y138_DLUT (
.I0(CLBLM_L_X8Y136_SLICE_X11Y136_AQ),
.I1(CLBLM_R_X7Y138_SLICE_X8Y138_CQ),
.I2(CLBLM_L_X8Y138_SLICE_X10Y138_CQ),
.I3(CLBLM_R_X5Y139_SLICE_X7Y139_BQ),
.I4(CLBLM_R_X7Y138_SLICE_X8Y138_BQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X7Y138_SLICE_X8Y138_DO5),
.O6(CLBLM_R_X7Y138_SLICE_X8Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8888888888dddd88)
  ) CLBLM_R_X7Y138_SLICE_X8Y138_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y139_SLICE_X7Y139_BQ),
.I2(1'b1),
.I3(CLBLM_R_X7Y135_SLICE_X9Y135_CO6),
.I4(CLBLM_L_X8Y140_SLICE_X10Y140_DQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X7Y138_SLICE_X8Y138_CO5),
.O6(CLBLM_R_X7Y138_SLICE_X8Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf101f101f202f202)
  ) CLBLM_R_X7Y138_SLICE_X8Y138_BLUT (
.I0(CLBLM_R_X7Y136_SLICE_X9Y136_BO5),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X11Y139_SLICE_X15Y139_A5Q),
.I4(1'b1),
.I5(CLBLM_R_X5Y138_SLICE_X6Y138_CQ),
.O5(CLBLM_R_X7Y138_SLICE_X8Y138_BO5),
.O6(CLBLM_R_X7Y138_SLICE_X8Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff44f4000044f4)
  ) CLBLM_R_X7Y138_SLICE_X8Y138_ALUT (
.I0(CLBLM_R_X7Y138_SLICE_X8Y138_DO6),
.I1(CLBLM_R_X7Y138_SLICE_X9Y138_BO6),
.I2(CLBLM_R_X7Y138_SLICE_X8Y138_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X12Y138_SLICE_X16Y138_BQ),
.O5(CLBLM_R_X7Y138_SLICE_X8Y138_AO5),
.O6(CLBLM_R_X7Y138_SLICE_X8Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y138_SLICE_X9Y138_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y138_SLICE_X9Y138_AO6),
.Q(CLBLM_R_X7Y138_SLICE_X9Y138_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffafffa)
  ) CLBLM_R_X7Y138_SLICE_X9Y138_DLUT (
.I0(CLBLM_R_X7Y134_SLICE_X9Y134_AQ),
.I1(1'b1),
.I2(CLBLM_L_X8Y140_SLICE_X10Y140_DQ),
.I3(CLBLM_R_X5Y138_SLICE_X6Y138_CQ),
.I4(1'b1),
.I5(CLBLM_R_X7Y138_SLICE_X9Y138_AQ),
.O5(CLBLM_R_X7Y138_SLICE_X9Y138_DO5),
.O6(CLBLM_R_X7Y138_SLICE_X9Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h4040000040400000)
  ) CLBLM_R_X7Y138_SLICE_X9Y138_CLUT (
.I0(CLBLM_L_X8Y138_SLICE_X10Y138_AQ),
.I1(CLBLM_R_X7Y137_SLICE_X8Y137_CQ),
.I2(CLBLM_R_X7Y140_SLICE_X9Y140_BQ),
.I3(1'b1),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y138_SLICE_X9Y138_CO5),
.O6(CLBLM_R_X7Y138_SLICE_X9Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000040000000)
  ) CLBLM_R_X7Y138_SLICE_X9Y138_BLUT (
.I0(CLBLM_R_X7Y138_SLICE_X9Y138_DO6),
.I1(CLBLM_R_X7Y134_SLICE_X8Y134_AQ),
.I2(CLBLL_L_X4Y138_SLICE_X5Y138_BQ),
.I3(CLBLM_L_X10Y134_SLICE_X13Y134_BQ),
.I4(CLBLM_R_X11Y137_SLICE_X14Y137_AQ),
.I5(CLBLM_L_X8Y140_SLICE_X11Y140_CO6),
.O5(CLBLM_R_X7Y138_SLICE_X9Y138_BO5),
.O6(CLBLM_R_X7Y138_SLICE_X9Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0faf500000a05)
  ) CLBLM_R_X7Y138_SLICE_X9Y138_ALUT (
.I0(CLBLM_L_X8Y138_SLICE_X10Y138_CQ),
.I1(1'b1),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y138_SLICE_X11Y138_CO5),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X11Y138_SLICE_X14Y138_DQ),
.O5(CLBLM_R_X7Y138_SLICE_X9Y138_AO5),
.O6(CLBLM_R_X7Y138_SLICE_X9Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y139_SLICE_X8Y139_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y139_SLICE_X8Y139_CO6),
.Q(CLBLM_R_X7Y139_SLICE_X8Y139_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y139_SLICE_X8Y139_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y139_SLICE_X8Y139_AO6),
.Q(CLBLM_R_X7Y139_SLICE_X8Y139_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y139_SLICE_X8Y139_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y139_SLICE_X8Y139_BO6),
.Q(CLBLM_R_X7Y139_SLICE_X8Y139_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000080008000)
  ) CLBLM_R_X7Y139_SLICE_X8Y139_DLUT (
.I0(CLBLM_R_X11Y136_SLICE_X14Y136_AQ),
.I1(CLBLM_R_X7Y139_SLICE_X8Y139_AQ),
.I2(CLBLM_R_X7Y139_SLICE_X9Y139_BO6),
.I3(CLBLM_R_X11Y138_SLICE_X14Y138_BQ),
.I4(CLBLM_L_X8Y142_SLICE_X10Y142_DQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y139_SLICE_X8Y139_DO5),
.O6(CLBLM_R_X7Y139_SLICE_X8Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0aa00c0c0c0c0)
  ) CLBLM_R_X7Y139_SLICE_X8Y139_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X7Y139_SLICE_X8Y139_AQ),
.I2(CLBLM_L_X8Y142_SLICE_X10Y142_DQ),
.I3(CLBLM_R_X11Y138_SLICE_X15Y138_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y139_SLICE_X8Y139_CO5),
.O6(CLBLM_R_X7Y139_SLICE_X8Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafaf0f00a0a0000)
  ) CLBLM_R_X7Y139_SLICE_X8Y139_BLUT (
.I0(CLBLM_R_X7Y139_SLICE_X9Y139_A5Q),
.I1(1'b1),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X7Y144_SLICE_X9Y144_AQ),
.O5(CLBLM_R_X7Y139_SLICE_X8Y139_BO5),
.O6(CLBLM_R_X7Y139_SLICE_X8Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00000f0f000ee)
  ) CLBLM_R_X7Y139_SLICE_X8Y139_ALUT (
.I0(CLBLM_R_X7Y139_SLICE_X8Y139_AQ),
.I1(CLBLM_R_X7Y140_SLICE_X8Y140_BO6),
.I2(CLBLM_L_X12Y135_SLICE_X17Y135_AQ),
.I3(CLBLM_R_X7Y139_SLICE_X8Y139_DO5),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X11Y135_SLICE_X14Y135_AQ),
.O5(CLBLM_R_X7Y139_SLICE_X8Y139_AO5),
.O6(CLBLM_R_X7Y139_SLICE_X8Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y139_SLICE_X9Y139_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y139_SLICE_X9Y139_AO5),
.Q(CLBLM_R_X7Y139_SLICE_X9Y139_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y139_SLICE_X9Y139_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y139_SLICE_X9Y139_AO6),
.Q(CLBLM_R_X7Y139_SLICE_X9Y139_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccddddddccffffff)
  ) CLBLM_R_X7Y139_SLICE_X9Y139_DLUT (
.I0(CLBLM_R_X5Y142_SLICE_X6Y142_CO6),
.I1(CLBLM_R_X11Y138_SLICE_X14Y138_DQ),
.I2(1'b1),
.I3(CLBLL_L_X4Y141_SLICE_X4Y141_DO6),
.I4(CLBLM_R_X3Y140_SLICE_X2Y140_DO6),
.I5(CLBLL_L_X4Y142_SLICE_X4Y142_BO6),
.O5(CLBLM_R_X7Y139_SLICE_X9Y139_DO5),
.O6(CLBLM_R_X7Y139_SLICE_X9Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ffa00000a0a0)
  ) CLBLM_R_X7Y139_SLICE_X9Y139_CLUT (
.I0(CLBLL_L_X4Y142_SLICE_X5Y142_DO6),
.I1(1'b1),
.I2(CLBLM_R_X5Y141_SLICE_X7Y141_DO6),
.I3(CLBLL_L_X4Y139_SLICE_X4Y139_BO6),
.I4(CLBLM_R_X7Y139_SLICE_X9Y139_DO6),
.I5(CLBLM_R_X5Y140_SLICE_X6Y140_AO6),
.O5(CLBLM_R_X7Y139_SLICE_X9Y139_CO5),
.O6(CLBLM_R_X7Y139_SLICE_X9Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0800000000000000)
  ) CLBLM_R_X7Y139_SLICE_X9Y139_BLUT (
.I0(CLBLM_R_X7Y140_SLICE_X9Y140_BQ),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_L_X8Y138_SLICE_X10Y138_AQ),
.I3(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I4(CLBLM_L_X8Y138_SLICE_X10Y138_BQ),
.I5(CLBLM_R_X7Y137_SLICE_X8Y137_CQ),
.O5(CLBLM_R_X7Y139_SLICE_X9Y139_BO5),
.O6(CLBLM_R_X7Y139_SLICE_X9Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccff00aaaa0c0c)
  ) CLBLM_R_X7Y139_SLICE_X9Y139_ALUT (
.I0(CLBLL_L_X4Y139_SLICE_X5Y139_AQ),
.I1(CLBLM_R_X11Y136_SLICE_X15Y136_BQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_L_X10Y139_SLICE_X12Y139_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y139_SLICE_X9Y139_AO5),
.O6(CLBLM_R_X7Y139_SLICE_X9Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y140_SLICE_X8Y140_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y140_SLICE_X8Y140_AO6),
.Q(CLBLM_R_X7Y140_SLICE_X8Y140_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h1333200033330000)
  ) CLBLM_R_X7Y140_SLICE_X8Y140_DLUT (
.I0(CLBLM_R_X7Y139_SLICE_X8Y139_AQ),
.I1(CLBLM_R_X11Y135_SLICE_X14Y135_AQ),
.I2(CLBLM_R_X7Y139_SLICE_X9Y139_BO6),
.I3(CLBLM_R_X11Y138_SLICE_X14Y138_BQ),
.I4(CLBLM_L_X8Y142_SLICE_X10Y142_DQ),
.I5(CLBLM_R_X11Y136_SLICE_X14Y136_AQ),
.O5(CLBLM_R_X7Y140_SLICE_X8Y140_DO5),
.O6(CLBLM_R_X7Y140_SLICE_X8Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0040000000000000)
  ) CLBLM_R_X7Y140_SLICE_X8Y140_CLUT (
.I0(CLBLL_L_X4Y143_SLICE_X5Y143_AO6),
.I1(CLBLM_L_X8Y137_SLICE_X10Y137_DO6),
.I2(CLBLM_R_X5Y132_SLICE_X7Y132_DO6),
.I3(CLBLL_L_X4Y142_SLICE_X4Y142_DO6),
.I4(CLBLM_R_X13Y141_SLICE_X18Y141_AO5),
.I5(CLBLM_L_X10Y141_SLICE_X13Y141_CQ),
.O5(CLBLM_R_X7Y140_SLICE_X8Y140_CO5),
.O6(CLBLM_R_X7Y140_SLICE_X8Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8800880033ff33ff)
  ) CLBLM_R_X7Y140_SLICE_X8Y140_BLUT (
.I0(CLBLM_R_X7Y139_SLICE_X9Y139_BO6),
.I1(CLBLM_R_X11Y138_SLICE_X14Y138_BQ),
.I2(1'b1),
.I3(CLBLM_R_X11Y136_SLICE_X14Y136_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y140_SLICE_X8Y140_BO5),
.O6(CLBLM_R_X7Y140_SLICE_X8Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc50facccc5050)
  ) CLBLM_R_X7Y140_SLICE_X8Y140_ALUT (
.I0(CLBLL_L_X4Y138_SLICE_X5Y138_CO5),
.I1(CLBLM_L_X8Y137_SLICE_X11Y137_BQ),
.I2(CLBLM_R_X7Y140_SLICE_X8Y140_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X5Y141_SLICE_X7Y141_DO6),
.O5(CLBLM_R_X7Y140_SLICE_X8Y140_AO5),
.O6(CLBLM_R_X7Y140_SLICE_X8Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y140_SLICE_X9Y140_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y140_SLICE_X9Y140_AO6),
.Q(CLBLM_R_X7Y140_SLICE_X9Y140_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y140_SLICE_X9Y140_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y140_SLICE_X9Y140_BO6),
.Q(CLBLM_R_X7Y140_SLICE_X9Y140_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y140_SLICE_X9Y140_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y140_SLICE_X9Y140_CO6),
.Q(CLBLM_R_X7Y140_SLICE_X9Y140_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h4444ffff44444444)
  ) CLBLM_R_X7Y140_SLICE_X9Y140_DLUT (
.I0(CLBLM_R_X7Y142_SLICE_X9Y142_CO5),
.I1(CLBLM_L_X8Y141_SLICE_X11Y141_CQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X5Y143_SLICE_X6Y143_AO5),
.I5(CLBLM_L_X10Y140_SLICE_X12Y140_AQ),
.O5(CLBLM_R_X7Y140_SLICE_X9Y140_DO5),
.O6(CLBLM_R_X7Y140_SLICE_X9Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hbfefbeee15451444)
  ) CLBLM_R_X7Y140_SLICE_X9Y140_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y140_SLICE_X8Y140_CO6),
.I2(CLBLM_L_X8Y143_SLICE_X10Y143_DO5),
.I3(CLBLM_L_X12Y139_SLICE_X16Y139_A5Q),
.I4(CLBLM_R_X7Y140_SLICE_X9Y140_CQ),
.I5(CLBLM_R_X11Y137_SLICE_X14Y137_AQ),
.O5(CLBLM_R_X7Y140_SLICE_X9Y140_CO5),
.O6(CLBLM_R_X7Y140_SLICE_X9Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaffffaaaac3cc)
  ) CLBLM_R_X7Y140_SLICE_X9Y140_BLUT (
.I0(CLBLM_L_X10Y140_SLICE_X13Y140_DQ),
.I1(CLBLM_R_X7Y140_SLICE_X9Y140_BQ),
.I2(CLBLM_L_X8Y138_SLICE_X10Y138_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X11Y135_SLICE_X14Y135_AQ),
.O5(CLBLM_R_X7Y140_SLICE_X9Y140_BO5),
.O6(CLBLM_R_X7Y140_SLICE_X9Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccf5f5cccca0a0)
  ) CLBLM_R_X7Y140_SLICE_X9Y140_ALUT (
.I0(CLBLM_L_X8Y143_SLICE_X10Y143_DO6),
.I1(CLBLM_R_X5Y140_SLICE_X7Y140_BQ),
.I2(CLBLM_R_X7Y140_SLICE_X9Y140_AQ),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X10Y140_SLICE_X13Y140_DQ),
.O5(CLBLM_R_X7Y140_SLICE_X9Y140_AO5),
.O6(CLBLM_R_X7Y140_SLICE_X9Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y141_SLICE_X8Y141_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y141_SLICE_X8Y141_AO6),
.Q(CLBLM_R_X7Y141_SLICE_X8Y141_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000880000008800)
  ) CLBLM_R_X7Y141_SLICE_X8Y141_DLUT (
.I0(CLBLM_R_X5Y139_SLICE_X7Y139_AQ),
.I1(CLBLM_L_X8Y138_SLICE_X10Y138_D5Q),
.I2(1'b1),
.I3(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I4(CLBLM_L_X8Y138_SLICE_X10Y138_BQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y141_SLICE_X8Y141_DO5),
.O6(CLBLM_R_X7Y141_SLICE_X8Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000a8fc88cc)
  ) CLBLM_R_X7Y141_SLICE_X8Y141_CLUT (
.I0(CLBLM_R_X7Y139_SLICE_X8Y139_CO5),
.I1(CLBLM_R_X7Y141_SLICE_X8Y141_BO5),
.I2(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I3(CLBLM_R_X7Y140_SLICE_X8Y140_BO5),
.I4(CLBLM_L_X8Y138_SLICE_X10Y138_BQ),
.I5(CLBLM_R_X11Y138_SLICE_X14Y138_DQ),
.O5(CLBLM_R_X7Y141_SLICE_X8Y141_CO5),
.O6(CLBLM_R_X7Y141_SLICE_X8Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fff7fffcc00cc00)
  ) CLBLM_R_X7Y141_SLICE_X8Y141_BLUT (
.I0(CLBLM_R_X7Y139_SLICE_X8Y139_AQ),
.I1(CLBLM_R_X7Y140_SLICE_X9Y140_BQ),
.I2(CLBLM_L_X8Y142_SLICE_X10Y142_DQ),
.I3(CLBLM_R_X7Y137_SLICE_X8Y137_CQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y141_SLICE_X8Y141_BO5),
.O6(CLBLM_R_X7Y141_SLICE_X8Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0c0cac0c0)
  ) CLBLM_R_X7Y141_SLICE_X8Y141_ALUT (
.I0(CLBLM_R_X7Y141_SLICE_X8Y141_DO6),
.I1(CLBLM_R_X7Y143_SLICE_X8Y143_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y141_SLICE_X8Y141_BO6),
.I4(CLBLM_R_X11Y138_SLICE_X14Y138_DQ),
.I5(CLBLM_R_X7Y140_SLICE_X8Y140_BO5),
.O5(CLBLM_R_X7Y141_SLICE_X8Y141_AO5),
.O6(CLBLM_R_X7Y141_SLICE_X8Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y141_SLICE_X9Y141_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y141_SLICE_X9Y141_AO6),
.Q(CLBLM_R_X7Y141_SLICE_X9Y141_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y141_SLICE_X9Y141_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y141_SLICE_X9Y141_BO6),
.Q(CLBLM_R_X7Y141_SLICE_X9Y141_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7f775f553f330f00)
  ) CLBLM_R_X7Y141_SLICE_X9Y141_DLUT (
.I0(CLBLM_R_X5Y143_SLICE_X6Y143_AO5),
.I1(CLBLL_L_X4Y143_SLICE_X5Y143_AO5),
.I2(CLBLM_R_X7Y142_SLICE_X9Y142_CO6),
.I3(CLBLM_R_X7Y142_SLICE_X9Y142_BQ),
.I4(CLBLM_R_X7Y141_SLICE_X9Y141_AQ),
.I5(CLBLM_R_X11Y141_SLICE_X15Y141_BQ),
.O5(CLBLM_R_X7Y141_SLICE_X9Y141_DO5),
.O6(CLBLM_R_X7Y141_SLICE_X9Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0302000200000000)
  ) CLBLM_R_X7Y141_SLICE_X9Y141_CLUT (
.I0(CLBLM_L_X12Y141_SLICE_X17Y141_AQ),
.I1(CLBLM_R_X3Y143_SLICE_X2Y143_AO5),
.I2(CLBLM_R_X7Y143_SLICE_X9Y143_DO6),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(CLBLM_L_X12Y136_SLICE_X16Y136_C5Q),
.I5(RIOB33_X105Y131_IOB_X1Y132_I),
.O5(CLBLM_R_X7Y141_SLICE_X9Y141_CO5),
.O6(CLBLM_R_X7Y141_SLICE_X9Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hafae0504ffee5544)
  ) CLBLM_R_X7Y141_SLICE_X9Y141_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y141_SLICE_X9Y141_BQ),
.I2(CLBLM_L_X10Y139_SLICE_X13Y139_B5Q),
.I3(CLBLM_R_X7Y140_SLICE_X9Y140_BQ),
.I4(CLBLM_R_X7Y140_SLICE_X9Y140_AQ),
.I5(CLBLM_L_X12Y134_SLICE_X17Y134_AO6),
.O5(CLBLM_R_X7Y141_SLICE_X9Y141_BO5),
.O6(CLBLM_R_X7Y141_SLICE_X9Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3fff2fa030f020a)
  ) CLBLM_R_X7Y141_SLICE_X9Y141_ALUT (
.I0(CLBLM_R_X7Y141_SLICE_X9Y141_AQ),
.I1(CLBLL_L_X4Y137_SLICE_X4Y137_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X12Y135_SLICE_X17Y135_AQ),
.I4(CLBLM_L_X8Y142_SLICE_X10Y142_DQ),
.I5(CLBLM_L_X8Y138_SLICE_X10Y138_D5Q),
.O5(CLBLM_R_X7Y141_SLICE_X9Y141_AO5),
.O6(CLBLM_R_X7Y141_SLICE_X9Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y142_SLICE_X8Y142_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y142_SLICE_X8Y142_AO6),
.Q(CLBLM_R_X7Y142_SLICE_X8Y142_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffff73ffffff50)
  ) CLBLM_R_X7Y142_SLICE_X8Y142_DLUT (
.I0(CLBLM_R_X3Y142_SLICE_X3Y142_AO6),
.I1(CLBLM_R_X7Y142_SLICE_X9Y142_CO6),
.I2(CLBLM_R_X7Y140_SLICE_X8Y140_AQ),
.I3(CLBLM_R_X7Y142_SLICE_X8Y142_CO6),
.I4(CLBLM_R_X7Y144_SLICE_X8Y144_DO6),
.I5(CLBLM_L_X12Y140_SLICE_X16Y140_AQ),
.O5(CLBLM_R_X7Y142_SLICE_X8Y142_DO5),
.O6(CLBLM_R_X7Y142_SLICE_X8Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000004000)
  ) CLBLM_R_X7Y142_SLICE_X8Y142_CLUT (
.I0(CLBLM_R_X3Y143_SLICE_X2Y143_AO5),
.I1(CLBLM_R_X7Y138_SLICE_X8Y138_AQ),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(RIOB33_X105Y131_IOB_X1Y132_I),
.I4(RIOB33_X105Y133_IOB_X1Y134_I),
.I5(RIOB33_X105Y133_IOB_X1Y133_I),
.O5(CLBLM_R_X7Y142_SLICE_X8Y142_CO5),
.O6(CLBLM_R_X7Y142_SLICE_X8Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'heeeeffeefefefffe)
  ) CLBLM_R_X7Y142_SLICE_X8Y142_BLUT (
.I0(CLBLM_R_X7Y143_SLICE_X8Y143_DO6),
.I1(CLBLM_R_X7Y142_SLICE_X9Y142_DO6),
.I2(CLBLM_L_X8Y141_SLICE_X11Y141_BQ),
.I3(CLBLM_R_X5Y138_SLICE_X7Y138_CQ),
.I4(CLBLM_R_X3Y142_SLICE_X3Y142_AO6),
.I5(CLBLL_L_X4Y143_SLICE_X5Y143_AO5),
.O5(CLBLM_R_X7Y142_SLICE_X8Y142_BO5),
.O6(CLBLM_R_X7Y142_SLICE_X8Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfaeefaee50445044)
  ) CLBLM_R_X7Y142_SLICE_X8Y142_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y135_SLICE_X7Y135_A5Q),
.I2(CLBLM_R_X7Y142_SLICE_X8Y142_AQ),
.I3(CLBLL_L_X4Y133_SLICE_X5Y133_BO6),
.I4(1'b1),
.I5(CLBLM_L_X12Y144_SLICE_X17Y144_AQ),
.O5(CLBLM_R_X7Y142_SLICE_X8Y142_AO5),
.O6(CLBLM_R_X7Y142_SLICE_X8Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y142_SLICE_X9Y142_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y142_SLICE_X9Y142_AO6),
.Q(CLBLM_R_X7Y142_SLICE_X9Y142_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y142_SLICE_X9Y142_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y142_SLICE_X9Y142_BO6),
.Q(CLBLM_R_X7Y142_SLICE_X9Y142_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000010000000000)
  ) CLBLM_R_X7Y142_SLICE_X9Y142_DLUT (
.I0(CLBLM_R_X3Y143_SLICE_X2Y143_AO5),
.I1(RIOB33_X105Y131_IOB_X1Y132_I),
.I2(RIOB33_X105Y133_IOB_X1Y134_I),
.I3(CLBLM_L_X8Y141_SLICE_X10Y141_BQ),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(RIOB33_X105Y133_IOB_X1Y133_I),
.O5(CLBLM_R_X7Y142_SLICE_X9Y142_DO5),
.O6(CLBLM_R_X7Y142_SLICE_X9Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffefffffffffb)
  ) CLBLM_R_X7Y142_SLICE_X9Y142_CLUT (
.I0(CLBLM_R_X3Y143_SLICE_X2Y143_AO5),
.I1(RIOB33_X105Y131_IOB_X1Y132_I),
.I2(RIOB33_X105Y133_IOB_X1Y134_I),
.I3(RIOB33_X105Y133_IOB_X1Y133_I),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y142_SLICE_X9Y142_CO5),
.O6(CLBLM_R_X7Y142_SLICE_X9Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fff0ccf000f000)
  ) CLBLM_R_X7Y142_SLICE_X9Y142_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y142_SLICE_X9Y142_BQ),
.I2(CLBLL_L_X4Y137_SLICE_X4Y137_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X11Y141_SLICE_X14Y141_AQ),
.I5(CLBLM_L_X8Y143_SLICE_X10Y143_DO6),
.O5(CLBLM_R_X7Y142_SLICE_X9Y142_BO5),
.O6(CLBLM_R_X7Y142_SLICE_X9Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00ff33cc00)
  ) CLBLM_R_X7Y142_SLICE_X9Y142_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(1'b1),
.I3(CLBLM_L_X12Y140_SLICE_X16Y140_AQ),
.I4(CLBLM_R_X7Y144_SLICE_X9Y144_AQ),
.I5(CLBLM_L_X10Y144_SLICE_X12Y144_AO5),
.O5(CLBLM_R_X7Y142_SLICE_X9Y142_AO5),
.O6(CLBLM_R_X7Y142_SLICE_X9Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y143_SLICE_X8Y143_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y143_SLICE_X8Y143_BO6),
.Q(CLBLM_R_X7Y143_SLICE_X8Y143_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y143_SLICE_X8Y143_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y143_SLICE_X8Y143_AO6),
.Q(CLBLM_R_X7Y143_SLICE_X8Y143_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y143_SLICE_X8Y143_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y143_SLICE_X8Y143_CO6),
.Q(CLBLM_R_X7Y143_SLICE_X8Y143_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000004000000000)
  ) CLBLM_R_X7Y143_SLICE_X8Y143_DLUT (
.I0(CLBLM_R_X3Y143_SLICE_X2Y143_AO5),
.I1(CLBLM_R_X7Y143_SLICE_X8Y143_AQ),
.I2(RIOB33_X105Y133_IOB_X1Y133_I),
.I3(RIOB33_X105Y133_IOB_X1Y134_I),
.I4(RIOB33_X105Y131_IOB_X1Y132_I),
.I5(RIOB33_X105Y131_IOB_X1Y131_I),
.O5(CLBLM_R_X7Y143_SLICE_X8Y143_DO5),
.O6(CLBLM_R_X7Y143_SLICE_X8Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hee44ee44fa50fa50)
  ) CLBLM_R_X7Y143_SLICE_X8Y143_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y143_SLICE_X8Y143_CQ),
.I2(CLBLM_R_X5Y135_SLICE_X6Y135_DQ),
.I3(CLBLM_L_X12Y141_SLICE_X16Y141_AQ),
.I4(1'b1),
.I5(CLBLL_L_X4Y133_SLICE_X5Y133_BO6),
.O5(CLBLM_R_X7Y143_SLICE_X8Y143_CO5),
.O6(CLBLM_R_X7Y143_SLICE_X8Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hd5d5c0c033003300)
  ) CLBLM_R_X7Y143_SLICE_X8Y143_BLUT (
.I0(CLBLM_R_X7Y133_SLICE_X8Y133_DO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y142_SLICE_X12Y142_BQ),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(CLBLM_R_X7Y143_SLICE_X8Y143_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X7Y143_SLICE_X8Y143_BO5),
.O6(CLBLM_R_X7Y143_SLICE_X8Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffe400e4ffe400e4)
  ) CLBLM_R_X7Y143_SLICE_X8Y143_ALUT (
.I0(CLBLM_L_X8Y143_SLICE_X10Y143_DO6),
.I1(CLBLM_L_X12Y144_SLICE_X17Y144_AQ),
.I2(CLBLM_R_X7Y143_SLICE_X8Y143_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y143_SLICE_X9Y143_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y143_SLICE_X8Y143_AO5),
.O6(CLBLM_R_X7Y143_SLICE_X8Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y143_SLICE_X9Y143_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y143_SLICE_X9Y143_AO6),
.Q(CLBLM_R_X7Y143_SLICE_X9Y143_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y143_SLICE_X9Y143_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y143_SLICE_X9Y143_BO6),
.Q(CLBLM_R_X7Y143_SLICE_X9Y143_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y143_SLICE_X9Y143_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y143_SLICE_X9Y143_CO6),
.Q(CLBLM_R_X7Y143_SLICE_X9Y143_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffff00ff00)
  ) CLBLM_R_X7Y143_SLICE_X9Y143_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(RIOB33_X105Y133_IOB_X1Y133_I),
.I4(1'b1),
.I5(RIOB33_X105Y133_IOB_X1Y134_I),
.O5(CLBLM_R_X7Y143_SLICE_X9Y143_DO5),
.O6(CLBLM_R_X7Y143_SLICE_X9Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00e4e4e4e4)
  ) CLBLM_R_X7Y143_SLICE_X9Y143_CLUT (
.I0(CLBLM_L_X8Y143_SLICE_X10Y143_DO5),
.I1(CLBLM_R_X7Y143_SLICE_X9Y143_CQ),
.I2(CLBLM_R_X7Y135_SLICE_X8Y135_AQ),
.I3(CLBLM_L_X12Y143_SLICE_X16Y143_BQ),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X7Y143_SLICE_X9Y143_CO5),
.O6(CLBLM_R_X7Y143_SLICE_X9Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0acacacac)
  ) CLBLM_R_X7Y143_SLICE_X9Y143_BLUT (
.I0(CLBLM_R_X3Y137_SLICE_X3Y137_CQ),
.I1(CLBLM_L_X8Y142_SLICE_X11Y142_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X10Y144_SLICE_X12Y144_AO5),
.O5(CLBLM_R_X7Y143_SLICE_X9Y143_BO5),
.O6(CLBLM_R_X7Y143_SLICE_X9Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hafafafafacacacac)
  ) CLBLM_R_X7Y143_SLICE_X9Y143_ALUT (
.I0(CLBLM_L_X10Y140_SLICE_X13Y140_C5Q),
.I1(CLBLM_R_X7Y143_SLICE_X9Y143_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X10Y144_SLICE_X12Y144_AO5),
.O5(CLBLM_R_X7Y143_SLICE_X9Y143_AO5),
.O6(CLBLM_R_X7Y143_SLICE_X9Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y144_SLICE_X8Y144_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y144_SLICE_X8Y144_AO6),
.Q(CLBLM_R_X7Y144_SLICE_X8Y144_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y144_SLICE_X8Y144_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y144_SLICE_X8Y144_BO6),
.Q(CLBLM_R_X7Y144_SLICE_X8Y144_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y144_SLICE_X8Y144_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y144_SLICE_X8Y144_CO6),
.Q(CLBLM_R_X7Y144_SLICE_X8Y144_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000400)
  ) CLBLM_R_X7Y144_SLICE_X8Y144_DLUT (
.I0(CLBLM_R_X3Y143_SLICE_X2Y143_AO5),
.I1(CLBLM_R_X7Y144_SLICE_X8Y144_CQ),
.I2(RIOB33_X105Y133_IOB_X1Y134_I),
.I3(RIOB33_X105Y131_IOB_X1Y132_I),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(RIOB33_X105Y133_IOB_X1Y133_I),
.O5(CLBLM_R_X7Y144_SLICE_X8Y144_DO5),
.O6(CLBLM_R_X7Y144_SLICE_X8Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffce00ceff000000)
  ) CLBLM_R_X7Y144_SLICE_X8Y144_CLUT (
.I0(CLBLM_R_X11Y136_SLICE_X14Y136_DQ),
.I1(CLBLM_R_X7Y144_SLICE_X8Y144_CQ),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y140_SLICE_X8Y140_AQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X7Y144_SLICE_X8Y144_CO5),
.O6(CLBLM_R_X7Y144_SLICE_X8Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f033cc0000)
  ) CLBLM_R_X7Y144_SLICE_X8Y144_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y144_SLICE_X8Y144_BQ),
.I2(CLBLM_L_X8Y143_SLICE_X10Y143_BQ),
.I3(CLBLM_R_X7Y143_SLICE_X9Y143_BQ),
.I4(CLBLM_L_X8Y144_SLICE_X11Y144_BO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X7Y144_SLICE_X8Y144_BO5),
.O6(CLBLM_R_X7Y144_SLICE_X8Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff90a0000090a0)
  ) CLBLM_R_X7Y144_SLICE_X8Y144_ALUT (
.I0(CLBLM_R_X7Y144_SLICE_X8Y144_AQ),
.I1(CLBLM_R_X7Y144_SLICE_X8Y144_BQ),
.I2(CLBLM_L_X8Y144_SLICE_X11Y144_BO6),
.I3(CLBLM_R_X7Y143_SLICE_X9Y143_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y140_SLICE_X10Y140_CQ),
.O5(CLBLM_R_X7Y144_SLICE_X8Y144_AO5),
.O6(CLBLM_R_X7Y144_SLICE_X8Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y144_SLICE_X9Y144_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y144_SLICE_X9Y144_AO6),
.Q(CLBLM_R_X7Y144_SLICE_X9Y144_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y144_SLICE_X9Y144_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y144_SLICE_X9Y144_DO5),
.O6(CLBLM_R_X7Y144_SLICE_X9Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y144_SLICE_X9Y144_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y144_SLICE_X9Y144_CO5),
.O6(CLBLM_R_X7Y144_SLICE_X9Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff000000af0000)
  ) CLBLM_R_X7Y144_SLICE_X9Y144_BLUT (
.I0(RIOB33_X105Y121_IOB_X1Y121_I),
.I1(1'b1),
.I2(CLBLM_R_X11Y136_SLICE_X14Y136_DQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X7Y144_SLICE_X8Y144_CQ),
.O5(CLBLM_R_X7Y144_SLICE_X9Y144_BO5),
.O6(CLBLM_R_X7Y144_SLICE_X9Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f033003300)
  ) CLBLM_R_X7Y144_SLICE_X9Y144_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y144_SLICE_X12Y144_AO5),
.I2(CLBLM_R_X7Y131_SLICE_X9Y131_BQ),
.I3(CLBLM_R_X7Y143_SLICE_X9Y143_AQ),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X7Y144_SLICE_X9Y144_AO5),
.O6(CLBLM_R_X7Y144_SLICE_X9Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y146_SLICE_X8Y146_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y146_SLICE_X12Y146_AO6),
.Q(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y146_SLICE_X8Y146_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y146_SLICE_X8Y146_DO5),
.O6(CLBLM_R_X7Y146_SLICE_X8Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y146_SLICE_X8Y146_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y146_SLICE_X8Y146_CO5),
.O6(CLBLM_R_X7Y146_SLICE_X8Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y146_SLICE_X8Y146_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y146_SLICE_X8Y146_BO5),
.O6(CLBLM_R_X7Y146_SLICE_X8Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y146_SLICE_X8Y146_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y146_SLICE_X8Y146_AO5),
.O6(CLBLM_R_X7Y146_SLICE_X8Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y146_SLICE_X9Y146_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y146_SLICE_X9Y146_DO5),
.O6(CLBLM_R_X7Y146_SLICE_X9Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y146_SLICE_X9Y146_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y146_SLICE_X9Y146_CO5),
.O6(CLBLM_R_X7Y146_SLICE_X9Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y146_SLICE_X9Y146_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y146_SLICE_X9Y146_BO5),
.O6(CLBLM_R_X7Y146_SLICE_X9Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y146_SLICE_X9Y146_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y146_SLICE_X9Y146_AO5),
.O6(CLBLM_R_X7Y146_SLICE_X9Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y131_SLICE_X14Y131_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y131_SLICE_X14Y131_BO6),
.Q(CLBLM_R_X11Y131_SLICE_X14Y131_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000272700007227)
  ) CLBLM_R_X11Y131_SLICE_X14Y131_DLUT (
.I0(CLBLM_R_X5Y132_SLICE_X7Y132_DO6),
.I1(CLBLM_R_X11Y146_SLICE_X14Y146_AQ),
.I2(CLBLM_L_X8Y131_SLICE_X10Y131_A5Q),
.I3(CLBLM_R_X11Y131_SLICE_X14Y131_AO5),
.I4(CLBLM_R_X11Y131_SLICE_X14Y131_BQ),
.I5(CLBLM_L_X10Y130_SLICE_X13Y130_AO5),
.O5(CLBLM_R_X11Y131_SLICE_X14Y131_DO5),
.O6(CLBLM_R_X11Y131_SLICE_X14Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff06f6ff00f606)
  ) CLBLM_R_X11Y131_SLICE_X14Y131_CLUT (
.I0(CLBLM_R_X11Y131_SLICE_X15Y131_AO6),
.I1(CLBLM_R_X11Y131_SLICE_X15Y131_CO6),
.I2(CLBLM_R_X5Y133_SLICE_X7Y133_CO6),
.I3(CLBLM_L_X10Y137_SLICE_X12Y137_BQ),
.I4(CLBLM_R_X3Y139_SLICE_X3Y139_BO6),
.I5(CLBLM_R_X13Y137_SLICE_X18Y137_A5Q),
.O5(CLBLM_R_X11Y131_SLICE_X14Y131_CO5),
.O6(CLBLM_R_X11Y131_SLICE_X14Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hd1d1c0d1d1d1c0d1)
  ) CLBLM_R_X11Y131_SLICE_X14Y131_BLUT (
.I0(CLBLM_R_X11Y131_SLICE_X14Y131_DO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X7Y141_SLICE_X9Y141_AQ),
.I3(RIOB33_X105Y141_IOB_X1Y142_I),
.I4(CLBLM_R_X7Y131_SLICE_X9Y131_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y131_SLICE_X14Y131_BO5),
.O6(CLBLM_R_X11Y131_SLICE_X14Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccc600005555)
  ) CLBLM_R_X11Y131_SLICE_X14Y131_ALUT (
.I0(CLBLL_L_X4Y135_SLICE_X5Y135_CQ),
.I1(CLBLM_R_X7Y131_SLICE_X9Y131_BQ),
.I2(CLBLM_L_X10Y130_SLICE_X12Y130_AQ),
.I3(CLBLM_R_X11Y131_SLICE_X15Y131_BQ),
.I4(CLBLM_L_X10Y131_SLICE_X12Y131_BQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y131_SLICE_X14Y131_AO5),
.O6(CLBLM_R_X11Y131_SLICE_X14Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y131_SLICE_X15Y131_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y131_SLICE_X15Y131_BO6),
.Q(CLBLM_R_X11Y131_SLICE_X15Y131_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff8800ffff)
  ) CLBLM_R_X11Y131_SLICE_X15Y131_DLUT (
.I0(CLBLL_L_X4Y135_SLICE_X5Y135_CQ),
.I1(CLBLM_L_X10Y131_SLICE_X12Y131_BQ),
.I2(1'b1),
.I3(CLBLM_R_X11Y131_SLICE_X15Y131_BQ),
.I4(CLBLM_L_X10Y130_SLICE_X12Y130_AQ),
.I5(CLBLM_R_X5Y132_SLICE_X7Y132_DO6),
.O5(CLBLM_R_X11Y131_SLICE_X15Y131_DO5),
.O6(CLBLM_R_X11Y131_SLICE_X15Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccc6ccccccc6c)
  ) CLBLM_R_X11Y131_SLICE_X15Y131_CLUT (
.I0(CLBLL_L_X4Y135_SLICE_X5Y135_CQ),
.I1(CLBLM_R_X11Y133_SLICE_X15Y133_AQ),
.I2(CLBLM_R_X11Y131_SLICE_X15Y131_BQ),
.I3(CLBLM_L_X10Y131_SLICE_X12Y131_BQ),
.I4(CLBLM_L_X10Y130_SLICE_X12Y130_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y131_SLICE_X15Y131_CO5),
.O6(CLBLM_R_X11Y131_SLICE_X15Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f099f000f000)
  ) CLBLM_R_X11Y131_SLICE_X15Y131_BLUT (
.I0(CLBLM_R_X11Y131_SLICE_X15Y131_DO6),
.I1(CLBLM_R_X11Y131_SLICE_X15Y131_BQ),
.I2(CLBLM_R_X13Y140_SLICE_X18Y140_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X11Y140_SLICE_X15Y140_CQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X11Y131_SLICE_X15Y131_BO5),
.O6(CLBLM_R_X11Y131_SLICE_X15Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00f708fafaffff)
  ) CLBLM_R_X11Y131_SLICE_X15Y131_ALUT (
.I0(CLBLM_L_X10Y131_SLICE_X12Y131_BQ),
.I1(CLBLM_R_X11Y131_SLICE_X15Y131_BQ),
.I2(CLBLM_L_X10Y130_SLICE_X12Y130_AQ),
.I3(CLBLM_L_X10Y131_SLICE_X13Y131_CQ),
.I4(CLBLL_L_X4Y135_SLICE_X5Y135_CQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y131_SLICE_X15Y131_AO5),
.O6(CLBLM_R_X11Y131_SLICE_X15Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y132_SLICE_X14Y132_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y132_SLICE_X14Y132_AO6),
.Q(CLBLM_R_X11Y132_SLICE_X14Y132_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y132_SLICE_X14Y132_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y132_SLICE_X14Y132_BO6),
.Q(CLBLM_R_X11Y132_SLICE_X14Y132_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h000005050a0a0f0f)
  ) CLBLM_R_X11Y132_SLICE_X14Y132_DLUT (
.I0(CLBLM_R_X5Y132_SLICE_X7Y132_DO6),
.I1(1'b1),
.I2(CLBLM_R_X11Y132_SLICE_X14Y132_BQ),
.I3(1'b1),
.I4(CLBLM_L_X10Y130_SLICE_X13Y130_AO6),
.I5(CLBLM_L_X10Y137_SLICE_X12Y137_B5Q),
.O5(CLBLM_R_X11Y132_SLICE_X14Y132_DO5),
.O6(CLBLM_R_X11Y132_SLICE_X14Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffffef)
  ) CLBLM_R_X11Y132_SLICE_X14Y132_CLUT (
.I0(CLBLM_R_X11Y133_SLICE_X15Y133_AQ),
.I1(CLBLM_R_X11Y133_SLICE_X14Y133_BQ),
.I2(CLBLM_L_X8Y131_SLICE_X10Y131_BO5),
.I3(CLBLM_R_X11Y133_SLICE_X14Y133_AQ),
.I4(CLBLM_R_X7Y131_SLICE_X9Y131_BQ),
.I5(CLBLM_R_X11Y133_SLICE_X15Y133_BQ),
.O5(CLBLM_R_X11Y132_SLICE_X14Y132_CO5),
.O6(CLBLM_R_X11Y132_SLICE_X14Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc50555055)
  ) CLBLM_R_X11Y132_SLICE_X14Y132_BLUT (
.I0(CLBLM_R_X11Y132_SLICE_X14Y132_DO6),
.I1(CLBLM_R_X11Y133_SLICE_X14Y133_CQ),
.I2(CLBLM_R_X7Y131_SLICE_X9Y131_AQ),
.I3(RIOB33_X105Y141_IOB_X1Y142_I),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y132_SLICE_X14Y132_BO5),
.O6(CLBLM_R_X11Y132_SLICE_X14Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff000000fcfc)
  ) CLBLM_R_X11Y132_SLICE_X14Y132_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y131_SLICE_X13Y131_BQ),
.I2(CLBLM_R_X11Y132_SLICE_X14Y132_AQ),
.I3(CLBLM_R_X11Y134_SLICE_X14Y134_BQ),
.I4(CLBLM_R_X5Y132_SLICE_X7Y132_DO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y132_SLICE_X14Y132_AO5),
.O6(CLBLM_R_X11Y132_SLICE_X14Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffcfc)
  ) CLBLM_R_X11Y132_SLICE_X15Y132_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y133_SLICE_X15Y133_CQ),
.I2(CLBLM_R_X11Y134_SLICE_X15Y134_CQ),
.I3(1'b1),
.I4(CLBLM_L_X8Y134_SLICE_X11Y134_BQ),
.I5(CLBLM_L_X10Y134_SLICE_X12Y134_AQ),
.O5(CLBLM_R_X11Y132_SLICE_X15Y132_DO5),
.O6(CLBLM_R_X11Y132_SLICE_X15Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5b5a5b5a5b5a5b5a)
  ) CLBLM_R_X11Y132_SLICE_X15Y132_CLUT (
.I0(CLBLM_L_X12Y132_SLICE_X16Y132_BQ),
.I1(CLBLM_R_X11Y132_SLICE_X14Y132_CO6),
.I2(CLBLM_L_X12Y136_SLICE_X16Y136_DQ),
.I3(CLBLM_L_X10Y133_SLICE_X13Y133_CO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y132_SLICE_X15Y132_CO5),
.O6(CLBLM_R_X11Y132_SLICE_X15Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0005010450555154)
  ) CLBLM_R_X11Y132_SLICE_X15Y132_BLUT (
.I0(CLBLM_L_X12Y132_SLICE_X16Y132_CQ),
.I1(CLBLM_R_X11Y131_SLICE_X15Y131_BQ),
.I2(CLBLM_R_X5Y132_SLICE_X7Y132_DO6),
.I3(CLBLM_R_X7Y131_SLICE_X9Y131_BQ),
.I4(CLBLM_R_X11Y131_SLICE_X15Y131_AO5),
.I5(CLBLM_L_X12Y136_SLICE_X16Y136_B5Q),
.O5(CLBLM_R_X11Y132_SLICE_X15Y132_BO5),
.O6(CLBLM_R_X11Y132_SLICE_X15Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h20002000ffef0010)
  ) CLBLM_R_X11Y132_SLICE_X15Y132_ALUT (
.I0(CLBLL_L_X4Y135_SLICE_X5Y135_CQ),
.I1(CLBLM_L_X10Y131_SLICE_X12Y131_BQ),
.I2(CLBLM_L_X10Y130_SLICE_X12Y130_AQ),
.I3(CLBLM_R_X11Y131_SLICE_X15Y131_BQ),
.I4(CLBLM_R_X11Y132_SLICE_X15Y132_CO6),
.I5(1'b1),
.O5(CLBLM_R_X11Y132_SLICE_X15Y132_AO5),
.O6(CLBLM_R_X11Y132_SLICE_X15Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y133_SLICE_X14Y133_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y133_SLICE_X14Y133_AO6),
.Q(CLBLM_R_X11Y133_SLICE_X14Y133_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y133_SLICE_X14Y133_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y133_SLICE_X14Y133_BO6),
.Q(CLBLM_R_X11Y133_SLICE_X14Y133_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y133_SLICE_X14Y133_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y133_SLICE_X14Y133_CO6),
.Q(CLBLM_R_X11Y133_SLICE_X14Y133_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h000003f3000009f9)
  ) CLBLM_R_X11Y133_SLICE_X14Y133_DLUT (
.I0(CLBLM_R_X11Y131_SLICE_X15Y131_BQ),
.I1(CLBLM_L_X10Y131_SLICE_X13Y131_CQ),
.I2(CLBLM_R_X5Y132_SLICE_X7Y132_DO6),
.I3(CLBLM_L_X10Y137_SLICE_X12Y137_BQ),
.I4(CLBLM_R_X11Y133_SLICE_X15Y133_DQ),
.I5(CLBLM_L_X10Y133_SLICE_X12Y133_DO6),
.O5(CLBLM_R_X11Y133_SLICE_X14Y133_DO5),
.O6(CLBLM_R_X11Y133_SLICE_X14Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcf0fcf00c000c00)
  ) CLBLM_R_X11Y133_SLICE_X14Y133_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y133_SLICE_X14Y133_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(1'b1),
.I5(CLBLM_R_X7Y134_SLICE_X8Y134_AQ),
.O5(CLBLM_R_X11Y133_SLICE_X14Y133_CO5),
.O6(CLBLM_R_X11Y133_SLICE_X14Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fff0fc000f000c)
  ) CLBLM_R_X11Y133_SLICE_X14Y133_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y133_SLICE_X14Y133_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X5Y134_SLICE_X7Y134_DO6),
.I4(CLBLM_R_X11Y132_SLICE_X14Y132_AQ),
.I5(CLBLM_R_X11Y140_SLICE_X14Y140_AQ),
.O5(CLBLM_R_X11Y133_SLICE_X14Y133_BO5),
.O6(CLBLM_R_X11Y133_SLICE_X14Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000000fc00fc)
  ) CLBLM_R_X11Y133_SLICE_X14Y133_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y133_SLICE_X14Y133_BQ),
.I2(CLBLM_R_X11Y133_SLICE_X14Y133_AQ),
.I3(CLBLM_R_X5Y134_SLICE_X7Y134_DO6),
.I4(CLBLM_L_X10Y142_SLICE_X13Y142_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y133_SLICE_X14Y133_AO5),
.O6(CLBLM_R_X11Y133_SLICE_X14Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y133_SLICE_X15Y133_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y133_SLICE_X15Y133_AO6),
.Q(CLBLM_R_X11Y133_SLICE_X15Y133_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y133_SLICE_X15Y133_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y133_SLICE_X15Y133_BO6),
.Q(CLBLM_R_X11Y133_SLICE_X15Y133_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y133_SLICE_X15Y133_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y133_SLICE_X15Y133_CO6),
.Q(CLBLM_R_X11Y133_SLICE_X15Y133_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y133_SLICE_X15Y133_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y133_SLICE_X15Y133_DO6),
.Q(CLBLM_R_X11Y133_SLICE_X15Y133_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0a0fcccc0a0f)
  ) CLBLM_R_X11Y133_SLICE_X15Y133_DLUT (
.I0(CLBLM_R_X7Y131_SLICE_X9Y131_AQ),
.I1(CLBLM_L_X12Y133_SLICE_X17Y133_BQ),
.I2(CLBLM_R_X11Y133_SLICE_X14Y133_DO6),
.I3(RIOB33_X105Y141_IOB_X1Y142_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y133_SLICE_X15Y133_DO5),
.O6(CLBLM_R_X11Y133_SLICE_X15Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00fe54aa00fe54)
  ) CLBLM_R_X11Y133_SLICE_X15Y133_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X11Y133_SLICE_X15Y133_CQ),
.I2(CLBLM_R_X11Y134_SLICE_X15Y134_CQ),
.I3(CLBLM_R_X11Y140_SLICE_X15Y140_BQ),
.I4(CLBLM_R_X5Y132_SLICE_X7Y132_DO6),
.I5(1'b1),
.O5(CLBLM_R_X11Y133_SLICE_X15Y133_CO5),
.O6(CLBLM_R_X11Y133_SLICE_X15Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaaee00550044)
  ) CLBLM_R_X11Y133_SLICE_X15Y133_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X11Y133_SLICE_X15Y133_BQ),
.I2(1'b1),
.I3(CLBLM_R_X5Y134_SLICE_X7Y134_DO6),
.I4(CLBLM_R_X7Y131_SLICE_X9Y131_BQ),
.I5(CLBLM_L_X12Y136_SLICE_X17Y136_CQ),
.O5(CLBLM_R_X11Y133_SLICE_X15Y133_BO5),
.O6(CLBLM_R_X11Y133_SLICE_X15Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haafeaafe00540054)
  ) CLBLM_R_X11Y133_SLICE_X15Y133_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X11Y133_SLICE_X15Y133_BQ),
.I2(CLBLM_R_X11Y133_SLICE_X15Y133_AQ),
.I3(CLBLM_R_X5Y133_SLICE_X7Y133_DO6),
.I4(1'b1),
.I5(CLBLM_L_X10Y140_SLICE_X12Y140_A5Q),
.O5(CLBLM_R_X11Y133_SLICE_X15Y133_AO5),
.O6(CLBLM_R_X11Y133_SLICE_X15Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y134_SLICE_X14Y134_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y134_SLICE_X14Y134_AO6),
.Q(CLBLM_R_X11Y134_SLICE_X14Y134_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y134_SLICE_X14Y134_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y134_SLICE_X14Y134_BO6),
.Q(CLBLM_R_X11Y134_SLICE_X14Y134_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y134_SLICE_X14Y134_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y134_SLICE_X14Y134_CO6),
.Q(CLBLM_R_X11Y134_SLICE_X14Y134_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y134_SLICE_X14Y134_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y134_SLICE_X14Y134_DO6),
.Q(CLBLM_R_X11Y134_SLICE_X14Y134_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0022222222)
  ) CLBLM_R_X11Y134_SLICE_X14Y134_DLUT (
.I0(CLBLM_R_X11Y136_SLICE_X15Y136_AQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(1'b1),
.I3(CLBLM_L_X10Y131_SLICE_X12Y131_BQ),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y134_SLICE_X14Y134_DO5),
.O6(CLBLM_R_X11Y134_SLICE_X14Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff00008f808f80)
  ) CLBLM_R_X11Y134_SLICE_X14Y134_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X11Y134_SLICE_X14Y134_CQ),
.I2(CLBLM_L_X10Y135_SLICE_X12Y135_DO6),
.I3(CLBLM_R_X13Y134_SLICE_X19Y134_AQ),
.I4(CLBLM_L_X10Y138_SLICE_X13Y138_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y134_SLICE_X14Y134_CO5),
.O6(CLBLM_R_X11Y134_SLICE_X14Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffd800d8ff500050)
  ) CLBLM_R_X11Y134_SLICE_X14Y134_BLUT (
.I0(CLBLM_L_X10Y135_SLICE_X12Y135_DO6),
.I1(CLBLM_R_X11Y134_SLICE_X14Y134_BQ),
.I2(CLBLM_R_X11Y134_SLICE_X14Y134_CQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLL_L_X4Y138_SLICE_X5Y138_BQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X11Y134_SLICE_X14Y134_BO5),
.O6(CLBLM_R_X11Y134_SLICE_X14Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdec3120ddcc1100)
  ) CLBLM_R_X11Y134_SLICE_X14Y134_ALUT (
.I0(CLBLM_L_X10Y135_SLICE_X12Y135_DO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X11Y134_SLICE_X14Y134_AQ),
.I3(CLBLM_L_X12Y135_SLICE_X16Y135_BQ),
.I4(CLBLM_R_X5Y136_SLICE_X7Y136_BQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X11Y134_SLICE_X14Y134_AO5),
.O6(CLBLM_R_X11Y134_SLICE_X14Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y134_SLICE_X15Y134_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y134_SLICE_X15Y134_AO6),
.Q(CLBLM_R_X11Y134_SLICE_X15Y134_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y134_SLICE_X15Y134_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y134_SLICE_X15Y134_BO6),
.Q(CLBLM_R_X11Y134_SLICE_X15Y134_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y134_SLICE_X15Y134_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y134_SLICE_X15Y134_CO6),
.Q(CLBLM_R_X11Y134_SLICE_X15Y134_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6699669999669966)
  ) CLBLM_R_X11Y134_SLICE_X15Y134_DLUT (
.I0(CLBLM_L_X8Y132_SLICE_X11Y132_BQ),
.I1(CLBLM_R_X11Y139_SLICE_X14Y139_AQ),
.I2(1'b1),
.I3(CLBLM_L_X8Y134_SLICE_X11Y134_AQ),
.I4(1'b1),
.I5(CLBLM_R_X7Y133_SLICE_X9Y133_AQ),
.O5(CLBLM_R_X11Y134_SLICE_X15Y134_DO5),
.O6(CLBLM_R_X11Y134_SLICE_X15Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f055554444)
  ) CLBLM_R_X11Y134_SLICE_X15Y134_CLUT (
.I0(CLBLM_R_X5Y133_SLICE_X7Y133_DO6),
.I1(CLBLM_R_X11Y134_SLICE_X15Y134_CQ),
.I2(CLBLM_L_X12Y138_SLICE_X17Y138_AQ),
.I3(1'b1),
.I4(CLBLM_L_X10Y134_SLICE_X12Y134_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y134_SLICE_X15Y134_CO5),
.O6(CLBLM_R_X11Y134_SLICE_X15Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000aaacaaac)
  ) CLBLM_R_X11Y134_SLICE_X15Y134_BLUT (
.I0(CLBLM_L_X8Y134_SLICE_X11Y134_CQ),
.I1(CLBLM_R_X11Y134_SLICE_X15Y134_BQ),
.I2(RIOB33_X105Y117_IOB_X1Y118_I),
.I3(CLBLM_L_X8Y138_SLICE_X10Y138_AQ),
.I4(CLBLM_R_X11Y139_SLICE_X15Y139_BQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y134_SLICE_X15Y134_BO5),
.O6(CLBLM_R_X11Y134_SLICE_X15Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffcc00ccf0cc00)
  ) CLBLM_R_X11Y134_SLICE_X15Y134_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y133_SLICE_X11Y133_BQ),
.I2(CLBLM_R_X11Y134_SLICE_X15Y134_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y143_SLICE_X10Y143_DO6),
.I5(CLBLM_L_X8Y140_SLICE_X11Y140_AQ),
.O5(CLBLM_R_X11Y134_SLICE_X15Y134_AO5),
.O6(CLBLM_R_X11Y134_SLICE_X15Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y135_SLICE_X14Y135_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y135_SLICE_X14Y135_AO6),
.Q(CLBLM_R_X11Y135_SLICE_X14Y135_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y135_SLICE_X14Y135_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y135_SLICE_X14Y135_BO6),
.Q(CLBLM_R_X11Y135_SLICE_X14Y135_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y135_SLICE_X14Y135_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y135_SLICE_X14Y135_CO6),
.Q(CLBLM_R_X11Y135_SLICE_X14Y135_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y135_SLICE_X14Y135_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y135_SLICE_X14Y135_DO6),
.Q(CLBLM_R_X11Y135_SLICE_X14Y135_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaaf0aaccaac0)
  ) CLBLM_R_X11Y135_SLICE_X14Y135_DLUT (
.I0(CLBLM_R_X11Y133_SLICE_X14Y133_AQ),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_R_X11Y135_SLICE_X14Y135_DQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y135_SLICE_X13Y135_CO6),
.I5(CLBLM_L_X8Y138_SLICE_X10Y138_AQ),
.O5(CLBLM_R_X11Y135_SLICE_X14Y135_DO5),
.O6(CLBLM_R_X11Y135_SLICE_X14Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf033f022f000f000)
  ) CLBLM_R_X11Y135_SLICE_X14Y135_CLUT (
.I0(CLBLM_R_X11Y132_SLICE_X14Y132_BQ),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_L_X8Y136_SLICE_X11Y136_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X11Y135_SLICE_X14Y135_CQ),
.I5(CLBLM_L_X8Y138_SLICE_X10Y138_AQ),
.O5(CLBLM_R_X11Y135_SLICE_X14Y135_CO5),
.O6(CLBLM_R_X11Y135_SLICE_X14Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000aaacaaac)
  ) CLBLM_R_X11Y135_SLICE_X14Y135_BLUT (
.I0(CLBLM_R_X11Y135_SLICE_X14Y135_CQ),
.I1(CLBLM_R_X11Y135_SLICE_X14Y135_BQ),
.I2(RIOB33_X105Y117_IOB_X1Y118_I),
.I3(CLBLM_L_X8Y138_SLICE_X10Y138_AQ),
.I4(CLBLM_L_X10Y144_SLICE_X12Y144_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y135_SLICE_X14Y135_BO5),
.O6(CLBLM_R_X11Y135_SLICE_X14Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haafcaafcaafcaa00)
  ) CLBLM_R_X11Y135_SLICE_X14Y135_ALUT (
.I0(CLBLM_R_X11Y135_SLICE_X14Y135_CQ),
.I1(CLBLM_R_X11Y138_SLICE_X14Y138_D5Q),
.I2(CLBLM_R_X11Y135_SLICE_X14Y135_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLM_L_X8Y138_SLICE_X10Y138_AQ),
.O5(CLBLM_R_X11Y135_SLICE_X14Y135_AO5),
.O6(CLBLM_R_X11Y135_SLICE_X14Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y135_SLICE_X15Y135_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y135_SLICE_X15Y135_AO6),
.Q(CLBLM_R_X11Y135_SLICE_X15Y135_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y135_SLICE_X15Y135_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y135_SLICE_X15Y135_BO6),
.Q(CLBLM_R_X11Y135_SLICE_X15Y135_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h010004050b0a0e0f)
  ) CLBLM_R_X11Y135_SLICE_X15Y135_DLUT (
.I0(CLBLM_R_X5Y132_SLICE_X7Y132_DO6),
.I1(CLBLM_R_X11Y131_SLICE_X15Y131_AO5),
.I2(CLBLM_L_X10Y139_SLICE_X13Y139_CQ),
.I3(CLBLM_R_X11Y131_SLICE_X15Y131_BQ),
.I4(CLBLM_R_X11Y133_SLICE_X15Y133_AQ),
.I5(CLBLM_R_X13Y137_SLICE_X18Y137_A5Q),
.O5(CLBLM_R_X11Y135_SLICE_X15Y135_DO5),
.O6(CLBLM_R_X11Y135_SLICE_X15Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f07030000ff00)
  ) CLBLM_R_X11Y135_SLICE_X15Y135_CLUT (
.I0(CLBLL_L_X4Y139_SLICE_X4Y139_BO6),
.I1(CLBLM_L_X10Y134_SLICE_X12Y134_CQ),
.I2(CLBLM_L_X12Y135_SLICE_X17Y135_A5Q),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLL_L_X4Y134_SLICE_X4Y134_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y135_SLICE_X15Y135_CO5),
.O6(CLBLM_R_X11Y135_SLICE_X15Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff008888ff008888)
  ) CLBLM_R_X11Y135_SLICE_X15Y135_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X8Y133_SLICE_X11Y133_BQ),
.I2(1'b1),
.I3(CLBLM_L_X10Y136_SLICE_X12Y136_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y135_SLICE_X15Y135_BO5),
.O6(CLBLM_R_X11Y135_SLICE_X15Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdddc1110cccc0000)
  ) CLBLM_R_X11Y135_SLICE_X15Y135_ALUT (
.I0(CLBLM_R_X11Y136_SLICE_X14Y136_DQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X11Y135_SLICE_X15Y135_AQ),
.I3(CLBLM_L_X8Y135_SLICE_X11Y135_CQ),
.I4(CLBLM_R_X13Y137_SLICE_X19Y137_AQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X11Y135_SLICE_X15Y135_AO5),
.O6(CLBLM_R_X11Y135_SLICE_X15Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y136_SLICE_X14Y136_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y136_SLICE_X14Y136_AO6),
.Q(CLBLM_R_X11Y136_SLICE_X14Y136_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y136_SLICE_X14Y136_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y136_SLICE_X14Y136_BO6),
.Q(CLBLM_R_X11Y136_SLICE_X14Y136_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y136_SLICE_X14Y136_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y136_SLICE_X14Y136_DO6),
.Q(CLBLM_R_X11Y136_SLICE_X14Y136_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00ba10aa00)
  ) CLBLM_R_X11Y136_SLICE_X14Y136_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X13Y137_SLICE_X18Y137_AQ),
.I3(CLBLM_R_X11Y136_SLICE_X14Y136_BQ),
.I4(CLBLM_R_X11Y135_SLICE_X15Y135_AQ),
.I5(CLBLM_L_X10Y136_SLICE_X13Y136_AO6),
.O5(CLBLM_R_X11Y136_SLICE_X14Y136_DO5),
.O6(CLBLM_R_X11Y136_SLICE_X14Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hee44ea40ccccc0c0)
  ) CLBLM_R_X11Y136_SLICE_X14Y136_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y121_IOB_X1Y121_I),
.I2(CLBLM_L_X10Y141_SLICE_X13Y141_BQ),
.I3(CLBLM_R_X11Y133_SLICE_X15Y133_DQ),
.I4(CLBLM_L_X12Y136_SLICE_X17Y136_CQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y136_SLICE_X14Y136_CO5),
.O6(CLBLM_R_X11Y136_SLICE_X14Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc0cf404fc0cf404)
  ) CLBLM_R_X11Y136_SLICE_X14Y136_BLUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_R_X11Y136_SLICE_X14Y136_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X11Y138_SLICE_X14Y138_D5Q),
.I4(CLBLM_L_X8Y138_SLICE_X10Y138_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y136_SLICE_X14Y136_BO5),
.O6(CLBLM_R_X11Y136_SLICE_X14Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00de12cc00de12)
  ) CLBLM_R_X11Y136_SLICE_X14Y136_ALUT (
.I0(CLBLM_R_X7Y139_SLICE_X9Y139_BO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X11Y136_SLICE_X14Y136_AQ),
.I3(CLBLM_R_X13Y136_SLICE_X18Y136_AQ),
.I4(CLBLM_R_X11Y135_SLICE_X14Y135_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y136_SLICE_X14Y136_AO5),
.O6(CLBLM_R_X11Y136_SLICE_X14Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y136_SLICE_X15Y136_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y136_SLICE_X15Y136_AO5),
.Q(CLBLM_R_X11Y136_SLICE_X15Y136_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y136_SLICE_X15Y136_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y136_SLICE_X15Y136_BO5),
.Q(CLBLM_R_X11Y136_SLICE_X15Y136_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y136_SLICE_X15Y136_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y136_SLICE_X15Y136_AO6),
.Q(CLBLM_R_X11Y136_SLICE_X15Y136_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y136_SLICE_X15Y136_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y136_SLICE_X15Y136_BO6),
.Q(CLBLM_R_X11Y136_SLICE_X15Y136_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffeeffee)
  ) CLBLM_R_X11Y136_SLICE_X15Y136_DLUT (
.I0(CLBLM_L_X8Y136_SLICE_X10Y136_CQ),
.I1(CLBLM_L_X8Y135_SLICE_X11Y135_A5Q),
.I2(1'b1),
.I3(CLBLM_R_X13Y136_SLICE_X18Y136_CQ),
.I4(1'b1),
.I5(CLBLM_R_X11Y135_SLICE_X15Y135_BQ),
.O5(CLBLM_R_X11Y136_SLICE_X15Y136_DO5),
.O6(CLBLM_R_X11Y136_SLICE_X15Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hc8dd0000ccdd0000)
  ) CLBLM_R_X11Y136_SLICE_X15Y136_CLUT (
.I0(CLBLL_L_X4Y134_SLICE_X4Y134_AQ),
.I1(CLBLM_R_X11Y137_SLICE_X14Y137_CO5),
.I2(CLBLM_R_X5Y141_SLICE_X7Y141_DO6),
.I3(CLBLM_L_X10Y134_SLICE_X12Y134_CQ),
.I4(CLBLM_L_X12Y135_SLICE_X17Y135_BO5),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X11Y136_SLICE_X15Y136_CO5),
.O6(CLBLM_R_X11Y136_SLICE_X15Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haca0aca0cfcfc0c0)
  ) CLBLM_R_X11Y136_SLICE_X15Y136_BLUT (
.I0(CLBLM_L_X8Y132_SLICE_X10Y132_AQ),
.I1(CLBLM_R_X11Y136_SLICE_X15Y136_A5Q),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_L_X10Y141_SLICE_X13Y141_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y136_SLICE_X15Y136_BO5),
.O6(CLBLM_R_X11Y136_SLICE_X15Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf022f022aa33aa00)
  ) CLBLM_R_X11Y136_SLICE_X15Y136_ALUT (
.I0(CLBLM_R_X13Y136_SLICE_X18Y136_CQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_L_X10Y139_SLICE_X13Y139_CQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X5Y140_SLICE_X7Y140_BQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y136_SLICE_X15Y136_AO5),
.O6(CLBLM_R_X11Y136_SLICE_X15Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y137_SLICE_X14Y137_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y137_SLICE_X14Y137_AO6),
.Q(CLBLM_R_X11Y137_SLICE_X14Y137_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hee40ee0000000000)
  ) CLBLM_R_X11Y137_SLICE_X14Y137_DLUT (
.I0(CLBLL_L_X4Y134_SLICE_X4Y134_AQ),
.I1(CLBLM_L_X10Y134_SLICE_X12Y134_CQ),
.I2(CLBLL_L_X4Y142_SLICE_X5Y142_DO6),
.I3(CLBLM_R_X11Y137_SLICE_X14Y137_CO6),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_L_X12Y135_SLICE_X17Y135_BO5),
.O5(CLBLM_R_X11Y137_SLICE_X14Y137_DO5),
.O6(CLBLM_R_X11Y137_SLICE_X14Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfc0000ff00aaaa)
  ) CLBLM_R_X11Y137_SLICE_X14Y137_CLUT (
.I0(CLBLM_R_X11Y138_SLICE_X14Y138_AQ),
.I1(CLBLM_R_X7Y139_SLICE_X8Y139_A5Q),
.I2(CLBLM_L_X10Y138_SLICE_X13Y138_AQ),
.I3(CLBLM_L_X10Y141_SLICE_X13Y141_BQ),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y137_SLICE_X14Y137_CO5),
.O6(CLBLM_R_X11Y137_SLICE_X14Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbb88888fff00000)
  ) CLBLM_R_X11Y137_SLICE_X14Y137_BLUT (
.I0(CLBLM_R_X11Y133_SLICE_X15Y133_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X7Y136_SLICE_X9Y136_AQ),
.I3(CLBLM_L_X8Y135_SLICE_X11Y135_A5Q),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y137_SLICE_X14Y137_BO5),
.O6(CLBLM_R_X11Y137_SLICE_X14Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a3a3a3a3a0a0)
  ) CLBLM_R_X11Y137_SLICE_X14Y137_ALUT (
.I0(CLBLM_L_X12Y137_SLICE_X16Y137_A5Q),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(CLBLM_R_X11Y137_SLICE_X14Y137_CO5),
.I5(CLBLM_R_X7Y134_SLICE_X8Y134_AQ),
.O5(CLBLM_R_X11Y137_SLICE_X14Y137_AO5),
.O6(CLBLM_R_X11Y137_SLICE_X14Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y137_SLICE_X15Y137_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y137_SLICE_X15Y137_AO6),
.Q(CLBLM_R_X11Y137_SLICE_X15Y137_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffefffefffefffe)
  ) CLBLM_R_X11Y137_SLICE_X15Y137_DLUT (
.I0(CLBLM_R_X11Y136_SLICE_X15Y136_A5Q),
.I1(CLBLM_L_X12Y139_SLICE_X16Y139_CQ),
.I2(CLBLM_R_X11Y138_SLICE_X15Y138_CQ),
.I3(CLBLM_L_X8Y139_SLICE_X11Y139_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y137_SLICE_X15Y137_DO5),
.O6(CLBLM_R_X11Y137_SLICE_X15Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffffcc)
  ) CLBLM_R_X11Y137_SLICE_X15Y137_CLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y135_SLICE_X12Y135_BQ),
.I2(1'b1),
.I3(CLBLM_R_X5Y140_SLICE_X7Y140_BQ),
.I4(CLBLM_L_X12Y136_SLICE_X16Y136_AQ),
.I5(CLBLM_R_X7Y139_SLICE_X8Y139_BQ),
.O5(CLBLM_R_X11Y137_SLICE_X15Y137_CO5),
.O6(CLBLM_R_X11Y137_SLICE_X15Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_R_X11Y137_SLICE_X15Y137_BLUT (
.I0(CLBLM_R_X11Y136_SLICE_X15Y136_DO6),
.I1(CLBLM_R_X11Y138_SLICE_X15Y138_AQ),
.I2(CLBLM_R_X5Y137_SLICE_X7Y137_CQ),
.I3(CLBLM_R_X11Y137_SLICE_X15Y137_DO6),
.I4(CLBLM_R_X11Y136_SLICE_X15Y136_AQ),
.I5(CLBLM_R_X11Y137_SLICE_X15Y137_CO6),
.O5(CLBLM_R_X11Y137_SLICE_X15Y137_BO5),
.O6(CLBLM_R_X11Y137_SLICE_X15Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffccfff0ffccffa0)
  ) CLBLM_R_X11Y137_SLICE_X15Y137_ALUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_L_X10Y137_SLICE_X12Y137_CQ),
.I2(CLBLM_R_X11Y137_SLICE_X15Y137_AQ),
.I3(CLBLM_R_X11Y137_SLICE_X14Y137_DO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y138_SLICE_X10Y138_AQ),
.O5(CLBLM_R_X11Y137_SLICE_X15Y137_AO5),
.O6(CLBLM_R_X11Y137_SLICE_X15Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y138_SLICE_X14Y138_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y138_SLICE_X14Y138_DO5),
.Q(CLBLM_R_X11Y138_SLICE_X14Y138_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y138_SLICE_X14Y138_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y138_SLICE_X14Y138_AO6),
.Q(CLBLM_R_X11Y138_SLICE_X14Y138_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y138_SLICE_X14Y138_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y138_SLICE_X14Y138_BO6),
.Q(CLBLM_R_X11Y138_SLICE_X14Y138_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y138_SLICE_X14Y138_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y138_SLICE_X14Y138_CO6),
.Q(CLBLM_R_X11Y138_SLICE_X14Y138_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y138_SLICE_X14Y138_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y138_SLICE_X14Y138_DO6),
.Q(CLBLM_R_X11Y138_SLICE_X14Y138_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc0fcc00aaccaaff)
  ) CLBLM_R_X11Y138_SLICE_X14Y138_DLUT (
.I0(CLBLM_R_X5Y135_SLICE_X6Y135_BQ),
.I1(CLBLM_L_X8Y138_SLICE_X10Y138_DQ),
.I2(CLBLM_R_X11Y138_SLICE_X14Y138_DQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y119_IOB_X1Y119_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y138_SLICE_X14Y138_DO5),
.O6(CLBLM_R_X11Y138_SLICE_X14Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f055f055f000)
  ) CLBLM_R_X11Y138_SLICE_X14Y138_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(1'b1),
.I2(CLBLM_R_X11Y136_SLICE_X14Y136_DQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X11Y140_SLICE_X15Y140_DQ),
.I5(CLBLM_L_X10Y135_SLICE_X13Y135_AO5),
.O5(CLBLM_R_X11Y138_SLICE_X14Y138_CO5),
.O6(CLBLM_R_X11Y138_SLICE_X14Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0006600cc)
  ) CLBLM_R_X11Y138_SLICE_X14Y138_BLUT (
.I0(CLBLM_R_X7Y139_SLICE_X9Y139_BO6),
.I1(CLBLM_R_X11Y138_SLICE_X14Y138_BQ),
.I2(CLBLM_R_X11Y138_SLICE_X14Y138_AQ),
.I3(CLBLM_R_X11Y135_SLICE_X14Y135_AQ),
.I4(CLBLM_R_X11Y136_SLICE_X14Y136_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y138_SLICE_X14Y138_BO5),
.O6(CLBLM_R_X11Y138_SLICE_X14Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8888bbbb88b8bbb8)
  ) CLBLM_R_X11Y138_SLICE_X14Y138_ALUT (
.I0(CLBLM_L_X12Y139_SLICE_X17Y139_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X11Y138_SLICE_X14Y138_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_L_X10Y138_SLICE_X12Y138_BO6),
.I5(CLBLM_L_X8Y138_SLICE_X10Y138_AQ),
.O5(CLBLM_R_X11Y138_SLICE_X14Y138_AO5),
.O6(CLBLM_R_X11Y138_SLICE_X14Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y138_SLICE_X15Y138_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y138_SLICE_X15Y138_BO5),
.Q(CLBLM_R_X11Y138_SLICE_X15Y138_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y138_SLICE_X15Y138_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y138_SLICE_X15Y138_DO5),
.Q(CLBLM_R_X11Y138_SLICE_X15Y138_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y138_SLICE_X15Y138_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y138_SLICE_X15Y138_AO6),
.Q(CLBLM_R_X11Y138_SLICE_X15Y138_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y138_SLICE_X15Y138_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y138_SLICE_X15Y138_BO6),
.Q(CLBLM_R_X11Y138_SLICE_X15Y138_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y138_SLICE_X15Y138_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y138_SLICE_X15Y138_CO6),
.Q(CLBLM_R_X11Y138_SLICE_X15Y138_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y138_SLICE_X15Y138_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y138_SLICE_X15Y138_DO6),
.Q(CLBLM_R_X11Y138_SLICE_X15Y138_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3c0f3c0bbbb8888)
  ) CLBLM_R_X11Y138_SLICE_X15Y138_DLUT (
.I0(CLBLM_L_X8Y136_SLICE_X10Y136_DQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X11Y142_SLICE_X15Y142_AQ),
.I3(CLBLM_L_X10Y141_SLICE_X13Y141_A5Q),
.I4(RIOB33_X105Y103_IOB_X1Y103_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y138_SLICE_X15Y138_DO5),
.O6(CLBLM_R_X11Y138_SLICE_X15Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00ee22ee22)
  ) CLBLM_R_X11Y138_SLICE_X15Y138_CLUT (
.I0(CLBLM_R_X5Y137_SLICE_X7Y137_CQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(1'b1),
.I3(CLBLM_L_X12Y135_SLICE_X17Y135_A5Q),
.I4(1'b1),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X11Y138_SLICE_X15Y138_CO5),
.O6(CLBLM_R_X11Y138_SLICE_X15Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff33cc00cece0202)
  ) CLBLM_R_X11Y138_SLICE_X15Y138_BLUT (
.I0(CLBLM_R_X11Y138_SLICE_X15Y138_B5Q),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X11Y138_SLICE_X15Y138_D5Q),
.I4(CLBLM_L_X12Y138_SLICE_X16Y138_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y138_SLICE_X15Y138_BO5),
.O6(CLBLM_R_X11Y138_SLICE_X15Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0f00cccc0f00)
  ) CLBLM_R_X11Y138_SLICE_X15Y138_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y138_SLICE_X15Y138_BQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_L_X10Y141_SLICE_X13Y141_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y138_SLICE_X15Y138_AO5),
.O6(CLBLM_R_X11Y138_SLICE_X15Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y139_SLICE_X14Y139_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y139_SLICE_X14Y139_BO5),
.Q(CLBLM_R_X11Y139_SLICE_X14Y139_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y139_SLICE_X14Y139_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y139_SLICE_X14Y139_AO6),
.Q(CLBLM_R_X11Y139_SLICE_X14Y139_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y139_SLICE_X14Y139_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y139_SLICE_X14Y139_BO6),
.Q(CLBLM_R_X11Y139_SLICE_X14Y139_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y139_SLICE_X14Y139_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y139_SLICE_X14Y139_CO6),
.Q(CLBLM_R_X11Y139_SLICE_X14Y139_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000ff00ff00)
  ) CLBLM_R_X11Y139_SLICE_X14Y139_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X11Y139_SLICE_X15Y139_CQ),
.I4(1'b1),
.I5(CLBLM_L_X10Y139_SLICE_X13Y139_AQ),
.O5(CLBLM_R_X11Y139_SLICE_X14Y139_DO5),
.O6(CLBLM_R_X11Y139_SLICE_X14Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haafeaaaa00540000)
  ) CLBLM_R_X11Y139_SLICE_X14Y139_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X11Y139_SLICE_X14Y139_CQ),
.I2(CLBLM_L_X8Y137_SLICE_X11Y137_CO6),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_L_X8Y138_SLICE_X10Y138_AQ),
.I5(CLBLM_L_X10Y138_SLICE_X13Y138_BQ),
.O5(CLBLM_R_X11Y139_SLICE_X14Y139_CO5),
.O6(CLBLM_R_X11Y139_SLICE_X14Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hea40ea40dddd8888)
  ) CLBLM_R_X11Y139_SLICE_X14Y139_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X11Y139_SLICE_X14Y139_BQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_L_X12Y133_SLICE_X16Y133_BQ),
.I4(CLBLM_R_X7Y141_SLICE_X8Y141_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y139_SLICE_X14Y139_BO5),
.O6(CLBLM_R_X11Y139_SLICE_X14Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heeee2222eefc2230)
  ) CLBLM_R_X11Y139_SLICE_X14Y139_ALUT (
.I0(CLBLM_R_X11Y140_SLICE_X14Y140_CQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X11Y139_SLICE_X14Y139_AQ),
.I3(CLBLM_L_X8Y138_SLICE_X10Y138_AQ),
.I4(CLBLM_R_X7Y136_SLICE_X9Y136_AQ),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_R_X11Y139_SLICE_X14Y139_AO5),
.O6(CLBLM_R_X11Y139_SLICE_X14Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y139_SLICE_X15Y139_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y139_SLICE_X15Y139_AO5),
.Q(CLBLM_R_X11Y139_SLICE_X15Y139_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y139_SLICE_X15Y139_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y139_SLICE_X15Y139_AO6),
.Q(CLBLM_R_X11Y139_SLICE_X15Y139_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y139_SLICE_X15Y139_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y139_SLICE_X15Y139_BO6),
.Q(CLBLM_R_X11Y139_SLICE_X15Y139_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y139_SLICE_X15Y139_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y139_SLICE_X15Y139_CO6),
.Q(CLBLM_R_X11Y139_SLICE_X15Y139_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y139_SLICE_X15Y139_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y139_SLICE_X15Y139_DO6),
.Q(CLBLM_R_X11Y139_SLICE_X15Y139_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0011114444)
  ) CLBLM_R_X11Y139_SLICE_X15Y139_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X12Y139_SLICE_X16Y139_DO5),
.I2(1'b1),
.I3(CLBLM_R_X11Y138_SLICE_X15Y138_AQ),
.I4(CLBLM_R_X11Y140_SLICE_X15Y140_BQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y139_SLICE_X15Y139_DO5),
.O6(CLBLM_R_X11Y139_SLICE_X15Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaee0044aaaa0000)
  ) CLBLM_R_X11Y139_SLICE_X15Y139_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X11Y139_SLICE_X15Y139_CQ),
.I2(1'b1),
.I3(CLBLM_R_X7Y139_SLICE_X9Y139_AQ),
.I4(CLBLM_R_X11Y139_SLICE_X15Y139_AQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X11Y139_SLICE_X15Y139_CO5),
.O6(CLBLM_R_X11Y139_SLICE_X15Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00fc30cc00fc30)
  ) CLBLM_R_X11Y139_SLICE_X15Y139_BLUT (
.I0(1'b1),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X11Y139_SLICE_X15Y139_AQ),
.I3(CLBLM_R_X11Y139_SLICE_X15Y139_DQ),
.I4(CLBLM_R_X13Y141_SLICE_X18Y141_AO6),
.I5(1'b1),
.O5(CLBLM_R_X11Y139_SLICE_X15Y139_BO5),
.O6(CLBLM_R_X11Y139_SLICE_X15Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0acacfa0afa0a)
  ) CLBLM_R_X11Y139_SLICE_X15Y139_ALUT (
.I0(CLBLM_R_X11Y138_SLICE_X15Y138_DQ),
.I1(CLBLM_L_X12Y140_SLICE_X16Y140_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y135_SLICE_X12Y135_BQ),
.I4(CLBLM_R_X13Y141_SLICE_X18Y141_AO6),
.I5(1'b1),
.O5(CLBLM_R_X11Y139_SLICE_X15Y139_AO5),
.O6(CLBLM_R_X11Y139_SLICE_X15Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y140_SLICE_X14Y140_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y140_SLICE_X14Y140_AO6),
.Q(CLBLM_R_X11Y140_SLICE_X14Y140_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y140_SLICE_X14Y140_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y140_SLICE_X14Y140_BO6),
.Q(CLBLM_R_X11Y140_SLICE_X14Y140_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y140_SLICE_X14Y140_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y140_SLICE_X14Y140_CO6),
.Q(CLBLM_R_X11Y140_SLICE_X14Y140_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffff55)
  ) CLBLM_R_X11Y140_SLICE_X14Y140_DLUT (
.I0(CLBLM_L_X10Y140_SLICE_X13Y140_DQ),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_L_X12Y138_SLICE_X16Y138_DQ),
.I4(CLBLM_R_X11Y140_SLICE_X15Y140_DQ),
.I5(CLBLM_R_X11Y138_SLICE_X14Y138_CQ),
.O5(CLBLM_R_X11Y140_SLICE_X14Y140_DO5),
.O6(CLBLM_R_X11Y140_SLICE_X14Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff504000005040)
  ) CLBLM_R_X11Y140_SLICE_X14Y140_CLUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_R_X11Y140_SLICE_X14Y140_CQ),
.I2(CLBLM_L_X8Y138_SLICE_X10Y138_AQ),
.I3(CLBLM_L_X10Y139_SLICE_X13Y139_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X11Y142_SLICE_X14Y142_BQ),
.O5(CLBLM_R_X11Y140_SLICE_X14Y140_CO5),
.O6(CLBLM_R_X11Y140_SLICE_X14Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf044f0fff044f000)
  ) CLBLM_R_X11Y140_SLICE_X14Y140_BLUT (
.I0(CLBLM_R_X13Y143_SLICE_X18Y143_AO6),
.I1(CLBLM_R_X11Y140_SLICE_X14Y140_BQ),
.I2(CLBLM_R_X11Y136_SLICE_X14Y136_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X12Y143_SLICE_X17Y143_CO5),
.I5(CLBLM_L_X12Y140_SLICE_X17Y140_CQ),
.O5(CLBLM_R_X11Y140_SLICE_X14Y140_BO5),
.O6(CLBLM_R_X11Y140_SLICE_X14Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff50cc000050cc)
  ) CLBLM_R_X11Y140_SLICE_X14Y140_ALUT (
.I0(CLBLM_R_X13Y143_SLICE_X18Y143_AO6),
.I1(CLBLM_R_X11Y140_SLICE_X14Y140_BQ),
.I2(CLBLM_R_X11Y140_SLICE_X14Y140_AQ),
.I3(CLBLM_L_X12Y143_SLICE_X17Y143_CO5),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y140_SLICE_X9Y140_CQ),
.O5(CLBLM_R_X11Y140_SLICE_X14Y140_AO5),
.O6(CLBLM_R_X11Y140_SLICE_X14Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y140_SLICE_X15Y140_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y140_SLICE_X15Y140_CO5),
.Q(CLBLM_R_X11Y140_SLICE_X15Y140_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y140_SLICE_X15Y140_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y140_SLICE_X15Y140_BO6),
.Q(CLBLM_R_X11Y140_SLICE_X15Y140_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y140_SLICE_X15Y140_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y140_SLICE_X15Y140_CO6),
.Q(CLBLM_R_X11Y140_SLICE_X15Y140_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y140_SLICE_X15Y140_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y140_SLICE_X15Y140_DO6),
.Q(CLBLM_R_X11Y140_SLICE_X15Y140_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h888888888b8bb8b8)
  ) CLBLM_R_X11Y140_SLICE_X15Y140_DLUT (
.I0(CLBLM_L_X12Y142_SLICE_X17Y142_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y140_SLICE_X12Y140_A5Q),
.I3(1'b1),
.I4(CLBLM_L_X12Y136_SLICE_X17Y136_BO5),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X11Y140_SLICE_X15Y140_DO5),
.O6(CLBLM_R_X11Y140_SLICE_X15Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaa00ccf0ccf0)
  ) CLBLM_R_X11Y140_SLICE_X15Y140_CLUT (
.I0(CLBLM_R_X11Y132_SLICE_X14Y132_BQ),
.I1(CLBLM_L_X12Y138_SLICE_X16Y138_DQ),
.I2(CLBLM_R_X11Y143_SLICE_X14Y143_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X12Y143_SLICE_X16Y143_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y140_SLICE_X15Y140_CO5),
.O6(CLBLM_R_X11Y140_SLICE_X15Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00af05aa00fa50)
  ) CLBLM_R_X11Y140_SLICE_X15Y140_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(1'b1),
.I2(CLBLM_L_X10Y140_SLICE_X13Y140_DQ),
.I3(CLBLM_L_X8Y142_SLICE_X11Y142_CQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X11Y140_SLICE_X15Y140_AO5),
.O5(CLBLM_R_X11Y140_SLICE_X15Y140_BO5),
.O6(CLBLM_R_X11Y140_SLICE_X15Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffc800c8c8c8c8c8)
  ) CLBLM_R_X11Y140_SLICE_X15Y140_ALUT (
.I0(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.I1(RIOB33_X105Y121_IOB_X1Y121_I),
.I2(CLBLM_R_X11Y136_SLICE_X15Y136_BQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X11Y140_SLICE_X15Y140_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X11Y140_SLICE_X15Y140_AO5),
.O6(CLBLM_R_X11Y140_SLICE_X15Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y141_SLICE_X14Y141_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y141_SLICE_X14Y141_AO6),
.Q(CLBLM_R_X11Y141_SLICE_X14Y141_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y141_SLICE_X14Y141_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y141_SLICE_X14Y141_BO6),
.Q(CLBLM_R_X11Y141_SLICE_X14Y141_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0ff0f00f0ff0f0)
  ) CLBLM_R_X11Y141_SLICE_X14Y141_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_L_X12Y144_SLICE_X17Y144_AQ),
.I3(1'b1),
.I4(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y141_SLICE_X14Y141_DO5),
.O6(CLBLM_R_X11Y141_SLICE_X14Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0e0e0e0e0f0f0f00)
  ) CLBLM_R_X11Y141_SLICE_X14Y141_CLUT (
.I0(CLBLM_R_X11Y141_SLICE_X14Y141_BQ),
.I1(CLBLM_R_X7Y133_SLICE_X9Y133_CQ),
.I2(CLBLM_R_X11Y138_SLICE_X14Y138_DQ),
.I3(CLBLM_R_X11Y139_SLICE_X14Y139_CQ),
.I4(CLBLM_L_X8Y133_SLICE_X11Y133_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y141_SLICE_X14Y141_CO5),
.O6(CLBLM_R_X11Y141_SLICE_X14Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f0f4f005000400)
  ) CLBLM_R_X11Y141_SLICE_X14Y141_BLUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_L_X10Y135_SLICE_X13Y135_CO6),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y138_SLICE_X10Y138_AQ),
.I4(CLBLM_R_X11Y141_SLICE_X14Y141_BQ),
.I5(CLBLM_R_X11Y143_SLICE_X15Y143_BQ),
.O5(CLBLM_R_X11Y141_SLICE_X14Y141_BO5),
.O6(CLBLM_R_X11Y141_SLICE_X14Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa0300c03c)
  ) CLBLM_R_X11Y141_SLICE_X14Y141_ALUT (
.I0(CLBLM_L_X10Y141_SLICE_X13Y141_AQ),
.I1(CLBLM_L_X12Y140_SLICE_X16Y140_DQ),
.I2(CLBLM_R_X11Y141_SLICE_X14Y141_AQ),
.I3(CLBLM_R_X11Y141_SLICE_X14Y141_DO6),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y141_SLICE_X14Y141_AO5),
.O6(CLBLM_R_X11Y141_SLICE_X14Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y141_SLICE_X15Y141_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y141_SLICE_X15Y141_AO6),
.Q(CLBLM_R_X11Y141_SLICE_X15Y141_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y141_SLICE_X15Y141_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y141_SLICE_X15Y141_BO6),
.Q(CLBLM_R_X11Y141_SLICE_X15Y141_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y141_SLICE_X15Y141_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y141_SLICE_X15Y141_CO6),
.Q(CLBLM_R_X11Y141_SLICE_X15Y141_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y141_SLICE_X15Y141_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y141_SLICE_X15Y141_DO6),
.Q(CLBLM_R_X11Y141_SLICE_X15Y141_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0000009999)
  ) CLBLM_R_X11Y141_SLICE_X15Y141_DLUT (
.I0(CLBLM_L_X10Y140_SLICE_X13Y140_BQ),
.I1(CLBLM_L_X12Y137_SLICE_X17Y137_BO5),
.I2(1'b1),
.I3(CLBLM_R_X11Y143_SLICE_X15Y143_AQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y141_SLICE_X15Y141_DO5),
.O6(CLBLM_R_X11Y141_SLICE_X15Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000c0cff00aaaa)
  ) CLBLM_R_X11Y141_SLICE_X15Y141_CLUT (
.I0(CLBLM_R_X11Y140_SLICE_X14Y140_AQ),
.I1(CLBLM_R_X11Y141_SLICE_X15Y141_CQ),
.I2(CLBLM_R_X13Y143_SLICE_X18Y143_AO6),
.I3(CLBLM_R_X11Y139_SLICE_X14Y139_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X12Y143_SLICE_X17Y143_CO5),
.O5(CLBLM_R_X11Y141_SLICE_X15Y141_CO5),
.O6(CLBLM_R_X11Y141_SLICE_X15Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00f0f0cccc)
  ) CLBLM_R_X11Y141_SLICE_X15Y141_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y141_SLICE_X15Y141_BQ),
.I2(CLBLM_R_X11Y140_SLICE_X15Y140_BQ),
.I3(CLBLM_R_X11Y141_SLICE_X14Y141_BQ),
.I4(CLBLM_L_X8Y143_SLICE_X10Y143_DO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y141_SLICE_X15Y141_BO5),
.O6(CLBLM_R_X11Y141_SLICE_X15Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00a2a2a0a0)
  ) CLBLM_R_X11Y141_SLICE_X15Y141_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(RIOB33_X105Y121_IOB_X1Y121_I),
.I2(CLBLM_R_X11Y141_SLICE_X15Y141_AQ),
.I3(CLBLM_L_X10Y131_SLICE_X13Y131_CQ),
.I4(CLBLM_R_X11Y136_SLICE_X14Y136_DQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y141_SLICE_X15Y141_AO5),
.O6(CLBLM_R_X11Y141_SLICE_X15Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y142_SLICE_X14Y142_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y142_SLICE_X14Y142_AO6),
.Q(CLBLM_R_X11Y142_SLICE_X14Y142_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y142_SLICE_X14Y142_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y142_SLICE_X14Y142_BO6),
.Q(CLBLM_R_X11Y142_SLICE_X14Y142_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_R_X11Y142_SLICE_X14Y142_DLUT (
.I0(CLBLM_R_X11Y142_SLICE_X15Y142_DQ),
.I1(CLBLM_R_X11Y144_SLICE_X14Y144_CO6),
.I2(CLBLM_L_X10Y143_SLICE_X12Y143_CQ),
.I3(CLBLM_R_X11Y142_SLICE_X15Y142_CQ),
.I4(CLBLM_R_X11Y143_SLICE_X15Y143_BQ),
.I5(CLBLM_L_X10Y142_SLICE_X13Y142_CQ),
.O5(CLBLM_R_X11Y142_SLICE_X14Y142_DO5),
.O6(CLBLM_R_X11Y142_SLICE_X14Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hc3c3c3c3c9c9c9c3)
  ) CLBLM_R_X11Y142_SLICE_X14Y142_CLUT (
.I0(CLBLM_R_X11Y142_SLICE_X15Y142_AQ),
.I1(CLBLM_R_X11Y142_SLICE_X14Y142_AQ),
.I2(CLBLM_L_X10Y144_SLICE_X13Y144_DO6),
.I3(CLBLM_R_X11Y143_SLICE_X15Y143_CO6),
.I4(CLBLM_R_X11Y142_SLICE_X14Y142_DO6),
.I5(CLBLM_L_X10Y145_SLICE_X12Y145_CO6),
.O5(CLBLM_R_X11Y142_SLICE_X14Y142_CO5),
.O6(CLBLM_R_X11Y142_SLICE_X14Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff004444f0f0)
  ) CLBLM_R_X11Y142_SLICE_X14Y142_BLUT (
.I0(CLBLM_R_X13Y143_SLICE_X18Y143_AO6),
.I1(CLBLM_R_X11Y142_SLICE_X14Y142_BQ),
.I2(CLBLM_R_X11Y141_SLICE_X15Y141_CQ),
.I3(CLBLL_L_X4Y134_SLICE_X5Y134_CQ),
.I4(CLBLM_L_X12Y143_SLICE_X17Y143_CO5),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y142_SLICE_X14Y142_BO5),
.O6(CLBLM_R_X11Y142_SLICE_X14Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h55055505dd0ddd0d)
  ) CLBLM_R_X11Y142_SLICE_X14Y142_ALUT (
.I0(CLBLM_R_X11Y144_SLICE_X14Y144_DO6),
.I1(CLBLM_L_X10Y144_SLICE_X12Y144_AO6),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X12Y136_SLICE_X17Y136_A5Q),
.I4(1'b1),
.I5(CLBLM_R_X11Y142_SLICE_X14Y142_CO6),
.O5(CLBLM_R_X11Y142_SLICE_X14Y142_AO5),
.O6(CLBLM_R_X11Y142_SLICE_X14Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y142_SLICE_X15Y142_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y142_SLICE_X15Y142_AO6),
.Q(CLBLM_R_X11Y142_SLICE_X15Y142_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y142_SLICE_X15Y142_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y142_SLICE_X15Y142_BO6),
.Q(CLBLM_R_X11Y142_SLICE_X15Y142_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y142_SLICE_X15Y142_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y142_SLICE_X15Y142_CO6),
.Q(CLBLM_R_X11Y142_SLICE_X15Y142_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y142_SLICE_X15Y142_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y142_SLICE_X15Y142_DO6),
.Q(CLBLM_R_X11Y142_SLICE_X15Y142_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8400cccca500ffff)
  ) CLBLM_R_X11Y142_SLICE_X15Y142_DLUT (
.I0(CLBLM_R_X11Y144_SLICE_X15Y144_CO6),
.I1(CLBLM_R_X11Y135_SLICE_X14Y135_DQ),
.I2(CLBLM_R_X11Y142_SLICE_X15Y142_DQ),
.I3(CLBLM_L_X10Y144_SLICE_X12Y144_AO6),
.I4(CLBLM_R_X11Y144_SLICE_X14Y144_DO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y142_SLICE_X15Y142_DO5),
.O6(CLBLM_R_X11Y142_SLICE_X15Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h2a0a2a0a3f0f3f0f)
  ) CLBLM_R_X11Y142_SLICE_X15Y142_CLUT (
.I0(CLBLM_R_X11Y137_SLICE_X15Y137_AQ),
.I1(CLBLM_L_X10Y143_SLICE_X13Y143_CO6),
.I2(CLBLM_R_X11Y144_SLICE_X14Y144_DO6),
.I3(CLBLM_L_X10Y144_SLICE_X12Y144_AO6),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y142_SLICE_X15Y142_CO5),
.O6(CLBLM_R_X11Y142_SLICE_X15Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff005050ff00d8d8)
  ) CLBLM_R_X11Y142_SLICE_X15Y142_BLUT (
.I0(CLBLM_L_X8Y144_SLICE_X11Y144_CO6),
.I1(CLBLM_R_X11Y142_SLICE_X15Y142_BQ),
.I2(CLBLM_L_X10Y142_SLICE_X12Y142_BQ),
.I3(CLBLM_L_X8Y138_SLICE_X10Y138_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X10Y145_SLICE_X13Y145_BO6),
.O5(CLBLM_R_X11Y142_SLICE_X15Y142_BO5),
.O6(CLBLM_R_X11Y142_SLICE_X15Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd11cc00fd31ec20)
  ) CLBLM_R_X11Y142_SLICE_X15Y142_ALUT (
.I0(CLBLM_L_X8Y144_SLICE_X11Y144_CO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X11Y142_SLICE_X15Y142_AQ),
.I3(CLBLM_L_X10Y135_SLICE_X13Y135_BQ),
.I4(CLBLM_R_X11Y143_SLICE_X15Y143_AQ),
.I5(CLBLM_L_X10Y145_SLICE_X13Y145_BO6),
.O5(CLBLM_R_X11Y142_SLICE_X15Y142_AO5),
.O6(CLBLM_R_X11Y142_SLICE_X15Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y143_SLICE_X14Y143_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y143_SLICE_X14Y143_AO6),
.Q(CLBLM_R_X11Y143_SLICE_X14Y143_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ac0c00000c0c)
  ) CLBLM_R_X11Y143_SLICE_X14Y143_DLUT (
.I0(CLBLM_R_X11Y143_SLICE_X15Y143_BQ),
.I1(CLBLM_R_X11Y143_SLICE_X15Y143_CO6),
.I2(CLBLM_R_X11Y142_SLICE_X14Y142_AQ),
.I3(CLBLM_R_X11Y143_SLICE_X14Y143_CO6),
.I4(CLBLM_L_X10Y145_SLICE_X12Y145_CO6),
.I5(CLBLM_R_X11Y142_SLICE_X15Y142_DQ),
.O5(CLBLM_R_X11Y143_SLICE_X14Y143_DO5),
.O6(CLBLM_R_X11Y143_SLICE_X14Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0000000f000f000)
  ) CLBLM_R_X11Y143_SLICE_X14Y143_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y142_SLICE_X15Y142_CQ),
.I2(CLBLM_L_X10Y142_SLICE_X13Y142_CQ),
.I3(CLBLM_R_X11Y144_SLICE_X14Y144_CO6),
.I4(CLBLM_L_X10Y143_SLICE_X12Y143_CQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y143_SLICE_X14Y143_CO5),
.O6(CLBLM_R_X11Y143_SLICE_X14Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0000aaa000000f0)
  ) CLBLM_R_X11Y143_SLICE_X14Y143_BLUT (
.I0(CLBLM_R_X11Y143_SLICE_X14Y143_DO6),
.I1(1'b1),
.I2(CLBLM_L_X10Y142_SLICE_X12Y142_CQ),
.I3(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.I4(CLBLM_R_X11Y144_SLICE_X14Y144_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y143_SLICE_X14Y143_BO5),
.O6(CLBLM_R_X11Y143_SLICE_X14Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccf0f0aaff)
  ) CLBLM_R_X11Y143_SLICE_X14Y143_ALUT (
.I0(CLBLM_R_X11Y143_SLICE_X14Y143_BO5),
.I1(CLBLM_L_X12Y142_SLICE_X16Y142_BQ),
.I2(CLBLM_L_X8Y141_SLICE_X11Y141_DO5),
.I3(CLBLM_L_X10Y144_SLICE_X12Y144_BO6),
.I4(CLBLM_L_X10Y145_SLICE_X13Y145_BO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y143_SLICE_X14Y143_AO5),
.O6(CLBLM_R_X11Y143_SLICE_X14Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y143_SLICE_X15Y143_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y143_SLICE_X15Y143_AO6),
.Q(CLBLM_R_X11Y143_SLICE_X15Y143_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y143_SLICE_X15Y143_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y143_SLICE_X15Y143_BO6),
.Q(CLBLM_R_X11Y143_SLICE_X15Y143_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0fef00f0f010f)
  ) CLBLM_R_X11Y143_SLICE_X15Y143_DLUT (
.I0(CLBLM_R_X11Y143_SLICE_X15Y143_CO5),
.I1(CLBLM_R_X11Y143_SLICE_X14Y143_CO6),
.I2(CLBLM_L_X10Y144_SLICE_X13Y144_DO6),
.I3(CLBLM_R_X11Y142_SLICE_X15Y142_BQ),
.I4(CLBLM_L_X10Y145_SLICE_X12Y145_CO6),
.I5(CLBLM_R_X11Y143_SLICE_X15Y143_BQ),
.O5(CLBLM_R_X11Y143_SLICE_X15Y143_DO5),
.O6(CLBLM_R_X11Y143_SLICE_X15Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000010000000f00)
  ) CLBLM_R_X11Y143_SLICE_X15Y143_CLUT (
.I0(CLBLM_R_X11Y143_SLICE_X15Y143_BQ),
.I1(CLBLM_R_X11Y142_SLICE_X15Y142_DQ),
.I2(CLBLM_L_X10Y143_SLICE_X12Y143_CQ),
.I3(CLBLM_L_X10Y143_SLICE_X13Y143_DO6),
.I4(CLBLM_R_X11Y142_SLICE_X15Y142_CQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y143_SLICE_X15Y143_CO5),
.O6(CLBLM_R_X11Y143_SLICE_X15Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5f0f13035f0f1303)
  ) CLBLM_R_X11Y143_SLICE_X15Y143_BLUT (
.I0(CLBLM_R_X11Y143_SLICE_X15Y143_DO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X11Y144_SLICE_X14Y144_DO6),
.I3(CLBLM_L_X10Y144_SLICE_X12Y144_AO6),
.I4(CLBLM_L_X12Y143_SLICE_X17Y143_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y143_SLICE_X15Y143_BO5),
.O6(CLBLM_R_X11Y143_SLICE_X15Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00fc30ee22ee22)
  ) CLBLM_R_X11Y143_SLICE_X15Y143_ALUT (
.I0(CLBLM_R_X11Y142_SLICE_X15Y142_BQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X11Y143_SLICE_X15Y143_AQ),
.I3(CLBLM_L_X8Y143_SLICE_X10Y143_CQ),
.I4(CLBLM_L_X10Y145_SLICE_X13Y145_BO6),
.I5(CLBLM_L_X8Y144_SLICE_X11Y144_CO6),
.O5(CLBLM_R_X11Y143_SLICE_X15Y143_AO5),
.O6(CLBLM_R_X11Y143_SLICE_X15Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y144_SLICE_X14Y144_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y144_SLICE_X14Y144_AO6),
.Q(CLBLM_R_X11Y144_SLICE_X14Y144_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5500550055555555)
  ) CLBLM_R_X11Y144_SLICE_X14Y144_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X11Y145_SLICE_X14Y145_AO5),
.I4(1'b1),
.I5(CLBLM_R_X11Y143_SLICE_X14Y143_DO6),
.O5(CLBLM_R_X11Y144_SLICE_X14Y144_DO5),
.O6(CLBLM_R_X11Y144_SLICE_X14Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h10f0000000000000)
  ) CLBLM_R_X11Y144_SLICE_X14Y144_CLUT (
.I0(CLBLM_L_X10Y142_SLICE_X12Y142_CQ),
.I1(CLBLM_R_X11Y144_SLICE_X14Y144_AQ),
.I2(CLBLM_L_X10Y143_SLICE_X12Y143_AQ),
.I3(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.I4(CLBLM_R_X11Y144_SLICE_X15Y144_BQ),
.I5(CLBLM_L_X10Y144_SLICE_X13Y144_AQ),
.O5(CLBLM_R_X11Y144_SLICE_X14Y144_CO5),
.O6(CLBLM_R_X11Y144_SLICE_X14Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0eeeef0fff0ff)
  ) CLBLM_R_X11Y144_SLICE_X14Y144_BLUT (
.I0(CLBLM_L_X10Y144_SLICE_X12Y144_AQ),
.I1(CLBLM_L_X8Y140_SLICE_X10Y140_DQ),
.I2(CLBLM_L_X10Y143_SLICE_X13Y143_AQ),
.I3(RIOB33_X105Y143_IOB_X1Y143_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y144_SLICE_X14Y144_BO5),
.O6(CLBLM_R_X11Y144_SLICE_X14Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8888d88d8888d8d8)
  ) CLBLM_R_X11Y144_SLICE_X14Y144_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X11Y141_SLICE_X14Y141_AQ),
.I2(CLBLM_R_X11Y144_SLICE_X14Y144_AQ),
.I3(CLBLM_R_X11Y145_SLICE_X14Y145_AO6),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(CLBLM_R_X11Y143_SLICE_X14Y143_DO6),
.O5(CLBLM_R_X11Y144_SLICE_X14Y144_AO5),
.O6(CLBLM_R_X11Y144_SLICE_X14Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y144_SLICE_X15Y144_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y144_SLICE_X15Y144_AO6),
.Q(CLBLM_R_X11Y144_SLICE_X15Y144_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y144_SLICE_X15Y144_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y144_SLICE_X15Y144_BO6),
.Q(CLBLM_R_X11Y144_SLICE_X15Y144_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha5a5f0a5a5a5f0a5)
  ) CLBLM_R_X11Y144_SLICE_X15Y144_DLUT (
.I0(CLBLM_L_X10Y144_SLICE_X13Y144_DO6),
.I1(1'b1),
.I2(CLBLM_R_X11Y144_SLICE_X15Y144_BQ),
.I3(CLBLM_L_X10Y145_SLICE_X13Y145_AQ),
.I4(CLBLM_L_X10Y145_SLICE_X12Y145_CO6),
.I5(1'b1),
.O5(CLBLM_R_X11Y144_SLICE_X15Y144_DO5),
.O6(CLBLM_R_X11Y144_SLICE_X15Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333033333331313)
  ) CLBLM_R_X11Y144_SLICE_X15Y144_CLUT (
.I0(CLBLM_R_X11Y143_SLICE_X15Y143_CO5),
.I1(CLBLM_L_X10Y144_SLICE_X13Y144_DO6),
.I2(CLBLM_R_X11Y143_SLICE_X15Y143_AQ),
.I3(CLBLM_R_X11Y143_SLICE_X14Y143_CO6),
.I4(CLBLM_L_X10Y145_SLICE_X12Y145_CO6),
.I5(CLBLM_R_X11Y143_SLICE_X15Y143_BQ),
.O5(CLBLM_R_X11Y144_SLICE_X15Y144_CO5),
.O6(CLBLM_R_X11Y144_SLICE_X15Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h44ff44ff040f040f)
  ) CLBLM_R_X11Y144_SLICE_X15Y144_BLUT (
.I0(CLBLM_R_X11Y144_SLICE_X15Y144_DO6),
.I1(CLBLM_L_X10Y144_SLICE_X12Y144_AO6),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X11Y144_SLICE_X14Y144_DO6),
.I4(1'b1),
.I5(CLBLM_L_X10Y141_SLICE_X13Y141_CQ),
.O5(CLBLM_R_X11Y144_SLICE_X15Y144_BO5),
.O6(CLBLM_R_X11Y144_SLICE_X15Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa50fa50fe54fe54)
  ) CLBLM_R_X11Y144_SLICE_X15Y144_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y141_IOB_X1Y142_I),
.I2(CLBLM_R_X11Y144_SLICE_X15Y144_AQ),
.I3(CLBLM_R_X11Y142_SLICE_X15Y142_DQ),
.I4(1'b1),
.I5(CLBLM_R_X7Y131_SLICE_X9Y131_AQ),
.O5(CLBLM_R_X11Y144_SLICE_X15Y144_AO5),
.O6(CLBLM_R_X11Y144_SLICE_X15Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y145_SLICE_X14Y145_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y145_SLICE_X14Y145_DO5),
.O6(CLBLM_R_X11Y145_SLICE_X14Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y145_SLICE_X14Y145_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y145_SLICE_X14Y145_CO5),
.O6(CLBLM_R_X11Y145_SLICE_X14Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y145_SLICE_X14Y145_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y145_SLICE_X14Y145_BO5),
.O6(CLBLM_R_X11Y145_SLICE_X14Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa5f22570f518fd9)
  ) CLBLM_R_X11Y145_SLICE_X14Y145_ALUT (
.I0(CLBLM_R_X11Y144_SLICE_X14Y144_AQ),
.I1(CLBLM_L_X8Y142_SLICE_X10Y142_D5Q),
.I2(CLBLM_L_X10Y142_SLICE_X12Y142_CQ),
.I3(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.I4(CLBLM_L_X10Y141_SLICE_X12Y141_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X11Y145_SLICE_X14Y145_AO5),
.O6(CLBLM_R_X11Y145_SLICE_X14Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y145_SLICE_X15Y145_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y145_SLICE_X15Y145_DO5),
.O6(CLBLM_R_X11Y145_SLICE_X15Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y145_SLICE_X15Y145_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y145_SLICE_X15Y145_CO5),
.O6(CLBLM_R_X11Y145_SLICE_X15Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y145_SLICE_X15Y145_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y145_SLICE_X15Y145_BO5),
.O6(CLBLM_R_X11Y145_SLICE_X15Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y145_SLICE_X15Y145_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y145_SLICE_X15Y145_AO5),
.O6(CLBLM_R_X11Y145_SLICE_X15Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y146_SLICE_X14Y146_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y146_SLICE_X16Y146_AO5),
.Q(CLBLM_R_X11Y146_SLICE_X14Y146_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y146_SLICE_X14Y146_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y146_SLICE_X14Y146_DO5),
.O6(CLBLM_R_X11Y146_SLICE_X14Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y146_SLICE_X14Y146_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y146_SLICE_X14Y146_CO5),
.O6(CLBLM_R_X11Y146_SLICE_X14Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y146_SLICE_X14Y146_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y146_SLICE_X14Y146_BO5),
.O6(CLBLM_R_X11Y146_SLICE_X14Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y146_SLICE_X14Y146_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y146_SLICE_X14Y146_AO5),
.O6(CLBLM_R_X11Y146_SLICE_X14Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y146_SLICE_X15Y146_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y146_SLICE_X15Y146_DO5),
.O6(CLBLM_R_X11Y146_SLICE_X15Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y146_SLICE_X15Y146_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y146_SLICE_X15Y146_CO5),
.O6(CLBLM_R_X11Y146_SLICE_X15Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y146_SLICE_X15Y146_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y146_SLICE_X15Y146_BO5),
.O6(CLBLM_R_X11Y146_SLICE_X15Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y146_SLICE_X15Y146_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y146_SLICE_X15Y146_AO5),
.O6(CLBLM_R_X11Y146_SLICE_X15Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y153_SLICE_X14Y153_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y153_SLICE_X14Y153_DO5),
.O6(CLBLM_R_X11Y153_SLICE_X14Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y153_SLICE_X14Y153_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y153_SLICE_X14Y153_CO5),
.O6(CLBLM_R_X11Y153_SLICE_X14Y153_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y153_SLICE_X14Y153_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y153_SLICE_X14Y153_BO5),
.O6(CLBLM_R_X11Y153_SLICE_X14Y153_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555555555555555)
  ) CLBLM_R_X11Y153_SLICE_X14Y153_ALUT (
.I0(CLBLM_R_X11Y139_SLICE_X14Y139_B5Q),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y153_SLICE_X14Y153_AO5),
.O6(CLBLM_R_X11Y153_SLICE_X14Y153_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y153_SLICE_X15Y153_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y153_SLICE_X15Y153_DO5),
.O6(CLBLM_R_X11Y153_SLICE_X15Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y153_SLICE_X15Y153_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y153_SLICE_X15Y153_CO5),
.O6(CLBLM_R_X11Y153_SLICE_X15Y153_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y153_SLICE_X15Y153_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y153_SLICE_X15Y153_BO5),
.O6(CLBLM_R_X11Y153_SLICE_X15Y153_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y153_SLICE_X15Y153_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y153_SLICE_X15Y153_AO5),
.O6(CLBLM_R_X11Y153_SLICE_X15Y153_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y133_SLICE_X18Y133_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y133_SLICE_X18Y133_AO6),
.Q(CLBLM_R_X13Y133_SLICE_X18Y133_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y133_SLICE_X18Y133_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y133_SLICE_X18Y133_BO6),
.Q(CLBLM_R_X13Y133_SLICE_X18Y133_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y133_SLICE_X18Y133_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y133_SLICE_X18Y133_DO5),
.O6(CLBLM_R_X13Y133_SLICE_X18Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y133_SLICE_X18Y133_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y133_SLICE_X18Y133_CO5),
.O6(CLBLM_R_X13Y133_SLICE_X18Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff005454ff000000)
  ) CLBLM_R_X13Y133_SLICE_X18Y133_BLUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_R_X13Y133_SLICE_X18Y133_BQ),
.I2(CLBLM_R_X11Y131_SLICE_X14Y131_BQ),
.I3(CLBLM_L_X12Y133_SLICE_X17Y133_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y138_SLICE_X10Y138_AQ),
.O5(CLBLM_R_X13Y133_SLICE_X18Y133_BO5),
.O6(CLBLM_R_X13Y133_SLICE_X18Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hec20ff33ec20cc00)
  ) CLBLM_R_X13Y133_SLICE_X18Y133_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X13Y133_SLICE_X18Y133_AQ),
.I3(CLBLM_L_X10Y142_SLICE_X13Y142_CQ),
.I4(CLBLM_L_X10Y135_SLICE_X12Y135_DO6),
.I5(CLBLM_R_X11Y134_SLICE_X14Y134_BQ),
.O5(CLBLM_R_X13Y133_SLICE_X18Y133_AO5),
.O6(CLBLM_R_X13Y133_SLICE_X18Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y133_SLICE_X19Y133_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y133_SLICE_X19Y133_DO5),
.O6(CLBLM_R_X13Y133_SLICE_X19Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y133_SLICE_X19Y133_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y133_SLICE_X19Y133_CO5),
.O6(CLBLM_R_X13Y133_SLICE_X19Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y133_SLICE_X19Y133_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y133_SLICE_X19Y133_BO5),
.O6(CLBLM_R_X13Y133_SLICE_X19Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y133_SLICE_X19Y133_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y133_SLICE_X19Y133_AO5),
.O6(CLBLM_R_X13Y133_SLICE_X19Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f00f0d0f0d)
  ) CLBLM_R_X13Y134_SLICE_X18Y134_DLUT (
.I0(CLBLM_L_X12Y134_SLICE_X17Y134_BO6),
.I1(CLBLM_R_X13Y135_SLICE_X18Y135_CO6),
.I2(CLBLM_R_X13Y135_SLICE_X18Y135_BQ),
.I3(CLBLM_R_X13Y134_SLICE_X18Y134_AO5),
.I4(1'b1),
.I5(CLBLM_L_X12Y133_SLICE_X17Y133_AQ),
.O5(CLBLM_R_X13Y134_SLICE_X18Y134_DO5),
.O6(CLBLM_R_X13Y134_SLICE_X18Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hddf0ddf088f088f0)
  ) CLBLM_R_X13Y134_SLICE_X18Y134_CLUT (
.I0(CLBLM_L_X12Y133_SLICE_X17Y133_AQ),
.I1(CLBLM_R_X13Y135_SLICE_X18Y135_BQ),
.I2(CLBLM_L_X12Y133_SLICE_X16Y133_DO6),
.I3(CLBLM_L_X12Y138_SLICE_X17Y138_BO5),
.I4(1'b1),
.I5(CLBLM_R_X13Y134_SLICE_X18Y134_BO6),
.O5(CLBLM_R_X13Y134_SLICE_X18Y134_CO5),
.O6(CLBLM_R_X13Y134_SLICE_X18Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555555555555545)
  ) CLBLM_R_X13Y134_SLICE_X18Y134_BLUT (
.I0(CLBLM_R_X13Y135_SLICE_X18Y135_BQ),
.I1(CLBLM_L_X12Y139_SLICE_X17Y139_CQ),
.I2(CLBLM_L_X12Y134_SLICE_X17Y134_BO6),
.I3(CLBLM_L_X12Y133_SLICE_X16Y133_BQ),
.I4(CLBLM_R_X13Y133_SLICE_X18Y133_AQ),
.I5(CLBLM_R_X13Y135_SLICE_X18Y135_CO6),
.O5(CLBLM_R_X13Y134_SLICE_X18Y134_BO5),
.O6(CLBLM_R_X13Y134_SLICE_X18Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5a0f5a0fffffcfc)
  ) CLBLM_R_X13Y134_SLICE_X18Y134_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X12Y139_SLICE_X17Y139_CQ),
.I2(CLBLM_R_X13Y133_SLICE_X18Y133_AQ),
.I3(CLBLM_L_X12Y134_SLICE_X17Y134_AO6),
.I4(CLBLM_L_X12Y133_SLICE_X16Y133_BQ),
.I5(1'b1),
.O5(CLBLM_R_X13Y134_SLICE_X18Y134_AO5),
.O6(CLBLM_R_X13Y134_SLICE_X18Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y134_SLICE_X19Y134_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y134_SLICE_X19Y134_AO6),
.Q(CLBLM_R_X13Y134_SLICE_X19Y134_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y134_SLICE_X19Y134_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y134_SLICE_X19Y134_BO6),
.Q(CLBLM_R_X13Y134_SLICE_X19Y134_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y134_SLICE_X19Y134_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y134_SLICE_X19Y134_CO6),
.Q(CLBLM_R_X13Y134_SLICE_X19Y134_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y134_SLICE_X19Y134_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y134_SLICE_X19Y134_DO6),
.Q(CLBLM_R_X13Y134_SLICE_X19Y134_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaccccccf0)
  ) CLBLM_R_X13Y134_SLICE_X19Y134_DLUT (
.I0(CLBLM_R_X13Y139_SLICE_X19Y139_AQ),
.I1(CLBLM_R_X13Y133_SLICE_X18Y133_BQ),
.I2(CLBLM_R_X13Y134_SLICE_X19Y134_DQ),
.I3(CLBLM_L_X8Y138_SLICE_X10Y138_AQ),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X13Y134_SLICE_X19Y134_DO5),
.O6(CLBLM_R_X13Y134_SLICE_X19Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa0afa0afa0afc0c)
  ) CLBLM_R_X13Y134_SLICE_X19Y134_CLUT (
.I0(CLBLM_L_X8Y134_SLICE_X10Y134_AQ),
.I1(CLBLM_R_X13Y134_SLICE_X19Y134_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X12Y140_SLICE_X16Y140_BQ),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLM_L_X8Y138_SLICE_X10Y138_AQ),
.O5(CLBLM_R_X13Y134_SLICE_X19Y134_CO5),
.O6(CLBLM_R_X13Y134_SLICE_X19Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'he4e4f5f5e4e4e4e4)
  ) CLBLM_R_X13Y134_SLICE_X19Y134_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X13Y134_SLICE_X19Y134_BQ),
.I2(CLBLM_L_X12Y136_SLICE_X16Y136_B5Q),
.I3(1'b1),
.I4(CLBLM_R_X7Y131_SLICE_X9Y131_AQ),
.I5(RIOB33_X105Y141_IOB_X1Y142_I),
.O5(CLBLM_R_X13Y134_SLICE_X19Y134_BO5),
.O6(CLBLM_R_X13Y134_SLICE_X19Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hd8888888d8dd88dd)
  ) CLBLM_R_X13Y134_SLICE_X19Y134_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X13Y134_SLICE_X19Y134_BQ),
.I2(CLBLM_R_X13Y134_SLICE_X19Y134_AQ),
.I3(CLBLM_L_X10Y135_SLICE_X12Y135_DO6),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X13Y134_SLICE_X18Y134_CO6),
.O5(CLBLM_R_X13Y134_SLICE_X19Y134_AO5),
.O6(CLBLM_R_X13Y134_SLICE_X19Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y135_SLICE_X18Y135_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y135_SLICE_X18Y135_AO6),
.Q(CLBLM_R_X13Y135_SLICE_X18Y135_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y135_SLICE_X18Y135_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y135_SLICE_X18Y135_BO6),
.Q(CLBLM_R_X13Y135_SLICE_X18Y135_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y135_SLICE_X18Y135_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y135_SLICE_X18Y135_DO5),
.O6(CLBLM_R_X13Y135_SLICE_X18Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffffaa)
  ) CLBLM_R_X13Y135_SLICE_X18Y135_CLUT (
.I0(CLBLM_R_X11Y134_SLICE_X14Y134_AQ),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X11Y134_SLICE_X14Y134_BQ),
.I4(CLBLM_L_X12Y135_SLICE_X16Y135_CQ),
.I5(CLBLM_R_X13Y136_SLICE_X18Y136_AQ),
.O5(CLBLM_R_X13Y135_SLICE_X18Y135_CO5),
.O6(CLBLM_R_X13Y135_SLICE_X18Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'heeaa4400fafa5050)
  ) CLBLM_R_X13Y135_SLICE_X18Y135_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X13Y135_SLICE_X18Y135_BQ),
.I2(CLBLM_R_X13Y135_SLICE_X18Y135_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X11Y134_SLICE_X15Y134_AQ),
.I5(CLBLM_L_X10Y135_SLICE_X12Y135_DO6),
.O5(CLBLM_R_X13Y135_SLICE_X18Y135_BO5),
.O6(CLBLM_R_X13Y135_SLICE_X18Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hd8ddd88888dd8888)
  ) CLBLM_R_X13Y135_SLICE_X18Y135_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y136_SLICE_X11Y136_BQ),
.I2(CLBLM_R_X13Y135_SLICE_X18Y135_AQ),
.I3(CLBLM_L_X10Y135_SLICE_X12Y135_DO6),
.I4(CLBLM_L_X12Y133_SLICE_X16Y133_AQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X13Y135_SLICE_X18Y135_AO5),
.O6(CLBLM_R_X13Y135_SLICE_X18Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y135_SLICE_X19Y135_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y135_SLICE_X19Y135_DO5),
.O6(CLBLM_R_X13Y135_SLICE_X19Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y135_SLICE_X19Y135_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y135_SLICE_X19Y135_CO5),
.O6(CLBLM_R_X13Y135_SLICE_X19Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y135_SLICE_X19Y135_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y135_SLICE_X19Y135_BO5),
.O6(CLBLM_R_X13Y135_SLICE_X19Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y135_SLICE_X19Y135_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y135_SLICE_X19Y135_AO5),
.O6(CLBLM_R_X13Y135_SLICE_X19Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y136_SLICE_X18Y136_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y136_SLICE_X18Y136_AO6),
.Q(CLBLM_R_X13Y136_SLICE_X18Y136_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y136_SLICE_X18Y136_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y136_SLICE_X18Y136_BO6),
.Q(CLBLM_R_X13Y136_SLICE_X18Y136_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y136_SLICE_X18Y136_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y136_SLICE_X18Y136_CO6),
.Q(CLBLM_R_X13Y136_SLICE_X18Y136_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y136_SLICE_X18Y136_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y136_SLICE_X18Y136_DO5),
.O6(CLBLM_R_X13Y136_SLICE_X18Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0cfc0cfc0c0c0c0)
  ) CLBLM_R_X13Y136_SLICE_X18Y136_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X13Y137_SLICE_X18Y137_A5Q),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(1'b1),
.I5(CLBLM_R_X11Y135_SLICE_X15Y135_BQ),
.O5(CLBLM_R_X13Y136_SLICE_X18Y136_CO5),
.O6(CLBLM_R_X13Y136_SLICE_X18Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000baee1044)
  ) CLBLM_R_X13Y136_SLICE_X18Y136_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X13Y136_SLICE_X18Y136_BQ),
.I2(CLBLM_R_X13Y137_SLICE_X19Y137_CQ),
.I3(CLBLM_R_X13Y137_SLICE_X18Y137_BO5),
.I4(CLBLM_R_X13Y133_SLICE_X18Y133_BQ),
.I5(CLBLM_R_X13Y143_SLICE_X18Y143_AO6),
.O5(CLBLM_R_X13Y136_SLICE_X18Y136_BO5),
.O6(CLBLM_R_X13Y136_SLICE_X18Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbbbeaaa51114000)
  ) CLBLM_R_X13Y136_SLICE_X18Y136_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y135_SLICE_X12Y135_DO6),
.I2(CLBLM_R_X13Y136_SLICE_X18Y136_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_L_X12Y135_SLICE_X16Y135_CQ),
.I5(CLBLM_R_X13Y140_SLICE_X19Y140_BQ),
.O5(CLBLM_R_X13Y136_SLICE_X18Y136_AO5),
.O6(CLBLM_R_X13Y136_SLICE_X18Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y136_SLICE_X19Y136_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y136_SLICE_X19Y136_DO5),
.O6(CLBLM_R_X13Y136_SLICE_X19Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y136_SLICE_X19Y136_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y136_SLICE_X19Y136_CO5),
.O6(CLBLM_R_X13Y136_SLICE_X19Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y136_SLICE_X19Y136_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y136_SLICE_X19Y136_BO5),
.O6(CLBLM_R_X13Y136_SLICE_X19Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y136_SLICE_X19Y136_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y136_SLICE_X19Y136_AO5),
.O6(CLBLM_R_X13Y136_SLICE_X19Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y137_SLICE_X18Y137_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y137_SLICE_X18Y137_BO6),
.Q(CLBLM_R_X13Y137_SLICE_X18Y137_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y137_SLICE_X18Y137_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y137_SLICE_X18Y137_AO6),
.Q(CLBLM_R_X13Y137_SLICE_X18Y137_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffcff3cff3)
  ) CLBLM_R_X13Y137_SLICE_X18Y137_DLUT (
.I0(1'b1),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X13Y137_SLICE_X18Y137_AQ),
.I3(CLBLM_L_X12Y137_SLICE_X17Y137_DO6),
.I4(1'b1),
.I5(CLBLM_R_X11Y135_SLICE_X15Y135_BQ),
.O5(CLBLM_R_X13Y137_SLICE_X18Y137_DO5),
.O6(CLBLM_R_X13Y137_SLICE_X18Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000101000000010)
  ) CLBLM_R_X13Y137_SLICE_X18Y137_CLUT (
.I0(CLBLM_R_X13Y136_SLICE_X18Y136_BQ),
.I1(CLBLM_R_X13Y137_SLICE_X19Y137_BQ),
.I2(CLBLM_R_X11Y139_SLICE_X15Y139_BQ),
.I3(CLBLM_R_X13Y137_SLICE_X19Y137_CQ),
.I4(CLBLM_L_X12Y137_SLICE_X16Y137_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X13Y137_SLICE_X18Y137_CO5),
.O6(CLBLM_R_X13Y137_SLICE_X18Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hee44ee44000f0000)
  ) CLBLM_R_X13Y137_SLICE_X18Y137_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X12Y137_SLICE_X17Y137_A5Q),
.I2(CLBLM_L_X12Y137_SLICE_X16Y137_A5Q),
.I3(CLBLM_R_X13Y137_SLICE_X19Y137_BQ),
.I4(CLBLM_R_X11Y139_SLICE_X15Y139_BQ),
.I5(1'b1),
.O5(CLBLM_R_X13Y137_SLICE_X18Y137_BO5),
.O6(CLBLM_R_X13Y137_SLICE_X18Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haabe0014abea0140)
  ) CLBLM_R_X13Y137_SLICE_X18Y137_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X11Y135_SLICE_X15Y135_BQ),
.I2(CLBLM_R_X13Y137_SLICE_X18Y137_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X11Y138_SLICE_X15Y138_B5Q),
.I5(CLBLM_L_X12Y137_SLICE_X17Y137_DO6),
.O5(CLBLM_R_X13Y137_SLICE_X18Y137_AO5),
.O6(CLBLM_R_X13Y137_SLICE_X18Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y137_SLICE_X19Y137_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y137_SLICE_X19Y137_AO6),
.Q(CLBLM_R_X13Y137_SLICE_X19Y137_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y137_SLICE_X19Y137_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y137_SLICE_X19Y137_BO6),
.Q(CLBLM_R_X13Y137_SLICE_X19Y137_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y137_SLICE_X19Y137_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y137_SLICE_X19Y137_CO6),
.Q(CLBLM_R_X13Y137_SLICE_X19Y137_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y137_SLICE_X19Y137_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y137_SLICE_X19Y137_DO5),
.O6(CLBLM_R_X13Y137_SLICE_X19Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00f3f3ff00fcfc)
  ) CLBLM_R_X13Y137_SLICE_X19Y137_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X13Y137_SLICE_X18Y137_CO6),
.I2(CLBLM_R_X13Y143_SLICE_X18Y143_AO6),
.I3(CLBLM_R_X5Y136_SLICE_X7Y136_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X13Y137_SLICE_X19Y137_CQ),
.O5(CLBLM_R_X13Y137_SLICE_X19Y137_CO5),
.O6(CLBLM_R_X13Y137_SLICE_X19Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8888888d888d8888)
  ) CLBLM_R_X13Y137_SLICE_X19Y137_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X12Y134_SLICE_X16Y134_AQ),
.I2(CLBLM_R_X13Y137_SLICE_X18Y137_CO5),
.I3(CLBLM_R_X13Y143_SLICE_X18Y143_AO6),
.I4(CLBLM_L_X12Y137_SLICE_X16Y137_BO5),
.I5(CLBLM_R_X13Y137_SLICE_X19Y137_BQ),
.O5(CLBLM_R_X13Y137_SLICE_X19Y137_BO5),
.O6(CLBLM_R_X13Y137_SLICE_X19Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffd8d8ffffd888)
  ) CLBLM_R_X13Y137_SLICE_X19Y137_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X15Y142_SLICE_X20Y142_AQ),
.I2(CLBLM_R_X13Y137_SLICE_X19Y137_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_L_X10Y136_SLICE_X13Y136_BO6),
.I5(CLBLM_L_X8Y138_SLICE_X10Y138_AQ),
.O5(CLBLM_R_X13Y137_SLICE_X19Y137_AO5),
.O6(CLBLM_R_X13Y137_SLICE_X19Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y138_SLICE_X18Y138_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y138_SLICE_X18Y138_AO6),
.Q(CLBLM_R_X13Y138_SLICE_X18Y138_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y138_SLICE_X18Y138_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y138_SLICE_X18Y138_DO5),
.O6(CLBLM_R_X13Y138_SLICE_X18Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y138_SLICE_X18Y138_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y138_SLICE_X18Y138_CO5),
.O6(CLBLM_R_X13Y138_SLICE_X18Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000010101010)
  ) CLBLM_R_X13Y138_SLICE_X18Y138_BLUT (
.I0(RIOB33_X105Y135_IOB_X1Y135_I),
.I1(CLBLM_R_X13Y139_SLICE_X18Y139_BO6),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(1'b1),
.I4(1'b1),
.I5(RIOB33_X105Y135_IOB_X1Y136_I),
.O5(CLBLM_R_X13Y138_SLICE_X18Y138_BO5),
.O6(CLBLM_R_X13Y138_SLICE_X18Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heceea0aaeccea00a)
  ) CLBLM_R_X13Y138_SLICE_X18Y138_ALUT (
.I0(CLBLM_L_X12Y139_SLICE_X17Y139_BO5),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X13Y138_SLICE_X18Y138_AQ),
.I3(CLBLM_L_X10Y135_SLICE_X12Y135_DO6),
.I4(CLBLM_R_X13Y140_SLICE_X18Y140_CQ),
.I5(CLBLM_L_X12Y138_SLICE_X17Y138_BO5),
.O5(CLBLM_R_X13Y138_SLICE_X18Y138_AO5),
.O6(CLBLM_R_X13Y138_SLICE_X18Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y138_SLICE_X19Y138_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y138_SLICE_X19Y138_DO5),
.O6(CLBLM_R_X13Y138_SLICE_X19Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y138_SLICE_X19Y138_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y138_SLICE_X19Y138_CO5),
.O6(CLBLM_R_X13Y138_SLICE_X19Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y138_SLICE_X19Y138_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y138_SLICE_X19Y138_BO5),
.O6(CLBLM_R_X13Y138_SLICE_X19Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y138_SLICE_X19Y138_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y138_SLICE_X19Y138_AO5),
.O6(CLBLM_R_X13Y138_SLICE_X19Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y139_SLICE_X18Y139_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y139_SLICE_X18Y139_AO6),
.Q(CLBLM_R_X13Y139_SLICE_X18Y139_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y139_SLICE_X18Y139_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y139_SLICE_X18Y139_DO5),
.O6(CLBLM_R_X13Y139_SLICE_X18Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y139_SLICE_X18Y139_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y139_SLICE_X18Y139_CO5),
.O6(CLBLM_R_X13Y139_SLICE_X18Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_R_X13Y139_SLICE_X18Y139_BLUT (
.I0(RIOB33_X105Y127_IOB_X1Y128_I),
.I1(RIOB33_X105Y131_IOB_X1Y132_I),
.I2(RIOB33_X105Y129_IOB_X1Y130_I),
.I3(RIOB33_X105Y137_IOB_X1Y137_I),
.I4(RIOB33_X105Y133_IOB_X1Y134_I),
.I5(RIOB33_X105Y133_IOB_X1Y133_I),
.O5(CLBLM_R_X13Y139_SLICE_X18Y139_BO5),
.O6(CLBLM_R_X13Y139_SLICE_X18Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000babebabe)
  ) CLBLM_R_X13Y139_SLICE_X18Y139_ALUT (
.I0(CLBLM_R_X13Y143_SLICE_X18Y143_AO6),
.I1(CLBLM_R_X13Y137_SLICE_X18Y137_CO5),
.I2(CLBLM_R_X13Y139_SLICE_X18Y139_AQ),
.I3(CLBLM_R_X13Y141_SLICE_X18Y141_BO6),
.I4(CLBLM_R_X7Y132_SLICE_X9Y132_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X13Y139_SLICE_X18Y139_AO5),
.O6(CLBLM_R_X13Y139_SLICE_X18Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y139_SLICE_X19Y139_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y139_SLICE_X19Y139_AO6),
.Q(CLBLM_R_X13Y139_SLICE_X19Y139_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y139_SLICE_X19Y139_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y139_SLICE_X19Y139_DO5),
.O6(CLBLM_R_X13Y139_SLICE_X19Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y139_SLICE_X19Y139_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y139_SLICE_X19Y139_CO5),
.O6(CLBLM_R_X13Y139_SLICE_X19Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y139_SLICE_X19Y139_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y139_SLICE_X19Y139_BO5),
.O6(CLBLM_R_X13Y139_SLICE_X19Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccf0f0fafa)
  ) CLBLM_R_X13Y139_SLICE_X19Y139_ALUT (
.I0(RIOB33_X105Y141_IOB_X1Y142_I),
.I1(CLBLM_L_X8Y139_SLICE_X11Y139_AQ),
.I2(CLBLM_R_X13Y139_SLICE_X19Y139_AQ),
.I3(1'b1),
.I4(CLBLM_R_X7Y131_SLICE_X9Y131_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X13Y139_SLICE_X19Y139_AO5),
.O6(CLBLM_R_X13Y139_SLICE_X19Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y140_SLICE_X18Y140_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y140_SLICE_X18Y140_AO6),
.Q(CLBLM_R_X13Y140_SLICE_X18Y140_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y140_SLICE_X18Y140_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y140_SLICE_X18Y140_BO6),
.Q(CLBLM_R_X13Y140_SLICE_X18Y140_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y140_SLICE_X18Y140_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y140_SLICE_X18Y140_CO6),
.Q(CLBLM_R_X13Y140_SLICE_X18Y140_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccfccc33330333)
  ) CLBLM_R_X13Y140_SLICE_X18Y140_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X13Y144_SLICE_X18Y144_CO6),
.I2(CLBLM_R_X11Y142_SLICE_X14Y142_BQ),
.I3(CLBLM_R_X13Y143_SLICE_X18Y143_BO6),
.I4(CLBLM_R_X13Y141_SLICE_X18Y141_BO5),
.I5(CLBLM_R_X13Y140_SLICE_X19Y140_BQ),
.O5(CLBLM_R_X13Y140_SLICE_X18Y140_DO5),
.O6(CLBLM_R_X13Y140_SLICE_X18Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hafacafaca3a0a3a0)
  ) CLBLM_R_X13Y140_SLICE_X18Y140_CLUT (
.I0(CLBLM_R_X13Y141_SLICE_X19Y141_AQ),
.I1(CLBLM_R_X13Y143_SLICE_X18Y143_AO6),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X12Y141_SLICE_X17Y141_CO6),
.I4(1'b1),
.I5(CLBLM_R_X5Y137_SLICE_X7Y137_DO6),
.O5(CLBLM_R_X13Y140_SLICE_X18Y140_CO5),
.O6(CLBLM_R_X13Y140_SLICE_X18Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f022aaf0f02288)
  ) CLBLM_R_X13Y140_SLICE_X18Y140_BLUT (
.I0(RIOB33_X105Y121_IOB_X1Y121_I),
.I1(CLBLM_R_X13Y140_SLICE_X18Y140_BQ),
.I2(CLBLM_R_X13Y138_SLICE_X18Y138_AQ),
.I3(CLBLM_R_X13Y141_SLICE_X18Y141_DO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X13Y143_SLICE_X18Y143_AO6),
.O5(CLBLM_R_X13Y140_SLICE_X18Y140_BO5),
.O6(CLBLM_R_X13Y140_SLICE_X18Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h21ff000021ff21ff)
  ) CLBLM_R_X13Y140_SLICE_X18Y140_ALUT (
.I0(CLBLM_R_X13Y140_SLICE_X18Y140_AQ),
.I1(CLBLM_R_X13Y141_SLICE_X18Y141_AO5),
.I2(CLBLM_R_X13Y142_SLICE_X18Y142_AO6),
.I3(CLBLM_L_X12Y143_SLICE_X17Y143_DO6),
.I4(CLBLM_L_X8Y141_SLICE_X11Y141_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X13Y140_SLICE_X18Y140_AO5),
.O6(CLBLM_R_X13Y140_SLICE_X18Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y140_SLICE_X19Y140_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y140_SLICE_X19Y140_AO6),
.Q(CLBLM_R_X13Y140_SLICE_X19Y140_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y140_SLICE_X19Y140_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y140_SLICE_X19Y140_BO6),
.Q(CLBLM_R_X13Y140_SLICE_X19Y140_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y140_SLICE_X19Y140_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y140_SLICE_X19Y140_DO5),
.O6(CLBLM_R_X13Y140_SLICE_X19Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcfcfcfcfcfcfcf)
  ) CLBLM_R_X13Y140_SLICE_X19Y140_CLUT (
.I0(1'b1),
.I1(CLBLM_L_X12Y143_SLICE_X17Y143_CO5),
.I2(CLBLM_L_X12Y142_SLICE_X16Y142_CQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y140_SLICE_X19Y140_CO5),
.O6(CLBLM_R_X13Y140_SLICE_X19Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333111133ff1155)
  ) CLBLM_R_X13Y140_SLICE_X19Y140_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X12Y143_SLICE_X17Y143_DO6),
.I2(1'b1),
.I3(CLBLM_R_X13Y141_SLICE_X18Y141_AO5),
.I4(CLBLM_R_X7Y133_SLICE_X9Y133_BQ),
.I5(CLBLM_R_X13Y140_SLICE_X18Y140_DO6),
.O5(CLBLM_R_X13Y140_SLICE_X19Y140_BO5),
.O6(CLBLM_R_X13Y140_SLICE_X19Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff540054ff050005)
  ) CLBLM_R_X13Y140_SLICE_X19Y140_ALUT (
.I0(RIOB33_X105Y121_IOB_X1Y121_I),
.I1(CLBLM_R_X13Y143_SLICE_X18Y143_AO5),
.I2(CLBLM_R_X13Y140_SLICE_X19Y140_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.I5(CLBLM_R_X13Y140_SLICE_X19Y140_CO6),
.O5(CLBLM_R_X13Y140_SLICE_X19Y140_AO5),
.O6(CLBLM_R_X13Y140_SLICE_X19Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hdc0050007300dc00)
  ) CLBLM_R_X13Y141_SLICE_X18Y141_DLUT (
.I0(CLBLM_L_X12Y143_SLICE_X17Y143_AQ),
.I1(CLBLM_R_X13Y140_SLICE_X18Y140_BQ),
.I2(CLBLM_L_X12Y142_SLICE_X17Y142_CO5),
.I3(CLBLM_R_X13Y141_SLICE_X19Y141_CO5),
.I4(CLBLM_L_X12Y142_SLICE_X16Y142_BQ),
.I5(CLBLM_R_X13Y144_SLICE_X18Y144_AQ),
.O5(CLBLM_R_X13Y141_SLICE_X18Y141_DO5),
.O6(CLBLM_R_X13Y141_SLICE_X18Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8a8a9bdff0c0f0c0)
  ) CLBLM_R_X13Y141_SLICE_X18Y141_CLUT (
.I0(CLBLM_R_X13Y139_SLICE_X18Y139_AQ),
.I1(CLBLM_R_X13Y144_SLICE_X18Y144_AQ),
.I2(CLBLM_L_X12Y142_SLICE_X16Y142_BQ),
.I3(CLBLM_R_X13Y140_SLICE_X18Y140_BQ),
.I4(CLBLM_L_X12Y143_SLICE_X17Y143_BQ),
.I5(1'b1),
.O5(CLBLM_R_X13Y141_SLICE_X18Y141_CO5),
.O6(CLBLM_R_X13Y141_SLICE_X18Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h003300330515ffff)
  ) CLBLM_R_X13Y141_SLICE_X18Y141_BLUT (
.I0(CLBLM_L_X12Y142_SLICE_X17Y142_CO5),
.I1(CLBLM_L_X12Y142_SLICE_X16Y142_BQ),
.I2(CLBLM_R_X13Y139_SLICE_X18Y139_AQ),
.I3(CLBLM_R_X13Y140_SLICE_X18Y140_BQ),
.I4(CLBLM_R_X13Y137_SLICE_X18Y137_CO5),
.I5(1'b1),
.O5(CLBLM_R_X13Y141_SLICE_X18Y141_BO5),
.O6(CLBLM_R_X13Y141_SLICE_X18Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00aa00bb0f0f0f0e)
  ) CLBLM_R_X13Y141_SLICE_X18Y141_ALUT (
.I0(CLBLM_L_X12Y143_SLICE_X17Y143_BQ),
.I1(CLBLM_L_X12Y142_SLICE_X16Y142_BQ),
.I2(CLBLM_R_X13Y141_SLICE_X19Y141_CO5),
.I3(CLBLM_R_X13Y144_SLICE_X18Y144_AQ),
.I4(CLBLM_R_X13Y140_SLICE_X18Y140_BQ),
.I5(1'b1),
.O5(CLBLM_R_X13Y141_SLICE_X18Y141_AO5),
.O6(CLBLM_R_X13Y141_SLICE_X18Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y141_SLICE_X19Y141_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y141_SLICE_X19Y141_AO6),
.Q(CLBLM_R_X13Y141_SLICE_X19Y141_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y141_SLICE_X19Y141_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y141_SLICE_X19Y141_BO6),
.Q(CLBLM_R_X13Y141_SLICE_X19Y141_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcecececc31313133)
  ) CLBLM_R_X13Y141_SLICE_X19Y141_DLUT (
.I0(CLBLM_L_X12Y142_SLICE_X16Y142_CQ),
.I1(CLBLM_R_X13Y144_SLICE_X18Y144_CO6),
.I2(CLBLM_R_X13Y141_SLICE_X18Y141_BO5),
.I3(CLBLM_R_X13Y142_SLICE_X19Y142_CO6),
.I4(CLBLM_R_X13Y142_SLICE_X19Y142_DO6),
.I5(CLBLM_R_X13Y141_SLICE_X19Y141_AQ),
.O5(CLBLM_R_X13Y141_SLICE_X19Y141_DO5),
.O6(CLBLM_R_X13Y141_SLICE_X19Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0c03000f0c0300)
  ) CLBLM_R_X13Y141_SLICE_X19Y141_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X13Y141_SLICE_X19Y141_AQ),
.I2(CLBLM_R_X13Y141_SLICE_X18Y141_BO5),
.I3(CLBLM_R_X13Y142_SLICE_X19Y142_CO6),
.I4(CLBLM_R_X13Y142_SLICE_X19Y142_DO6),
.I5(1'b1),
.O5(CLBLM_R_X13Y141_SLICE_X19Y141_CO5),
.O6(CLBLM_R_X13Y141_SLICE_X19Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff000c0c0c0c)
  ) CLBLM_R_X13Y141_SLICE_X19Y141_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X13Y141_SLICE_X19Y141_BQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_L_X12Y142_SLICE_X17Y142_BQ),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X13Y141_SLICE_X19Y141_BO5),
.O6(CLBLM_R_X13Y141_SLICE_X19Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0404cccc0505ffff)
  ) CLBLM_R_X13Y141_SLICE_X19Y141_ALUT (
.I0(CLBLM_R_X13Y141_SLICE_X19Y141_DO6),
.I1(CLBLM_R_X13Y144_SLICE_X18Y144_AQ),
.I2(CLBLM_R_X13Y141_SLICE_X18Y141_AO5),
.I3(1'b1),
.I4(CLBLM_L_X12Y143_SLICE_X17Y143_DO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X13Y141_SLICE_X19Y141_AO5),
.O6(CLBLM_R_X13Y141_SLICE_X19Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffd)
  ) CLBLM_R_X13Y142_SLICE_X18Y142_DLUT (
.I0(CLBLM_R_X13Y141_SLICE_X18Y141_CO5),
.I1(CLBLM_R_X13Y140_SLICE_X18Y140_AQ),
.I2(CLBLM_L_X12Y141_SLICE_X16Y141_AQ),
.I3(CLBLM_L_X12Y140_SLICE_X17Y140_AQ),
.I4(CLBLM_L_X12Y142_SLICE_X17Y142_AQ),
.I5(CLBLM_L_X12Y142_SLICE_X16Y142_AQ),
.O5(CLBLM_R_X13Y142_SLICE_X18Y142_DO5),
.O6(CLBLM_R_X13Y142_SLICE_X18Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hbfffffffffffffff)
  ) CLBLM_R_X13Y142_SLICE_X18Y142_CLUT (
.I0(CLBLM_R_X13Y141_SLICE_X18Y141_CO5),
.I1(CLBLM_R_X13Y140_SLICE_X18Y140_AQ),
.I2(CLBLM_L_X12Y141_SLICE_X16Y141_AQ),
.I3(CLBLM_L_X12Y140_SLICE_X17Y140_AQ),
.I4(CLBLM_L_X12Y142_SLICE_X17Y142_AQ),
.I5(CLBLM_L_X12Y142_SLICE_X16Y142_AQ),
.O5(CLBLM_R_X13Y142_SLICE_X18Y142_CO5),
.O6(CLBLM_R_X13Y142_SLICE_X18Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0e0f0f0f020f0f)
  ) CLBLM_R_X13Y142_SLICE_X18Y142_BLUT (
.I0(CLBLM_R_X13Y142_SLICE_X18Y142_DO6),
.I1(CLBLM_R_X13Y140_SLICE_X19Y140_BQ),
.I2(CLBLM_R_X13Y144_SLICE_X18Y144_CO6),
.I3(CLBLM_R_X13Y141_SLICE_X18Y141_BO5),
.I4(CLBLM_L_X12Y143_SLICE_X16Y143_CQ),
.I5(CLBLM_R_X13Y142_SLICE_X18Y142_CO6),
.O5(CLBLM_R_X13Y142_SLICE_X18Y142_BO5),
.O6(CLBLM_R_X13Y142_SLICE_X18Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00ff003700f7)
  ) CLBLM_R_X13Y142_SLICE_X18Y142_ALUT (
.I0(CLBLM_R_X13Y143_SLICE_X18Y143_DO6),
.I1(CLBLM_R_X11Y141_SLICE_X15Y141_CQ),
.I2(CLBLM_L_X12Y141_SLICE_X16Y141_AQ),
.I3(CLBLM_R_X13Y144_SLICE_X18Y144_CO6),
.I4(CLBLM_R_X13Y143_SLICE_X18Y143_CO6),
.I5(CLBLM_R_X13Y141_SLICE_X18Y141_BO5),
.O5(CLBLM_R_X13Y142_SLICE_X18Y142_AO5),
.O6(CLBLM_R_X13Y142_SLICE_X18Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y142_SLICE_X19Y142_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y142_SLICE_X19Y142_AO6),
.Q(CLBLM_R_X13Y142_SLICE_X19Y142_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_R_X13Y142_SLICE_X19Y142_DLUT (
.I0(CLBLM_R_X13Y143_SLICE_X18Y143_CO6),
.I1(CLBLM_L_X12Y142_SLICE_X17Y142_BQ),
.I2(CLBLM_R_X13Y140_SLICE_X19Y140_BQ),
.I3(CLBLM_R_X13Y140_SLICE_X18Y140_AQ),
.I4(CLBLM_L_X12Y141_SLICE_X16Y141_AQ),
.I5(CLBLM_R_X13Y142_SLICE_X19Y142_AQ),
.O5(CLBLM_R_X13Y142_SLICE_X19Y142_DO5),
.O6(CLBLM_R_X13Y142_SLICE_X19Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000010)
  ) CLBLM_R_X13Y142_SLICE_X19Y142_CLUT (
.I0(CLBLM_R_X13Y140_SLICE_X19Y140_BQ),
.I1(CLBLM_L_X12Y141_SLICE_X16Y141_AQ),
.I2(CLBLM_R_X13Y143_SLICE_X18Y143_DO6),
.I3(CLBLM_L_X12Y142_SLICE_X17Y142_BQ),
.I4(CLBLM_R_X13Y140_SLICE_X18Y140_AQ),
.I5(CLBLM_R_X13Y142_SLICE_X19Y142_AQ),
.O5(CLBLM_R_X13Y142_SLICE_X19Y142_CO5),
.O6(CLBLM_R_X13Y142_SLICE_X19Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0040bfff0050af)
  ) CLBLM_R_X13Y142_SLICE_X19Y142_BLUT (
.I0(CLBLM_R_X13Y141_SLICE_X18Y141_BO5),
.I1(CLBLM_R_X13Y143_SLICE_X19Y143_BO6),
.I2(CLBLM_L_X12Y140_SLICE_X16Y140_BQ),
.I3(CLBLM_R_X13Y142_SLICE_X19Y142_AQ),
.I4(CLBLM_R_X13Y144_SLICE_X18Y144_CO6),
.I5(CLBLM_R_X13Y143_SLICE_X19Y143_AO6),
.O5(CLBLM_R_X13Y142_SLICE_X19Y142_BO5),
.O6(CLBLM_R_X13Y142_SLICE_X19Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5070507055775577)
  ) CLBLM_R_X13Y142_SLICE_X19Y142_ALUT (
.I0(CLBLM_L_X12Y143_SLICE_X17Y143_DO6),
.I1(CLBLM_R_X13Y141_SLICE_X18Y141_AO5),
.I2(CLBLM_L_X12Y137_SLICE_X17Y137_AQ),
.I3(CLBLM_R_X13Y142_SLICE_X19Y142_BO6),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X13Y142_SLICE_X19Y142_AO5),
.O6(CLBLM_R_X13Y142_SLICE_X19Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y143_SLICE_X18Y143_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y77_IOB_X0Y77_I),
.D(CLBLM_R_X13Y140_SLICE_X18Y140_BQ),
.Q(CLBLM_R_X13Y143_SLICE_X18Y143_AQ),
.R(CLBLM_L_X12Y144_SLICE_X16Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y143_SLICE_X18Y143_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y77_IOB_X0Y77_I),
.D(CLBLM_L_X12Y143_SLICE_X16Y143_CQ),
.Q(CLBLM_R_X13Y143_SLICE_X18Y143_BQ),
.R(CLBLM_L_X12Y144_SLICE_X16Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000500040)
  ) CLBLM_R_X13Y143_SLICE_X18Y143_DLUT (
.I0(CLBLM_L_X12Y142_SLICE_X17Y142_AQ),
.I1(CLBLM_R_X13Y140_SLICE_X18Y140_BQ),
.I2(CLBLM_L_X12Y142_SLICE_X16Y142_BQ),
.I3(CLBLM_L_X12Y140_SLICE_X17Y140_AQ),
.I4(CLBLM_R_X13Y144_SLICE_X18Y144_AQ),
.I5(CLBLM_L_X12Y142_SLICE_X16Y142_AQ),
.O5(CLBLM_R_X13Y143_SLICE_X18Y143_DO5),
.O6(CLBLM_R_X13Y143_SLICE_X18Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0a0000002a000000)
  ) CLBLM_R_X13Y143_SLICE_X18Y143_CLUT (
.I0(CLBLM_L_X12Y142_SLICE_X17Y142_AQ),
.I1(CLBLM_R_X13Y140_SLICE_X18Y140_BQ),
.I2(CLBLM_L_X12Y142_SLICE_X16Y142_BQ),
.I3(CLBLM_L_X12Y140_SLICE_X17Y140_AQ),
.I4(CLBLM_L_X12Y142_SLICE_X16Y142_AQ),
.I5(CLBLM_R_X13Y144_SLICE_X18Y144_AQ),
.O5(CLBLM_R_X13Y143_SLICE_X18Y143_CO5),
.O6(CLBLM_R_X13Y143_SLICE_X18Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000800000010000)
  ) CLBLM_R_X13Y143_SLICE_X18Y143_BLUT (
.I0(CLBLM_L_X12Y141_SLICE_X16Y141_AQ),
.I1(CLBLM_L_X12Y142_SLICE_X16Y142_AQ),
.I2(CLBLM_L_X12Y142_SLICE_X17Y142_AQ),
.I3(CLBLM_R_X13Y140_SLICE_X18Y140_AQ),
.I4(CLBLM_R_X13Y141_SLICE_X18Y141_CO5),
.I5(CLBLM_L_X12Y140_SLICE_X17Y140_AQ),
.O5(CLBLM_R_X13Y143_SLICE_X18Y143_BO5),
.O6(CLBLM_R_X13Y143_SLICE_X18Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000300000200)
  ) CLBLM_R_X13Y143_SLICE_X18Y143_ALUT (
.I0(CLBLM_R_X13Y137_SLICE_X18Y137_CO5),
.I1(CLBLM_R_X13Y140_SLICE_X18Y140_BQ),
.I2(CLBLM_L_X12Y142_SLICE_X16Y142_BQ),
.I3(CLBLM_R_X13Y144_SLICE_X18Y144_AQ),
.I4(CLBLM_L_X12Y143_SLICE_X17Y143_BQ),
.I5(1'b1),
.O5(CLBLM_R_X13Y143_SLICE_X18Y143_AO5),
.O6(CLBLM_R_X13Y143_SLICE_X18Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y143_SLICE_X19Y143_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y143_SLICE_X19Y143_DO5),
.O6(CLBLM_R_X13Y143_SLICE_X19Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y143_SLICE_X19Y143_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y143_SLICE_X19Y143_CO5),
.O6(CLBLM_R_X13Y143_SLICE_X19Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000010000000100)
  ) CLBLM_R_X13Y143_SLICE_X19Y143_BLUT (
.I0(CLBLM_L_X12Y141_SLICE_X16Y141_AQ),
.I1(CLBLM_R_X13Y140_SLICE_X18Y140_AQ),
.I2(CLBLM_R_X13Y140_SLICE_X19Y140_BQ),
.I3(CLBLM_R_X13Y143_SLICE_X18Y143_DO6),
.I4(CLBLM_L_X12Y142_SLICE_X17Y142_BQ),
.I5(1'b1),
.O5(CLBLM_R_X13Y143_SLICE_X19Y143_BO5),
.O6(CLBLM_R_X13Y143_SLICE_X19Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fffffff7fffffff)
  ) CLBLM_R_X13Y143_SLICE_X19Y143_ALUT (
.I0(CLBLM_L_X12Y141_SLICE_X16Y141_AQ),
.I1(CLBLM_R_X13Y140_SLICE_X18Y140_AQ),
.I2(CLBLM_R_X13Y140_SLICE_X19Y140_BQ),
.I3(CLBLM_R_X13Y143_SLICE_X18Y143_CO6),
.I4(CLBLM_L_X12Y142_SLICE_X17Y142_BQ),
.I5(1'b1),
.O5(CLBLM_R_X13Y143_SLICE_X19Y143_AO5),
.O6(CLBLM_R_X13Y143_SLICE_X19Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y144_SLICE_X18Y144_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y144_SLICE_X18Y144_AO6),
.Q(CLBLM_R_X13Y144_SLICE_X18Y144_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y144_SLICE_X18Y144_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y144_SLICE_X18Y144_DO5),
.O6(CLBLM_R_X13Y144_SLICE_X18Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00efffffffff)
  ) CLBLM_R_X13Y144_SLICE_X18Y144_CLUT (
.I0(CLBLM_L_X12Y142_SLICE_X16Y142_BQ),
.I1(CLBLM_L_X12Y143_SLICE_X17Y143_BQ),
.I2(CLBLM_R_X13Y144_SLICE_X18Y144_AQ),
.I3(CLBLM_R_X13Y140_SLICE_X19Y140_AQ),
.I4(CLBLM_R_X13Y140_SLICE_X18Y140_BQ),
.I5(CLBLM_R_X13Y137_SLICE_X18Y137_CO5),
.O5(CLBLM_R_X13Y144_SLICE_X18Y144_CO5),
.O6(CLBLM_R_X13Y144_SLICE_X18Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00c001c1f0305f1f)
  ) CLBLM_R_X13Y144_SLICE_X18Y144_BLUT (
.I0(CLBLM_R_X13Y140_SLICE_X18Y140_BQ),
.I1(CLBLM_L_X12Y143_SLICE_X17Y143_BQ),
.I2(CLBLM_R_X13Y144_SLICE_X18Y144_AQ),
.I3(CLBLM_R_X13Y140_SLICE_X19Y140_AQ),
.I4(CLBLM_L_X12Y142_SLICE_X16Y142_BQ),
.I5(1'b1),
.O5(CLBLM_R_X13Y144_SLICE_X18Y144_BO5),
.O6(CLBLM_R_X13Y144_SLICE_X18Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000041504150)
  ) CLBLM_R_X13Y144_SLICE_X18Y144_ALUT (
.I0(RIOB33_X105Y121_IOB_X1Y121_I),
.I1(CLBLM_R_X13Y144_SLICE_X18Y144_BO5),
.I2(CLBLM_R_X13Y144_SLICE_X18Y144_AQ),
.I3(CLBLM_R_X13Y141_SLICE_X19Y141_CO5),
.I4(CLBLM_L_X12Y143_SLICE_X16Y143_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X13Y144_SLICE_X18Y144_AO5),
.O6(CLBLM_R_X13Y144_SLICE_X18Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y144_SLICE_X19Y144_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y144_SLICE_X19Y144_AO6),
.Q(CLBLM_R_X13Y144_SLICE_X19Y144_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y144_SLICE_X19Y144_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y144_SLICE_X19Y144_DO5),
.O6(CLBLM_R_X13Y144_SLICE_X19Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y144_SLICE_X19Y144_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y144_SLICE_X19Y144_CO5),
.O6(CLBLM_R_X13Y144_SLICE_X19Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y144_SLICE_X19Y144_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y144_SLICE_X19Y144_BO5),
.O6(CLBLM_R_X13Y144_SLICE_X19Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaf0aaf0aafcaafc)
  ) CLBLM_R_X13Y144_SLICE_X19Y144_ALUT (
.I0(CLBLM_L_X10Y145_SLICE_X13Y145_AQ),
.I1(RIOB33_X105Y141_IOB_X1Y142_I),
.I2(CLBLM_R_X13Y144_SLICE_X19Y144_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLM_R_X7Y131_SLICE_X9Y131_AQ),
.O5(CLBLM_R_X13Y144_SLICE_X19Y144_AO5),
.O6(CLBLM_R_X13Y144_SLICE_X19Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y142_SLICE_X20Y142_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X15Y142_SLICE_X20Y142_AO6),
.Q(CLBLM_R_X15Y142_SLICE_X20Y142_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y142_SLICE_X20Y142_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y142_SLICE_X20Y142_DO5),
.O6(CLBLM_R_X15Y142_SLICE_X20Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y142_SLICE_X20Y142_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y142_SLICE_X20Y142_CO5),
.O6(CLBLM_R_X15Y142_SLICE_X20Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y142_SLICE_X20Y142_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y142_SLICE_X20Y142_BO5),
.O6(CLBLM_R_X15Y142_SLICE_X20Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000f3f0f3f0)
  ) CLBLM_R_X15Y142_SLICE_X20Y142_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y131_SLICE_X9Y131_AQ),
.I2(CLBLM_R_X15Y142_SLICE_X20Y142_AQ),
.I3(RIOB33_X105Y141_IOB_X1Y142_I),
.I4(CLBLM_R_X13Y142_SLICE_X19Y142_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X15Y142_SLICE_X20Y142_AO5),
.O6(CLBLM_R_X15Y142_SLICE_X20Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y142_SLICE_X21Y142_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y142_SLICE_X21Y142_DO5),
.O6(CLBLM_R_X15Y142_SLICE_X21Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y142_SLICE_X21Y142_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y142_SLICE_X21Y142_CO5),
.O6(CLBLM_R_X15Y142_SLICE_X21Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y142_SLICE_X21Y142_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y142_SLICE_X21Y142_BO5),
.O6(CLBLM_R_X15Y142_SLICE_X21Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y142_SLICE_X21Y142_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y142_SLICE_X21Y142_AO5),
.O6(CLBLM_R_X15Y142_SLICE_X21Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X37Y138_SLICE_X56Y138_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X37Y138_SLICE_X56Y138_DO5),
.O6(CLBLM_R_X37Y138_SLICE_X56Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X37Y138_SLICE_X56Y138_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X37Y138_SLICE_X56Y138_CO5),
.O6(CLBLM_R_X37Y138_SLICE_X56Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X37Y138_SLICE_X56Y138_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X37Y138_SLICE_X56Y138_BO5),
.O6(CLBLM_R_X37Y138_SLICE_X56Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000022222222)
  ) CLBLM_R_X37Y138_SLICE_X56Y138_ALUT (
.I0(RIOB33_X105Y119_IOB_X1Y119_I),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X8Y138_SLICE_X10Y138_DQ),
.O5(CLBLM_R_X37Y138_SLICE_X56Y138_AO5),
.O6(CLBLM_R_X37Y138_SLICE_X56Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X37Y138_SLICE_X57Y138_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X37Y138_SLICE_X57Y138_DO5),
.O6(CLBLM_R_X37Y138_SLICE_X57Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X37Y138_SLICE_X57Y138_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X37Y138_SLICE_X57Y138_CO5),
.O6(CLBLM_R_X37Y138_SLICE_X57Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X37Y138_SLICE_X57Y138_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X37Y138_SLICE_X57Y138_BO5),
.O6(CLBLM_R_X37Y138_SLICE_X57Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X37Y138_SLICE_X57Y138_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X37Y138_SLICE_X57Y138_AO5),
.O6(CLBLM_R_X37Y138_SLICE_X57Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y140_SLICE_X162Y140_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y140_SLICE_X162Y140_DO5),
.O6(CLBLM_R_X103Y140_SLICE_X162Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y140_SLICE_X162Y140_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y140_SLICE_X162Y140_CO5),
.O6(CLBLM_R_X103Y140_SLICE_X162Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y140_SLICE_X162Y140_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y140_SLICE_X162Y140_BO5),
.O6(CLBLM_R_X103Y140_SLICE_X162Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y140_SLICE_X162Y140_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y140_SLICE_X162Y140_AO5),
.O6(CLBLM_R_X103Y140_SLICE_X162Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y140_SLICE_X163Y140_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y140_SLICE_X163Y140_DO5),
.O6(CLBLM_R_X103Y140_SLICE_X163Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y140_SLICE_X163Y140_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y140_SLICE_X163Y140_CO5),
.O6(CLBLM_R_X103Y140_SLICE_X163Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y140_SLICE_X163Y140_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y140_SLICE_X163Y140_BO5),
.O6(CLBLM_R_X103Y140_SLICE_X163Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc000c00088880000)
  ) CLBLM_R_X103Y140_SLICE_X163Y140_ALUT (
.I0(RIOB33_X105Y141_IOB_X1Y141_I),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(RIOB33_X105Y137_IOB_X1Y138_I),
.I3(RIOB33_X105Y139_IOB_X1Y139_I),
.I4(RIOB33_X105Y139_IOB_X1Y140_I),
.I5(1'b1),
.O5(CLBLM_R_X103Y140_SLICE_X163Y140_AO5),
.O6(CLBLM_R_X103Y140_SLICE_X163Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y169_SLICE_X162Y169_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y169_SLICE_X162Y169_DO5),
.O6(CLBLM_R_X103Y169_SLICE_X162Y169_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y169_SLICE_X162Y169_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y169_SLICE_X162Y169_CO5),
.O6(CLBLM_R_X103Y169_SLICE_X162Y169_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y169_SLICE_X162Y169_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y169_SLICE_X162Y169_BO5),
.O6(CLBLM_R_X103Y169_SLICE_X162Y169_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y169_SLICE_X162Y169_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y169_SLICE_X162Y169_AO5),
.O6(CLBLM_R_X103Y169_SLICE_X162Y169_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y169_SLICE_X163Y169_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y169_SLICE_X163Y169_DO5),
.O6(CLBLM_R_X103Y169_SLICE_X163Y169_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y169_SLICE_X163Y169_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y169_SLICE_X163Y169_CO5),
.O6(CLBLM_R_X103Y169_SLICE_X163Y169_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y169_SLICE_X163Y169_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y169_SLICE_X163Y169_BO5),
.O6(CLBLM_R_X103Y169_SLICE_X163Y169_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hafafafafafafafaf)
  ) CLBLM_R_X103Y169_SLICE_X163Y169_ALUT (
.I0(CLBLM_L_X12Y134_SLICE_X16Y134_AQ),
.I1(1'b1),
.I2(RIOB33_X105Y143_IOB_X1Y143_I),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y169_SLICE_X163Y169_AO5),
.O6(CLBLM_R_X103Y169_SLICE_X163Y169_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y170_SLICE_X162Y170_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y170_SLICE_X162Y170_DO5),
.O6(CLBLM_R_X103Y170_SLICE_X162Y170_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y170_SLICE_X162Y170_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y170_SLICE_X162Y170_CO5),
.O6(CLBLM_R_X103Y170_SLICE_X162Y170_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y170_SLICE_X162Y170_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y170_SLICE_X162Y170_BO5),
.O6(CLBLM_R_X103Y170_SLICE_X162Y170_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y170_SLICE_X162Y170_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y170_SLICE_X162Y170_AO5),
.O6(CLBLM_R_X103Y170_SLICE_X162Y170_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y170_SLICE_X163Y170_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y170_SLICE_X163Y170_DO5),
.O6(CLBLM_R_X103Y170_SLICE_X163Y170_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y170_SLICE_X163Y170_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y170_SLICE_X163Y170_CO5),
.O6(CLBLM_R_X103Y170_SLICE_X163Y170_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y170_SLICE_X163Y170_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y170_SLICE_X163Y170_BO5),
.O6(CLBLM_R_X103Y170_SLICE_X163Y170_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaafffff0f0ffff)
  ) CLBLM_R_X103Y170_SLICE_X163Y170_ALUT (
.I0(CLBLM_R_X11Y144_SLICE_X15Y144_AQ),
.I1(1'b1),
.I2(CLBLM_R_X15Y142_SLICE_X20Y142_AQ),
.I3(1'b1),
.I4(RIOB33_X105Y143_IOB_X1Y143_I),
.I5(1'b1),
.O5(CLBLM_R_X103Y170_SLICE_X163Y170_AO5),
.O6(CLBLM_R_X103Y170_SLICE_X163Y170_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y173_SLICE_X162Y173_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y173_SLICE_X162Y173_DO5),
.O6(CLBLM_R_X103Y173_SLICE_X162Y173_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y173_SLICE_X162Y173_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y173_SLICE_X162Y173_CO5),
.O6(CLBLM_R_X103Y173_SLICE_X162Y173_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y173_SLICE_X162Y173_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y173_SLICE_X162Y173_BO5),
.O6(CLBLM_R_X103Y173_SLICE_X162Y173_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y173_SLICE_X162Y173_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y173_SLICE_X162Y173_AO5),
.O6(CLBLM_R_X103Y173_SLICE_X162Y173_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y173_SLICE_X163Y173_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y173_SLICE_X163Y173_DO5),
.O6(CLBLM_R_X103Y173_SLICE_X163Y173_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y173_SLICE_X163Y173_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y173_SLICE_X163Y173_CO5),
.O6(CLBLM_R_X103Y173_SLICE_X163Y173_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y173_SLICE_X163Y173_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y173_SLICE_X163Y173_BO5),
.O6(CLBLM_R_X103Y173_SLICE_X163Y173_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ffffccccffff)
  ) CLBLM_R_X103Y173_SLICE_X163Y173_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X13Y144_SLICE_X19Y144_AQ),
.I2(1'b1),
.I3(CLBLM_R_X13Y134_SLICE_X19Y134_BQ),
.I4(RIOB33_X105Y143_IOB_X1Y143_I),
.I5(1'b1),
.O5(CLBLM_R_X103Y173_SLICE_X163Y173_AO5),
.O6(CLBLM_R_X103Y173_SLICE_X163Y173_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y175_SLICE_X162Y175_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y175_SLICE_X162Y175_DO5),
.O6(CLBLM_R_X103Y175_SLICE_X162Y175_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y175_SLICE_X162Y175_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y175_SLICE_X162Y175_CO5),
.O6(CLBLM_R_X103Y175_SLICE_X162Y175_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y175_SLICE_X162Y175_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y175_SLICE_X162Y175_BO5),
.O6(CLBLM_R_X103Y175_SLICE_X162Y175_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y175_SLICE_X162Y175_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y175_SLICE_X162Y175_AO5),
.O6(CLBLM_R_X103Y175_SLICE_X162Y175_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y175_SLICE_X163Y175_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y175_SLICE_X163Y175_DO5),
.O6(CLBLM_R_X103Y175_SLICE_X163Y175_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y175_SLICE_X163Y175_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y175_SLICE_X163Y175_CO5),
.O6(CLBLM_R_X103Y175_SLICE_X163Y175_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y175_SLICE_X163Y175_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y175_SLICE_X163Y175_BO5),
.O6(CLBLM_R_X103Y175_SLICE_X163Y175_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffccffcc)
  ) CLBLM_R_X103Y175_SLICE_X163Y175_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y127_IOB_X1Y128_I),
.I2(1'b1),
.I3(RIOB33_X105Y129_IOB_X1Y129_I),
.I4(1'b1),
.I5(RIOB33_X105Y129_IOB_X1Y130_I),
.O5(CLBLM_R_X103Y175_SLICE_X163Y175_AO5),
.O6(CLBLM_R_X103Y175_SLICE_X163Y175_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y177_SLICE_X162Y177_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X162Y177_DO5),
.O6(CLBLM_R_X103Y177_SLICE_X162Y177_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y177_SLICE_X162Y177_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X162Y177_CO5),
.O6(CLBLM_R_X103Y177_SLICE_X162Y177_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y177_SLICE_X162Y177_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X162Y177_BO5),
.O6(CLBLM_R_X103Y177_SLICE_X162Y177_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y177_SLICE_X162Y177_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X162Y177_AO5),
.O6(CLBLM_R_X103Y177_SLICE_X162Y177_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y177_SLICE_X163Y177_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X163Y177_DO5),
.O6(CLBLM_R_X103Y177_SLICE_X163Y177_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y177_SLICE_X163Y177_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X163Y177_CO5),
.O6(CLBLM_R_X103Y177_SLICE_X163Y177_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y177_SLICE_X163Y177_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X163Y177_BO5),
.O6(CLBLM_R_X103Y177_SLICE_X163Y177_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0fff0fcfcfcfcf)
  ) CLBLM_R_X103Y177_SLICE_X163Y177_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X13Y143_SLICE_X18Y143_BQ),
.I2(RIOB33_X105Y143_IOB_X1Y143_I),
.I3(CLBLM_R_X13Y139_SLICE_X19Y139_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X163Y177_AO5),
.O6(CLBLM_R_X103Y177_SLICE_X163Y177_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFGCTRL" *)
  BUFGCTRL #(
    .INIT_OUT(0),
    .IS_CE0_INVERTED(0),
    .IS_CE1_INVERTED(1),
    .IS_IGNORE0_INVERTED(1),
    .IS_IGNORE1_INVERTED(0),
    .IS_S0_INVERTED(0),
    .IS_S1_INVERTED(1),
    .PRESELECT_I0("TRUE"),
    .PRESELECT_I1("FALSE")
  ) CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_BUFGCTRL (
.CE0(1'b1),
.CE1(1'b1),
.I0(LIOB33_X0Y77_IOB_X0Y78_I),
.I1(1'b1),
.IGNORE0(1'b1),
.IGNORE1(1'b1),
.O(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.S0(1'b1),
.S1(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFHCE" *)
  BUFHCE #(
    .CE_TYPE("SYNC"),
    .INIT_OUT(0),
    .IS_CE_INVERTED(0)
  ) CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_BUFHCE (
.CE(1'b1),
.I(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.O(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y51_IOB_X0Y51_IBUF (
.I(LIOB33_X0Y51_IOB_X0Y51_IPAD),
.O(LIOB33_X0Y51_IOB_X0Y51_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y51_IOB_X0Y52_IBUF (
.I(LIOB33_X0Y51_IOB_X0Y52_IPAD),
.O(LIOB33_X0Y51_IOB_X0Y52_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y53_IOB_X0Y53_IBUF (
.I(LIOB33_X0Y53_IOB_X0Y53_IPAD),
.O(LIOB33_X0Y53_IOB_X0Y53_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y53_IOB_X0Y54_IBUF (
.I(LIOB33_X0Y53_IOB_X0Y54_IPAD),
.O(LIOB33_X0Y53_IOB_X0Y54_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y55_IOB_X0Y55_IBUF (
.I(LIOB33_X0Y55_IOB_X0Y55_IPAD),
.O(LIOB33_X0Y55_IOB_X0Y55_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y55_IOB_X0Y56_IBUF (
.I(LIOB33_X0Y55_IOB_X0Y56_IPAD),
.O(LIOB33_X0Y55_IOB_X0Y56_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y57_IOB_X0Y57_IBUF (
.I(LIOB33_X0Y57_IOB_X0Y57_IPAD),
.O(LIOB33_X0Y57_IOB_X0Y57_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y57_IOB_X0Y58_IBUF (
.I(LIOB33_X0Y57_IOB_X0Y58_IPAD),
.O(LIOB33_X0Y57_IOB_X0Y58_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y59_IOB_X0Y59_IBUF (
.I(LIOB33_X0Y59_IOB_X0Y59_IPAD),
.O(LIOB33_X0Y59_IOB_X0Y59_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y59_IOB_X0Y60_IBUF (
.I(LIOB33_X0Y59_IOB_X0Y60_IPAD),
.O(LIOB33_X0Y59_IOB_X0Y60_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y61_IOB_X0Y61_IBUF (
.I(LIOB33_X0Y61_IOB_X0Y61_IPAD),
.O(LIOB33_X0Y61_IOB_X0Y61_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y61_IOB_X0Y62_IBUF (
.I(LIOB33_X0Y61_IOB_X0Y62_IPAD),
.O(LIOB33_X0Y61_IOB_X0Y62_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y63_IOB_X0Y63_IBUF (
.I(LIOB33_X0Y63_IOB_X0Y63_IPAD),
.O(LIOB33_X0Y63_IOB_X0Y63_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y63_IOB_X0Y64_IBUF (
.I(LIOB33_X0Y63_IOB_X0Y64_IPAD),
.O(LIOB33_X0Y63_IOB_X0Y64_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y65_IOB_X0Y65_IBUF (
.I(LIOB33_X0Y65_IOB_X0Y65_IPAD),
.O(LIOB33_X0Y65_IOB_X0Y65_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y65_IOB_X0Y66_IBUF (
.I(LIOB33_X0Y65_IOB_X0Y66_IPAD),
.O(LIOB33_X0Y65_IOB_X0Y66_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y67_IOB_X0Y67_IBUF (
.I(LIOB33_X0Y67_IOB_X0Y67_IPAD),
.O(LIOB33_X0Y67_IOB_X0Y67_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y67_IOB_X0Y68_IBUF (
.I(LIOB33_X0Y67_IOB_X0Y68_IPAD),
.O(LIOB33_X0Y67_IOB_X0Y68_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y69_IOB_X0Y69_IBUF (
.I(LIOB33_X0Y69_IOB_X0Y69_IPAD),
.O(LIOB33_X0Y69_IOB_X0Y69_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y69_IOB_X0Y70_IBUF (
.I(LIOB33_X0Y69_IOB_X0Y70_IPAD),
.O(LIOB33_X0Y69_IOB_X0Y70_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y71_IOB_X0Y71_IBUF (
.I(LIOB33_X0Y71_IOB_X0Y71_IPAD),
.O(LIOB33_X0Y71_IOB_X0Y71_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y71_IOB_X0Y72_IBUF (
.I(LIOB33_X0Y71_IOB_X0Y72_IPAD),
.O(LIOB33_X0Y71_IOB_X0Y72_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y73_IOB_X0Y73_IBUF (
.I(LIOB33_X0Y73_IOB_X0Y73_IPAD),
.O(LIOB33_X0Y73_IOB_X0Y73_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y73_IOB_X0Y74_IBUF (
.I(LIOB33_X0Y73_IOB_X0Y74_IPAD),
.O(LIOB33_X0Y73_IOB_X0Y74_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y75_IOB_X0Y75_IBUF (
.I(LIOB33_X0Y75_IOB_X0Y75_IPAD),
.O(LIOB33_X0Y75_IOB_X0Y75_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y75_IOB_X0Y76_IBUF (
.I(LIOB33_X0Y75_IOB_X0Y76_IPAD),
.O(LIOB33_X0Y75_IOB_X0Y76_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y77_IOB_X0Y77_IBUF (
.I(LIOB33_X0Y77_IOB_X0Y77_IPAD),
.O(LIOB33_X0Y77_IOB_X0Y77_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y77_IOB_X0Y78_IBUF (
.I(LIOB33_X0Y77_IOB_X0Y78_IPAD),
.O(LIOB33_X0Y77_IOB_X0Y78_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y79_IOB_X0Y79_IBUF (
.I(LIOB33_X0Y79_IOB_X0Y79_IPAD),
.O(LIOB33_X0Y79_IOB_X0Y79_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y79_IOB_X0Y80_OBUF (
.I(CLBLL_L_X2Y133_SLICE_X0Y133_AO6),
.O(LIOB33_X0Y79_IOB_X0Y80_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y101_IOB_X0Y101_OBUF (
.I(CLBLM_R_X3Y133_SLICE_X2Y133_AO6),
.O(LIOB33_X0Y101_IOB_X0Y101_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y101_IOB_X0Y102_OBUF (
.I(CLBLM_R_X3Y133_SLICE_X2Y133_AO5),
.O(LIOB33_X0Y101_IOB_X0Y102_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y103_IOB_X0Y103_OBUF (
.I(CLBLL_L_X2Y133_SLICE_X0Y133_AO5),
.O(LIOB33_X0Y103_IOB_X0Y103_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y103_IOB_X0Y104_OBUF (
.I(CLBLL_L_X2Y133_SLICE_X0Y133_CO6),
.O(LIOB33_X0Y103_IOB_X0Y104_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y105_IOB_X0Y105_OBUF (
.I(CLBLL_L_X2Y133_SLICE_X0Y133_BO5),
.O(LIOB33_X0Y105_IOB_X0Y105_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y105_IOB_X0Y106_OBUF (
.I(CLBLL_L_X4Y138_SLICE_X5Y138_DO6),
.O(LIOB33_X0Y105_IOB_X0Y106_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y107_IOB_X0Y107_OBUF (
.I(CLBLL_L_X2Y108_SLICE_X0Y108_AO6),
.O(LIOB33_X0Y107_IOB_X0Y107_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y107_IOB_X0Y108_OBUF (
.I(CLBLL_L_X2Y133_SLICE_X0Y133_CO5),
.O(LIOB33_X0Y107_IOB_X0Y108_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y109_IOB_X0Y109_OBUF (
.I(CLBLL_L_X2Y127_SLICE_X0Y127_AO6),
.O(LIOB33_X0Y109_IOB_X0Y109_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y109_IOB_X0Y110_OBUF (
.I(CLBLL_L_X2Y127_SLICE_X0Y127_AO5),
.O(LIOB33_X0Y109_IOB_X0Y110_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y111_IOB_X0Y111_OBUF (
.I(1'b0),
.O(LIOB33_X0Y111_IOB_X0Y111_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y111_IOB_X0Y112_OBUF (
.I(CLBLM_L_X12Y133_SLICE_X16Y133_C5Q),
.O(LIOB33_X0Y111_IOB_X0Y112_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y113_IOB_X0Y113_OBUF (
.I(RIOB33_X105Y121_IOB_X1Y121_I),
.O(LIOB33_X0Y113_IOB_X0Y113_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y113_IOB_X0Y114_OBUF (
.I(CLBLM_R_X7Y132_SLICE_X9Y132_DQ),
.O(LIOB33_X0Y113_IOB_X0Y114_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y115_IOB_X0Y115_OBUF (
.I(CLBLM_L_X12Y133_SLICE_X16Y133_CQ),
.O(LIOB33_X0Y115_IOB_X0Y115_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y115_IOB_X0Y116_OBUF (
.I(CLBLM_L_X8Y135_SLICE_X11Y135_BQ),
.O(LIOB33_X0Y115_IOB_X0Y116_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y117_IOB_X0Y117_OBUF (
.I(CLBLM_R_X5Y136_SLICE_X6Y136_D5Q),
.O(LIOB33_X0Y117_IOB_X0Y117_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y117_IOB_X0Y118_OBUF (
.I(CLBLL_L_X4Y135_SLICE_X5Y135_DQ),
.O(LIOB33_X0Y117_IOB_X0Y118_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y119_IOB_X0Y119_OBUF (
.I(CLBLM_L_X10Y135_SLICE_X13Y135_BQ),
.O(LIOB33_X0Y119_IOB_X0Y119_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y119_IOB_X0Y120_OBUF (
.I(CLBLM_L_X12Y136_SLICE_X16Y136_BQ),
.O(LIOB33_X0Y119_IOB_X0Y120_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y121_IOB_X0Y121_OBUF (
.I(CLBLM_L_X8Y135_SLICE_X11Y135_B5Q),
.O(LIOB33_X0Y121_IOB_X0Y121_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y121_IOB_X0Y122_OBUF (
.I(CLBLL_L_X4Y133_SLICE_X5Y133_A5Q),
.O(LIOB33_X0Y121_IOB_X0Y122_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y123_IOB_X0Y123_OBUF (
.I(CLBLM_R_X7Y132_SLICE_X9Y132_D5Q),
.O(LIOB33_X0Y123_IOB_X0Y123_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y123_IOB_X0Y124_OBUF (
.I(CLBLL_L_X4Y135_SLICE_X5Y135_D5Q),
.O(LIOB33_X0Y123_IOB_X0Y124_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y125_IOB_X0Y125_OBUF (
.I(CLBLM_R_X11Y138_SLICE_X15Y138_D5Q),
.O(LIOB33_X0Y125_IOB_X0Y125_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y125_IOB_X0Y126_OBUF (
.I(CLBLM_R_X3Y136_SLICE_X3Y136_CQ),
.O(LIOB33_X0Y125_IOB_X0Y126_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y127_IOB_X0Y127_OBUF (
.I(CLBLM_R_X5Y137_SLICE_X6Y137_BQ),
.O(LIOB33_X0Y127_IOB_X0Y127_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y127_IOB_X0Y128_OBUF (
.I(CLBLL_L_X4Y134_SLICE_X5Y134_A5Q),
.O(LIOB33_X0Y127_IOB_X0Y128_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y129_IOB_X0Y129_OBUF (
.I(CLBLM_R_X5Y136_SLICE_X6Y136_CQ),
.O(LIOB33_X0Y129_IOB_X0Y129_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y129_IOB_X0Y130_OBUF (
.I(CLBLL_L_X52Y126_SLICE_X78Y126_AO6),
.O(LIOB33_X0Y129_IOB_X0Y130_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y131_IOB_X0Y131_OBUF (
.I(CLBLM_R_X7Y131_SLICE_X9Y131_AO5),
.O(LIOB33_X0Y131_IOB_X0Y131_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y131_IOB_X0Y132_OBUF (
.I(CLBLM_R_X7Y131_SLICE_X9Y131_AQ),
.O(LIOB33_X0Y131_IOB_X0Y132_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y133_IOB_X0Y133_OBUF (
.I(CLBLM_R_X3Y137_SLICE_X3Y137_AQ),
.O(LIOB33_X0Y133_IOB_X0Y133_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y133_IOB_X0Y134_OBUF (
.I(CLBLM_R_X3Y133_SLICE_X3Y133_AQ),
.O(LIOB33_X0Y133_IOB_X0Y134_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y135_IOB_X0Y135_OBUF (
.I(CLBLM_R_X3Y136_SLICE_X3Y136_AQ),
.O(LIOB33_X0Y135_IOB_X0Y135_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y135_IOB_X0Y136_OBUF (
.I(CLBLM_R_X3Y135_SLICE_X3Y135_AQ),
.O(LIOB33_X0Y135_IOB_X0Y136_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y137_IOB_X0Y137_OBUF (
.I(CLBLM_R_X3Y137_SLICE_X2Y137_BQ),
.O(LIOB33_X0Y137_IOB_X0Y137_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y137_IOB_X0Y138_OBUF (
.I(CLBLM_R_X3Y136_SLICE_X3Y136_DQ),
.O(LIOB33_X0Y137_IOB_X0Y138_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y139_IOB_X0Y139_OBUF (
.I(CLBLM_R_X3Y137_SLICE_X2Y137_AQ),
.O(LIOB33_X0Y139_IOB_X0Y139_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y139_IOB_X0Y140_OBUF (
.I(CLBLM_R_X3Y136_SLICE_X2Y136_AQ),
.O(LIOB33_X0Y139_IOB_X0Y140_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y141_IOB_X0Y141_OBUF (
.I(CLBLM_R_X3Y136_SLICE_X3Y136_BQ),
.O(LIOB33_X0Y141_IOB_X0Y141_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y141_IOB_X0Y142_OBUF (
.I(LIOB33_X0Y53_IOB_X0Y54_I),
.O(LIOB33_X0Y141_IOB_X0Y142_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y143_IOB_X0Y143_OBUF (
.I(LIOB33_X0Y55_IOB_X0Y55_I),
.O(LIOB33_X0Y143_IOB_X0Y143_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y145_IOB_X0Y145_OBUF (
.I(LIOB33_X0Y57_IOB_X0Y58_I),
.O(LIOB33_X0Y145_IOB_X0Y145_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y145_IOB_X0Y146_OBUF (
.I(LIOB33_X0Y59_IOB_X0Y59_I),
.O(LIOB33_X0Y145_IOB_X0Y146_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y147_IOB_X0Y147_OBUF (
.I(LIOB33_X0Y71_IOB_X0Y71_I),
.O(LIOB33_X0Y147_IOB_X0Y147_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y147_IOB_X0Y148_OBUF (
.I(LIOB33_X0Y61_IOB_X0Y61_I),
.O(LIOB33_X0Y147_IOB_X0Y148_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y151_IOB_X0Y151_OBUF (
.I(LIOB33_X0Y65_IOB_X0Y65_I),
.O(LIOB33_X0Y151_IOB_X0Y151_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y151_IOB_X0Y152_OBUF (
.I(LIOB33_X0Y65_IOB_X0Y66_I),
.O(LIOB33_X0Y151_IOB_X0Y152_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y153_IOB_X0Y153_OBUF (
.I(LIOB33_X0Y67_IOB_X0Y67_I),
.O(LIOB33_X0Y153_IOB_X0Y153_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y153_IOB_X0Y154_OBUF (
.I(LIOB33_X0Y67_IOB_X0Y68_I),
.O(LIOB33_X0Y153_IOB_X0Y154_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y155_IOB_X0Y155_OBUF (
.I(LIOB33_X0Y69_IOB_X0Y70_I),
.O(LIOB33_X0Y155_IOB_X0Y155_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y155_IOB_X0Y156_OBUF (
.I(RIOB33_X105Y105_IOB_X1Y106_I),
.O(LIOB33_X0Y155_IOB_X0Y156_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y157_IOB_X0Y157_OBUF (
.I(RIOB33_X105Y115_IOB_X1Y115_I),
.O(LIOB33_X0Y157_IOB_X0Y157_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y157_IOB_X0Y158_OBUF (
.I(RIOB33_X105Y115_IOB_X1Y116_I),
.O(LIOB33_X0Y157_IOB_X0Y158_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y159_IOB_X0Y159_OBUF (
.I(RIOB33_X105Y117_IOB_X1Y117_I),
.O(LIOB33_X0Y159_IOB_X0Y159_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y159_IOB_X0Y160_OBUF (
.I(RIOB33_X105Y107_IOB_X1Y107_I),
.O(LIOB33_X0Y159_IOB_X0Y160_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y161_IOB_X0Y161_OBUF (
.I(RIOB33_X105Y107_IOB_X1Y108_I),
.O(LIOB33_X0Y161_IOB_X0Y161_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y161_IOB_X0Y162_OBUF (
.I(RIOB33_X105Y109_IOB_X1Y109_I),
.O(LIOB33_X0Y161_IOB_X0Y162_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y163_IOB_X0Y163_OBUF (
.I(RIOB33_X105Y109_IOB_X1Y110_I),
.O(LIOB33_X0Y163_IOB_X0Y163_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y163_IOB_X0Y164_OBUF (
.I(RIOB33_X105Y111_IOB_X1Y111_I),
.O(LIOB33_X0Y163_IOB_X0Y164_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y165_IOB_X0Y165_OBUF (
.I(RIOB33_X105Y111_IOB_X1Y112_I),
.O(LIOB33_X0Y165_IOB_X0Y165_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y165_IOB_X0Y166_OBUF (
.I(RIOB33_X105Y113_IOB_X1Y113_I),
.O(LIOB33_X0Y165_IOB_X0Y166_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y167_IOB_X0Y167_OBUF (
.I(RIOB33_X105Y113_IOB_X1Y114_I),
.O(LIOB33_X0Y167_IOB_X0Y167_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y167_IOB_X0Y168_OBUF (
.I(RIOB33_X105Y123_IOB_X1Y123_I),
.O(LIOB33_X0Y167_IOB_X0Y168_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y169_IOB_X0Y169_OBUF (
.I(RIOB33_X105Y121_IOB_X1Y122_I),
.O(LIOB33_X0Y169_IOB_X0Y169_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y169_IOB_X0Y170_OBUF (
.I(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.O(LIOB33_X0Y169_IOB_X0Y170_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y171_IOB_X0Y171_OBUF (
.I(LIOB33_SING_X0Y50_IOB_X0Y50_I),
.O(LIOB33_X0Y171_IOB_X0Y171_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y171_IOB_X0Y172_OBUF (
.I(CLBLM_R_X103Y140_SLICE_X163Y140_AO6),
.O(LIOB33_X0Y171_IOB_X0Y172_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y173_IOB_X0Y173_OBUF (
.I(CLBLM_R_X103Y140_SLICE_X163Y140_AO5),
.O(LIOB33_X0Y173_IOB_X0Y173_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y173_IOB_X0Y174_OBUF (
.I(CLBLM_R_X11Y153_SLICE_X14Y153_AO6),
.O(LIOB33_X0Y173_IOB_X0Y174_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y175_IOB_X0Y175_OBUF (
.I(RIOB33_X105Y127_IOB_X1Y127_I),
.O(LIOB33_X0Y175_IOB_X0Y175_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y175_IOB_X0Y176_OBUF (
.I(RIOB33_X105Y127_IOB_X1Y128_I),
.O(LIOB33_X0Y175_IOB_X0Y176_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y177_IOB_X0Y177_OBUF (
.I(RIOB33_X105Y129_IOB_X1Y129_I),
.O(LIOB33_X0Y177_IOB_X0Y177_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y177_IOB_X0Y178_OBUF (
.I(RIOB33_X105Y129_IOB_X1Y130_I),
.O(LIOB33_X0Y177_IOB_X0Y178_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y179_IOB_X0Y179_OBUF (
.I(RIOB33_X105Y131_IOB_X1Y131_I),
.O(LIOB33_X0Y179_IOB_X0Y179_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y179_IOB_X0Y180_OBUF (
.I(RIOB33_X105Y131_IOB_X1Y132_I),
.O(LIOB33_X0Y179_IOB_X0Y180_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y181_IOB_X0Y181_OBUF (
.I(RIOB33_X105Y133_IOB_X1Y133_I),
.O(LIOB33_X0Y181_IOB_X0Y181_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y181_IOB_X0Y182_OBUF (
.I(RIOB33_X105Y133_IOB_X1Y134_I),
.O(LIOB33_X0Y181_IOB_X0Y182_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y183_IOB_X0Y183_OBUF (
.I(RIOB33_X105Y135_IOB_X1Y135_I),
.O(LIOB33_X0Y183_IOB_X0Y183_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y183_IOB_X0Y184_OBUF (
.I(RIOB33_X105Y135_IOB_X1Y136_I),
.O(LIOB33_X0Y183_IOB_X0Y184_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y185_IOB_X0Y185_OBUF (
.I(RIOB33_X105Y137_IOB_X1Y137_I),
.O(LIOB33_X0Y185_IOB_X0Y185_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y185_IOB_X0Y186_OBUF (
.I(RIOB33_X105Y143_IOB_X1Y143_I),
.O(LIOB33_X0Y185_IOB_X0Y186_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y187_IOB_X0Y187_OBUF (
.I(RIOB33_X105Y143_IOB_X1Y144_I),
.O(LIOB33_X0Y187_IOB_X0Y187_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y187_IOB_X0Y188_OBUF (
.I(RIOB33_X105Y145_IOB_X1Y145_I),
.O(LIOB33_X0Y187_IOB_X0Y188_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y189_IOB_X0Y189_OBUF (
.I(RIOB33_X105Y145_IOB_X1Y146_I),
.O(LIOB33_X0Y189_IOB_X0Y189_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y189_IOB_X0Y190_OBUF (
.I(RIOB33_X105Y147_IOB_X1Y147_I),
.O(LIOB33_X0Y189_IOB_X0Y190_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y191_IOB_X0Y191_OBUF (
.I(RIOB33_X105Y147_IOB_X1Y148_I),
.O(LIOB33_X0Y191_IOB_X0Y191_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y191_IOB_X0Y192_OBUF (
.I(LIOB33_X0Y51_IOB_X0Y52_I),
.O(LIOB33_X0Y191_IOB_X0Y192_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y193_IOB_X0Y193_OBUF (
.I(LIOB33_X0Y55_IOB_X0Y56_I),
.O(LIOB33_X0Y193_IOB_X0Y193_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y193_IOB_X0Y194_OBUF (
.I(LIOB33_X0Y59_IOB_X0Y60_I),
.O(LIOB33_X0Y193_IOB_X0Y194_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y195_IOB_X0Y195_OBUF (
.I(LIOB33_X0Y63_IOB_X0Y64_I),
.O(LIOB33_X0Y195_IOB_X0Y195_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y195_IOB_X0Y196_OBUF (
.I(LIOB33_X0Y69_IOB_X0Y69_I),
.O(LIOB33_X0Y195_IOB_X0Y196_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y197_IOB_X0Y197_OBUF (
.I(LIOB33_X0Y71_IOB_X0Y72_I),
.O(LIOB33_X0Y197_IOB_X0Y197_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y197_IOB_X0Y198_OBUF (
.I(LIOB33_X0Y73_IOB_X0Y73_I),
.O(LIOB33_X0Y197_IOB_X0Y198_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_SING_X0Y50_IOB_X0Y50_IBUF (
.I(LIOB33_SING_X0Y50_IOB_X0Y50_IPAD),
.O(LIOB33_SING_X0Y50_IOB_X0Y50_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y100_IOB_X0Y100_OBUF (
.I(CLBLL_L_X2Y133_SLICE_X0Y133_BO6),
.O(LIOB33_SING_X0Y100_IOB_X0Y100_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y149_IOB_X0Y149_OBUF (
.I(LIOB33_X0Y61_IOB_X0Y62_I),
.O(LIOB33_SING_X0Y149_IOB_X0Y149_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y150_IOB_X0Y150_OBUF (
.I(LIOB33_X0Y63_IOB_X0Y63_I),
.O(LIOB33_SING_X0Y150_IOB_X0Y150_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y199_IOB_X0Y199_OBUF (
.I(LIOB33_X0Y73_IOB_X0Y74_I),
.O(LIOB33_SING_X0Y199_IOB_X0Y199_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y101_IOB_X1Y101_IBUF (
.I(RIOB33_X105Y101_IOB_X1Y101_IPAD),
.O(RIOB33_X105Y101_IOB_X1Y101_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y101_IOB_X1Y102_IBUF (
.I(RIOB33_X105Y101_IOB_X1Y102_IPAD),
.O(RIOB33_X105Y101_IOB_X1Y102_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y103_IOB_X1Y103_IBUF (
.I(RIOB33_X105Y103_IOB_X1Y103_IPAD),
.O(RIOB33_X105Y103_IOB_X1Y103_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y103_IOB_X1Y104_IBUF (
.I(RIOB33_X105Y103_IOB_X1Y104_IPAD),
.O(RIOB33_X105Y103_IOB_X1Y104_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y105_IOB_X1Y105_IBUF (
.I(RIOB33_X105Y105_IOB_X1Y105_IPAD),
.O(RIOB33_X105Y105_IOB_X1Y105_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y105_IOB_X1Y106_IBUF (
.I(RIOB33_X105Y105_IOB_X1Y106_IPAD),
.O(RIOB33_X105Y105_IOB_X1Y106_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y107_IOB_X1Y107_IBUF (
.I(RIOB33_X105Y107_IOB_X1Y107_IPAD),
.O(RIOB33_X105Y107_IOB_X1Y107_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y107_IOB_X1Y108_IBUF (
.I(RIOB33_X105Y107_IOB_X1Y108_IPAD),
.O(RIOB33_X105Y107_IOB_X1Y108_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y109_IOB_X1Y109_IBUF (
.I(RIOB33_X105Y109_IOB_X1Y109_IPAD),
.O(RIOB33_X105Y109_IOB_X1Y109_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y109_IOB_X1Y110_IBUF (
.I(RIOB33_X105Y109_IOB_X1Y110_IPAD),
.O(RIOB33_X105Y109_IOB_X1Y110_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y111_IOB_X1Y111_IBUF (
.I(RIOB33_X105Y111_IOB_X1Y111_IPAD),
.O(RIOB33_X105Y111_IOB_X1Y111_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y111_IOB_X1Y112_IBUF (
.I(RIOB33_X105Y111_IOB_X1Y112_IPAD),
.O(RIOB33_X105Y111_IOB_X1Y112_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y113_IOB_X1Y113_IBUF (
.I(RIOB33_X105Y113_IOB_X1Y113_IPAD),
.O(RIOB33_X105Y113_IOB_X1Y113_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y113_IOB_X1Y114_IBUF (
.I(RIOB33_X105Y113_IOB_X1Y114_IPAD),
.O(RIOB33_X105Y113_IOB_X1Y114_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y115_IOB_X1Y115_IBUF (
.I(RIOB33_X105Y115_IOB_X1Y115_IPAD),
.O(RIOB33_X105Y115_IOB_X1Y115_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y115_IOB_X1Y116_IBUF (
.I(RIOB33_X105Y115_IOB_X1Y116_IPAD),
.O(RIOB33_X105Y115_IOB_X1Y116_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y117_IOB_X1Y117_IBUF (
.I(RIOB33_X105Y117_IOB_X1Y117_IPAD),
.O(RIOB33_X105Y117_IOB_X1Y117_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y117_IOB_X1Y118_IBUF (
.I(RIOB33_X105Y117_IOB_X1Y118_IPAD),
.O(RIOB33_X105Y117_IOB_X1Y118_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y119_IOB_X1Y119_IBUF (
.I(RIOB33_X105Y119_IOB_X1Y119_IPAD),
.O(RIOB33_X105Y119_IOB_X1Y119_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y119_IOB_X1Y120_IBUF (
.I(RIOB33_X105Y119_IOB_X1Y120_IPAD),
.O(RIOB33_X105Y119_IOB_X1Y120_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y121_IOB_X1Y121_IBUF (
.I(RIOB33_X105Y121_IOB_X1Y121_IPAD),
.O(RIOB33_X105Y121_IOB_X1Y121_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y121_IOB_X1Y122_IBUF (
.I(RIOB33_X105Y121_IOB_X1Y122_IPAD),
.O(RIOB33_X105Y121_IOB_X1Y122_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y123_IOB_X1Y123_IBUF (
.I(RIOB33_X105Y123_IOB_X1Y123_IPAD),
.O(RIOB33_X105Y123_IOB_X1Y123_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y123_IOB_X1Y124_IBUF (
.I(RIOB33_X105Y123_IOB_X1Y124_IPAD),
.O(RIOB33_X105Y123_IOB_X1Y124_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y125_IOB_X1Y125_IBUF (
.I(RIOB33_X105Y125_IOB_X1Y125_IPAD),
.O(RIOB33_X105Y125_IOB_X1Y125_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y125_IOB_X1Y126_IBUF (
.I(RIOB33_X105Y125_IOB_X1Y126_IPAD),
.O(RIOB33_X105Y125_IOB_X1Y126_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y127_IOB_X1Y127_IBUF (
.I(RIOB33_X105Y127_IOB_X1Y127_IPAD),
.O(RIOB33_X105Y127_IOB_X1Y127_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y127_IOB_X1Y128_IBUF (
.I(RIOB33_X105Y127_IOB_X1Y128_IPAD),
.O(RIOB33_X105Y127_IOB_X1Y128_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y129_IOB_X1Y129_IBUF (
.I(RIOB33_X105Y129_IOB_X1Y129_IPAD),
.O(RIOB33_X105Y129_IOB_X1Y129_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y129_IOB_X1Y130_IBUF (
.I(RIOB33_X105Y129_IOB_X1Y130_IPAD),
.O(RIOB33_X105Y129_IOB_X1Y130_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y131_IOB_X1Y131_IBUF (
.I(RIOB33_X105Y131_IOB_X1Y131_IPAD),
.O(RIOB33_X105Y131_IOB_X1Y131_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y131_IOB_X1Y132_IBUF (
.I(RIOB33_X105Y131_IOB_X1Y132_IPAD),
.O(RIOB33_X105Y131_IOB_X1Y132_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y133_IOB_X1Y133_IBUF (
.I(RIOB33_X105Y133_IOB_X1Y133_IPAD),
.O(RIOB33_X105Y133_IOB_X1Y133_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y133_IOB_X1Y134_IBUF (
.I(RIOB33_X105Y133_IOB_X1Y134_IPAD),
.O(RIOB33_X105Y133_IOB_X1Y134_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y135_IOB_X1Y135_IBUF (
.I(RIOB33_X105Y135_IOB_X1Y135_IPAD),
.O(RIOB33_X105Y135_IOB_X1Y135_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y135_IOB_X1Y136_IBUF (
.I(RIOB33_X105Y135_IOB_X1Y136_IPAD),
.O(RIOB33_X105Y135_IOB_X1Y136_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y137_IOB_X1Y137_IBUF (
.I(RIOB33_X105Y137_IOB_X1Y137_IPAD),
.O(RIOB33_X105Y137_IOB_X1Y137_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y137_IOB_X1Y138_IBUF (
.I(RIOB33_X105Y137_IOB_X1Y138_IPAD),
.O(RIOB33_X105Y137_IOB_X1Y138_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y139_IOB_X1Y139_IBUF (
.I(RIOB33_X105Y139_IOB_X1Y139_IPAD),
.O(RIOB33_X105Y139_IOB_X1Y139_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y139_IOB_X1Y140_IBUF (
.I(RIOB33_X105Y139_IOB_X1Y140_IPAD),
.O(RIOB33_X105Y139_IOB_X1Y140_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y141_IOB_X1Y141_IBUF (
.I(RIOB33_X105Y141_IOB_X1Y141_IPAD),
.O(RIOB33_X105Y141_IOB_X1Y141_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y141_IOB_X1Y142_IBUF (
.I(RIOB33_X105Y141_IOB_X1Y142_IPAD),
.O(RIOB33_X105Y141_IOB_X1Y142_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y143_IOB_X1Y143_IBUF (
.I(RIOB33_X105Y143_IOB_X1Y143_IPAD),
.O(RIOB33_X105Y143_IOB_X1Y143_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y143_IOB_X1Y144_IBUF (
.I(RIOB33_X105Y143_IOB_X1Y144_IPAD),
.O(RIOB33_X105Y143_IOB_X1Y144_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y145_IOB_X1Y145_IBUF (
.I(RIOB33_X105Y145_IOB_X1Y145_IPAD),
.O(RIOB33_X105Y145_IOB_X1Y145_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y145_IOB_X1Y146_IBUF (
.I(RIOB33_X105Y145_IOB_X1Y146_IPAD),
.O(RIOB33_X105Y145_IOB_X1Y146_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y147_IOB_X1Y147_IBUF (
.I(RIOB33_X105Y147_IOB_X1Y147_IPAD),
.O(RIOB33_X105Y147_IOB_X1Y147_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y147_IOB_X1Y148_IBUF (
.I(RIOB33_X105Y147_IOB_X1Y148_IPAD),
.O(RIOB33_X105Y147_IOB_X1Y148_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y151_IOB_X1Y151_OBUF (
.I(LIOB33_X0Y75_IOB_X0Y76_I),
.O(RIOB33_X105Y151_IOB_X1Y151_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y151_IOB_X1Y152_OBUF (
.I(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.O(RIOB33_X105Y151_IOB_X1Y152_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y153_IOB_X1Y153_OBUF (
.I(RIOB33_X105Y101_IOB_X1Y101_I),
.O(RIOB33_X105Y153_IOB_X1Y153_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y153_IOB_X1Y154_OBUF (
.I(RIOB33_X105Y101_IOB_X1Y102_I),
.O(RIOB33_X105Y153_IOB_X1Y154_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y155_IOB_X1Y155_OBUF (
.I(RIOB33_X105Y103_IOB_X1Y103_I),
.O(RIOB33_X105Y155_IOB_X1Y155_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y155_IOB_X1Y156_OBUF (
.I(RIOB33_X105Y103_IOB_X1Y104_I),
.O(RIOB33_X105Y155_IOB_X1Y156_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y157_IOB_X1Y157_OBUF (
.I(RIOB33_X105Y125_IOB_X1Y126_I),
.O(RIOB33_X105Y157_IOB_X1Y157_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y157_IOB_X1Y158_OBUF (
.I(CLBLM_R_X37Y138_SLICE_X56Y138_AO6),
.O(RIOB33_X105Y157_IOB_X1Y158_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y159_IOB_X1Y159_OBUF (
.I(CLBLM_L_X12Y138_SLICE_X17Y138_DO6),
.O(RIOB33_X105Y159_IOB_X1Y159_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y159_IOB_X1Y160_OBUF (
.I(CLBLM_L_X12Y138_SLICE_X17Y138_DO5),
.O(RIOB33_X105Y159_IOB_X1Y160_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y161_IOB_X1Y161_OBUF (
.I(CLBLM_R_X11Y141_SLICE_X14Y141_CO6),
.O(RIOB33_X105Y161_IOB_X1Y161_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y161_IOB_X1Y162_OBUF (
.I(CLBLM_R_X11Y141_SLICE_X14Y141_CO5),
.O(RIOB33_X105Y161_IOB_X1Y162_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y163_IOB_X1Y163_OBUF (
.I(CLBLM_L_X12Y139_SLICE_X17Y139_DO6),
.O(RIOB33_X105Y163_IOB_X1Y163_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y163_IOB_X1Y164_OBUF (
.I(CLBLM_L_X12Y139_SLICE_X17Y139_DO5),
.O(RIOB33_X105Y163_IOB_X1Y164_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y165_IOB_X1Y165_OBUF (
.I(RIOB33_X105Y125_IOB_X1Y125_I),
.O(RIOB33_X105Y165_IOB_X1Y165_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y165_IOB_X1Y166_OBUF (
.I(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.O(RIOB33_X105Y165_IOB_X1Y166_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y167_IOB_X1Y167_OBUF (
.I(LIOB33_SING_X0Y50_IOB_X0Y50_I),
.O(RIOB33_X105Y167_IOB_X1Y167_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y167_IOB_X1Y168_OBUF (
.I(CLBLM_R_X11Y153_SLICE_X14Y153_AO6),
.O(RIOB33_X105Y167_IOB_X1Y168_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y169_IOB_X1Y169_OBUF (
.I(CLBLM_R_X103Y169_SLICE_X163Y169_AO6),
.O(RIOB33_X105Y169_IOB_X1Y169_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y169_IOB_X1Y170_OBUF (
.I(CLBLM_R_X103Y170_SLICE_X163Y170_AO6),
.O(RIOB33_X105Y169_IOB_X1Y170_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y171_IOB_X1Y171_OBUF (
.I(CLBLM_L_X10Y146_SLICE_X12Y146_AO5),
.O(RIOB33_X105Y171_IOB_X1Y171_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y171_IOB_X1Y172_OBUF (
.I(CLBLM_R_X103Y170_SLICE_X163Y170_AO5),
.O(RIOB33_X105Y171_IOB_X1Y172_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y173_IOB_X1Y173_OBUF (
.I(CLBLM_R_X11Y144_SLICE_X14Y144_BO5),
.O(RIOB33_X105Y173_IOB_X1Y173_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y173_IOB_X1Y174_OBUF (
.I(CLBLM_R_X103Y173_SLICE_X163Y173_AO6),
.O(RIOB33_X105Y173_IOB_X1Y174_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y175_IOB_X1Y175_OBUF (
.I(CLBLM_L_X12Y146_SLICE_X16Y146_AO6),
.O(RIOB33_X105Y175_IOB_X1Y175_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y175_IOB_X1Y176_OBUF (
.I(CLBLM_R_X103Y173_SLICE_X163Y173_AO5),
.O(RIOB33_X105Y175_IOB_X1Y176_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y177_IOB_X1Y177_OBUF (
.I(CLBLM_R_X103Y177_SLICE_X163Y177_AO6),
.O(RIOB33_X105Y177_IOB_X1Y177_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y177_IOB_X1Y178_OBUF (
.I(CLBLM_R_X103Y177_SLICE_X163Y177_AO5),
.O(RIOB33_X105Y177_IOB_X1Y178_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y179_IOB_X1Y179_OBUF (
.I(CLBLM_L_X12Y144_SLICE_X17Y144_AO5),
.O(RIOB33_X105Y179_IOB_X1Y179_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y179_IOB_X1Y180_OBUF (
.I(CLBLM_L_X12Y138_SLICE_X17Y138_DO6),
.O(RIOB33_X105Y179_IOB_X1Y180_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y181_IOB_X1Y181_OBUF (
.I(CLBLM_L_X12Y138_SLICE_X17Y138_DO5),
.O(RIOB33_X105Y181_IOB_X1Y181_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y181_IOB_X1Y182_OBUF (
.I(CLBLM_R_X11Y141_SLICE_X14Y141_CO6),
.O(RIOB33_X105Y181_IOB_X1Y182_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y183_IOB_X1Y183_OBUF (
.I(CLBLM_R_X11Y141_SLICE_X14Y141_CO5),
.O(RIOB33_X105Y183_IOB_X1Y183_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y183_IOB_X1Y184_OBUF (
.I(CLBLM_L_X12Y139_SLICE_X17Y139_DO6),
.O(RIOB33_X105Y183_IOB_X1Y184_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y185_IOB_X1Y185_OBUF (
.I(CLBLM_L_X12Y139_SLICE_X17Y139_DO5),
.O(RIOB33_X105Y185_IOB_X1Y185_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y185_IOB_X1Y186_OBUF (
.I(CLBLM_R_X13Y139_SLICE_X19Y139_AQ),
.O(RIOB33_X105Y185_IOB_X1Y186_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y187_IOB_X1Y187_OBUF (
.I(CLBLM_L_X12Y134_SLICE_X16Y134_AQ),
.O(RIOB33_X105Y187_IOB_X1Y187_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y187_IOB_X1Y188_OBUF (
.I(CLBLM_R_X11Y144_SLICE_X15Y144_AQ),
.O(RIOB33_X105Y187_IOB_X1Y188_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y189_IOB_X1Y189_OBUF (
.I(CLBLM_L_X10Y143_SLICE_X13Y143_BQ),
.O(RIOB33_X105Y189_IOB_X1Y189_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y189_IOB_X1Y190_OBUF (
.I(CLBLM_R_X15Y142_SLICE_X20Y142_AQ),
.O(RIOB33_X105Y189_IOB_X1Y190_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y191_IOB_X1Y191_OBUF (
.I(CLBLM_L_X10Y143_SLICE_X13Y143_AQ),
.O(RIOB33_X105Y191_IOB_X1Y191_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y191_IOB_X1Y192_OBUF (
.I(CLBLM_R_X13Y134_SLICE_X19Y134_BQ),
.O(RIOB33_X105Y191_IOB_X1Y192_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y193_IOB_X1Y193_OBUF (
.I(CLBLM_L_X12Y144_SLICE_X16Y144_AQ),
.O(RIOB33_X105Y193_IOB_X1Y193_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y193_IOB_X1Y194_OBUF (
.I(CLBLM_R_X13Y144_SLICE_X19Y144_AQ),
.O(RIOB33_X105Y193_IOB_X1Y194_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y195_IOB_X1Y195_OBUF (
.I(CLBLM_R_X13Y143_SLICE_X18Y143_BQ),
.O(RIOB33_X105Y195_IOB_X1Y195_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y195_IOB_X1Y196_OBUF (
.I(CLBLM_R_X13Y143_SLICE_X18Y143_AQ),
.O(RIOB33_X105Y195_IOB_X1Y196_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y197_IOB_X1Y197_OBUF (
.I(CLBLM_R_X103Y175_SLICE_X163Y175_AO6),
.O(RIOB33_X105Y197_IOB_X1Y197_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y197_IOB_X1Y198_OBUF (
.I(CLBLM_R_X103Y175_SLICE_X163Y175_AO6),
.O(RIOB33_X105Y197_IOB_X1Y198_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_SING_X105Y100_IOB_X1Y100_IBUF (
.I(RIOB33_SING_X105Y100_IOB_X1Y100_IPAD),
.O(RIOB33_SING_X105Y100_IOB_X1Y100_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_SING_X105Y149_IOB_X1Y149_IBUF (
.I(RIOB33_SING_X105Y149_IOB_X1Y149_IPAD),
.O(RIOB33_SING_X105Y149_IOB_X1Y149_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_SING_X105Y150_IOB_X1Y150_OBUF (
.I(LIOB33_X0Y75_IOB_X0Y75_I),
.O(RIOB33_SING_X105Y150_IOB_X1Y150_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_SING_X105Y199_IOB_X1Y199_OBUF (
.I(CLBLM_R_X13Y144_SLICE_X19Y144_AQ),
.O(RIOB33_SING_X105Y199_IOB_X1Y199_OPAD)
  );
  assign CLBLL_L_X2Y108_SLICE_X0Y108_A = CLBLL_L_X2Y108_SLICE_X0Y108_AO6;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_B = CLBLL_L_X2Y108_SLICE_X0Y108_BO6;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_C = CLBLL_L_X2Y108_SLICE_X0Y108_CO6;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_D = CLBLL_L_X2Y108_SLICE_X0Y108_DO6;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_A = CLBLL_L_X2Y108_SLICE_X1Y108_AO6;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_B = CLBLL_L_X2Y108_SLICE_X1Y108_BO6;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_C = CLBLL_L_X2Y108_SLICE_X1Y108_CO6;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_D = CLBLL_L_X2Y108_SLICE_X1Y108_DO6;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_A = CLBLL_L_X2Y127_SLICE_X0Y127_AO6;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_B = CLBLL_L_X2Y127_SLICE_X0Y127_BO6;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_C = CLBLL_L_X2Y127_SLICE_X0Y127_CO6;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_D = CLBLL_L_X2Y127_SLICE_X0Y127_DO6;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_AMUX = CLBLL_L_X2Y127_SLICE_X0Y127_AO5;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_A = CLBLL_L_X2Y127_SLICE_X1Y127_AO6;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_B = CLBLL_L_X2Y127_SLICE_X1Y127_BO6;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_C = CLBLL_L_X2Y127_SLICE_X1Y127_CO6;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_D = CLBLL_L_X2Y127_SLICE_X1Y127_DO6;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_A = CLBLL_L_X2Y133_SLICE_X0Y133_AO6;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_B = CLBLL_L_X2Y133_SLICE_X0Y133_BO6;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_C = CLBLL_L_X2Y133_SLICE_X0Y133_CO6;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_D = CLBLL_L_X2Y133_SLICE_X0Y133_DO6;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_AMUX = CLBLL_L_X2Y133_SLICE_X0Y133_AO5;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_BMUX = CLBLL_L_X2Y133_SLICE_X0Y133_BO5;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_CMUX = CLBLL_L_X2Y133_SLICE_X0Y133_CO5;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_A = CLBLL_L_X2Y133_SLICE_X1Y133_AO6;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_B = CLBLL_L_X2Y133_SLICE_X1Y133_BO6;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_C = CLBLL_L_X2Y133_SLICE_X1Y133_CO6;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_D = CLBLL_L_X2Y133_SLICE_X1Y133_DO6;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_A = CLBLL_L_X2Y140_SLICE_X0Y140_AO6;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_B = CLBLL_L_X2Y140_SLICE_X0Y140_BO6;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_C = CLBLL_L_X2Y140_SLICE_X0Y140_CO6;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_D = CLBLL_L_X2Y140_SLICE_X0Y140_DO6;
  assign CLBLL_L_X2Y140_SLICE_X1Y140_A = CLBLL_L_X2Y140_SLICE_X1Y140_AO6;
  assign CLBLL_L_X2Y140_SLICE_X1Y140_B = CLBLL_L_X2Y140_SLICE_X1Y140_BO6;
  assign CLBLL_L_X2Y140_SLICE_X1Y140_C = CLBLL_L_X2Y140_SLICE_X1Y140_CO6;
  assign CLBLL_L_X2Y140_SLICE_X1Y140_D = CLBLL_L_X2Y140_SLICE_X1Y140_DO6;
  assign CLBLL_L_X2Y140_SLICE_X1Y140_AMUX = CLBLL_L_X2Y140_SLICE_X1Y140_AO5;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_A = CLBLL_L_X2Y141_SLICE_X0Y141_AO6;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_B = CLBLL_L_X2Y141_SLICE_X0Y141_BO6;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_C = CLBLL_L_X2Y141_SLICE_X0Y141_CO6;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_D = CLBLL_L_X2Y141_SLICE_X0Y141_DO6;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_AMUX = CLBLL_L_X2Y141_SLICE_X0Y141_AO6;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_A = CLBLL_L_X2Y141_SLICE_X1Y141_AO6;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_B = CLBLL_L_X2Y141_SLICE_X1Y141_BO6;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_C = CLBLL_L_X2Y141_SLICE_X1Y141_CO6;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_D = CLBLL_L_X2Y141_SLICE_X1Y141_DO6;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_AMUX = CLBLL_L_X2Y141_SLICE_X1Y141_AO5;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_BMUX = CLBLL_L_X2Y141_SLICE_X1Y141_BO5;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_A = CLBLL_L_X4Y132_SLICE_X4Y132_AO6;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_B = CLBLL_L_X4Y132_SLICE_X4Y132_BO6;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_C = CLBLL_L_X4Y132_SLICE_X4Y132_CO6;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_D = CLBLL_L_X4Y132_SLICE_X4Y132_DO6;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_A = CLBLL_L_X4Y132_SLICE_X5Y132_AO6;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_B = CLBLL_L_X4Y132_SLICE_X5Y132_BO6;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_C = CLBLL_L_X4Y132_SLICE_X5Y132_CO6;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_D = CLBLL_L_X4Y132_SLICE_X5Y132_DO6;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_A = CLBLL_L_X4Y133_SLICE_X4Y133_AO6;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_B = CLBLL_L_X4Y133_SLICE_X4Y133_BO6;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_C = CLBLL_L_X4Y133_SLICE_X4Y133_CO6;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_D = CLBLL_L_X4Y133_SLICE_X4Y133_DO6;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_BMUX = CLBLL_L_X4Y133_SLICE_X4Y133_BO5;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_A = CLBLL_L_X4Y133_SLICE_X5Y133_AO6;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_B = CLBLL_L_X4Y133_SLICE_X5Y133_BO6;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_C = CLBLL_L_X4Y133_SLICE_X5Y133_CO6;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_D = CLBLL_L_X4Y133_SLICE_X5Y133_DO6;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_AMUX = CLBLL_L_X4Y133_SLICE_X5Y133_A5Q;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_A = CLBLL_L_X4Y134_SLICE_X4Y134_AO6;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_B = CLBLL_L_X4Y134_SLICE_X4Y134_BO6;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_C = CLBLL_L_X4Y134_SLICE_X4Y134_CO6;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_D = CLBLL_L_X4Y134_SLICE_X4Y134_DO6;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_BMUX = CLBLL_L_X4Y134_SLICE_X4Y134_B5Q;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_A = CLBLL_L_X4Y134_SLICE_X5Y134_AO6;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_B = CLBLL_L_X4Y134_SLICE_X5Y134_BO6;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_C = CLBLL_L_X4Y134_SLICE_X5Y134_CO6;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_D = CLBLL_L_X4Y134_SLICE_X5Y134_DO6;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_AMUX = CLBLL_L_X4Y134_SLICE_X5Y134_A5Q;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_DMUX = CLBLL_L_X4Y134_SLICE_X5Y134_DO5;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_A = CLBLL_L_X4Y135_SLICE_X4Y135_AO6;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_B = CLBLL_L_X4Y135_SLICE_X4Y135_BO6;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_C = CLBLL_L_X4Y135_SLICE_X4Y135_CO6;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_D = CLBLL_L_X4Y135_SLICE_X4Y135_DO6;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_AMUX = CLBLL_L_X4Y135_SLICE_X4Y135_A5Q;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_DMUX = CLBLL_L_X4Y135_SLICE_X4Y135_DO5;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_A = CLBLL_L_X4Y135_SLICE_X5Y135_AO6;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_B = CLBLL_L_X4Y135_SLICE_X5Y135_BO6;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_C = CLBLL_L_X4Y135_SLICE_X5Y135_CO6;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_D = CLBLL_L_X4Y135_SLICE_X5Y135_DO6;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_CMUX = CLBLL_L_X4Y135_SLICE_X5Y135_C5Q;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_DMUX = CLBLL_L_X4Y135_SLICE_X5Y135_D5Q;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_A = CLBLL_L_X4Y136_SLICE_X4Y136_AO6;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_B = CLBLL_L_X4Y136_SLICE_X4Y136_BO6;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_C = CLBLL_L_X4Y136_SLICE_X4Y136_CO6;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_D = CLBLL_L_X4Y136_SLICE_X4Y136_DO6;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_AMUX = CLBLL_L_X4Y136_SLICE_X4Y136_AO5;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_DMUX = CLBLL_L_X4Y136_SLICE_X4Y136_D5Q;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_A = CLBLL_L_X4Y136_SLICE_X5Y136_AO6;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_B = CLBLL_L_X4Y136_SLICE_X5Y136_BO6;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_C = CLBLL_L_X4Y136_SLICE_X5Y136_CO6;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_D = CLBLL_L_X4Y136_SLICE_X5Y136_DO6;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_AMUX = CLBLL_L_X4Y136_SLICE_X5Y136_A5Q;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_DMUX = CLBLL_L_X4Y136_SLICE_X5Y136_DO5;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_A = CLBLL_L_X4Y137_SLICE_X4Y137_AO6;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_B = CLBLL_L_X4Y137_SLICE_X4Y137_BO6;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_C = CLBLL_L_X4Y137_SLICE_X4Y137_CO6;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_D = CLBLL_L_X4Y137_SLICE_X4Y137_DO6;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_AMUX = CLBLL_L_X4Y137_SLICE_X4Y137_A5Q;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_DMUX = CLBLL_L_X4Y137_SLICE_X4Y137_D5Q;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_A = CLBLL_L_X4Y137_SLICE_X5Y137_AO6;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_B = CLBLL_L_X4Y137_SLICE_X5Y137_BO6;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_C = CLBLL_L_X4Y137_SLICE_X5Y137_CO6;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_D = CLBLL_L_X4Y137_SLICE_X5Y137_DO6;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_AMUX = CLBLL_L_X4Y137_SLICE_X5Y137_AO5;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_A = CLBLL_L_X4Y138_SLICE_X4Y138_AO6;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_B = CLBLL_L_X4Y138_SLICE_X4Y138_BO6;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_C = CLBLL_L_X4Y138_SLICE_X4Y138_CO6;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_D = CLBLL_L_X4Y138_SLICE_X4Y138_DO6;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_A = CLBLL_L_X4Y138_SLICE_X5Y138_AO6;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_B = CLBLL_L_X4Y138_SLICE_X5Y138_BO6;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_C = CLBLL_L_X4Y138_SLICE_X5Y138_CO6;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_D = CLBLL_L_X4Y138_SLICE_X5Y138_DO6;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_AMUX = CLBLL_L_X4Y138_SLICE_X5Y138_A5Q;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_BMUX = CLBLL_L_X4Y138_SLICE_X5Y138_B5Q;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_CMUX = CLBLL_L_X4Y138_SLICE_X5Y138_CO5;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_DMUX = CLBLL_L_X4Y138_SLICE_X5Y138_DO5;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_A = CLBLL_L_X4Y139_SLICE_X4Y139_AO6;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_B = CLBLL_L_X4Y139_SLICE_X4Y139_BO6;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_C = CLBLL_L_X4Y139_SLICE_X4Y139_CO6;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_D = CLBLL_L_X4Y139_SLICE_X4Y139_DO6;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_A = CLBLL_L_X4Y139_SLICE_X5Y139_AO6;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_B = CLBLL_L_X4Y139_SLICE_X5Y139_BO6;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_C = CLBLL_L_X4Y139_SLICE_X5Y139_CO6;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_D = CLBLL_L_X4Y139_SLICE_X5Y139_DO6;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_A = CLBLL_L_X4Y140_SLICE_X4Y140_AO6;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_B = CLBLL_L_X4Y140_SLICE_X4Y140_BO6;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_C = CLBLL_L_X4Y140_SLICE_X4Y140_CO6;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_D = CLBLL_L_X4Y140_SLICE_X4Y140_DO6;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_CMUX = CLBLL_L_X4Y140_SLICE_X4Y140_CO6;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_A = CLBLL_L_X4Y140_SLICE_X5Y140_AO6;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_B = CLBLL_L_X4Y140_SLICE_X5Y140_BO6;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_C = CLBLL_L_X4Y140_SLICE_X5Y140_CO6;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_D = CLBLL_L_X4Y140_SLICE_X5Y140_DO6;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_DMUX = CLBLL_L_X4Y140_SLICE_X5Y140_DO6;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_A = CLBLL_L_X4Y141_SLICE_X4Y141_AO6;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_B = CLBLL_L_X4Y141_SLICE_X4Y141_BO6;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_C = CLBLL_L_X4Y141_SLICE_X4Y141_CO6;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_D = CLBLL_L_X4Y141_SLICE_X4Y141_DO6;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_A = CLBLL_L_X4Y141_SLICE_X5Y141_AO6;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_B = CLBLL_L_X4Y141_SLICE_X5Y141_BO6;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_C = CLBLL_L_X4Y141_SLICE_X5Y141_CO6;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_D = CLBLL_L_X4Y141_SLICE_X5Y141_DO6;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_A = CLBLL_L_X4Y142_SLICE_X4Y142_AO6;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_B = CLBLL_L_X4Y142_SLICE_X4Y142_BO6;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_C = CLBLL_L_X4Y142_SLICE_X4Y142_CO6;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_D = CLBLL_L_X4Y142_SLICE_X4Y142_DO6;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_A = CLBLL_L_X4Y142_SLICE_X5Y142_AO6;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_B = CLBLL_L_X4Y142_SLICE_X5Y142_BO6;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_C = CLBLL_L_X4Y142_SLICE_X5Y142_CO6;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_D = CLBLL_L_X4Y142_SLICE_X5Y142_DO6;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_A = CLBLL_L_X4Y143_SLICE_X4Y143_AO6;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_B = CLBLL_L_X4Y143_SLICE_X4Y143_BO6;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_C = CLBLL_L_X4Y143_SLICE_X4Y143_CO6;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_D = CLBLL_L_X4Y143_SLICE_X4Y143_DO6;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_AMUX = CLBLL_L_X4Y143_SLICE_X4Y143_AO5;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_BMUX = CLBLL_L_X4Y143_SLICE_X4Y143_BO5;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_A = CLBLL_L_X4Y143_SLICE_X5Y143_AO6;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_B = CLBLL_L_X4Y143_SLICE_X5Y143_BO6;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_C = CLBLL_L_X4Y143_SLICE_X5Y143_CO6;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_D = CLBLL_L_X4Y143_SLICE_X5Y143_DO6;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_AMUX = CLBLL_L_X4Y143_SLICE_X5Y143_AO5;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_BMUX = CLBLL_L_X4Y143_SLICE_X5Y143_BO5;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_CMUX = CLBLL_L_X4Y143_SLICE_X5Y143_CO5;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_A = CLBLL_L_X4Y144_SLICE_X4Y144_AO6;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_B = CLBLL_L_X4Y144_SLICE_X4Y144_BO6;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_C = CLBLL_L_X4Y144_SLICE_X4Y144_CO6;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_D = CLBLL_L_X4Y144_SLICE_X4Y144_DO6;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_A = CLBLL_L_X4Y144_SLICE_X5Y144_AO6;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_B = CLBLL_L_X4Y144_SLICE_X5Y144_BO6;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_C = CLBLL_L_X4Y144_SLICE_X5Y144_CO6;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_D = CLBLL_L_X4Y144_SLICE_X5Y144_DO6;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_A = CLBLL_L_X52Y126_SLICE_X78Y126_AO6;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_B = CLBLL_L_X52Y126_SLICE_X78Y126_BO6;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_C = CLBLL_L_X52Y126_SLICE_X78Y126_CO6;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_D = CLBLL_L_X52Y126_SLICE_X78Y126_DO6;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_A = CLBLL_L_X52Y126_SLICE_X79Y126_AO6;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_B = CLBLL_L_X52Y126_SLICE_X79Y126_BO6;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_C = CLBLL_L_X52Y126_SLICE_X79Y126_CO6;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_D = CLBLL_L_X52Y126_SLICE_X79Y126_DO6;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_A = CLBLM_L_X8Y131_SLICE_X10Y131_AO6;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_B = CLBLM_L_X8Y131_SLICE_X10Y131_BO6;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_C = CLBLM_L_X8Y131_SLICE_X10Y131_CO6;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_D = CLBLM_L_X8Y131_SLICE_X10Y131_DO6;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_AMUX = CLBLM_L_X8Y131_SLICE_X10Y131_A5Q;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_BMUX = CLBLM_L_X8Y131_SLICE_X10Y131_BO5;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_A = CLBLM_L_X8Y131_SLICE_X11Y131_AO6;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_B = CLBLM_L_X8Y131_SLICE_X11Y131_BO6;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_C = CLBLM_L_X8Y131_SLICE_X11Y131_CO6;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_D = CLBLM_L_X8Y131_SLICE_X11Y131_DO6;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_A = CLBLM_L_X8Y132_SLICE_X10Y132_AO6;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_B = CLBLM_L_X8Y132_SLICE_X10Y132_BO6;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_C = CLBLM_L_X8Y132_SLICE_X10Y132_CO6;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_D = CLBLM_L_X8Y132_SLICE_X10Y132_DO6;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_CMUX = CLBLM_L_X8Y132_SLICE_X10Y132_CO6;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_A = CLBLM_L_X8Y132_SLICE_X11Y132_AO6;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_B = CLBLM_L_X8Y132_SLICE_X11Y132_BO6;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_C = CLBLM_L_X8Y132_SLICE_X11Y132_CO6;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_D = CLBLM_L_X8Y132_SLICE_X11Y132_DO6;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_DMUX = CLBLM_L_X8Y132_SLICE_X11Y132_DO6;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_A = CLBLM_L_X8Y133_SLICE_X10Y133_AO6;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_B = CLBLM_L_X8Y133_SLICE_X10Y133_BO6;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_C = CLBLM_L_X8Y133_SLICE_X10Y133_CO6;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_D = CLBLM_L_X8Y133_SLICE_X10Y133_DO6;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_A = CLBLM_L_X8Y133_SLICE_X11Y133_AO6;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_B = CLBLM_L_X8Y133_SLICE_X11Y133_BO6;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_C = CLBLM_L_X8Y133_SLICE_X11Y133_CO6;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_D = CLBLM_L_X8Y133_SLICE_X11Y133_DO6;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_A = CLBLM_L_X8Y134_SLICE_X10Y134_AO6;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_B = CLBLM_L_X8Y134_SLICE_X10Y134_BO6;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_C = CLBLM_L_X8Y134_SLICE_X10Y134_CO6;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_D = CLBLM_L_X8Y134_SLICE_X10Y134_DO6;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_AMUX = CLBLM_L_X8Y134_SLICE_X10Y134_A5Q;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_BMUX = CLBLM_L_X8Y134_SLICE_X10Y134_BO5;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_A = CLBLM_L_X8Y134_SLICE_X11Y134_AO6;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_B = CLBLM_L_X8Y134_SLICE_X11Y134_BO6;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_C = CLBLM_L_X8Y134_SLICE_X11Y134_CO6;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_D = CLBLM_L_X8Y134_SLICE_X11Y134_DO6;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_A = CLBLM_L_X8Y135_SLICE_X10Y135_AO6;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_B = CLBLM_L_X8Y135_SLICE_X10Y135_BO6;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_C = CLBLM_L_X8Y135_SLICE_X10Y135_CO6;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_D = CLBLM_L_X8Y135_SLICE_X10Y135_DO6;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_AMUX = CLBLM_L_X8Y135_SLICE_X10Y135_A5Q;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_CMUX = CLBLM_L_X8Y135_SLICE_X10Y135_CO5;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_A = CLBLM_L_X8Y135_SLICE_X11Y135_AO6;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_B = CLBLM_L_X8Y135_SLICE_X11Y135_BO6;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_C = CLBLM_L_X8Y135_SLICE_X11Y135_CO6;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_D = CLBLM_L_X8Y135_SLICE_X11Y135_DO6;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_AMUX = CLBLM_L_X8Y135_SLICE_X11Y135_A5Q;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_BMUX = CLBLM_L_X8Y135_SLICE_X11Y135_B5Q;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_DMUX = CLBLM_L_X8Y135_SLICE_X11Y135_DO5;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_A = CLBLM_L_X8Y136_SLICE_X10Y136_AO6;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_B = CLBLM_L_X8Y136_SLICE_X10Y136_BO6;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_C = CLBLM_L_X8Y136_SLICE_X10Y136_CO6;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_D = CLBLM_L_X8Y136_SLICE_X10Y136_DO6;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_A = CLBLM_L_X8Y136_SLICE_X11Y136_AO6;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_B = CLBLM_L_X8Y136_SLICE_X11Y136_BO6;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_C = CLBLM_L_X8Y136_SLICE_X11Y136_CO6;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_D = CLBLM_L_X8Y136_SLICE_X11Y136_DO6;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_DMUX = CLBLM_L_X8Y136_SLICE_X11Y136_DO5;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_A = CLBLM_L_X8Y137_SLICE_X10Y137_AO6;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_B = CLBLM_L_X8Y137_SLICE_X10Y137_BO6;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_C = CLBLM_L_X8Y137_SLICE_X10Y137_CO6;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_D = CLBLM_L_X8Y137_SLICE_X10Y137_DO6;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_BMUX = CLBLM_L_X8Y137_SLICE_X10Y137_BO5;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_A = CLBLM_L_X8Y137_SLICE_X11Y137_AO6;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_B = CLBLM_L_X8Y137_SLICE_X11Y137_BO6;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_C = CLBLM_L_X8Y137_SLICE_X11Y137_CO6;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_D = CLBLM_L_X8Y137_SLICE_X11Y137_DO6;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_CMUX = CLBLM_L_X8Y137_SLICE_X11Y137_CO5;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_A = CLBLM_L_X8Y138_SLICE_X10Y138_AO6;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_B = CLBLM_L_X8Y138_SLICE_X10Y138_BO6;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_C = CLBLM_L_X8Y138_SLICE_X10Y138_CO6;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_D = CLBLM_L_X8Y138_SLICE_X10Y138_DO6;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_DMUX = CLBLM_L_X8Y138_SLICE_X10Y138_D5Q;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_A = CLBLM_L_X8Y138_SLICE_X11Y138_AO6;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_B = CLBLM_L_X8Y138_SLICE_X11Y138_BO6;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_C = CLBLM_L_X8Y138_SLICE_X11Y138_CO6;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_D = CLBLM_L_X8Y138_SLICE_X11Y138_DO6;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_CMUX = CLBLM_L_X8Y138_SLICE_X11Y138_CO5;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_A = CLBLM_L_X8Y139_SLICE_X10Y139_AO6;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_B = CLBLM_L_X8Y139_SLICE_X10Y139_BO6;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_C = CLBLM_L_X8Y139_SLICE_X10Y139_CO6;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_D = CLBLM_L_X8Y139_SLICE_X10Y139_DO6;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_A = CLBLM_L_X8Y139_SLICE_X11Y139_AO6;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_B = CLBLM_L_X8Y139_SLICE_X11Y139_BO6;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_C = CLBLM_L_X8Y139_SLICE_X11Y139_CO6;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_D = CLBLM_L_X8Y139_SLICE_X11Y139_DO6;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_CMUX = CLBLM_L_X8Y139_SLICE_X11Y139_CO6;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_A = CLBLM_L_X8Y140_SLICE_X10Y140_AO6;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_B = CLBLM_L_X8Y140_SLICE_X10Y140_BO6;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_C = CLBLM_L_X8Y140_SLICE_X10Y140_CO6;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_D = CLBLM_L_X8Y140_SLICE_X10Y140_DO6;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_AMUX = CLBLM_L_X8Y140_SLICE_X10Y140_A5Q;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_A = CLBLM_L_X8Y140_SLICE_X11Y140_AO6;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_B = CLBLM_L_X8Y140_SLICE_X11Y140_BO6;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_C = CLBLM_L_X8Y140_SLICE_X11Y140_CO6;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_D = CLBLM_L_X8Y140_SLICE_X11Y140_DO6;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_AMUX = CLBLM_L_X8Y140_SLICE_X11Y140_A5Q;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_CMUX = CLBLM_L_X8Y140_SLICE_X11Y140_CO5;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_A = CLBLM_L_X8Y141_SLICE_X10Y141_AO6;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_B = CLBLM_L_X8Y141_SLICE_X10Y141_BO6;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_C = CLBLM_L_X8Y141_SLICE_X10Y141_CO6;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_D = CLBLM_L_X8Y141_SLICE_X10Y141_DO6;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_A = CLBLM_L_X8Y141_SLICE_X11Y141_AO6;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_B = CLBLM_L_X8Y141_SLICE_X11Y141_BO6;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_C = CLBLM_L_X8Y141_SLICE_X11Y141_CO6;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_D = CLBLM_L_X8Y141_SLICE_X11Y141_DO6;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_DMUX = CLBLM_L_X8Y141_SLICE_X11Y141_DO5;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_A = CLBLM_L_X8Y142_SLICE_X10Y142_AO6;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_B = CLBLM_L_X8Y142_SLICE_X10Y142_BO6;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_C = CLBLM_L_X8Y142_SLICE_X10Y142_CO6;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_D = CLBLM_L_X8Y142_SLICE_X10Y142_DO6;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_DMUX = CLBLM_L_X8Y142_SLICE_X10Y142_D5Q;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_A = CLBLM_L_X8Y142_SLICE_X11Y142_AO6;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_B = CLBLM_L_X8Y142_SLICE_X11Y142_BO6;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_C = CLBLM_L_X8Y142_SLICE_X11Y142_CO6;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_D = CLBLM_L_X8Y142_SLICE_X11Y142_DO6;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_A = CLBLM_L_X8Y143_SLICE_X10Y143_AO6;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_B = CLBLM_L_X8Y143_SLICE_X10Y143_BO6;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_C = CLBLM_L_X8Y143_SLICE_X10Y143_CO6;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_D = CLBLM_L_X8Y143_SLICE_X10Y143_DO6;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_DMUX = CLBLM_L_X8Y143_SLICE_X10Y143_DO5;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_A = CLBLM_L_X8Y143_SLICE_X11Y143_AO6;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_B = CLBLM_L_X8Y143_SLICE_X11Y143_BO6;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_C = CLBLM_L_X8Y143_SLICE_X11Y143_CO6;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_D = CLBLM_L_X8Y143_SLICE_X11Y143_DO6;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_A = CLBLM_L_X8Y144_SLICE_X10Y144_AO6;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_B = CLBLM_L_X8Y144_SLICE_X10Y144_BO6;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_C = CLBLM_L_X8Y144_SLICE_X10Y144_CO6;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_D = CLBLM_L_X8Y144_SLICE_X10Y144_DO6;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_A = CLBLM_L_X8Y144_SLICE_X11Y144_AO6;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_B = CLBLM_L_X8Y144_SLICE_X11Y144_BO6;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_C = CLBLM_L_X8Y144_SLICE_X11Y144_CO6;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_D = CLBLM_L_X8Y144_SLICE_X11Y144_DO6;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_BMUX = CLBLM_L_X8Y144_SLICE_X11Y144_BO5;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_A = CLBLM_L_X10Y130_SLICE_X12Y130_AO6;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_B = CLBLM_L_X10Y130_SLICE_X12Y130_BO6;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_C = CLBLM_L_X10Y130_SLICE_X12Y130_CO6;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_D = CLBLM_L_X10Y130_SLICE_X12Y130_DO6;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_BMUX = CLBLM_L_X10Y130_SLICE_X12Y130_BO5;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_A = CLBLM_L_X10Y130_SLICE_X13Y130_AO6;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_B = CLBLM_L_X10Y130_SLICE_X13Y130_BO6;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_C = CLBLM_L_X10Y130_SLICE_X13Y130_CO6;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_D = CLBLM_L_X10Y130_SLICE_X13Y130_DO6;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_AMUX = CLBLM_L_X10Y130_SLICE_X13Y130_AO5;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_A = CLBLM_L_X10Y131_SLICE_X12Y131_AO6;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_B = CLBLM_L_X10Y131_SLICE_X12Y131_BO6;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_C = CLBLM_L_X10Y131_SLICE_X12Y131_CO6;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_D = CLBLM_L_X10Y131_SLICE_X12Y131_DO6;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_AMUX = CLBLM_L_X10Y131_SLICE_X12Y131_AO5;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_CMUX = CLBLM_L_X10Y131_SLICE_X12Y131_CO5;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_A = CLBLM_L_X10Y131_SLICE_X13Y131_AO6;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_B = CLBLM_L_X10Y131_SLICE_X13Y131_BO6;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_C = CLBLM_L_X10Y131_SLICE_X13Y131_CO6;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_D = CLBLM_L_X10Y131_SLICE_X13Y131_DO6;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_A = CLBLM_L_X10Y132_SLICE_X12Y132_AO6;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_B = CLBLM_L_X10Y132_SLICE_X12Y132_BO6;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_C = CLBLM_L_X10Y132_SLICE_X12Y132_CO6;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_D = CLBLM_L_X10Y132_SLICE_X12Y132_DO6;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_CMUX = CLBLM_L_X10Y132_SLICE_X12Y132_CO6;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_A = CLBLM_L_X10Y132_SLICE_X13Y132_AO6;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_B = CLBLM_L_X10Y132_SLICE_X13Y132_BO6;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_C = CLBLM_L_X10Y132_SLICE_X13Y132_CO6;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_D = CLBLM_L_X10Y132_SLICE_X13Y132_DO6;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_A = CLBLM_L_X10Y133_SLICE_X12Y133_AO6;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_B = CLBLM_L_X10Y133_SLICE_X12Y133_BO6;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_C = CLBLM_L_X10Y133_SLICE_X12Y133_CO6;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_D = CLBLM_L_X10Y133_SLICE_X12Y133_DO6;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_DMUX = CLBLM_L_X10Y133_SLICE_X12Y133_DO5;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_A = CLBLM_L_X10Y133_SLICE_X13Y133_AO6;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_B = CLBLM_L_X10Y133_SLICE_X13Y133_BO6;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_C = CLBLM_L_X10Y133_SLICE_X13Y133_CO6;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_D = CLBLM_L_X10Y133_SLICE_X13Y133_DO6;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_A = CLBLM_L_X10Y134_SLICE_X12Y134_AO6;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_B = CLBLM_L_X10Y134_SLICE_X12Y134_BO6;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_C = CLBLM_L_X10Y134_SLICE_X12Y134_CO6;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_D = CLBLM_L_X10Y134_SLICE_X12Y134_DO6;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_A = CLBLM_L_X10Y134_SLICE_X13Y134_AO6;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_B = CLBLM_L_X10Y134_SLICE_X13Y134_BO6;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_C = CLBLM_L_X10Y134_SLICE_X13Y134_CO6;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_D = CLBLM_L_X10Y134_SLICE_X13Y134_DO6;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_AMUX = CLBLM_L_X10Y134_SLICE_X13Y134_A5Q;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_BMUX = CLBLM_L_X10Y134_SLICE_X13Y134_B5Q;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_CMUX = CLBLM_L_X10Y134_SLICE_X13Y134_CO5;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_A = CLBLM_L_X10Y135_SLICE_X12Y135_AO6;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_B = CLBLM_L_X10Y135_SLICE_X12Y135_BO6;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_C = CLBLM_L_X10Y135_SLICE_X12Y135_CO6;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_D = CLBLM_L_X10Y135_SLICE_X12Y135_DO6;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_BMUX = CLBLM_L_X10Y135_SLICE_X12Y135_B5Q;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_A = CLBLM_L_X10Y135_SLICE_X13Y135_AO6;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_B = CLBLM_L_X10Y135_SLICE_X13Y135_BO6;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_C = CLBLM_L_X10Y135_SLICE_X13Y135_CO6;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_D = CLBLM_L_X10Y135_SLICE_X13Y135_DO6;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_AMUX = CLBLM_L_X10Y135_SLICE_X13Y135_AO5;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_BMUX = CLBLM_L_X10Y135_SLICE_X13Y135_B5Q;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_A = CLBLM_L_X10Y136_SLICE_X12Y136_AO6;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_B = CLBLM_L_X10Y136_SLICE_X12Y136_BO6;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_C = CLBLM_L_X10Y136_SLICE_X12Y136_CO6;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_D = CLBLM_L_X10Y136_SLICE_X12Y136_DO6;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_AMUX = CLBLM_L_X10Y136_SLICE_X12Y136_A5Q;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_CMUX = CLBLM_L_X10Y136_SLICE_X12Y136_CO5;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_A = CLBLM_L_X10Y136_SLICE_X13Y136_AO6;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_B = CLBLM_L_X10Y136_SLICE_X13Y136_BO6;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_C = CLBLM_L_X10Y136_SLICE_X13Y136_CO6;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_D = CLBLM_L_X10Y136_SLICE_X13Y136_DO6;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_A = CLBLM_L_X10Y137_SLICE_X12Y137_AO6;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_B = CLBLM_L_X10Y137_SLICE_X12Y137_BO6;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_C = CLBLM_L_X10Y137_SLICE_X12Y137_CO6;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_D = CLBLM_L_X10Y137_SLICE_X12Y137_DO6;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_BMUX = CLBLM_L_X10Y137_SLICE_X12Y137_B5Q;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_A = CLBLM_L_X10Y137_SLICE_X13Y137_AO6;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_B = CLBLM_L_X10Y137_SLICE_X13Y137_BO6;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_C = CLBLM_L_X10Y137_SLICE_X13Y137_CO6;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_D = CLBLM_L_X10Y137_SLICE_X13Y137_DO6;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_A = CLBLM_L_X10Y138_SLICE_X12Y138_AO6;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_B = CLBLM_L_X10Y138_SLICE_X12Y138_BO6;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_C = CLBLM_L_X10Y138_SLICE_X12Y138_CO6;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_D = CLBLM_L_X10Y138_SLICE_X12Y138_DO6;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_AMUX = CLBLM_L_X10Y138_SLICE_X12Y138_A5Q;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_BMUX = CLBLM_L_X10Y138_SLICE_X12Y138_BO5;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_A = CLBLM_L_X10Y138_SLICE_X13Y138_AO6;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_B = CLBLM_L_X10Y138_SLICE_X13Y138_BO6;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_C = CLBLM_L_X10Y138_SLICE_X13Y138_CO6;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_D = CLBLM_L_X10Y138_SLICE_X13Y138_DO6;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_A = CLBLM_L_X10Y139_SLICE_X12Y139_AO6;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_B = CLBLM_L_X10Y139_SLICE_X12Y139_BO6;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_C = CLBLM_L_X10Y139_SLICE_X12Y139_CO6;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_D = CLBLM_L_X10Y139_SLICE_X12Y139_DO6;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_A = CLBLM_L_X10Y139_SLICE_X13Y139_AO6;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_B = CLBLM_L_X10Y139_SLICE_X13Y139_BO6;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_C = CLBLM_L_X10Y139_SLICE_X13Y139_CO6;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_D = CLBLM_L_X10Y139_SLICE_X13Y139_DO6;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_BMUX = CLBLM_L_X10Y139_SLICE_X13Y139_B5Q;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_A = CLBLM_L_X10Y140_SLICE_X12Y140_AO6;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_B = CLBLM_L_X10Y140_SLICE_X12Y140_BO6;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_C = CLBLM_L_X10Y140_SLICE_X12Y140_CO6;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_D = CLBLM_L_X10Y140_SLICE_X12Y140_DO6;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_AMUX = CLBLM_L_X10Y140_SLICE_X12Y140_A5Q;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_BMUX = CLBLM_L_X10Y140_SLICE_X12Y140_BO5;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_A = CLBLM_L_X10Y140_SLICE_X13Y140_AO6;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_B = CLBLM_L_X10Y140_SLICE_X13Y140_BO6;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_C = CLBLM_L_X10Y140_SLICE_X13Y140_CO6;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_D = CLBLM_L_X10Y140_SLICE_X13Y140_DO6;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_AMUX = CLBLM_L_X10Y140_SLICE_X13Y140_AO5;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_CMUX = CLBLM_L_X10Y140_SLICE_X13Y140_C5Q;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_A = CLBLM_L_X10Y141_SLICE_X12Y141_AO6;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_B = CLBLM_L_X10Y141_SLICE_X12Y141_BO6;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_C = CLBLM_L_X10Y141_SLICE_X12Y141_CO6;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_D = CLBLM_L_X10Y141_SLICE_X12Y141_DO6;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_BMUX = CLBLM_L_X10Y141_SLICE_X12Y141_BO5;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_CMUX = CLBLM_L_X10Y141_SLICE_X12Y141_C5Q;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_A = CLBLM_L_X10Y141_SLICE_X13Y141_AO6;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_B = CLBLM_L_X10Y141_SLICE_X13Y141_BO6;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_C = CLBLM_L_X10Y141_SLICE_X13Y141_CO6;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_D = CLBLM_L_X10Y141_SLICE_X13Y141_DO6;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_AMUX = CLBLM_L_X10Y141_SLICE_X13Y141_A5Q;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_A = CLBLM_L_X10Y142_SLICE_X12Y142_AO6;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_B = CLBLM_L_X10Y142_SLICE_X12Y142_BO6;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_C = CLBLM_L_X10Y142_SLICE_X12Y142_CO6;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_D = CLBLM_L_X10Y142_SLICE_X12Y142_DO6;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_A = CLBLM_L_X10Y142_SLICE_X13Y142_AO6;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_B = CLBLM_L_X10Y142_SLICE_X13Y142_BO6;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_C = CLBLM_L_X10Y142_SLICE_X13Y142_CO6;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_D = CLBLM_L_X10Y142_SLICE_X13Y142_DO6;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_A = CLBLM_L_X10Y143_SLICE_X12Y143_AO6;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_B = CLBLM_L_X10Y143_SLICE_X12Y143_BO6;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_C = CLBLM_L_X10Y143_SLICE_X12Y143_CO6;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_D = CLBLM_L_X10Y143_SLICE_X12Y143_DO6;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_A = CLBLM_L_X10Y143_SLICE_X13Y143_AO6;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_B = CLBLM_L_X10Y143_SLICE_X13Y143_BO6;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_C = CLBLM_L_X10Y143_SLICE_X13Y143_CO6;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_D = CLBLM_L_X10Y143_SLICE_X13Y143_DO6;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_BMUX = CLBLM_L_X10Y143_SLICE_X13Y143_BO6;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_A = CLBLM_L_X10Y144_SLICE_X12Y144_AO6;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_B = CLBLM_L_X10Y144_SLICE_X12Y144_BO6;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_C = CLBLM_L_X10Y144_SLICE_X12Y144_CO6;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_D = CLBLM_L_X10Y144_SLICE_X12Y144_DO6;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_AMUX = CLBLM_L_X10Y144_SLICE_X12Y144_AO5;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_A = CLBLM_L_X10Y144_SLICE_X13Y144_AO6;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_B = CLBLM_L_X10Y144_SLICE_X13Y144_BO6;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_C = CLBLM_L_X10Y144_SLICE_X13Y144_CO6;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_D = CLBLM_L_X10Y144_SLICE_X13Y144_DO6;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_A = CLBLM_L_X10Y145_SLICE_X12Y145_AO6;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_B = CLBLM_L_X10Y145_SLICE_X12Y145_BO6;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_C = CLBLM_L_X10Y145_SLICE_X12Y145_CO6;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_D = CLBLM_L_X10Y145_SLICE_X12Y145_DO6;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_AMUX = CLBLM_L_X10Y145_SLICE_X12Y145_AO5;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_BMUX = CLBLM_L_X10Y145_SLICE_X12Y145_BO5;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_A = CLBLM_L_X10Y145_SLICE_X13Y145_AO6;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_B = CLBLM_L_X10Y145_SLICE_X13Y145_BO6;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_C = CLBLM_L_X10Y145_SLICE_X13Y145_CO6;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_D = CLBLM_L_X10Y145_SLICE_X13Y145_DO6;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_BMUX = CLBLM_L_X10Y145_SLICE_X13Y145_BO5;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_A = CLBLM_L_X10Y146_SLICE_X12Y146_AO6;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_B = CLBLM_L_X10Y146_SLICE_X12Y146_BO6;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_C = CLBLM_L_X10Y146_SLICE_X12Y146_CO6;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_D = CLBLM_L_X10Y146_SLICE_X12Y146_DO6;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_AMUX = CLBLM_L_X10Y146_SLICE_X12Y146_AO5;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_A = CLBLM_L_X10Y146_SLICE_X13Y146_AO6;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_B = CLBLM_L_X10Y146_SLICE_X13Y146_BO6;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_C = CLBLM_L_X10Y146_SLICE_X13Y146_CO6;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_D = CLBLM_L_X10Y146_SLICE_X13Y146_DO6;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_A = CLBLM_L_X12Y132_SLICE_X16Y132_AO6;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_B = CLBLM_L_X12Y132_SLICE_X16Y132_BO6;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_C = CLBLM_L_X12Y132_SLICE_X16Y132_CO6;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_D = CLBLM_L_X12Y132_SLICE_X16Y132_DO6;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_DMUX = CLBLM_L_X12Y132_SLICE_X16Y132_DO6;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_A = CLBLM_L_X12Y132_SLICE_X17Y132_AO6;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_B = CLBLM_L_X12Y132_SLICE_X17Y132_BO6;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_C = CLBLM_L_X12Y132_SLICE_X17Y132_CO6;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_D = CLBLM_L_X12Y132_SLICE_X17Y132_DO6;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_A = CLBLM_L_X12Y133_SLICE_X16Y133_AO6;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_B = CLBLM_L_X12Y133_SLICE_X16Y133_BO6;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_C = CLBLM_L_X12Y133_SLICE_X16Y133_CO6;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_D = CLBLM_L_X12Y133_SLICE_X16Y133_DO6;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_CMUX = CLBLM_L_X12Y133_SLICE_X16Y133_C5Q;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_DMUX = CLBLM_L_X12Y133_SLICE_X16Y133_DO5;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_A = CLBLM_L_X12Y133_SLICE_X17Y133_AO6;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_B = CLBLM_L_X12Y133_SLICE_X17Y133_BO6;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_C = CLBLM_L_X12Y133_SLICE_X17Y133_CO6;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_D = CLBLM_L_X12Y133_SLICE_X17Y133_DO6;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_A = CLBLM_L_X12Y134_SLICE_X16Y134_AO6;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_B = CLBLM_L_X12Y134_SLICE_X16Y134_BO6;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_C = CLBLM_L_X12Y134_SLICE_X16Y134_CO6;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_D = CLBLM_L_X12Y134_SLICE_X16Y134_DO6;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_A = CLBLM_L_X12Y134_SLICE_X17Y134_AO6;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_B = CLBLM_L_X12Y134_SLICE_X17Y134_BO6;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_C = CLBLM_L_X12Y134_SLICE_X17Y134_CO6;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_D = CLBLM_L_X12Y134_SLICE_X17Y134_DO6;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_DMUX = CLBLM_L_X12Y134_SLICE_X17Y134_DO6;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_A = CLBLM_L_X12Y135_SLICE_X16Y135_AO6;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_B = CLBLM_L_X12Y135_SLICE_X16Y135_BO6;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_C = CLBLM_L_X12Y135_SLICE_X16Y135_CO6;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_D = CLBLM_L_X12Y135_SLICE_X16Y135_DO6;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_A = CLBLM_L_X12Y135_SLICE_X17Y135_AO6;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_B = CLBLM_L_X12Y135_SLICE_X17Y135_BO6;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_C = CLBLM_L_X12Y135_SLICE_X17Y135_CO6;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_D = CLBLM_L_X12Y135_SLICE_X17Y135_DO6;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_AMUX = CLBLM_L_X12Y135_SLICE_X17Y135_A5Q;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_BMUX = CLBLM_L_X12Y135_SLICE_X17Y135_BO5;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_A = CLBLM_L_X12Y136_SLICE_X16Y136_AO6;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_B = CLBLM_L_X12Y136_SLICE_X16Y136_BO6;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_C = CLBLM_L_X12Y136_SLICE_X16Y136_CO6;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_D = CLBLM_L_X12Y136_SLICE_X16Y136_DO6;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_BMUX = CLBLM_L_X12Y136_SLICE_X16Y136_B5Q;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_CMUX = CLBLM_L_X12Y136_SLICE_X16Y136_C5Q;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_A = CLBLM_L_X12Y136_SLICE_X17Y136_AO6;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_B = CLBLM_L_X12Y136_SLICE_X17Y136_BO6;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_C = CLBLM_L_X12Y136_SLICE_X17Y136_CO6;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_D = CLBLM_L_X12Y136_SLICE_X17Y136_DO6;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_AMUX = CLBLM_L_X12Y136_SLICE_X17Y136_A5Q;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_BMUX = CLBLM_L_X12Y136_SLICE_X17Y136_BO5;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_A = CLBLM_L_X12Y137_SLICE_X16Y137_AO6;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_B = CLBLM_L_X12Y137_SLICE_X16Y137_BO6;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_C = CLBLM_L_X12Y137_SLICE_X16Y137_CO6;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_D = CLBLM_L_X12Y137_SLICE_X16Y137_DO6;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_AMUX = CLBLM_L_X12Y137_SLICE_X16Y137_A5Q;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_BMUX = CLBLM_L_X12Y137_SLICE_X16Y137_BO5;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_A = CLBLM_L_X12Y137_SLICE_X17Y137_AO6;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_B = CLBLM_L_X12Y137_SLICE_X17Y137_BO6;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_C = CLBLM_L_X12Y137_SLICE_X17Y137_CO6;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_D = CLBLM_L_X12Y137_SLICE_X17Y137_DO6;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_AMUX = CLBLM_L_X12Y137_SLICE_X17Y137_A5Q;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_BMUX = CLBLM_L_X12Y137_SLICE_X17Y137_BO5;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_A = CLBLM_L_X12Y138_SLICE_X16Y138_AO6;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_B = CLBLM_L_X12Y138_SLICE_X16Y138_BO6;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_C = CLBLM_L_X12Y138_SLICE_X16Y138_CO6;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_D = CLBLM_L_X12Y138_SLICE_X16Y138_DO6;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_A = CLBLM_L_X12Y138_SLICE_X17Y138_AO6;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_B = CLBLM_L_X12Y138_SLICE_X17Y138_BO6;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_C = CLBLM_L_X12Y138_SLICE_X17Y138_CO6;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_D = CLBLM_L_X12Y138_SLICE_X17Y138_DO6;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_AMUX = CLBLM_L_X12Y138_SLICE_X17Y138_A5Q;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_BMUX = CLBLM_L_X12Y138_SLICE_X17Y138_BO5;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_CMUX = CLBLM_L_X12Y138_SLICE_X17Y138_CO5;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_DMUX = CLBLM_L_X12Y138_SLICE_X17Y138_DO5;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_A = CLBLM_L_X12Y139_SLICE_X16Y139_AO6;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_B = CLBLM_L_X12Y139_SLICE_X16Y139_BO6;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_C = CLBLM_L_X12Y139_SLICE_X16Y139_CO6;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_D = CLBLM_L_X12Y139_SLICE_X16Y139_DO6;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_AMUX = CLBLM_L_X12Y139_SLICE_X16Y139_A5Q;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_BMUX = CLBLM_L_X12Y139_SLICE_X16Y139_BO5;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_DMUX = CLBLM_L_X12Y139_SLICE_X16Y139_DO5;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_A = CLBLM_L_X12Y139_SLICE_X17Y139_AO6;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_B = CLBLM_L_X12Y139_SLICE_X17Y139_BO6;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_C = CLBLM_L_X12Y139_SLICE_X17Y139_CO6;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_D = CLBLM_L_X12Y139_SLICE_X17Y139_DO6;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_BMUX = CLBLM_L_X12Y139_SLICE_X17Y139_BO5;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_DMUX = CLBLM_L_X12Y139_SLICE_X17Y139_DO5;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_A = CLBLM_L_X12Y140_SLICE_X16Y140_AO6;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_B = CLBLM_L_X12Y140_SLICE_X16Y140_BO6;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_C = CLBLM_L_X12Y140_SLICE_X16Y140_CO6;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_D = CLBLM_L_X12Y140_SLICE_X16Y140_DO6;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_A = CLBLM_L_X12Y140_SLICE_X17Y140_AO6;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_B = CLBLM_L_X12Y140_SLICE_X17Y140_BO6;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_C = CLBLM_L_X12Y140_SLICE_X17Y140_CO6;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_D = CLBLM_L_X12Y140_SLICE_X17Y140_DO6;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_A = CLBLM_L_X12Y141_SLICE_X16Y141_AO6;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_B = CLBLM_L_X12Y141_SLICE_X16Y141_BO6;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_C = CLBLM_L_X12Y141_SLICE_X16Y141_CO6;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_D = CLBLM_L_X12Y141_SLICE_X16Y141_DO6;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_A = CLBLM_L_X12Y141_SLICE_X17Y141_AO6;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_B = CLBLM_L_X12Y141_SLICE_X17Y141_BO6;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_C = CLBLM_L_X12Y141_SLICE_X17Y141_CO6;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_D = CLBLM_L_X12Y141_SLICE_X17Y141_DO6;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_BMUX = CLBLM_L_X12Y141_SLICE_X17Y141_BO5;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_DMUX = CLBLM_L_X12Y141_SLICE_X17Y141_DO6;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_A = CLBLM_L_X12Y142_SLICE_X16Y142_AO6;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_B = CLBLM_L_X12Y142_SLICE_X16Y142_BO6;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_C = CLBLM_L_X12Y142_SLICE_X16Y142_CO6;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_D = CLBLM_L_X12Y142_SLICE_X16Y142_DO6;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_AMUX = CLBLM_L_X12Y142_SLICE_X16Y142_A5Q;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_A = CLBLM_L_X12Y142_SLICE_X17Y142_AO6;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_B = CLBLM_L_X12Y142_SLICE_X17Y142_BO6;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_C = CLBLM_L_X12Y142_SLICE_X17Y142_CO6;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_D = CLBLM_L_X12Y142_SLICE_X17Y142_DO6;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_CMUX = CLBLM_L_X12Y142_SLICE_X17Y142_CO5;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_DMUX = CLBLM_L_X12Y142_SLICE_X17Y142_DO6;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_A = CLBLM_L_X12Y143_SLICE_X16Y143_AO6;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_B = CLBLM_L_X12Y143_SLICE_X16Y143_BO6;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_C = CLBLM_L_X12Y143_SLICE_X16Y143_CO6;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_D = CLBLM_L_X12Y143_SLICE_X16Y143_DO6;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_A = CLBLM_L_X12Y143_SLICE_X17Y143_AO6;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_B = CLBLM_L_X12Y143_SLICE_X17Y143_BO6;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_C = CLBLM_L_X12Y143_SLICE_X17Y143_CO6;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_D = CLBLM_L_X12Y143_SLICE_X17Y143_DO6;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_CMUX = CLBLM_L_X12Y143_SLICE_X17Y143_CO5;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_A = CLBLM_L_X12Y144_SLICE_X16Y144_AO6;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_B = CLBLM_L_X12Y144_SLICE_X16Y144_BO6;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_C = CLBLM_L_X12Y144_SLICE_X16Y144_CO6;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_D = CLBLM_L_X12Y144_SLICE_X16Y144_DO6;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_A = CLBLM_L_X12Y144_SLICE_X17Y144_AO6;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_B = CLBLM_L_X12Y144_SLICE_X17Y144_BO6;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_C = CLBLM_L_X12Y144_SLICE_X17Y144_CO6;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_D = CLBLM_L_X12Y144_SLICE_X17Y144_DO6;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_AMUX = CLBLM_L_X12Y144_SLICE_X17Y144_AO5;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_A = CLBLM_L_X12Y146_SLICE_X16Y146_AO6;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_B = CLBLM_L_X12Y146_SLICE_X16Y146_BO6;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_C = CLBLM_L_X12Y146_SLICE_X16Y146_CO6;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_D = CLBLM_L_X12Y146_SLICE_X16Y146_DO6;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_AMUX = CLBLM_L_X12Y146_SLICE_X16Y146_AO5;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_A = CLBLM_L_X12Y146_SLICE_X17Y146_AO6;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_B = CLBLM_L_X12Y146_SLICE_X17Y146_BO6;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_C = CLBLM_L_X12Y146_SLICE_X17Y146_CO6;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_D = CLBLM_L_X12Y146_SLICE_X17Y146_DO6;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_A = CLBLM_R_X3Y133_SLICE_X2Y133_AO6;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_B = CLBLM_R_X3Y133_SLICE_X2Y133_BO6;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_C = CLBLM_R_X3Y133_SLICE_X2Y133_CO6;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_D = CLBLM_R_X3Y133_SLICE_X2Y133_DO6;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_AMUX = CLBLM_R_X3Y133_SLICE_X2Y133_AO5;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_CMUX = CLBLM_R_X3Y133_SLICE_X2Y133_CO6;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_A = CLBLM_R_X3Y133_SLICE_X3Y133_AO6;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_B = CLBLM_R_X3Y133_SLICE_X3Y133_BO6;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_C = CLBLM_R_X3Y133_SLICE_X3Y133_CO6;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_D = CLBLM_R_X3Y133_SLICE_X3Y133_DO6;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_A = CLBLM_R_X3Y135_SLICE_X2Y135_AO6;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_B = CLBLM_R_X3Y135_SLICE_X2Y135_BO6;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_C = CLBLM_R_X3Y135_SLICE_X2Y135_CO6;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_D = CLBLM_R_X3Y135_SLICE_X2Y135_DO6;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_A = CLBLM_R_X3Y135_SLICE_X3Y135_AO6;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_B = CLBLM_R_X3Y135_SLICE_X3Y135_BO6;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_C = CLBLM_R_X3Y135_SLICE_X3Y135_CO6;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_D = CLBLM_R_X3Y135_SLICE_X3Y135_DO6;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_CMUX = CLBLM_R_X3Y135_SLICE_X3Y135_CO6;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_A = CLBLM_R_X3Y136_SLICE_X2Y136_AO6;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_B = CLBLM_R_X3Y136_SLICE_X2Y136_BO6;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_C = CLBLM_R_X3Y136_SLICE_X2Y136_CO6;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_D = CLBLM_R_X3Y136_SLICE_X2Y136_DO6;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_BMUX = CLBLM_R_X3Y136_SLICE_X2Y136_BO5;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_A = CLBLM_R_X3Y136_SLICE_X3Y136_AO6;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_B = CLBLM_R_X3Y136_SLICE_X3Y136_BO6;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_C = CLBLM_R_X3Y136_SLICE_X3Y136_CO6;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_D = CLBLM_R_X3Y136_SLICE_X3Y136_DO6;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_A = CLBLM_R_X3Y137_SLICE_X2Y137_AO6;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_B = CLBLM_R_X3Y137_SLICE_X2Y137_BO6;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_C = CLBLM_R_X3Y137_SLICE_X2Y137_CO6;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_D = CLBLM_R_X3Y137_SLICE_X2Y137_DO6;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_A = CLBLM_R_X3Y137_SLICE_X3Y137_AO6;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_B = CLBLM_R_X3Y137_SLICE_X3Y137_BO6;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_C = CLBLM_R_X3Y137_SLICE_X3Y137_CO6;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_D = CLBLM_R_X3Y137_SLICE_X3Y137_DO6;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_AMUX = CLBLM_R_X3Y137_SLICE_X3Y137_AO5;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_BMUX = CLBLM_R_X3Y137_SLICE_X3Y137_BO5;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_A = CLBLM_R_X3Y138_SLICE_X2Y138_AO6;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_B = CLBLM_R_X3Y138_SLICE_X2Y138_BO6;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_C = CLBLM_R_X3Y138_SLICE_X2Y138_CO6;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_D = CLBLM_R_X3Y138_SLICE_X2Y138_DO6;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_AMUX = CLBLM_R_X3Y138_SLICE_X2Y138_AO5;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_A = CLBLM_R_X3Y138_SLICE_X3Y138_AO6;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_B = CLBLM_R_X3Y138_SLICE_X3Y138_BO6;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_C = CLBLM_R_X3Y138_SLICE_X3Y138_CO6;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_D = CLBLM_R_X3Y138_SLICE_X3Y138_DO6;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_A = CLBLM_R_X3Y139_SLICE_X2Y139_AO6;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_B = CLBLM_R_X3Y139_SLICE_X2Y139_BO6;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_C = CLBLM_R_X3Y139_SLICE_X2Y139_CO6;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_D = CLBLM_R_X3Y139_SLICE_X2Y139_DO6;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_AMUX = CLBLM_R_X3Y139_SLICE_X2Y139_AO5;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_A = CLBLM_R_X3Y139_SLICE_X3Y139_AO6;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_B = CLBLM_R_X3Y139_SLICE_X3Y139_BO6;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_C = CLBLM_R_X3Y139_SLICE_X3Y139_CO6;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_D = CLBLM_R_X3Y139_SLICE_X3Y139_DO6;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_A = CLBLM_R_X3Y140_SLICE_X2Y140_AO6;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_B = CLBLM_R_X3Y140_SLICE_X2Y140_BO6;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_C = CLBLM_R_X3Y140_SLICE_X2Y140_CO6;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_D = CLBLM_R_X3Y140_SLICE_X2Y140_DO6;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_A = CLBLM_R_X3Y140_SLICE_X3Y140_AO6;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_B = CLBLM_R_X3Y140_SLICE_X3Y140_BO6;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_C = CLBLM_R_X3Y140_SLICE_X3Y140_CO6;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_D = CLBLM_R_X3Y140_SLICE_X3Y140_DO6;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_CMUX = CLBLM_R_X3Y140_SLICE_X3Y140_CO6;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_A = CLBLM_R_X3Y141_SLICE_X2Y141_AO6;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_B = CLBLM_R_X3Y141_SLICE_X2Y141_BO6;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_C = CLBLM_R_X3Y141_SLICE_X2Y141_CO6;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_D = CLBLM_R_X3Y141_SLICE_X2Y141_DO6;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_AMUX = CLBLM_R_X3Y141_SLICE_X2Y141_AO5;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_A = CLBLM_R_X3Y141_SLICE_X3Y141_AO6;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_B = CLBLM_R_X3Y141_SLICE_X3Y141_BO6;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_C = CLBLM_R_X3Y141_SLICE_X3Y141_CO6;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_D = CLBLM_R_X3Y141_SLICE_X3Y141_DO6;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_AMUX = CLBLM_R_X3Y141_SLICE_X3Y141_AO5;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_A = CLBLM_R_X3Y142_SLICE_X2Y142_AO6;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_B = CLBLM_R_X3Y142_SLICE_X2Y142_BO6;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_C = CLBLM_R_X3Y142_SLICE_X2Y142_CO6;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_D = CLBLM_R_X3Y142_SLICE_X2Y142_DO6;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_AMUX = CLBLM_R_X3Y142_SLICE_X2Y142_AO5;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_A = CLBLM_R_X3Y142_SLICE_X3Y142_AO6;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_B = CLBLM_R_X3Y142_SLICE_X3Y142_BO6;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_C = CLBLM_R_X3Y142_SLICE_X3Y142_CO6;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_D = CLBLM_R_X3Y142_SLICE_X3Y142_DO6;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_AMUX = CLBLM_R_X3Y142_SLICE_X3Y142_AO5;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_A = CLBLM_R_X3Y143_SLICE_X2Y143_AO6;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_B = CLBLM_R_X3Y143_SLICE_X2Y143_BO6;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_C = CLBLM_R_X3Y143_SLICE_X2Y143_CO6;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_D = CLBLM_R_X3Y143_SLICE_X2Y143_DO6;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_AMUX = CLBLM_R_X3Y143_SLICE_X2Y143_AO5;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_A = CLBLM_R_X3Y143_SLICE_X3Y143_AO6;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_B = CLBLM_R_X3Y143_SLICE_X3Y143_BO6;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_C = CLBLM_R_X3Y143_SLICE_X3Y143_CO6;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_D = CLBLM_R_X3Y143_SLICE_X3Y143_DO6;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_AMUX = CLBLM_R_X3Y143_SLICE_X3Y143_AO5;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_A = CLBLM_R_X5Y132_SLICE_X6Y132_AO6;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_B = CLBLM_R_X5Y132_SLICE_X6Y132_BO6;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_C = CLBLM_R_X5Y132_SLICE_X6Y132_CO6;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_D = CLBLM_R_X5Y132_SLICE_X6Y132_DO6;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_A = CLBLM_R_X5Y132_SLICE_X7Y132_AO6;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_B = CLBLM_R_X5Y132_SLICE_X7Y132_BO6;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_C = CLBLM_R_X5Y132_SLICE_X7Y132_CO6;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_D = CLBLM_R_X5Y132_SLICE_X7Y132_DO6;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_BMUX = CLBLM_R_X5Y132_SLICE_X7Y132_BO5;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_CMUX = CLBLM_R_X5Y132_SLICE_X7Y132_CO5;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_DMUX = CLBLM_R_X5Y132_SLICE_X7Y132_DO6;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_A = CLBLM_R_X5Y133_SLICE_X6Y133_AO6;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_B = CLBLM_R_X5Y133_SLICE_X6Y133_BO6;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_C = CLBLM_R_X5Y133_SLICE_X6Y133_CO6;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_D = CLBLM_R_X5Y133_SLICE_X6Y133_DO6;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_AMUX = CLBLM_R_X5Y133_SLICE_X6Y133_AO5;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_BMUX = CLBLM_R_X5Y133_SLICE_X6Y133_BO6;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_DMUX = CLBLM_R_X5Y133_SLICE_X6Y133_DO6;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_A = CLBLM_R_X5Y133_SLICE_X7Y133_AO6;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_B = CLBLM_R_X5Y133_SLICE_X7Y133_BO6;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_C = CLBLM_R_X5Y133_SLICE_X7Y133_CO6;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_D = CLBLM_R_X5Y133_SLICE_X7Y133_DO6;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_A = CLBLM_R_X5Y134_SLICE_X6Y134_AO6;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_B = CLBLM_R_X5Y134_SLICE_X6Y134_BO6;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_C = CLBLM_R_X5Y134_SLICE_X6Y134_CO6;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_D = CLBLM_R_X5Y134_SLICE_X6Y134_DO6;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_AMUX = CLBLM_R_X5Y134_SLICE_X6Y134_A5Q;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_BMUX = CLBLM_R_X5Y134_SLICE_X6Y134_BO5;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_CMUX = CLBLM_R_X5Y134_SLICE_X6Y134_CO5;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_A = CLBLM_R_X5Y134_SLICE_X7Y134_AO6;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_B = CLBLM_R_X5Y134_SLICE_X7Y134_BO6;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_C = CLBLM_R_X5Y134_SLICE_X7Y134_CO6;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_D = CLBLM_R_X5Y134_SLICE_X7Y134_DO6;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_AMUX = CLBLM_R_X5Y134_SLICE_X7Y134_AO5;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_DMUX = CLBLM_R_X5Y134_SLICE_X7Y134_DO6;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_A = CLBLM_R_X5Y135_SLICE_X6Y135_AO6;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_B = CLBLM_R_X5Y135_SLICE_X6Y135_BO6;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_C = CLBLM_R_X5Y135_SLICE_X6Y135_CO6;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_D = CLBLM_R_X5Y135_SLICE_X6Y135_DO6;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_DMUX = CLBLM_R_X5Y135_SLICE_X6Y135_D5Q;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_A = CLBLM_R_X5Y135_SLICE_X7Y135_AO6;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_B = CLBLM_R_X5Y135_SLICE_X7Y135_BO6;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_C = CLBLM_R_X5Y135_SLICE_X7Y135_CO6;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_D = CLBLM_R_X5Y135_SLICE_X7Y135_DO6;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_AMUX = CLBLM_R_X5Y135_SLICE_X7Y135_A5Q;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_BMUX = CLBLM_R_X5Y135_SLICE_X7Y135_BO5;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_CMUX = CLBLM_R_X5Y135_SLICE_X7Y135_CO5;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_A = CLBLM_R_X5Y136_SLICE_X6Y136_AO6;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_B = CLBLM_R_X5Y136_SLICE_X6Y136_BO6;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_C = CLBLM_R_X5Y136_SLICE_X6Y136_CO6;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_D = CLBLM_R_X5Y136_SLICE_X6Y136_DO6;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_DMUX = CLBLM_R_X5Y136_SLICE_X6Y136_D5Q;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_A = CLBLM_R_X5Y136_SLICE_X7Y136_AO6;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_B = CLBLM_R_X5Y136_SLICE_X7Y136_BO6;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_C = CLBLM_R_X5Y136_SLICE_X7Y136_CO6;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_D = CLBLM_R_X5Y136_SLICE_X7Y136_DO6;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_DMUX = CLBLM_R_X5Y136_SLICE_X7Y136_DO5;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_A = CLBLM_R_X5Y137_SLICE_X6Y137_AO6;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_B = CLBLM_R_X5Y137_SLICE_X6Y137_BO6;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_C = CLBLM_R_X5Y137_SLICE_X6Y137_CO6;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_D = CLBLM_R_X5Y137_SLICE_X6Y137_DO6;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_A = CLBLM_R_X5Y137_SLICE_X7Y137_AO6;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_B = CLBLM_R_X5Y137_SLICE_X7Y137_BO6;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_C = CLBLM_R_X5Y137_SLICE_X7Y137_CO6;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_D = CLBLM_R_X5Y137_SLICE_X7Y137_DO6;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_BMUX = CLBLM_R_X5Y137_SLICE_X7Y137_B5Q;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_CMUX = CLBLM_R_X5Y137_SLICE_X7Y137_C5Q;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_A = CLBLM_R_X5Y138_SLICE_X6Y138_AO6;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_B = CLBLM_R_X5Y138_SLICE_X6Y138_BO6;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_C = CLBLM_R_X5Y138_SLICE_X6Y138_CO6;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_D = CLBLM_R_X5Y138_SLICE_X6Y138_DO6;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_DMUX = CLBLM_R_X5Y138_SLICE_X6Y138_DO6;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_A = CLBLM_R_X5Y138_SLICE_X7Y138_AO6;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_B = CLBLM_R_X5Y138_SLICE_X7Y138_BO6;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_C = CLBLM_R_X5Y138_SLICE_X7Y138_CO6;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_D = CLBLM_R_X5Y138_SLICE_X7Y138_DO6;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_A = CLBLM_R_X5Y139_SLICE_X6Y139_AO6;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_B = CLBLM_R_X5Y139_SLICE_X6Y139_BO6;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_C = CLBLM_R_X5Y139_SLICE_X6Y139_CO6;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_D = CLBLM_R_X5Y139_SLICE_X6Y139_DO6;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_A = CLBLM_R_X5Y139_SLICE_X7Y139_AO6;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_B = CLBLM_R_X5Y139_SLICE_X7Y139_BO6;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_C = CLBLM_R_X5Y139_SLICE_X7Y139_CO6;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_D = CLBLM_R_X5Y139_SLICE_X7Y139_DO6;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_A = CLBLM_R_X5Y140_SLICE_X6Y140_AO6;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_B = CLBLM_R_X5Y140_SLICE_X6Y140_BO6;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_C = CLBLM_R_X5Y140_SLICE_X6Y140_CO6;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_D = CLBLM_R_X5Y140_SLICE_X6Y140_DO6;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_CMUX = CLBLM_R_X5Y140_SLICE_X6Y140_CO6;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_A = CLBLM_R_X5Y140_SLICE_X7Y140_AO6;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_B = CLBLM_R_X5Y140_SLICE_X7Y140_BO6;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_C = CLBLM_R_X5Y140_SLICE_X7Y140_CO6;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_D = CLBLM_R_X5Y140_SLICE_X7Y140_DO6;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_CMUX = CLBLM_R_X5Y140_SLICE_X7Y140_CO6;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_A = CLBLM_R_X5Y141_SLICE_X6Y141_AO6;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_B = CLBLM_R_X5Y141_SLICE_X6Y141_BO6;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_C = CLBLM_R_X5Y141_SLICE_X6Y141_CO6;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_D = CLBLM_R_X5Y141_SLICE_X6Y141_DO6;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_AMUX = CLBLM_R_X5Y141_SLICE_X6Y141_A5Q;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_A = CLBLM_R_X5Y141_SLICE_X7Y141_AO6;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_B = CLBLM_R_X5Y141_SLICE_X7Y141_BO6;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_C = CLBLM_R_X5Y141_SLICE_X7Y141_CO6;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_D = CLBLM_R_X5Y141_SLICE_X7Y141_DO6;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_A = CLBLM_R_X5Y142_SLICE_X6Y142_AO6;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_B = CLBLM_R_X5Y142_SLICE_X6Y142_BO6;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_C = CLBLM_R_X5Y142_SLICE_X6Y142_CO6;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_D = CLBLM_R_X5Y142_SLICE_X6Y142_DO6;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_A = CLBLM_R_X5Y142_SLICE_X7Y142_AO6;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_B = CLBLM_R_X5Y142_SLICE_X7Y142_BO6;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_C = CLBLM_R_X5Y142_SLICE_X7Y142_CO6;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_D = CLBLM_R_X5Y142_SLICE_X7Y142_DO6;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_A = CLBLM_R_X5Y143_SLICE_X6Y143_AO6;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_B = CLBLM_R_X5Y143_SLICE_X6Y143_BO6;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_C = CLBLM_R_X5Y143_SLICE_X6Y143_CO6;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_D = CLBLM_R_X5Y143_SLICE_X6Y143_DO6;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_AMUX = CLBLM_R_X5Y143_SLICE_X6Y143_AO5;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_BMUX = CLBLM_R_X5Y143_SLICE_X6Y143_BO5;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_A = CLBLM_R_X5Y143_SLICE_X7Y143_AO6;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_B = CLBLM_R_X5Y143_SLICE_X7Y143_BO6;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_C = CLBLM_R_X5Y143_SLICE_X7Y143_CO6;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_D = CLBLM_R_X5Y143_SLICE_X7Y143_DO6;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_A = CLBLM_R_X7Y131_SLICE_X8Y131_AO6;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_B = CLBLM_R_X7Y131_SLICE_X8Y131_BO6;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_C = CLBLM_R_X7Y131_SLICE_X8Y131_CO6;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_D = CLBLM_R_X7Y131_SLICE_X8Y131_DO6;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_A = CLBLM_R_X7Y131_SLICE_X9Y131_AO6;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_B = CLBLM_R_X7Y131_SLICE_X9Y131_BO6;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_C = CLBLM_R_X7Y131_SLICE_X9Y131_CO6;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_D = CLBLM_R_X7Y131_SLICE_X9Y131_DO6;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_AMUX = CLBLM_R_X7Y131_SLICE_X9Y131_AO5;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_A = CLBLM_R_X7Y132_SLICE_X8Y132_AO6;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_B = CLBLM_R_X7Y132_SLICE_X8Y132_BO6;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_C = CLBLM_R_X7Y132_SLICE_X8Y132_CO6;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_D = CLBLM_R_X7Y132_SLICE_X8Y132_DO6;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_AMUX = CLBLM_R_X7Y132_SLICE_X8Y132_AO5;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_A = CLBLM_R_X7Y132_SLICE_X9Y132_AO6;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_B = CLBLM_R_X7Y132_SLICE_X9Y132_BO6;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_C = CLBLM_R_X7Y132_SLICE_X9Y132_CO6;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_D = CLBLM_R_X7Y132_SLICE_X9Y132_DO6;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_DMUX = CLBLM_R_X7Y132_SLICE_X9Y132_D5Q;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_A = CLBLM_R_X7Y133_SLICE_X8Y133_AO6;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_B = CLBLM_R_X7Y133_SLICE_X8Y133_BO6;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_C = CLBLM_R_X7Y133_SLICE_X8Y133_CO6;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_D = CLBLM_R_X7Y133_SLICE_X8Y133_DO6;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_A = CLBLM_R_X7Y133_SLICE_X9Y133_AO6;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_B = CLBLM_R_X7Y133_SLICE_X9Y133_BO6;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_C = CLBLM_R_X7Y133_SLICE_X9Y133_CO6;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_D = CLBLM_R_X7Y133_SLICE_X9Y133_DO6;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_A = CLBLM_R_X7Y134_SLICE_X8Y134_AO6;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_B = CLBLM_R_X7Y134_SLICE_X8Y134_BO6;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_C = CLBLM_R_X7Y134_SLICE_X8Y134_CO6;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_D = CLBLM_R_X7Y134_SLICE_X8Y134_DO6;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_CMUX = CLBLM_R_X7Y134_SLICE_X8Y134_C5Q;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_DMUX = CLBLM_R_X7Y134_SLICE_X8Y134_DO5;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_A = CLBLM_R_X7Y134_SLICE_X9Y134_AO6;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_B = CLBLM_R_X7Y134_SLICE_X9Y134_BO6;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_C = CLBLM_R_X7Y134_SLICE_X9Y134_CO6;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_D = CLBLM_R_X7Y134_SLICE_X9Y134_DO6;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_A = CLBLM_R_X7Y135_SLICE_X8Y135_AO6;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_B = CLBLM_R_X7Y135_SLICE_X8Y135_BO6;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_C = CLBLM_R_X7Y135_SLICE_X8Y135_CO6;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_D = CLBLM_R_X7Y135_SLICE_X8Y135_DO6;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_DMUX = CLBLM_R_X7Y135_SLICE_X8Y135_DO5;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_A = CLBLM_R_X7Y135_SLICE_X9Y135_AO6;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_B = CLBLM_R_X7Y135_SLICE_X9Y135_BO6;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_C = CLBLM_R_X7Y135_SLICE_X9Y135_CO6;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_D = CLBLM_R_X7Y135_SLICE_X9Y135_DO6;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_AMUX = CLBLM_R_X7Y135_SLICE_X9Y135_A5Q;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_BMUX = CLBLM_R_X7Y135_SLICE_X9Y135_B5Q;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_CMUX = CLBLM_R_X7Y135_SLICE_X9Y135_CO5;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_A = CLBLM_R_X7Y136_SLICE_X8Y136_AO6;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_B = CLBLM_R_X7Y136_SLICE_X8Y136_BO6;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_C = CLBLM_R_X7Y136_SLICE_X8Y136_CO6;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_D = CLBLM_R_X7Y136_SLICE_X8Y136_DO6;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_DMUX = CLBLM_R_X7Y136_SLICE_X8Y136_DO6;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_A = CLBLM_R_X7Y136_SLICE_X9Y136_AO6;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_B = CLBLM_R_X7Y136_SLICE_X9Y136_BO6;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_C = CLBLM_R_X7Y136_SLICE_X9Y136_CO6;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_D = CLBLM_R_X7Y136_SLICE_X9Y136_DO6;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_BMUX = CLBLM_R_X7Y136_SLICE_X9Y136_BO5;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_A = CLBLM_R_X7Y137_SLICE_X8Y137_AO6;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_B = CLBLM_R_X7Y137_SLICE_X8Y137_BO6;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_C = CLBLM_R_X7Y137_SLICE_X8Y137_CO6;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_D = CLBLM_R_X7Y137_SLICE_X8Y137_DO6;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_DMUX = CLBLM_R_X7Y137_SLICE_X8Y137_DO6;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_A = CLBLM_R_X7Y137_SLICE_X9Y137_AO6;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_B = CLBLM_R_X7Y137_SLICE_X9Y137_BO6;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_C = CLBLM_R_X7Y137_SLICE_X9Y137_CO6;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_D = CLBLM_R_X7Y137_SLICE_X9Y137_DO6;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_A = CLBLM_R_X7Y138_SLICE_X8Y138_AO6;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_B = CLBLM_R_X7Y138_SLICE_X8Y138_BO6;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_C = CLBLM_R_X7Y138_SLICE_X8Y138_CO6;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_D = CLBLM_R_X7Y138_SLICE_X8Y138_DO6;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_A = CLBLM_R_X7Y138_SLICE_X9Y138_AO6;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_B = CLBLM_R_X7Y138_SLICE_X9Y138_BO6;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_C = CLBLM_R_X7Y138_SLICE_X9Y138_CO6;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_D = CLBLM_R_X7Y138_SLICE_X9Y138_DO6;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_A = CLBLM_R_X7Y139_SLICE_X8Y139_AO6;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_B = CLBLM_R_X7Y139_SLICE_X8Y139_BO6;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_C = CLBLM_R_X7Y139_SLICE_X8Y139_CO6;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_D = CLBLM_R_X7Y139_SLICE_X8Y139_DO6;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_AMUX = CLBLM_R_X7Y139_SLICE_X8Y139_A5Q;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_CMUX = CLBLM_R_X7Y139_SLICE_X8Y139_CO5;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_DMUX = CLBLM_R_X7Y139_SLICE_X8Y139_DO5;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_A = CLBLM_R_X7Y139_SLICE_X9Y139_AO6;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_B = CLBLM_R_X7Y139_SLICE_X9Y139_BO6;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_C = CLBLM_R_X7Y139_SLICE_X9Y139_CO6;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_D = CLBLM_R_X7Y139_SLICE_X9Y139_DO6;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_AMUX = CLBLM_R_X7Y139_SLICE_X9Y139_A5Q;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_BMUX = CLBLM_R_X7Y139_SLICE_X9Y139_BO6;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_A = CLBLM_R_X7Y140_SLICE_X8Y140_AO6;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_B = CLBLM_R_X7Y140_SLICE_X8Y140_BO6;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_C = CLBLM_R_X7Y140_SLICE_X8Y140_CO6;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_D = CLBLM_R_X7Y140_SLICE_X8Y140_DO6;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_BMUX = CLBLM_R_X7Y140_SLICE_X8Y140_BO5;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_A = CLBLM_R_X7Y140_SLICE_X9Y140_AO6;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_B = CLBLM_R_X7Y140_SLICE_X9Y140_BO6;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_C = CLBLM_R_X7Y140_SLICE_X9Y140_CO6;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_D = CLBLM_R_X7Y140_SLICE_X9Y140_DO6;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_A = CLBLM_R_X7Y141_SLICE_X8Y141_AO6;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_B = CLBLM_R_X7Y141_SLICE_X8Y141_BO6;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_C = CLBLM_R_X7Y141_SLICE_X8Y141_CO6;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_D = CLBLM_R_X7Y141_SLICE_X8Y141_DO6;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_BMUX = CLBLM_R_X7Y141_SLICE_X8Y141_BO5;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_A = CLBLM_R_X7Y141_SLICE_X9Y141_AO6;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_B = CLBLM_R_X7Y141_SLICE_X9Y141_BO6;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_C = CLBLM_R_X7Y141_SLICE_X9Y141_CO6;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_D = CLBLM_R_X7Y141_SLICE_X9Y141_DO6;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_A = CLBLM_R_X7Y142_SLICE_X8Y142_AO6;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_B = CLBLM_R_X7Y142_SLICE_X8Y142_BO6;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_C = CLBLM_R_X7Y142_SLICE_X8Y142_CO6;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_D = CLBLM_R_X7Y142_SLICE_X8Y142_DO6;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_A = CLBLM_R_X7Y142_SLICE_X9Y142_AO6;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_B = CLBLM_R_X7Y142_SLICE_X9Y142_BO6;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_C = CLBLM_R_X7Y142_SLICE_X9Y142_CO6;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_D = CLBLM_R_X7Y142_SLICE_X9Y142_DO6;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_CMUX = CLBLM_R_X7Y142_SLICE_X9Y142_CO5;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_DMUX = CLBLM_R_X7Y142_SLICE_X9Y142_DO6;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_A = CLBLM_R_X7Y143_SLICE_X8Y143_AO6;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_B = CLBLM_R_X7Y143_SLICE_X8Y143_BO6;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_C = CLBLM_R_X7Y143_SLICE_X8Y143_CO6;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_D = CLBLM_R_X7Y143_SLICE_X8Y143_DO6;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_AMUX = CLBLM_R_X7Y143_SLICE_X8Y143_A5Q;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_BMUX = CLBLM_R_X7Y143_SLICE_X8Y143_BO5;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_A = CLBLM_R_X7Y143_SLICE_X9Y143_AO6;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_B = CLBLM_R_X7Y143_SLICE_X9Y143_BO6;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_C = CLBLM_R_X7Y143_SLICE_X9Y143_CO6;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_D = CLBLM_R_X7Y143_SLICE_X9Y143_DO6;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_A = CLBLM_R_X7Y144_SLICE_X8Y144_AO6;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_B = CLBLM_R_X7Y144_SLICE_X8Y144_BO6;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_C = CLBLM_R_X7Y144_SLICE_X8Y144_CO6;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_D = CLBLM_R_X7Y144_SLICE_X8Y144_DO6;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_A = CLBLM_R_X7Y144_SLICE_X9Y144_AO6;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_B = CLBLM_R_X7Y144_SLICE_X9Y144_BO6;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_C = CLBLM_R_X7Y144_SLICE_X9Y144_CO6;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_D = CLBLM_R_X7Y144_SLICE_X9Y144_DO6;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_A = CLBLM_R_X7Y146_SLICE_X8Y146_AO6;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_B = CLBLM_R_X7Y146_SLICE_X8Y146_BO6;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_C = CLBLM_R_X7Y146_SLICE_X8Y146_CO6;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_D = CLBLM_R_X7Y146_SLICE_X8Y146_DO6;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_A = CLBLM_R_X7Y146_SLICE_X9Y146_AO6;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_B = CLBLM_R_X7Y146_SLICE_X9Y146_BO6;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_C = CLBLM_R_X7Y146_SLICE_X9Y146_CO6;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_D = CLBLM_R_X7Y146_SLICE_X9Y146_DO6;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_A = CLBLM_R_X11Y131_SLICE_X14Y131_AO6;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_B = CLBLM_R_X11Y131_SLICE_X14Y131_BO6;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_C = CLBLM_R_X11Y131_SLICE_X14Y131_CO6;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_D = CLBLM_R_X11Y131_SLICE_X14Y131_DO6;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_AMUX = CLBLM_R_X11Y131_SLICE_X14Y131_AO5;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_A = CLBLM_R_X11Y131_SLICE_X15Y131_AO6;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_B = CLBLM_R_X11Y131_SLICE_X15Y131_BO6;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_C = CLBLM_R_X11Y131_SLICE_X15Y131_CO6;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_D = CLBLM_R_X11Y131_SLICE_X15Y131_DO6;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_AMUX = CLBLM_R_X11Y131_SLICE_X15Y131_AO5;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_A = CLBLM_R_X11Y132_SLICE_X14Y132_AO6;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_B = CLBLM_R_X11Y132_SLICE_X14Y132_BO6;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_C = CLBLM_R_X11Y132_SLICE_X14Y132_CO6;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_D = CLBLM_R_X11Y132_SLICE_X14Y132_DO6;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_A = CLBLM_R_X11Y132_SLICE_X15Y132_AO6;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_B = CLBLM_R_X11Y132_SLICE_X15Y132_BO6;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_C = CLBLM_R_X11Y132_SLICE_X15Y132_CO6;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_D = CLBLM_R_X11Y132_SLICE_X15Y132_DO6;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_AMUX = CLBLM_R_X11Y132_SLICE_X15Y132_AO5;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_CMUX = CLBLM_R_X11Y132_SLICE_X15Y132_CO6;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_A = CLBLM_R_X11Y133_SLICE_X14Y133_AO6;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_B = CLBLM_R_X11Y133_SLICE_X14Y133_BO6;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_C = CLBLM_R_X11Y133_SLICE_X14Y133_CO6;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_D = CLBLM_R_X11Y133_SLICE_X14Y133_DO6;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_A = CLBLM_R_X11Y133_SLICE_X15Y133_AO6;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_B = CLBLM_R_X11Y133_SLICE_X15Y133_BO6;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_C = CLBLM_R_X11Y133_SLICE_X15Y133_CO6;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_D = CLBLM_R_X11Y133_SLICE_X15Y133_DO6;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_A = CLBLM_R_X11Y134_SLICE_X14Y134_AO6;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_B = CLBLM_R_X11Y134_SLICE_X14Y134_BO6;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_C = CLBLM_R_X11Y134_SLICE_X14Y134_CO6;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_D = CLBLM_R_X11Y134_SLICE_X14Y134_DO6;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_A = CLBLM_R_X11Y134_SLICE_X15Y134_AO6;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_B = CLBLM_R_X11Y134_SLICE_X15Y134_BO6;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_C = CLBLM_R_X11Y134_SLICE_X15Y134_CO6;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_D = CLBLM_R_X11Y134_SLICE_X15Y134_DO6;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_A = CLBLM_R_X11Y135_SLICE_X14Y135_AO6;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_B = CLBLM_R_X11Y135_SLICE_X14Y135_BO6;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_C = CLBLM_R_X11Y135_SLICE_X14Y135_CO6;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_D = CLBLM_R_X11Y135_SLICE_X14Y135_DO6;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_A = CLBLM_R_X11Y135_SLICE_X15Y135_AO6;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_B = CLBLM_R_X11Y135_SLICE_X15Y135_BO6;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_C = CLBLM_R_X11Y135_SLICE_X15Y135_CO6;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_D = CLBLM_R_X11Y135_SLICE_X15Y135_DO6;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_CMUX = CLBLM_R_X11Y135_SLICE_X15Y135_CO5;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_A = CLBLM_R_X11Y136_SLICE_X14Y136_AO6;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_B = CLBLM_R_X11Y136_SLICE_X14Y136_BO6;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_C = CLBLM_R_X11Y136_SLICE_X14Y136_CO6;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_D = CLBLM_R_X11Y136_SLICE_X14Y136_DO6;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_CMUX = CLBLM_R_X11Y136_SLICE_X14Y136_CO5;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_A = CLBLM_R_X11Y136_SLICE_X15Y136_AO6;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_B = CLBLM_R_X11Y136_SLICE_X15Y136_BO6;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_C = CLBLM_R_X11Y136_SLICE_X15Y136_CO6;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_D = CLBLM_R_X11Y136_SLICE_X15Y136_DO6;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_AMUX = CLBLM_R_X11Y136_SLICE_X15Y136_A5Q;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_BMUX = CLBLM_R_X11Y136_SLICE_X15Y136_B5Q;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_A = CLBLM_R_X11Y137_SLICE_X14Y137_AO6;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_B = CLBLM_R_X11Y137_SLICE_X14Y137_BO6;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_C = CLBLM_R_X11Y137_SLICE_X14Y137_CO6;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_D = CLBLM_R_X11Y137_SLICE_X14Y137_DO6;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_BMUX = CLBLM_R_X11Y137_SLICE_X14Y137_BO5;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_CMUX = CLBLM_R_X11Y137_SLICE_X14Y137_CO5;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_A = CLBLM_R_X11Y137_SLICE_X15Y137_AO6;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_B = CLBLM_R_X11Y137_SLICE_X15Y137_BO6;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_C = CLBLM_R_X11Y137_SLICE_X15Y137_CO6;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_D = CLBLM_R_X11Y137_SLICE_X15Y137_DO6;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_DMUX = CLBLM_R_X11Y137_SLICE_X15Y137_DO6;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_A = CLBLM_R_X11Y138_SLICE_X14Y138_AO6;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_B = CLBLM_R_X11Y138_SLICE_X14Y138_BO6;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_C = CLBLM_R_X11Y138_SLICE_X14Y138_CO6;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_D = CLBLM_R_X11Y138_SLICE_X14Y138_DO6;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_DMUX = CLBLM_R_X11Y138_SLICE_X14Y138_D5Q;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_A = CLBLM_R_X11Y138_SLICE_X15Y138_AO6;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_B = CLBLM_R_X11Y138_SLICE_X15Y138_BO6;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_C = CLBLM_R_X11Y138_SLICE_X15Y138_CO6;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_D = CLBLM_R_X11Y138_SLICE_X15Y138_DO6;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_BMUX = CLBLM_R_X11Y138_SLICE_X15Y138_B5Q;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_DMUX = CLBLM_R_X11Y138_SLICE_X15Y138_D5Q;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_A = CLBLM_R_X11Y139_SLICE_X14Y139_AO6;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_B = CLBLM_R_X11Y139_SLICE_X14Y139_BO6;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_C = CLBLM_R_X11Y139_SLICE_X14Y139_CO6;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_D = CLBLM_R_X11Y139_SLICE_X14Y139_DO6;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_BMUX = CLBLM_R_X11Y139_SLICE_X14Y139_B5Q;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_A = CLBLM_R_X11Y139_SLICE_X15Y139_AO6;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_B = CLBLM_R_X11Y139_SLICE_X15Y139_BO6;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_C = CLBLM_R_X11Y139_SLICE_X15Y139_CO6;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_D = CLBLM_R_X11Y139_SLICE_X15Y139_DO6;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_AMUX = CLBLM_R_X11Y139_SLICE_X15Y139_A5Q;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_A = CLBLM_R_X11Y140_SLICE_X14Y140_AO6;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_B = CLBLM_R_X11Y140_SLICE_X14Y140_BO6;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_C = CLBLM_R_X11Y140_SLICE_X14Y140_CO6;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_D = CLBLM_R_X11Y140_SLICE_X14Y140_DO6;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_A = CLBLM_R_X11Y140_SLICE_X15Y140_AO6;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_B = CLBLM_R_X11Y140_SLICE_X15Y140_BO6;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_C = CLBLM_R_X11Y140_SLICE_X15Y140_CO6;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_D = CLBLM_R_X11Y140_SLICE_X15Y140_DO6;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_AMUX = CLBLM_R_X11Y140_SLICE_X15Y140_AO5;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_CMUX = CLBLM_R_X11Y140_SLICE_X15Y140_C5Q;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_A = CLBLM_R_X11Y141_SLICE_X14Y141_AO6;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_B = CLBLM_R_X11Y141_SLICE_X14Y141_BO6;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_C = CLBLM_R_X11Y141_SLICE_X14Y141_CO6;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_D = CLBLM_R_X11Y141_SLICE_X14Y141_DO6;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_CMUX = CLBLM_R_X11Y141_SLICE_X14Y141_CO5;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_DMUX = CLBLM_R_X11Y141_SLICE_X14Y141_DO6;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_A = CLBLM_R_X11Y141_SLICE_X15Y141_AO6;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_B = CLBLM_R_X11Y141_SLICE_X15Y141_BO6;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_C = CLBLM_R_X11Y141_SLICE_X15Y141_CO6;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_D = CLBLM_R_X11Y141_SLICE_X15Y141_DO6;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_A = CLBLM_R_X11Y142_SLICE_X14Y142_AO6;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_B = CLBLM_R_X11Y142_SLICE_X14Y142_BO6;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_C = CLBLM_R_X11Y142_SLICE_X14Y142_CO6;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_D = CLBLM_R_X11Y142_SLICE_X14Y142_DO6;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_A = CLBLM_R_X11Y142_SLICE_X15Y142_AO6;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_B = CLBLM_R_X11Y142_SLICE_X15Y142_BO6;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_C = CLBLM_R_X11Y142_SLICE_X15Y142_CO6;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_D = CLBLM_R_X11Y142_SLICE_X15Y142_DO6;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_A = CLBLM_R_X11Y143_SLICE_X14Y143_AO6;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_B = CLBLM_R_X11Y143_SLICE_X14Y143_BO6;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_C = CLBLM_R_X11Y143_SLICE_X14Y143_CO6;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_D = CLBLM_R_X11Y143_SLICE_X14Y143_DO6;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_BMUX = CLBLM_R_X11Y143_SLICE_X14Y143_BO5;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_CMUX = CLBLM_R_X11Y143_SLICE_X14Y143_CO5;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_A = CLBLM_R_X11Y143_SLICE_X15Y143_AO6;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_B = CLBLM_R_X11Y143_SLICE_X15Y143_BO6;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_C = CLBLM_R_X11Y143_SLICE_X15Y143_CO6;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_D = CLBLM_R_X11Y143_SLICE_X15Y143_DO6;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_CMUX = CLBLM_R_X11Y143_SLICE_X15Y143_CO5;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_A = CLBLM_R_X11Y144_SLICE_X14Y144_AO6;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_B = CLBLM_R_X11Y144_SLICE_X14Y144_BO6;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_C = CLBLM_R_X11Y144_SLICE_X14Y144_CO6;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_D = CLBLM_R_X11Y144_SLICE_X14Y144_DO6;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_BMUX = CLBLM_R_X11Y144_SLICE_X14Y144_BO5;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_A = CLBLM_R_X11Y144_SLICE_X15Y144_AO6;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_B = CLBLM_R_X11Y144_SLICE_X15Y144_BO6;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_C = CLBLM_R_X11Y144_SLICE_X15Y144_CO6;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_D = CLBLM_R_X11Y144_SLICE_X15Y144_DO6;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_CMUX = CLBLM_R_X11Y144_SLICE_X15Y144_CO6;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_A = CLBLM_R_X11Y145_SLICE_X14Y145_AO6;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_B = CLBLM_R_X11Y145_SLICE_X14Y145_BO6;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_C = CLBLM_R_X11Y145_SLICE_X14Y145_CO6;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_D = CLBLM_R_X11Y145_SLICE_X14Y145_DO6;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_AMUX = CLBLM_R_X11Y145_SLICE_X14Y145_AO5;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_A = CLBLM_R_X11Y145_SLICE_X15Y145_AO6;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_B = CLBLM_R_X11Y145_SLICE_X15Y145_BO6;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_C = CLBLM_R_X11Y145_SLICE_X15Y145_CO6;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_D = CLBLM_R_X11Y145_SLICE_X15Y145_DO6;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_A = CLBLM_R_X11Y146_SLICE_X14Y146_AO6;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_B = CLBLM_R_X11Y146_SLICE_X14Y146_BO6;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_C = CLBLM_R_X11Y146_SLICE_X14Y146_CO6;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_D = CLBLM_R_X11Y146_SLICE_X14Y146_DO6;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_A = CLBLM_R_X11Y146_SLICE_X15Y146_AO6;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_B = CLBLM_R_X11Y146_SLICE_X15Y146_BO6;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_C = CLBLM_R_X11Y146_SLICE_X15Y146_CO6;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_D = CLBLM_R_X11Y146_SLICE_X15Y146_DO6;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_A = CLBLM_R_X11Y153_SLICE_X14Y153_AO6;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_B = CLBLM_R_X11Y153_SLICE_X14Y153_BO6;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_C = CLBLM_R_X11Y153_SLICE_X14Y153_CO6;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_D = CLBLM_R_X11Y153_SLICE_X14Y153_DO6;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_A = CLBLM_R_X11Y153_SLICE_X15Y153_AO6;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_B = CLBLM_R_X11Y153_SLICE_X15Y153_BO6;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_C = CLBLM_R_X11Y153_SLICE_X15Y153_CO6;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_D = CLBLM_R_X11Y153_SLICE_X15Y153_DO6;
  assign CLBLM_R_X13Y133_SLICE_X18Y133_A = CLBLM_R_X13Y133_SLICE_X18Y133_AO6;
  assign CLBLM_R_X13Y133_SLICE_X18Y133_B = CLBLM_R_X13Y133_SLICE_X18Y133_BO6;
  assign CLBLM_R_X13Y133_SLICE_X18Y133_C = CLBLM_R_X13Y133_SLICE_X18Y133_CO6;
  assign CLBLM_R_X13Y133_SLICE_X18Y133_D = CLBLM_R_X13Y133_SLICE_X18Y133_DO6;
  assign CLBLM_R_X13Y133_SLICE_X19Y133_A = CLBLM_R_X13Y133_SLICE_X19Y133_AO6;
  assign CLBLM_R_X13Y133_SLICE_X19Y133_B = CLBLM_R_X13Y133_SLICE_X19Y133_BO6;
  assign CLBLM_R_X13Y133_SLICE_X19Y133_C = CLBLM_R_X13Y133_SLICE_X19Y133_CO6;
  assign CLBLM_R_X13Y133_SLICE_X19Y133_D = CLBLM_R_X13Y133_SLICE_X19Y133_DO6;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_A = CLBLM_R_X13Y134_SLICE_X18Y134_AO6;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_B = CLBLM_R_X13Y134_SLICE_X18Y134_BO6;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_C = CLBLM_R_X13Y134_SLICE_X18Y134_CO6;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_D = CLBLM_R_X13Y134_SLICE_X18Y134_DO6;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_AMUX = CLBLM_R_X13Y134_SLICE_X18Y134_AO5;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_CMUX = CLBLM_R_X13Y134_SLICE_X18Y134_CO6;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_A = CLBLM_R_X13Y134_SLICE_X19Y134_AO6;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_B = CLBLM_R_X13Y134_SLICE_X19Y134_BO6;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_C = CLBLM_R_X13Y134_SLICE_X19Y134_CO6;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_D = CLBLM_R_X13Y134_SLICE_X19Y134_DO6;
  assign CLBLM_R_X13Y135_SLICE_X18Y135_A = CLBLM_R_X13Y135_SLICE_X18Y135_AO6;
  assign CLBLM_R_X13Y135_SLICE_X18Y135_B = CLBLM_R_X13Y135_SLICE_X18Y135_BO6;
  assign CLBLM_R_X13Y135_SLICE_X18Y135_C = CLBLM_R_X13Y135_SLICE_X18Y135_CO6;
  assign CLBLM_R_X13Y135_SLICE_X18Y135_D = CLBLM_R_X13Y135_SLICE_X18Y135_DO6;
  assign CLBLM_R_X13Y135_SLICE_X19Y135_A = CLBLM_R_X13Y135_SLICE_X19Y135_AO6;
  assign CLBLM_R_X13Y135_SLICE_X19Y135_B = CLBLM_R_X13Y135_SLICE_X19Y135_BO6;
  assign CLBLM_R_X13Y135_SLICE_X19Y135_C = CLBLM_R_X13Y135_SLICE_X19Y135_CO6;
  assign CLBLM_R_X13Y135_SLICE_X19Y135_D = CLBLM_R_X13Y135_SLICE_X19Y135_DO6;
  assign CLBLM_R_X13Y136_SLICE_X18Y136_A = CLBLM_R_X13Y136_SLICE_X18Y136_AO6;
  assign CLBLM_R_X13Y136_SLICE_X18Y136_B = CLBLM_R_X13Y136_SLICE_X18Y136_BO6;
  assign CLBLM_R_X13Y136_SLICE_X18Y136_C = CLBLM_R_X13Y136_SLICE_X18Y136_CO6;
  assign CLBLM_R_X13Y136_SLICE_X18Y136_D = CLBLM_R_X13Y136_SLICE_X18Y136_DO6;
  assign CLBLM_R_X13Y136_SLICE_X19Y136_A = CLBLM_R_X13Y136_SLICE_X19Y136_AO6;
  assign CLBLM_R_X13Y136_SLICE_X19Y136_B = CLBLM_R_X13Y136_SLICE_X19Y136_BO6;
  assign CLBLM_R_X13Y136_SLICE_X19Y136_C = CLBLM_R_X13Y136_SLICE_X19Y136_CO6;
  assign CLBLM_R_X13Y136_SLICE_X19Y136_D = CLBLM_R_X13Y136_SLICE_X19Y136_DO6;
  assign CLBLM_R_X13Y137_SLICE_X18Y137_A = CLBLM_R_X13Y137_SLICE_X18Y137_AO6;
  assign CLBLM_R_X13Y137_SLICE_X18Y137_B = CLBLM_R_X13Y137_SLICE_X18Y137_BO6;
  assign CLBLM_R_X13Y137_SLICE_X18Y137_C = CLBLM_R_X13Y137_SLICE_X18Y137_CO6;
  assign CLBLM_R_X13Y137_SLICE_X18Y137_D = CLBLM_R_X13Y137_SLICE_X18Y137_DO6;
  assign CLBLM_R_X13Y137_SLICE_X18Y137_AMUX = CLBLM_R_X13Y137_SLICE_X18Y137_A5Q;
  assign CLBLM_R_X13Y137_SLICE_X18Y137_BMUX = CLBLM_R_X13Y137_SLICE_X18Y137_BO5;
  assign CLBLM_R_X13Y137_SLICE_X18Y137_CMUX = CLBLM_R_X13Y137_SLICE_X18Y137_CO5;
  assign CLBLM_R_X13Y137_SLICE_X19Y137_A = CLBLM_R_X13Y137_SLICE_X19Y137_AO6;
  assign CLBLM_R_X13Y137_SLICE_X19Y137_B = CLBLM_R_X13Y137_SLICE_X19Y137_BO6;
  assign CLBLM_R_X13Y137_SLICE_X19Y137_C = CLBLM_R_X13Y137_SLICE_X19Y137_CO6;
  assign CLBLM_R_X13Y137_SLICE_X19Y137_D = CLBLM_R_X13Y137_SLICE_X19Y137_DO6;
  assign CLBLM_R_X13Y138_SLICE_X18Y138_A = CLBLM_R_X13Y138_SLICE_X18Y138_AO6;
  assign CLBLM_R_X13Y138_SLICE_X18Y138_B = CLBLM_R_X13Y138_SLICE_X18Y138_BO6;
  assign CLBLM_R_X13Y138_SLICE_X18Y138_C = CLBLM_R_X13Y138_SLICE_X18Y138_CO6;
  assign CLBLM_R_X13Y138_SLICE_X18Y138_D = CLBLM_R_X13Y138_SLICE_X18Y138_DO6;
  assign CLBLM_R_X13Y138_SLICE_X19Y138_A = CLBLM_R_X13Y138_SLICE_X19Y138_AO6;
  assign CLBLM_R_X13Y138_SLICE_X19Y138_B = CLBLM_R_X13Y138_SLICE_X19Y138_BO6;
  assign CLBLM_R_X13Y138_SLICE_X19Y138_C = CLBLM_R_X13Y138_SLICE_X19Y138_CO6;
  assign CLBLM_R_X13Y138_SLICE_X19Y138_D = CLBLM_R_X13Y138_SLICE_X19Y138_DO6;
  assign CLBLM_R_X13Y139_SLICE_X18Y139_A = CLBLM_R_X13Y139_SLICE_X18Y139_AO6;
  assign CLBLM_R_X13Y139_SLICE_X18Y139_B = CLBLM_R_X13Y139_SLICE_X18Y139_BO6;
  assign CLBLM_R_X13Y139_SLICE_X18Y139_C = CLBLM_R_X13Y139_SLICE_X18Y139_CO6;
  assign CLBLM_R_X13Y139_SLICE_X18Y139_D = CLBLM_R_X13Y139_SLICE_X18Y139_DO6;
  assign CLBLM_R_X13Y139_SLICE_X19Y139_A = CLBLM_R_X13Y139_SLICE_X19Y139_AO6;
  assign CLBLM_R_X13Y139_SLICE_X19Y139_B = CLBLM_R_X13Y139_SLICE_X19Y139_BO6;
  assign CLBLM_R_X13Y139_SLICE_X19Y139_C = CLBLM_R_X13Y139_SLICE_X19Y139_CO6;
  assign CLBLM_R_X13Y139_SLICE_X19Y139_D = CLBLM_R_X13Y139_SLICE_X19Y139_DO6;
  assign CLBLM_R_X13Y140_SLICE_X18Y140_A = CLBLM_R_X13Y140_SLICE_X18Y140_AO6;
  assign CLBLM_R_X13Y140_SLICE_X18Y140_B = CLBLM_R_X13Y140_SLICE_X18Y140_BO6;
  assign CLBLM_R_X13Y140_SLICE_X18Y140_C = CLBLM_R_X13Y140_SLICE_X18Y140_CO6;
  assign CLBLM_R_X13Y140_SLICE_X18Y140_D = CLBLM_R_X13Y140_SLICE_X18Y140_DO6;
  assign CLBLM_R_X13Y140_SLICE_X19Y140_A = CLBLM_R_X13Y140_SLICE_X19Y140_AO6;
  assign CLBLM_R_X13Y140_SLICE_X19Y140_B = CLBLM_R_X13Y140_SLICE_X19Y140_BO6;
  assign CLBLM_R_X13Y140_SLICE_X19Y140_C = CLBLM_R_X13Y140_SLICE_X19Y140_CO6;
  assign CLBLM_R_X13Y140_SLICE_X19Y140_D = CLBLM_R_X13Y140_SLICE_X19Y140_DO6;
  assign CLBLM_R_X13Y141_SLICE_X18Y141_A = CLBLM_R_X13Y141_SLICE_X18Y141_AO6;
  assign CLBLM_R_X13Y141_SLICE_X18Y141_B = CLBLM_R_X13Y141_SLICE_X18Y141_BO6;
  assign CLBLM_R_X13Y141_SLICE_X18Y141_C = CLBLM_R_X13Y141_SLICE_X18Y141_CO6;
  assign CLBLM_R_X13Y141_SLICE_X18Y141_D = CLBLM_R_X13Y141_SLICE_X18Y141_DO6;
  assign CLBLM_R_X13Y141_SLICE_X18Y141_AMUX = CLBLM_R_X13Y141_SLICE_X18Y141_AO5;
  assign CLBLM_R_X13Y141_SLICE_X18Y141_BMUX = CLBLM_R_X13Y141_SLICE_X18Y141_BO5;
  assign CLBLM_R_X13Y141_SLICE_X18Y141_CMUX = CLBLM_R_X13Y141_SLICE_X18Y141_CO5;
  assign CLBLM_R_X13Y141_SLICE_X18Y141_DMUX = CLBLM_R_X13Y141_SLICE_X18Y141_DO6;
  assign CLBLM_R_X13Y141_SLICE_X19Y141_A = CLBLM_R_X13Y141_SLICE_X19Y141_AO6;
  assign CLBLM_R_X13Y141_SLICE_X19Y141_B = CLBLM_R_X13Y141_SLICE_X19Y141_BO6;
  assign CLBLM_R_X13Y141_SLICE_X19Y141_C = CLBLM_R_X13Y141_SLICE_X19Y141_CO6;
  assign CLBLM_R_X13Y141_SLICE_X19Y141_D = CLBLM_R_X13Y141_SLICE_X19Y141_DO6;
  assign CLBLM_R_X13Y141_SLICE_X19Y141_CMUX = CLBLM_R_X13Y141_SLICE_X19Y141_CO5;
  assign CLBLM_R_X13Y142_SLICE_X18Y142_A = CLBLM_R_X13Y142_SLICE_X18Y142_AO6;
  assign CLBLM_R_X13Y142_SLICE_X18Y142_B = CLBLM_R_X13Y142_SLICE_X18Y142_BO6;
  assign CLBLM_R_X13Y142_SLICE_X18Y142_C = CLBLM_R_X13Y142_SLICE_X18Y142_CO6;
  assign CLBLM_R_X13Y142_SLICE_X18Y142_D = CLBLM_R_X13Y142_SLICE_X18Y142_DO6;
  assign CLBLM_R_X13Y142_SLICE_X19Y142_A = CLBLM_R_X13Y142_SLICE_X19Y142_AO6;
  assign CLBLM_R_X13Y142_SLICE_X19Y142_B = CLBLM_R_X13Y142_SLICE_X19Y142_BO6;
  assign CLBLM_R_X13Y142_SLICE_X19Y142_C = CLBLM_R_X13Y142_SLICE_X19Y142_CO6;
  assign CLBLM_R_X13Y142_SLICE_X19Y142_D = CLBLM_R_X13Y142_SLICE_X19Y142_DO6;
  assign CLBLM_R_X13Y143_SLICE_X18Y143_A = CLBLM_R_X13Y143_SLICE_X18Y143_AO6;
  assign CLBLM_R_X13Y143_SLICE_X18Y143_B = CLBLM_R_X13Y143_SLICE_X18Y143_BO6;
  assign CLBLM_R_X13Y143_SLICE_X18Y143_C = CLBLM_R_X13Y143_SLICE_X18Y143_CO6;
  assign CLBLM_R_X13Y143_SLICE_X18Y143_D = CLBLM_R_X13Y143_SLICE_X18Y143_DO6;
  assign CLBLM_R_X13Y143_SLICE_X18Y143_AMUX = CLBLM_R_X13Y143_SLICE_X18Y143_AO5;
  assign CLBLM_R_X13Y143_SLICE_X18Y143_CMUX = CLBLM_R_X13Y143_SLICE_X18Y143_CO6;
  assign CLBLM_R_X13Y143_SLICE_X19Y143_A = CLBLM_R_X13Y143_SLICE_X19Y143_AO6;
  assign CLBLM_R_X13Y143_SLICE_X19Y143_B = CLBLM_R_X13Y143_SLICE_X19Y143_BO6;
  assign CLBLM_R_X13Y143_SLICE_X19Y143_C = CLBLM_R_X13Y143_SLICE_X19Y143_CO6;
  assign CLBLM_R_X13Y143_SLICE_X19Y143_D = CLBLM_R_X13Y143_SLICE_X19Y143_DO6;
  assign CLBLM_R_X13Y144_SLICE_X18Y144_A = CLBLM_R_X13Y144_SLICE_X18Y144_AO6;
  assign CLBLM_R_X13Y144_SLICE_X18Y144_B = CLBLM_R_X13Y144_SLICE_X18Y144_BO6;
  assign CLBLM_R_X13Y144_SLICE_X18Y144_C = CLBLM_R_X13Y144_SLICE_X18Y144_CO6;
  assign CLBLM_R_X13Y144_SLICE_X18Y144_D = CLBLM_R_X13Y144_SLICE_X18Y144_DO6;
  assign CLBLM_R_X13Y144_SLICE_X18Y144_BMUX = CLBLM_R_X13Y144_SLICE_X18Y144_BO5;
  assign CLBLM_R_X13Y144_SLICE_X19Y144_A = CLBLM_R_X13Y144_SLICE_X19Y144_AO6;
  assign CLBLM_R_X13Y144_SLICE_X19Y144_B = CLBLM_R_X13Y144_SLICE_X19Y144_BO6;
  assign CLBLM_R_X13Y144_SLICE_X19Y144_C = CLBLM_R_X13Y144_SLICE_X19Y144_CO6;
  assign CLBLM_R_X13Y144_SLICE_X19Y144_D = CLBLM_R_X13Y144_SLICE_X19Y144_DO6;
  assign CLBLM_R_X15Y142_SLICE_X20Y142_A = CLBLM_R_X15Y142_SLICE_X20Y142_AO6;
  assign CLBLM_R_X15Y142_SLICE_X20Y142_B = CLBLM_R_X15Y142_SLICE_X20Y142_BO6;
  assign CLBLM_R_X15Y142_SLICE_X20Y142_C = CLBLM_R_X15Y142_SLICE_X20Y142_CO6;
  assign CLBLM_R_X15Y142_SLICE_X20Y142_D = CLBLM_R_X15Y142_SLICE_X20Y142_DO6;
  assign CLBLM_R_X15Y142_SLICE_X21Y142_A = CLBLM_R_X15Y142_SLICE_X21Y142_AO6;
  assign CLBLM_R_X15Y142_SLICE_X21Y142_B = CLBLM_R_X15Y142_SLICE_X21Y142_BO6;
  assign CLBLM_R_X15Y142_SLICE_X21Y142_C = CLBLM_R_X15Y142_SLICE_X21Y142_CO6;
  assign CLBLM_R_X15Y142_SLICE_X21Y142_D = CLBLM_R_X15Y142_SLICE_X21Y142_DO6;
  assign CLBLM_R_X37Y138_SLICE_X56Y138_A = CLBLM_R_X37Y138_SLICE_X56Y138_AO6;
  assign CLBLM_R_X37Y138_SLICE_X56Y138_B = CLBLM_R_X37Y138_SLICE_X56Y138_BO6;
  assign CLBLM_R_X37Y138_SLICE_X56Y138_C = CLBLM_R_X37Y138_SLICE_X56Y138_CO6;
  assign CLBLM_R_X37Y138_SLICE_X56Y138_D = CLBLM_R_X37Y138_SLICE_X56Y138_DO6;
  assign CLBLM_R_X37Y138_SLICE_X57Y138_A = CLBLM_R_X37Y138_SLICE_X57Y138_AO6;
  assign CLBLM_R_X37Y138_SLICE_X57Y138_B = CLBLM_R_X37Y138_SLICE_X57Y138_BO6;
  assign CLBLM_R_X37Y138_SLICE_X57Y138_C = CLBLM_R_X37Y138_SLICE_X57Y138_CO6;
  assign CLBLM_R_X37Y138_SLICE_X57Y138_D = CLBLM_R_X37Y138_SLICE_X57Y138_DO6;
  assign CLBLM_R_X103Y140_SLICE_X162Y140_A = CLBLM_R_X103Y140_SLICE_X162Y140_AO6;
  assign CLBLM_R_X103Y140_SLICE_X162Y140_B = CLBLM_R_X103Y140_SLICE_X162Y140_BO6;
  assign CLBLM_R_X103Y140_SLICE_X162Y140_C = CLBLM_R_X103Y140_SLICE_X162Y140_CO6;
  assign CLBLM_R_X103Y140_SLICE_X162Y140_D = CLBLM_R_X103Y140_SLICE_X162Y140_DO6;
  assign CLBLM_R_X103Y140_SLICE_X163Y140_A = CLBLM_R_X103Y140_SLICE_X163Y140_AO6;
  assign CLBLM_R_X103Y140_SLICE_X163Y140_B = CLBLM_R_X103Y140_SLICE_X163Y140_BO6;
  assign CLBLM_R_X103Y140_SLICE_X163Y140_C = CLBLM_R_X103Y140_SLICE_X163Y140_CO6;
  assign CLBLM_R_X103Y140_SLICE_X163Y140_D = CLBLM_R_X103Y140_SLICE_X163Y140_DO6;
  assign CLBLM_R_X103Y140_SLICE_X163Y140_AMUX = CLBLM_R_X103Y140_SLICE_X163Y140_AO5;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_A = CLBLM_R_X103Y169_SLICE_X162Y169_AO6;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_B = CLBLM_R_X103Y169_SLICE_X162Y169_BO6;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_C = CLBLM_R_X103Y169_SLICE_X162Y169_CO6;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_D = CLBLM_R_X103Y169_SLICE_X162Y169_DO6;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_A = CLBLM_R_X103Y169_SLICE_X163Y169_AO6;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_B = CLBLM_R_X103Y169_SLICE_X163Y169_BO6;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_C = CLBLM_R_X103Y169_SLICE_X163Y169_CO6;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_D = CLBLM_R_X103Y169_SLICE_X163Y169_DO6;
  assign CLBLM_R_X103Y170_SLICE_X162Y170_A = CLBLM_R_X103Y170_SLICE_X162Y170_AO6;
  assign CLBLM_R_X103Y170_SLICE_X162Y170_B = CLBLM_R_X103Y170_SLICE_X162Y170_BO6;
  assign CLBLM_R_X103Y170_SLICE_X162Y170_C = CLBLM_R_X103Y170_SLICE_X162Y170_CO6;
  assign CLBLM_R_X103Y170_SLICE_X162Y170_D = CLBLM_R_X103Y170_SLICE_X162Y170_DO6;
  assign CLBLM_R_X103Y170_SLICE_X163Y170_A = CLBLM_R_X103Y170_SLICE_X163Y170_AO6;
  assign CLBLM_R_X103Y170_SLICE_X163Y170_B = CLBLM_R_X103Y170_SLICE_X163Y170_BO6;
  assign CLBLM_R_X103Y170_SLICE_X163Y170_C = CLBLM_R_X103Y170_SLICE_X163Y170_CO6;
  assign CLBLM_R_X103Y170_SLICE_X163Y170_D = CLBLM_R_X103Y170_SLICE_X163Y170_DO6;
  assign CLBLM_R_X103Y170_SLICE_X163Y170_AMUX = CLBLM_R_X103Y170_SLICE_X163Y170_AO5;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_A = CLBLM_R_X103Y173_SLICE_X162Y173_AO6;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_B = CLBLM_R_X103Y173_SLICE_X162Y173_BO6;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_C = CLBLM_R_X103Y173_SLICE_X162Y173_CO6;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_D = CLBLM_R_X103Y173_SLICE_X162Y173_DO6;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_A = CLBLM_R_X103Y173_SLICE_X163Y173_AO6;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_B = CLBLM_R_X103Y173_SLICE_X163Y173_BO6;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_C = CLBLM_R_X103Y173_SLICE_X163Y173_CO6;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_D = CLBLM_R_X103Y173_SLICE_X163Y173_DO6;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_AMUX = CLBLM_R_X103Y173_SLICE_X163Y173_AO5;
  assign CLBLM_R_X103Y175_SLICE_X162Y175_A = CLBLM_R_X103Y175_SLICE_X162Y175_AO6;
  assign CLBLM_R_X103Y175_SLICE_X162Y175_B = CLBLM_R_X103Y175_SLICE_X162Y175_BO6;
  assign CLBLM_R_X103Y175_SLICE_X162Y175_C = CLBLM_R_X103Y175_SLICE_X162Y175_CO6;
  assign CLBLM_R_X103Y175_SLICE_X162Y175_D = CLBLM_R_X103Y175_SLICE_X162Y175_DO6;
  assign CLBLM_R_X103Y175_SLICE_X163Y175_A = CLBLM_R_X103Y175_SLICE_X163Y175_AO6;
  assign CLBLM_R_X103Y175_SLICE_X163Y175_B = CLBLM_R_X103Y175_SLICE_X163Y175_BO6;
  assign CLBLM_R_X103Y175_SLICE_X163Y175_C = CLBLM_R_X103Y175_SLICE_X163Y175_CO6;
  assign CLBLM_R_X103Y175_SLICE_X163Y175_D = CLBLM_R_X103Y175_SLICE_X163Y175_DO6;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_A = CLBLM_R_X103Y177_SLICE_X162Y177_AO6;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_B = CLBLM_R_X103Y177_SLICE_X162Y177_BO6;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_C = CLBLM_R_X103Y177_SLICE_X162Y177_CO6;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_D = CLBLM_R_X103Y177_SLICE_X162Y177_DO6;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_A = CLBLM_R_X103Y177_SLICE_X163Y177_AO6;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_B = CLBLM_R_X103Y177_SLICE_X163Y177_BO6;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_C = CLBLM_R_X103Y177_SLICE_X163Y177_CO6;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_D = CLBLM_R_X103Y177_SLICE_X163Y177_DO6;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_AMUX = CLBLM_R_X103Y177_SLICE_X163Y177_AO5;
  assign LIOI3_X0Y51_ILOGIC_X0Y52_O = LIOB33_X0Y51_IOB_X0Y52_I;
  assign LIOI3_X0Y51_ILOGIC_X0Y51_O = LIOB33_X0Y51_IOB_X0Y51_I;
  assign LIOI3_X0Y53_ILOGIC_X0Y54_O = LIOB33_X0Y53_IOB_X0Y54_I;
  assign LIOI3_X0Y53_ILOGIC_X0Y53_O = LIOB33_X0Y53_IOB_X0Y53_I;
  assign LIOI3_X0Y55_ILOGIC_X0Y56_O = LIOB33_X0Y55_IOB_X0Y56_I;
  assign LIOI3_X0Y55_ILOGIC_X0Y55_O = LIOB33_X0Y55_IOB_X0Y55_I;
  assign LIOI3_X0Y59_ILOGIC_X0Y60_O = LIOB33_X0Y59_IOB_X0Y60_I;
  assign LIOI3_X0Y59_ILOGIC_X0Y59_O = LIOB33_X0Y59_IOB_X0Y59_I;
  assign LIOI3_X0Y61_ILOGIC_X0Y62_O = LIOB33_X0Y61_IOB_X0Y62_I;
  assign LIOI3_X0Y61_ILOGIC_X0Y61_O = LIOB33_X0Y61_IOB_X0Y61_I;
  assign LIOI3_X0Y65_ILOGIC_X0Y66_O = LIOB33_X0Y65_IOB_X0Y66_I;
  assign LIOI3_X0Y65_ILOGIC_X0Y65_O = LIOB33_X0Y65_IOB_X0Y65_I;
  assign LIOI3_X0Y67_ILOGIC_X0Y68_O = LIOB33_X0Y67_IOB_X0Y68_I;
  assign LIOI3_X0Y67_ILOGIC_X0Y67_O = LIOB33_X0Y67_IOB_X0Y67_I;
  assign LIOI3_X0Y71_ILOGIC_X0Y72_O = LIOB33_X0Y71_IOB_X0Y72_I;
  assign LIOI3_X0Y71_ILOGIC_X0Y71_O = LIOB33_X0Y71_IOB_X0Y71_I;
  assign LIOI3_X0Y73_ILOGIC_X0Y74_O = LIOB33_X0Y73_IOB_X0Y74_I;
  assign LIOI3_X0Y73_ILOGIC_X0Y73_O = LIOB33_X0Y73_IOB_X0Y73_I;
  assign LIOI3_X0Y75_ILOGIC_X0Y76_O = LIOB33_X0Y75_IOB_X0Y76_I;
  assign LIOI3_X0Y75_ILOGIC_X0Y75_O = LIOB33_X0Y75_IOB_X0Y75_I;
  assign LIOI3_X0Y77_ILOGIC_X0Y78_O = LIOB33_X0Y77_IOB_X0Y78_I;
  assign LIOI3_X0Y77_ILOGIC_X0Y77_O = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOI3_X0Y79_ILOGIC_X0Y79_O = LIOB33_X0Y79_IOB_X0Y79_I;
  assign LIOI3_X0Y79_OLOGIC_X0Y80_OQ = CLBLL_L_X2Y133_SLICE_X0Y133_AO6;
  assign LIOI3_X0Y79_OLOGIC_X0Y80_TQ = 1'b1;
  assign LIOI3_X0Y101_OLOGIC_X0Y102_OQ = CLBLM_R_X3Y133_SLICE_X2Y133_AO5;
  assign LIOI3_X0Y101_OLOGIC_X0Y102_TQ = 1'b1;
  assign LIOI3_X0Y101_OLOGIC_X0Y101_OQ = CLBLM_R_X3Y133_SLICE_X2Y133_AO6;
  assign LIOI3_X0Y101_OLOGIC_X0Y101_TQ = 1'b1;
  assign LIOI3_X0Y103_OLOGIC_X0Y104_OQ = CLBLL_L_X2Y133_SLICE_X0Y133_CO6;
  assign LIOI3_X0Y103_OLOGIC_X0Y104_TQ = 1'b1;
  assign LIOI3_X0Y103_OLOGIC_X0Y103_OQ = CLBLL_L_X2Y133_SLICE_X0Y133_AO5;
  assign LIOI3_X0Y103_OLOGIC_X0Y103_TQ = 1'b1;
  assign LIOI3_X0Y105_OLOGIC_X0Y106_OQ = CLBLL_L_X4Y138_SLICE_X5Y138_DO6;
  assign LIOI3_X0Y105_OLOGIC_X0Y106_TQ = 1'b1;
  assign LIOI3_X0Y105_OLOGIC_X0Y105_OQ = CLBLL_L_X2Y133_SLICE_X0Y133_BO5;
  assign LIOI3_X0Y105_OLOGIC_X0Y105_TQ = 1'b1;
  assign LIOI3_X0Y109_OLOGIC_X0Y110_OQ = CLBLL_L_X2Y127_SLICE_X0Y127_AO5;
  assign LIOI3_X0Y109_OLOGIC_X0Y110_TQ = 1'b1;
  assign LIOI3_X0Y109_OLOGIC_X0Y109_OQ = CLBLL_L_X2Y127_SLICE_X0Y127_AO6;
  assign LIOI3_X0Y109_OLOGIC_X0Y109_TQ = 1'b1;
  assign LIOI3_X0Y111_OLOGIC_X0Y112_OQ = CLBLM_L_X12Y133_SLICE_X16Y133_C5Q;
  assign LIOI3_X0Y111_OLOGIC_X0Y112_TQ = 1'b1;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_OQ = 1'b0;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_TQ = 1'b1;
  assign LIOI3_X0Y115_OLOGIC_X0Y116_OQ = CLBLM_L_X8Y135_SLICE_X11Y135_BQ;
  assign LIOI3_X0Y115_OLOGIC_X0Y116_TQ = 1'b1;
  assign LIOI3_X0Y115_OLOGIC_X0Y115_OQ = CLBLM_L_X12Y133_SLICE_X16Y133_CQ;
  assign LIOI3_X0Y115_OLOGIC_X0Y115_TQ = 1'b1;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_OQ = CLBLL_L_X4Y135_SLICE_X5Y135_DQ;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_TQ = 1'b1;
  assign LIOI3_X0Y117_OLOGIC_X0Y117_OQ = CLBLM_R_X5Y136_SLICE_X6Y136_D5Q;
  assign LIOI3_X0Y117_OLOGIC_X0Y117_TQ = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_OQ = CLBLL_L_X4Y133_SLICE_X5Y133_A5Q;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_TQ = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_OQ = CLBLM_L_X8Y135_SLICE_X11Y135_B5Q;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_TQ = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_OQ = CLBLL_L_X4Y135_SLICE_X5Y135_D5Q;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_TQ = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_OQ = CLBLM_R_X7Y132_SLICE_X9Y132_D5Q;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_TQ = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_OQ = CLBLM_R_X3Y136_SLICE_X3Y136_CQ;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_TQ = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_OQ = CLBLM_R_X11Y138_SLICE_X15Y138_D5Q;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_TQ = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_OQ = CLBLL_L_X4Y134_SLICE_X5Y134_A5Q;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_TQ = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_OQ = CLBLM_R_X5Y137_SLICE_X6Y137_BQ;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_TQ = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_OQ = CLBLL_L_X52Y126_SLICE_X78Y126_AO6;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_TQ = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_OQ = CLBLM_R_X5Y136_SLICE_X6Y136_CQ;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_TQ = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_OQ = CLBLM_R_X3Y133_SLICE_X3Y133_AQ;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_TQ = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_OQ = CLBLM_R_X3Y137_SLICE_X3Y137_AQ;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_TQ = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_OQ = CLBLM_R_X3Y135_SLICE_X3Y135_AQ;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_TQ = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_OQ = CLBLM_R_X3Y136_SLICE_X3Y136_AQ;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_TQ = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_OQ = CLBLM_R_X3Y136_SLICE_X2Y136_AQ;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_TQ = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_OQ = CLBLM_R_X3Y137_SLICE_X2Y137_AQ;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_TQ = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_OQ = LIOB33_X0Y53_IOB_X0Y54_I;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_TQ = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_OQ = CLBLM_R_X3Y136_SLICE_X3Y136_BQ;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_TQ = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_OQ = LIOB33_X0Y59_IOB_X0Y59_I;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_TQ = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_OQ = LIOB33_X0Y57_IOB_X0Y58_I;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_TQ = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_OQ = LIOB33_X0Y61_IOB_X0Y61_I;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_TQ = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_OQ = LIOB33_X0Y71_IOB_X0Y71_I;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_TQ = 1'b1;
  assign LIOI3_X0Y151_OLOGIC_X0Y152_OQ = LIOB33_X0Y65_IOB_X0Y66_I;
  assign LIOI3_X0Y151_OLOGIC_X0Y152_TQ = 1'b1;
  assign LIOI3_X0Y151_OLOGIC_X0Y151_OQ = LIOB33_X0Y65_IOB_X0Y65_I;
  assign LIOI3_X0Y151_OLOGIC_X0Y151_TQ = 1'b1;
  assign LIOI3_X0Y153_OLOGIC_X0Y154_OQ = LIOB33_X0Y67_IOB_X0Y68_I;
  assign LIOI3_X0Y153_OLOGIC_X0Y154_TQ = 1'b1;
  assign LIOI3_X0Y153_OLOGIC_X0Y153_OQ = LIOB33_X0Y67_IOB_X0Y67_I;
  assign LIOI3_X0Y153_OLOGIC_X0Y153_TQ = 1'b1;
  assign LIOI3_X0Y155_OLOGIC_X0Y156_OQ = RIOB33_X105Y105_IOB_X1Y106_I;
  assign LIOI3_X0Y155_OLOGIC_X0Y156_TQ = 1'b1;
  assign LIOI3_X0Y155_OLOGIC_X0Y155_OQ = LIOB33_X0Y69_IOB_X0Y70_I;
  assign LIOI3_X0Y155_OLOGIC_X0Y155_TQ = 1'b1;
  assign LIOI3_X0Y159_OLOGIC_X0Y160_OQ = RIOB33_X105Y107_IOB_X1Y107_I;
  assign LIOI3_X0Y159_OLOGIC_X0Y160_TQ = 1'b1;
  assign LIOI3_X0Y159_OLOGIC_X0Y159_OQ = RIOB33_X105Y117_IOB_X1Y117_I;
  assign LIOI3_X0Y159_OLOGIC_X0Y159_TQ = 1'b1;
  assign LIOI3_X0Y161_OLOGIC_X0Y162_OQ = RIOB33_X105Y109_IOB_X1Y109_I;
  assign LIOI3_X0Y161_OLOGIC_X0Y162_TQ = 1'b1;
  assign LIOI3_X0Y161_OLOGIC_X0Y161_OQ = RIOB33_X105Y107_IOB_X1Y108_I;
  assign LIOI3_X0Y161_OLOGIC_X0Y161_TQ = 1'b1;
  assign LIOI3_X0Y165_OLOGIC_X0Y166_OQ = RIOB33_X105Y113_IOB_X1Y113_I;
  assign LIOI3_X0Y165_OLOGIC_X0Y166_TQ = 1'b1;
  assign LIOI3_X0Y165_OLOGIC_X0Y165_OQ = RIOB33_X105Y111_IOB_X1Y112_I;
  assign LIOI3_X0Y165_OLOGIC_X0Y165_TQ = 1'b1;
  assign LIOI3_X0Y167_OLOGIC_X0Y168_OQ = RIOB33_X105Y123_IOB_X1Y123_I;
  assign LIOI3_X0Y167_OLOGIC_X0Y168_TQ = 1'b1;
  assign LIOI3_X0Y167_OLOGIC_X0Y167_OQ = RIOB33_X105Y113_IOB_X1Y114_I;
  assign LIOI3_X0Y167_OLOGIC_X0Y167_TQ = 1'b1;
  assign LIOI3_X0Y171_OLOGIC_X0Y172_OQ = CLBLM_R_X103Y140_SLICE_X163Y140_AO6;
  assign LIOI3_X0Y171_OLOGIC_X0Y172_TQ = 1'b1;
  assign LIOI3_X0Y171_OLOGIC_X0Y171_OQ = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign LIOI3_X0Y171_OLOGIC_X0Y171_TQ = 1'b1;
  assign LIOI3_X0Y173_OLOGIC_X0Y174_OQ = CLBLM_R_X11Y153_SLICE_X14Y153_AO6;
  assign LIOI3_X0Y173_OLOGIC_X0Y174_TQ = 1'b1;
  assign LIOI3_X0Y173_OLOGIC_X0Y173_OQ = CLBLM_R_X103Y140_SLICE_X163Y140_AO5;
  assign LIOI3_X0Y173_OLOGIC_X0Y173_TQ = 1'b1;
  assign LIOI3_X0Y175_OLOGIC_X0Y176_OQ = RIOB33_X105Y127_IOB_X1Y128_I;
  assign LIOI3_X0Y175_OLOGIC_X0Y176_TQ = 1'b1;
  assign LIOI3_X0Y175_OLOGIC_X0Y175_OQ = RIOB33_X105Y127_IOB_X1Y127_I;
  assign LIOI3_X0Y175_OLOGIC_X0Y175_TQ = 1'b1;
  assign LIOI3_X0Y177_OLOGIC_X0Y178_OQ = RIOB33_X105Y129_IOB_X1Y130_I;
  assign LIOI3_X0Y177_OLOGIC_X0Y178_TQ = 1'b1;
  assign LIOI3_X0Y177_OLOGIC_X0Y177_OQ = RIOB33_X105Y129_IOB_X1Y129_I;
  assign LIOI3_X0Y177_OLOGIC_X0Y177_TQ = 1'b1;
  assign LIOI3_X0Y179_OLOGIC_X0Y180_OQ = RIOB33_X105Y131_IOB_X1Y132_I;
  assign LIOI3_X0Y179_OLOGIC_X0Y180_TQ = 1'b1;
  assign LIOI3_X0Y179_OLOGIC_X0Y179_OQ = RIOB33_X105Y131_IOB_X1Y131_I;
  assign LIOI3_X0Y179_OLOGIC_X0Y179_TQ = 1'b1;
  assign LIOI3_X0Y183_OLOGIC_X0Y184_OQ = RIOB33_X105Y135_IOB_X1Y136_I;
  assign LIOI3_X0Y183_OLOGIC_X0Y184_TQ = 1'b1;
  assign LIOI3_X0Y183_OLOGIC_X0Y183_OQ = RIOB33_X105Y135_IOB_X1Y135_I;
  assign LIOI3_X0Y183_OLOGIC_X0Y183_TQ = 1'b1;
  assign LIOI3_X0Y185_OLOGIC_X0Y186_OQ = RIOB33_X105Y143_IOB_X1Y143_I;
  assign LIOI3_X0Y185_OLOGIC_X0Y186_TQ = 1'b1;
  assign LIOI3_X0Y185_OLOGIC_X0Y185_OQ = RIOB33_X105Y137_IOB_X1Y137_I;
  assign LIOI3_X0Y185_OLOGIC_X0Y185_TQ = 1'b1;
  assign LIOI3_X0Y189_OLOGIC_X0Y190_OQ = RIOB33_X105Y147_IOB_X1Y147_I;
  assign LIOI3_X0Y189_OLOGIC_X0Y190_TQ = 1'b1;
  assign LIOI3_X0Y189_OLOGIC_X0Y189_OQ = RIOB33_X105Y145_IOB_X1Y146_I;
  assign LIOI3_X0Y189_OLOGIC_X0Y189_TQ = 1'b1;
  assign LIOI3_X0Y191_OLOGIC_X0Y192_OQ = LIOB33_X0Y51_IOB_X0Y52_I;
  assign LIOI3_X0Y191_OLOGIC_X0Y192_TQ = 1'b1;
  assign LIOI3_X0Y191_OLOGIC_X0Y191_OQ = RIOB33_X105Y147_IOB_X1Y148_I;
  assign LIOI3_X0Y191_OLOGIC_X0Y191_TQ = 1'b1;
  assign LIOI3_X0Y195_OLOGIC_X0Y196_OQ = LIOB33_X0Y69_IOB_X0Y69_I;
  assign LIOI3_X0Y195_OLOGIC_X0Y196_TQ = 1'b1;
  assign LIOI3_X0Y195_OLOGIC_X0Y195_OQ = LIOB33_X0Y63_IOB_X0Y64_I;
  assign LIOI3_X0Y195_OLOGIC_X0Y195_TQ = 1'b1;
  assign LIOI3_X0Y197_OLOGIC_X0Y198_OQ = LIOB33_X0Y73_IOB_X0Y73_I;
  assign LIOI3_X0Y197_OLOGIC_X0Y198_TQ = 1'b1;
  assign LIOI3_X0Y197_OLOGIC_X0Y197_OQ = LIOB33_X0Y71_IOB_X0Y72_I;
  assign LIOI3_X0Y197_OLOGIC_X0Y197_TQ = 1'b1;
  assign LIOI3_SING_X0Y50_ILOGIC_X0Y50_O = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign LIOI3_SING_X0Y100_OLOGIC_X0Y100_OQ = CLBLL_L_X2Y133_SLICE_X0Y133_BO6;
  assign LIOI3_SING_X0Y100_OLOGIC_X0Y100_TQ = 1'b1;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_OQ = LIOB33_X0Y61_IOB_X0Y62_I;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_TQ = 1'b1;
  assign LIOI3_SING_X0Y150_OLOGIC_X0Y150_OQ = LIOB33_X0Y63_IOB_X0Y63_I;
  assign LIOI3_SING_X0Y150_OLOGIC_X0Y150_TQ = 1'b1;
  assign LIOI3_SING_X0Y199_OLOGIC_X0Y199_OQ = LIOB33_X0Y73_IOB_X0Y74_I;
  assign LIOI3_SING_X0Y199_OLOGIC_X0Y199_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y58_O = LIOB33_X0Y57_IOB_X0Y58_I;
  assign LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y57_O = LIOB33_X0Y57_IOB_X0Y57_I;
  assign LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y70_O = LIOB33_X0Y69_IOB_X0Y70_I;
  assign LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y69_O = LIOB33_X0Y69_IOB_X0Y69_I;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_OQ = CLBLL_L_X2Y133_SLICE_X0Y133_CO5;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_OQ = CLBLL_L_X2Y108_SLICE_X0Y108_AO6;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_OQ = CLBLM_L_X12Y136_SLICE_X16Y136_BQ;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_OQ = CLBLM_L_X10Y135_SLICE_X13Y135_BQ;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_OQ = CLBLM_R_X7Y131_SLICE_X9Y131_AQ;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_OQ = CLBLM_R_X7Y131_SLICE_X9Y131_AO5;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_OQ = LIOB33_X0Y57_IOB_X0Y57_I;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_OQ = LIOB33_X0Y55_IOB_X0Y55_I;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_OQ = RIOB33_X105Y115_IOB_X1Y116_I;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_OQ = RIOB33_X105Y115_IOB_X1Y115_I;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_OQ = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_OQ = RIOB33_X105Y121_IOB_X1Y122_I;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_OQ = RIOB33_X105Y133_IOB_X1Y134_I;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_OQ = RIOB33_X105Y133_IOB_X1Y133_I;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_OQ = LIOB33_X0Y59_IOB_X0Y60_I;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_OQ = LIOB33_X0Y55_IOB_X0Y56_I;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y64_O = LIOB33_X0Y63_IOB_X0Y64_I;
  assign LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y63_O = LIOB33_X0Y63_IOB_X0Y63_I;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_OQ = CLBLM_R_X7Y132_SLICE_X9Y132_DQ;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_OQ = RIOB33_X105Y121_IOB_X1Y121_I;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_OQ = CLBLM_R_X3Y136_SLICE_X3Y136_DQ;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_OQ = CLBLM_R_X3Y137_SLICE_X2Y137_BQ;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_OQ = RIOB33_X105Y111_IOB_X1Y111_I;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_OQ = RIOB33_X105Y109_IOB_X1Y110_I;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_OQ = RIOB33_X105Y145_IOB_X1Y145_I;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_OQ = RIOB33_X105Y143_IOB_X1Y144_I;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_TQ = 1'b1;
  assign RIOI3_X105Y101_ILOGIC_X1Y102_O = RIOB33_X105Y101_IOB_X1Y102_I;
  assign RIOI3_X105Y101_ILOGIC_X1Y101_O = RIOB33_X105Y101_IOB_X1Y101_I;
  assign RIOI3_X105Y103_ILOGIC_X1Y104_O = RIOB33_X105Y103_IOB_X1Y104_I;
  assign RIOI3_X105Y103_ILOGIC_X1Y103_O = RIOB33_X105Y103_IOB_X1Y103_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y106_O = RIOB33_X105Y105_IOB_X1Y106_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y105_O = RIOB33_X105Y105_IOB_X1Y105_I;
  assign RIOI3_X105Y109_ILOGIC_X1Y110_O = RIOB33_X105Y109_IOB_X1Y110_I;
  assign RIOI3_X105Y109_ILOGIC_X1Y109_O = RIOB33_X105Y109_IOB_X1Y109_I;
  assign RIOI3_X105Y111_ILOGIC_X1Y112_O = RIOB33_X105Y111_IOB_X1Y112_I;
  assign RIOI3_X105Y111_ILOGIC_X1Y111_O = RIOB33_X105Y111_IOB_X1Y111_I;
  assign RIOI3_X105Y115_ILOGIC_X1Y116_O = RIOB33_X105Y115_IOB_X1Y116_I;
  assign RIOI3_X105Y115_ILOGIC_X1Y115_O = RIOB33_X105Y115_IOB_X1Y115_I;
  assign RIOI3_X105Y117_ILOGIC_X1Y118_O = RIOB33_X105Y117_IOB_X1Y118_I;
  assign RIOI3_X105Y117_ILOGIC_X1Y117_O = RIOB33_X105Y117_IOB_X1Y117_I;
  assign RIOI3_X105Y121_ILOGIC_X1Y122_O = RIOB33_X105Y121_IOB_X1Y122_I;
  assign RIOI3_X105Y121_ILOGIC_X1Y121_O = RIOB33_X105Y121_IOB_X1Y121_I;
  assign RIOI3_X105Y123_ILOGIC_X1Y124_O = RIOB33_X105Y123_IOB_X1Y124_I;
  assign RIOI3_X105Y123_ILOGIC_X1Y123_O = RIOB33_X105Y123_IOB_X1Y123_I;
  assign RIOI3_X105Y125_ILOGIC_X1Y126_O = RIOB33_X105Y125_IOB_X1Y126_I;
  assign RIOI3_X105Y125_ILOGIC_X1Y125_O = RIOB33_X105Y125_IOB_X1Y125_I;
  assign RIOI3_X105Y127_ILOGIC_X1Y128_O = RIOB33_X105Y127_IOB_X1Y128_I;
  assign RIOI3_X105Y127_ILOGIC_X1Y127_O = RIOB33_X105Y127_IOB_X1Y127_I;
  assign RIOI3_X105Y129_ILOGIC_X1Y130_O = RIOB33_X105Y129_IOB_X1Y130_I;
  assign RIOI3_X105Y129_ILOGIC_X1Y129_O = RIOB33_X105Y129_IOB_X1Y129_I;
  assign RIOI3_X105Y133_ILOGIC_X1Y134_O = RIOB33_X105Y133_IOB_X1Y134_I;
  assign RIOI3_X105Y133_ILOGIC_X1Y133_O = RIOB33_X105Y133_IOB_X1Y133_I;
  assign RIOI3_X105Y135_ILOGIC_X1Y136_O = RIOB33_X105Y135_IOB_X1Y136_I;
  assign RIOI3_X105Y135_ILOGIC_X1Y135_O = RIOB33_X105Y135_IOB_X1Y135_I;
  assign RIOI3_X105Y139_ILOGIC_X1Y140_O = RIOB33_X105Y139_IOB_X1Y140_I;
  assign RIOI3_X105Y139_ILOGIC_X1Y139_O = RIOB33_X105Y139_IOB_X1Y139_I;
  assign RIOI3_X105Y141_ILOGIC_X1Y142_O = RIOB33_X105Y141_IOB_X1Y142_I;
  assign RIOI3_X105Y141_ILOGIC_X1Y141_O = RIOB33_X105Y141_IOB_X1Y141_I;
  assign RIOI3_X105Y145_ILOGIC_X1Y146_O = RIOB33_X105Y145_IOB_X1Y146_I;
  assign RIOI3_X105Y145_ILOGIC_X1Y145_O = RIOB33_X105Y145_IOB_X1Y145_I;
  assign RIOI3_X105Y147_ILOGIC_X1Y148_O = RIOB33_X105Y147_IOB_X1Y148_I;
  assign RIOI3_X105Y147_ILOGIC_X1Y147_O = RIOB33_X105Y147_IOB_X1Y147_I;
  assign RIOI3_X105Y151_OLOGIC_X1Y152_OQ = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign RIOI3_X105Y151_OLOGIC_X1Y152_TQ = 1'b1;
  assign RIOI3_X105Y151_OLOGIC_X1Y151_OQ = LIOB33_X0Y75_IOB_X0Y76_I;
  assign RIOI3_X105Y151_OLOGIC_X1Y151_TQ = 1'b1;
  assign RIOI3_X105Y153_OLOGIC_X1Y154_OQ = RIOB33_X105Y101_IOB_X1Y102_I;
  assign RIOI3_X105Y153_OLOGIC_X1Y154_TQ = 1'b1;
  assign RIOI3_X105Y153_OLOGIC_X1Y153_OQ = RIOB33_X105Y101_IOB_X1Y101_I;
  assign RIOI3_X105Y153_OLOGIC_X1Y153_TQ = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y156_OQ = RIOB33_X105Y103_IOB_X1Y104_I;
  assign RIOI3_X105Y155_OLOGIC_X1Y156_TQ = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y155_OQ = RIOB33_X105Y103_IOB_X1Y103_I;
  assign RIOI3_X105Y155_OLOGIC_X1Y155_TQ = 1'b1;
  assign RIOI3_X105Y159_OLOGIC_X1Y160_OQ = CLBLM_L_X12Y138_SLICE_X17Y138_DO5;
  assign RIOI3_X105Y159_OLOGIC_X1Y160_TQ = 1'b1;
  assign RIOI3_X105Y159_OLOGIC_X1Y159_OQ = CLBLM_L_X12Y138_SLICE_X17Y138_DO6;
  assign RIOI3_X105Y159_OLOGIC_X1Y159_TQ = 1'b1;
  assign RIOI3_X105Y161_OLOGIC_X1Y162_OQ = CLBLM_R_X11Y141_SLICE_X14Y141_CO5;
  assign RIOI3_X105Y161_OLOGIC_X1Y162_TQ = 1'b1;
  assign RIOI3_X105Y161_OLOGIC_X1Y161_OQ = CLBLM_R_X11Y141_SLICE_X14Y141_CO6;
  assign RIOI3_X105Y161_OLOGIC_X1Y161_TQ = 1'b1;
  assign RIOI3_X105Y165_OLOGIC_X1Y166_OQ = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign RIOI3_X105Y165_OLOGIC_X1Y166_TQ = 1'b1;
  assign RIOI3_X105Y165_OLOGIC_X1Y165_OQ = RIOB33_X105Y125_IOB_X1Y125_I;
  assign RIOI3_X105Y165_OLOGIC_X1Y165_TQ = 1'b1;
  assign RIOI3_X105Y167_OLOGIC_X1Y168_OQ = CLBLM_R_X11Y153_SLICE_X14Y153_AO6;
  assign RIOI3_X105Y167_OLOGIC_X1Y168_TQ = 1'b1;
  assign RIOI3_X105Y167_OLOGIC_X1Y167_OQ = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign RIOI3_X105Y167_OLOGIC_X1Y167_TQ = 1'b1;
  assign RIOI3_X105Y171_OLOGIC_X1Y172_OQ = CLBLM_R_X103Y170_SLICE_X163Y170_AO5;
  assign RIOI3_X105Y171_OLOGIC_X1Y172_TQ = 1'b1;
  assign RIOI3_X105Y171_OLOGIC_X1Y171_OQ = CLBLM_L_X10Y146_SLICE_X12Y146_AO5;
  assign RIOI3_X105Y171_OLOGIC_X1Y171_TQ = 1'b1;
  assign RIOI3_X105Y173_OLOGIC_X1Y174_OQ = CLBLM_R_X103Y173_SLICE_X163Y173_AO6;
  assign RIOI3_X105Y173_OLOGIC_X1Y174_TQ = 1'b1;
  assign RIOI3_X105Y173_OLOGIC_X1Y173_OQ = CLBLM_R_X11Y144_SLICE_X14Y144_BO5;
  assign RIOI3_X105Y173_OLOGIC_X1Y173_TQ = 1'b1;
  assign RIOI3_X105Y175_OLOGIC_X1Y176_OQ = CLBLM_R_X103Y173_SLICE_X163Y173_AO5;
  assign RIOI3_X105Y175_OLOGIC_X1Y176_TQ = 1'b1;
  assign RIOI3_X105Y175_OLOGIC_X1Y175_OQ = CLBLM_L_X12Y146_SLICE_X16Y146_AO6;
  assign RIOI3_X105Y175_OLOGIC_X1Y175_TQ = 1'b1;
  assign RIOI3_X105Y177_OLOGIC_X1Y178_OQ = CLBLM_R_X103Y177_SLICE_X163Y177_AO5;
  assign RIOI3_X105Y177_OLOGIC_X1Y178_TQ = 1'b1;
  assign RIOI3_X105Y177_OLOGIC_X1Y177_OQ = CLBLM_R_X103Y177_SLICE_X163Y177_AO6;
  assign RIOI3_X105Y177_OLOGIC_X1Y177_TQ = 1'b1;
  assign RIOI3_X105Y179_OLOGIC_X1Y180_OQ = CLBLM_L_X12Y138_SLICE_X17Y138_DO6;
  assign RIOI3_X105Y179_OLOGIC_X1Y180_TQ = 1'b1;
  assign RIOI3_X105Y179_OLOGIC_X1Y179_OQ = CLBLM_L_X12Y144_SLICE_X17Y144_AO5;
  assign RIOI3_X105Y179_OLOGIC_X1Y179_TQ = 1'b1;
  assign RIOI3_X105Y183_OLOGIC_X1Y184_OQ = CLBLM_L_X12Y139_SLICE_X17Y139_DO6;
  assign RIOI3_X105Y183_OLOGIC_X1Y184_TQ = 1'b1;
  assign RIOI3_X105Y183_OLOGIC_X1Y183_OQ = CLBLM_R_X11Y141_SLICE_X14Y141_CO5;
  assign RIOI3_X105Y183_OLOGIC_X1Y183_TQ = 1'b1;
  assign RIOI3_X105Y185_OLOGIC_X1Y186_OQ = CLBLM_R_X13Y139_SLICE_X19Y139_AQ;
  assign RIOI3_X105Y185_OLOGIC_X1Y186_TQ = 1'b1;
  assign RIOI3_X105Y185_OLOGIC_X1Y185_OQ = CLBLM_L_X12Y139_SLICE_X17Y139_DO5;
  assign RIOI3_X105Y185_OLOGIC_X1Y185_TQ = 1'b1;
  assign RIOI3_X105Y189_OLOGIC_X1Y190_OQ = CLBLM_R_X15Y142_SLICE_X20Y142_AQ;
  assign RIOI3_X105Y189_OLOGIC_X1Y190_TQ = 1'b1;
  assign RIOI3_X105Y189_OLOGIC_X1Y189_OQ = CLBLM_L_X10Y143_SLICE_X13Y143_BQ;
  assign RIOI3_X105Y189_OLOGIC_X1Y189_TQ = 1'b1;
  assign RIOI3_X105Y191_OLOGIC_X1Y192_OQ = CLBLM_R_X13Y134_SLICE_X19Y134_BQ;
  assign RIOI3_X105Y191_OLOGIC_X1Y192_TQ = 1'b1;
  assign RIOI3_X105Y191_OLOGIC_X1Y191_OQ = CLBLM_L_X10Y143_SLICE_X13Y143_AQ;
  assign RIOI3_X105Y191_OLOGIC_X1Y191_TQ = 1'b1;
  assign RIOI3_X105Y195_OLOGIC_X1Y196_OQ = CLBLM_R_X13Y143_SLICE_X18Y143_AQ;
  assign RIOI3_X105Y195_OLOGIC_X1Y196_TQ = 1'b1;
  assign RIOI3_X105Y195_OLOGIC_X1Y195_OQ = CLBLM_R_X13Y143_SLICE_X18Y143_BQ;
  assign RIOI3_X105Y195_OLOGIC_X1Y195_TQ = 1'b1;
  assign RIOI3_X105Y197_OLOGIC_X1Y198_OQ = CLBLM_R_X103Y175_SLICE_X163Y175_AO6;
  assign RIOI3_X105Y197_OLOGIC_X1Y198_TQ = 1'b1;
  assign RIOI3_X105Y197_OLOGIC_X1Y197_OQ = CLBLM_R_X103Y175_SLICE_X163Y175_AO6;
  assign RIOI3_X105Y197_OLOGIC_X1Y197_TQ = 1'b1;
  assign RIOI3_SING_X105Y100_ILOGIC_X1Y100_O = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign RIOI3_SING_X105Y149_ILOGIC_X1Y149_O = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign RIOI3_SING_X105Y150_OLOGIC_X1Y150_OQ = LIOB33_X0Y75_IOB_X0Y75_I;
  assign RIOI3_SING_X105Y150_OLOGIC_X1Y150_TQ = 1'b1;
  assign RIOI3_SING_X105Y199_OLOGIC_X1Y199_OQ = CLBLM_R_X13Y144_SLICE_X19Y144_AQ;
  assign RIOI3_SING_X105Y199_OLOGIC_X1Y199_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_O = RIOB33_X105Y107_IOB_X1Y108_I;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_O = RIOB33_X105Y107_IOB_X1Y107_I;
  assign RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_O = RIOB33_X105Y119_IOB_X1Y119_I;
  assign RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y132_O = RIOB33_X105Y131_IOB_X1Y132_I;
  assign RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y131_O = RIOB33_X105Y131_IOB_X1Y131_I;
  assign RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y144_O = RIOB33_X105Y143_IOB_X1Y144_I;
  assign RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y143_O = RIOB33_X105Y143_IOB_X1Y143_I;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_OQ = CLBLM_R_X37Y138_SLICE_X56Y138_AO6;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_OQ = RIOB33_X105Y125_IOB_X1Y126_I;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_OQ = CLBLM_R_X103Y170_SLICE_X163Y170_AO6;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_OQ = CLBLM_R_X103Y169_SLICE_X163Y169_AO6;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_OQ = CLBLM_R_X11Y141_SLICE_X14Y141_CO6;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_OQ = CLBLM_L_X12Y138_SLICE_X17Y138_DO5;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_OQ = CLBLM_R_X13Y144_SLICE_X19Y144_AQ;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_OQ = CLBLM_L_X12Y144_SLICE_X16Y144_AQ;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y114_O = RIOB33_X105Y113_IOB_X1Y114_I;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_O = RIOB33_X105Y113_IOB_X1Y113_I;
  assign RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y138_O = RIOB33_X105Y137_IOB_X1Y138_I;
  assign RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y137_O = RIOB33_X105Y137_IOB_X1Y137_I;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_OQ = CLBLM_L_X12Y139_SLICE_X17Y139_DO5;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_OQ = CLBLM_L_X12Y139_SLICE_X17Y139_DO6;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_OQ = CLBLM_R_X11Y144_SLICE_X15Y144_AQ;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_OQ = CLBLM_L_X12Y134_SLICE_X16Y134_AQ;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_TQ = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_B5 = 1'b1;
  assign LIOB33_X0Y147_IOB_X0Y148_O = LIOB33_X0Y61_IOB_X0Y61_I;
  assign LIOB33_X0Y147_IOB_X0Y147_O = LIOB33_X0Y71_IOB_X0Y71_I;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_B5 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_C1 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_C2 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_C3 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_C4 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_C6 = 1'b1;
  assign LIOI3_X0Y155_OLOGIC_X0Y156_D1 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_A1 = CLBLL_L_X4Y139_SLICE_X5Y139_AQ;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_A2 = CLBLM_R_X11Y136_SLICE_X15Y136_BQ;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_A3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_A4 = CLBLM_L_X10Y139_SLICE_X12Y139_AQ;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_A6 = 1'b1;
  assign LIOI3_X0Y155_OLOGIC_X0Y156_T1 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_B1 = CLBLM_R_X7Y140_SLICE_X9Y140_BQ;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_B2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_B3 = CLBLM_L_X8Y138_SLICE_X10Y138_AQ;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_B4 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_B5 = CLBLM_L_X8Y138_SLICE_X10Y138_BQ;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_B6 = CLBLM_R_X7Y137_SLICE_X8Y137_CQ;
  assign LIOI3_X0Y155_OLOGIC_X0Y155_D1 = LIOB33_X0Y69_IOB_X0Y70_I;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_C1 = CLBLL_L_X4Y142_SLICE_X5Y142_DO6;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_C2 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_C3 = CLBLM_R_X5Y141_SLICE_X7Y141_DO6;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_C4 = CLBLL_L_X4Y139_SLICE_X4Y139_BO6;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_C5 = CLBLM_R_X7Y139_SLICE_X9Y139_DO6;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_C6 = CLBLM_R_X5Y140_SLICE_X6Y140_AO6;
  assign LIOB33_X0Y127_IOB_X0Y127_O = CLBLM_R_X5Y137_SLICE_X6Y137_BQ;
  assign LIOB33_X0Y127_IOB_X0Y128_O = CLBLL_L_X4Y134_SLICE_X5Y134_A5Q;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y155_OLOGIC_X0Y155_T1 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_D1 = CLBLM_R_X5Y142_SLICE_X6Y142_CO6;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_D2 = CLBLM_R_X11Y138_SLICE_X14Y138_DQ;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_D3 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_D4 = CLBLL_L_X4Y141_SLICE_X4Y141_DO6;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_D5 = CLBLM_R_X3Y140_SLICE_X2Y140_DO6;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_D6 = CLBLL_L_X4Y142_SLICE_X4Y142_BO6;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_A1 = CLBLM_R_X7Y139_SLICE_X8Y139_AQ;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_A2 = CLBLM_R_X7Y140_SLICE_X8Y140_BO6;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_A3 = CLBLM_L_X12Y135_SLICE_X17Y135_AQ;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_A4 = CLBLM_R_X7Y139_SLICE_X8Y139_DO5;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_A6 = CLBLM_R_X11Y135_SLICE_X14Y135_AQ;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_AX = CLBLM_R_X7Y139_SLICE_X8Y139_CO6;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_B1 = CLBLM_R_X7Y139_SLICE_X9Y139_A5Q;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_B2 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_B4 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_B6 = CLBLM_R_X7Y144_SLICE_X9Y144_AQ;
  assign RIOB33_SING_X105Y150_IOB_X1Y150_O = LIOB33_X0Y75_IOB_X0Y75_I;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_C2 = CLBLM_R_X7Y139_SLICE_X8Y139_AQ;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_C3 = CLBLM_L_X8Y142_SLICE_X10Y142_DQ;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_C4 = CLBLM_R_X11Y138_SLICE_X15Y138_AQ;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_C6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_D1 = CLBLM_R_X11Y141_SLICE_X14Y141_CO6;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_D1 = CLBLM_R_X11Y136_SLICE_X14Y136_AQ;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_D2 = CLBLM_R_X7Y139_SLICE_X8Y139_AQ;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_D3 = CLBLM_R_X7Y139_SLICE_X9Y139_BO6;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_D4 = CLBLM_R_X11Y138_SLICE_X14Y138_BQ;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_D5 = CLBLM_L_X8Y142_SLICE_X10Y142_DQ;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_D6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_D1 = CLBLM_L_X12Y138_SLICE_X17Y138_DO5;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_T1 = 1'b1;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_A3 = CLBLM_R_X7Y132_SLICE_X9Y132_BQ;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_A4 = CLBLM_R_X7Y132_SLICE_X9Y132_CQ;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_A5 = CLBLM_L_X8Y138_SLICE_X10Y138_AQ;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_A6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_B2 = CLBLM_L_X8Y134_SLICE_X11Y134_BQ;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_D6 = 1'b1;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_B5 = 1'b1;
  assign LIOI3_SING_X0Y199_OLOGIC_X0Y199_D1 = LIOB33_X0Y73_IOB_X0Y74_I;
  assign LIOB33_X0Y151_IOB_X0Y152_O = LIOB33_X0Y65_IOB_X0Y66_I;
  assign LIOB33_X0Y151_IOB_X0Y151_O = LIOB33_X0Y65_IOB_X0Y65_I;
  assign RIOB33_SING_X105Y199_IOB_X1Y199_O = CLBLM_R_X13Y144_SLICE_X19Y144_AQ;
  assign LIOI3_SING_X0Y199_OLOGIC_X0Y199_T1 = 1'b1;
  assign RIOI3_X105Y139_ILOGIC_X1Y140_D = RIOB33_X105Y139_IOB_X1Y140_I;
  assign RIOI3_X105Y139_ILOGIC_X1Y139_D = RIOB33_X105Y139_IOB_X1Y139_I;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_A1 = CLBLM_L_X8Y143_SLICE_X10Y143_DO6;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_A2 = CLBLM_R_X5Y140_SLICE_X7Y140_BQ;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_A3 = CLBLM_R_X7Y140_SLICE_X9Y140_AQ;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_A4 = 1'b1;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_A6 = CLBLM_L_X10Y140_SLICE_X13Y140_DQ;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_B1 = CLBLM_L_X10Y140_SLICE_X13Y140_DQ;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_B2 = CLBLM_R_X7Y140_SLICE_X9Y140_BQ;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_B3 = CLBLM_L_X8Y138_SLICE_X10Y138_AQ;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_B4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_B6 = CLBLM_R_X11Y135_SLICE_X14Y135_AQ;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_C2 = CLBLM_R_X7Y140_SLICE_X8Y140_CO6;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_C3 = CLBLM_L_X8Y143_SLICE_X10Y143_DO5;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_C4 = CLBLM_L_X12Y139_SLICE_X16Y139_A5Q;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_C5 = CLBLM_R_X7Y140_SLICE_X9Y140_CQ;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_C6 = CLBLM_R_X11Y137_SLICE_X14Y137_AQ;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y191_OLOGIC_X0Y192_D1 = LIOB33_X0Y51_IOB_X0Y52_I;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_D1 = CLBLM_R_X7Y142_SLICE_X9Y142_CO5;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_D2 = CLBLM_L_X8Y141_SLICE_X11Y141_CQ;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_D3 = 1'b1;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_D4 = 1'b1;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_D5 = CLBLM_R_X5Y143_SLICE_X6Y143_AO5;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_D6 = CLBLM_L_X10Y140_SLICE_X12Y140_AQ;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_A1 = CLBLL_L_X4Y138_SLICE_X5Y138_CO5;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_A2 = CLBLM_L_X8Y137_SLICE_X11Y137_BQ;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_A3 = CLBLM_R_X7Y140_SLICE_X8Y140_AQ;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_A6 = CLBLM_R_X5Y141_SLICE_X7Y141_DO6;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_B1 = CLBLM_R_X7Y139_SLICE_X9Y139_BO6;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_B2 = CLBLM_R_X11Y138_SLICE_X14Y138_BQ;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_B3 = 1'b1;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_B4 = CLBLM_R_X11Y136_SLICE_X14Y136_AQ;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_B5 = 1'b1;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_B6 = 1'b1;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_C1 = CLBLL_L_X4Y143_SLICE_X5Y143_AO6;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_C2 = CLBLM_L_X8Y137_SLICE_X10Y137_DO6;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_C3 = CLBLM_R_X5Y132_SLICE_X7Y132_DO6;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_C4 = CLBLL_L_X4Y142_SLICE_X4Y142_DO6;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_C5 = CLBLM_R_X13Y141_SLICE_X18Y141_AO5;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_C6 = CLBLM_L_X10Y141_SLICE_X13Y141_CQ;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_D1 = CLBLM_R_X7Y139_SLICE_X8Y139_AQ;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_D2 = CLBLM_R_X11Y135_SLICE_X14Y135_AQ;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_D3 = CLBLM_R_X7Y139_SLICE_X9Y139_BO6;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_D4 = CLBLM_R_X11Y138_SLICE_X14Y138_BQ;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_D5 = CLBLM_L_X8Y142_SLICE_X10Y142_DQ;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_D6 = CLBLM_R_X11Y136_SLICE_X14Y136_AQ;
  assign LIOB33_X0Y153_IOB_X0Y154_O = LIOB33_X0Y67_IOB_X0Y68_I;
  assign LIOB33_X0Y153_IOB_X0Y153_O = LIOB33_X0Y67_IOB_X0Y67_I;
  assign RIOI3_X105Y165_OLOGIC_X1Y165_D1 = RIOB33_X105Y125_IOB_X1Y125_I;
  assign CLBLM_R_X103Y175_SLICE_X163Y175_A1 = 1'b1;
  assign CLBLM_R_X103Y175_SLICE_X163Y175_A2 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLM_R_X103Y175_SLICE_X163Y175_A3 = 1'b1;
  assign CLBLM_R_X103Y175_SLICE_X163Y175_A4 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X103Y175_SLICE_X163Y175_A5 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_A1 = CLBLM_R_X7Y141_SLICE_X9Y141_AQ;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_A2 = CLBLL_L_X4Y137_SLICE_X4Y137_CQ;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_A4 = CLBLM_L_X12Y135_SLICE_X17Y135_AQ;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_A5 = CLBLM_L_X8Y142_SLICE_X10Y142_DQ;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_A6 = CLBLM_L_X8Y138_SLICE_X10Y138_D5Q;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_B2 = CLBLM_R_X7Y141_SLICE_X9Y141_BQ;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_B3 = CLBLM_L_X10Y139_SLICE_X13Y139_B5Q;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_B4 = CLBLM_R_X7Y140_SLICE_X9Y140_BQ;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_B5 = CLBLM_R_X7Y140_SLICE_X9Y140_AQ;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_B6 = CLBLM_L_X12Y134_SLICE_X17Y134_AO6;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_D6 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_C1 = CLBLM_L_X12Y141_SLICE_X17Y141_AQ;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_C2 = CLBLM_R_X3Y143_SLICE_X2Y143_AO5;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_C3 = CLBLM_R_X7Y143_SLICE_X9Y143_DO6;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_C4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_C5 = CLBLM_L_X12Y136_SLICE_X16Y136_C5Q;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_C6 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_D1 = CLBLM_R_X5Y143_SLICE_X6Y143_AO5;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_D2 = CLBLL_L_X4Y143_SLICE_X5Y143_AO5;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_D3 = CLBLM_R_X7Y142_SLICE_X9Y142_CO6;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_D4 = CLBLM_R_X7Y142_SLICE_X9Y142_BQ;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_D5 = CLBLM_R_X7Y141_SLICE_X9Y141_AQ;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_D6 = CLBLM_R_X11Y141_SLICE_X15Y141_BQ;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_A1 = CLBLM_R_X7Y141_SLICE_X8Y141_DO6;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_A2 = CLBLM_R_X7Y143_SLICE_X8Y143_CQ;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_A4 = CLBLM_R_X7Y141_SLICE_X8Y141_BO6;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_A5 = CLBLM_R_X11Y138_SLICE_X14Y138_DQ;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_A6 = CLBLM_R_X7Y140_SLICE_X8Y140_BO5;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_B1 = CLBLM_R_X7Y139_SLICE_X8Y139_AQ;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_B2 = CLBLM_R_X7Y140_SLICE_X9Y140_BQ;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_B3 = CLBLM_L_X8Y142_SLICE_X10Y142_DQ;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_B4 = CLBLM_R_X7Y137_SLICE_X8Y137_CQ;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_B5 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_B6 = 1'b1;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_BX = CLBLM_R_X11Y140_SLICE_X15Y140_AO6;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_C1 = CLBLM_R_X7Y139_SLICE_X8Y139_CO5;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_C2 = CLBLM_R_X7Y141_SLICE_X8Y141_BO5;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_C3 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_C4 = CLBLM_R_X7Y140_SLICE_X8Y140_BO5;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_C5 = CLBLM_L_X8Y138_SLICE_X10Y138_BQ;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_A1 = 1'b1;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_A2 = 1'b1;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_A3 = 1'b1;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_A4 = 1'b1;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_A5 = 1'b1;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_A6 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_C6 = CLBLM_R_X11Y138_SLICE_X14Y138_DQ;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_B1 = 1'b1;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_B2 = 1'b1;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_B3 = 1'b1;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_B4 = 1'b1;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_B5 = 1'b1;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_B6 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_D1 = CLBLM_R_X5Y139_SLICE_X7Y139_AQ;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_D2 = CLBLM_L_X8Y138_SLICE_X10Y138_D5Q;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_D3 = 1'b1;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_C1 = 1'b1;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_C2 = 1'b1;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_C3 = 1'b1;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_C4 = 1'b1;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_C5 = 1'b1;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_C6 = 1'b1;
  assign LIOI3_X0Y159_OLOGIC_X0Y160_D1 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_D1 = 1'b1;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_D2 = 1'b1;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_D3 = 1'b1;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_D4 = 1'b1;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_D5 = 1'b1;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_D6 = 1'b1;
  assign LIOI3_X0Y159_OLOGIC_X0Y160_T1 = 1'b1;
  assign LIOI3_X0Y159_OLOGIC_X0Y159_D1 = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLL_L_X2Y140_SLICE_X1Y140_A1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y140_SLICE_X1Y140_A2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y140_SLICE_X1Y140_A3 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y140_SLICE_X1Y140_A4 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y140_SLICE_X1Y140_A5 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLL_L_X2Y140_SLICE_X1Y140_A6 = 1'b1;
  assign LIOB33_X0Y155_IOB_X0Y155_O = LIOB33_X0Y69_IOB_X0Y70_I;
  assign LIOB33_X0Y155_IOB_X0Y156_O = RIOB33_X105Y105_IOB_X1Y106_I;
  assign LIOI3_X0Y159_OLOGIC_X0Y159_T1 = 1'b1;
  assign CLBLL_L_X2Y140_SLICE_X1Y140_B1 = 1'b1;
  assign CLBLL_L_X2Y140_SLICE_X1Y140_B2 = 1'b1;
  assign CLBLL_L_X2Y140_SLICE_X1Y140_B3 = 1'b1;
  assign CLBLL_L_X2Y140_SLICE_X1Y140_B4 = 1'b1;
  assign CLBLL_L_X2Y140_SLICE_X1Y140_B5 = 1'b1;
  assign CLBLL_L_X2Y140_SLICE_X1Y140_B6 = 1'b1;
  assign CLBLL_L_X2Y140_SLICE_X1Y140_C1 = 1'b1;
  assign CLBLL_L_X2Y140_SLICE_X1Y140_C2 = 1'b1;
  assign CLBLL_L_X2Y140_SLICE_X1Y140_C3 = 1'b1;
  assign CLBLL_L_X2Y140_SLICE_X1Y140_C4 = 1'b1;
  assign CLBLL_L_X2Y140_SLICE_X1Y140_C5 = 1'b1;
  assign CLBLL_L_X2Y140_SLICE_X1Y140_C6 = 1'b1;
  assign CLBLL_L_X2Y140_SLICE_X1Y140_D1 = 1'b1;
  assign CLBLL_L_X2Y140_SLICE_X1Y140_D2 = 1'b1;
  assign CLBLL_L_X2Y140_SLICE_X1Y140_D3 = 1'b1;
  assign CLBLL_L_X2Y140_SLICE_X1Y140_D4 = 1'b1;
  assign CLBLL_L_X2Y140_SLICE_X1Y140_D5 = 1'b1;
  assign CLBLL_L_X2Y140_SLICE_X1Y140_D6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_D1 = CLBLM_R_X13Y144_SLICE_X19Y144_AQ;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_D1 = CLBLM_L_X12Y144_SLICE_X16Y144_AQ;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_A3 = CLBLM_R_X7Y132_SLICE_X8Y132_AQ;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_T1 = 1'b1;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_A4 = CLBLM_L_X10Y132_SLICE_X12Y132_AO6;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_D1 = LIOB33_X0Y59_IOB_X0Y59_I;
  assign CLBLM_R_X103Y175_SLICE_X162Y175_B4 = 1'b1;
  assign CLBLM_R_X103Y175_SLICE_X162Y175_B6 = 1'b1;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_B1 = 1'b1;
  assign RIOB33_X105Y181_IOB_X1Y182_O = CLBLM_R_X11Y141_SLICE_X14Y141_CO6;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_C4 = CLBLM_L_X12Y136_SLICE_X17Y136_A5Q;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_C5 = CLBLM_L_X12Y141_SLICE_X17Y141_BO5;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_C6 = CLBLM_L_X12Y141_SLICE_X17Y141_DO6;
  assign CLBLM_R_X103Y175_SLICE_X162Y175_C3 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_A1 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_A3 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_A4 = CLBLM_L_X12Y140_SLICE_X16Y140_AQ;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_A5 = CLBLM_R_X7Y144_SLICE_X9Y144_AQ;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_A6 = CLBLM_L_X10Y144_SLICE_X12Y144_AO5;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_C1 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_B1 = 1'b1;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_C2 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_B2 = CLBLM_R_X7Y142_SLICE_X9Y142_BQ;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_B3 = CLBLL_L_X4Y137_SLICE_X4Y137_AQ;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_B5 = CLBLM_R_X11Y141_SLICE_X14Y141_AQ;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_B6 = CLBLM_L_X8Y143_SLICE_X10Y143_DO6;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_A1 = CLBLM_R_X7Y133_SLICE_X8Y133_AQ;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_A2 = CLBLM_R_X11Y138_SLICE_X15Y138_BQ;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_A3 = CLBLM_R_X5Y132_SLICE_X7Y132_AQ;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_A6 = CLBLM_R_X5Y132_SLICE_X7Y132_CO6;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_C1 = CLBLM_R_X3Y143_SLICE_X2Y143_AO5;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_C2 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_C3 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_B1 = CLBLL_L_X4Y133_SLICE_X4Y133_AQ;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_B2 = CLBLM_R_X5Y134_SLICE_X7Y134_DO6;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_B3 = CLBLM_R_X5Y132_SLICE_X7Y132_AQ;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_B4 = CLBLM_R_X7Y132_SLICE_X8Y132_CQ;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_B5 = CLBLM_R_X7Y132_SLICE_X8Y132_AQ;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_B6 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_D2 = CLBLM_L_X12Y143_SLICE_X17Y143_BQ;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_C1 = CLBLM_R_X7Y132_SLICE_X8Y132_AQ;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_C2 = CLBLM_R_X5Y132_SLICE_X7Y132_AQ;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_C3 = CLBLL_L_X4Y133_SLICE_X4Y133_AQ;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_C4 = CLBLM_R_X7Y132_SLICE_X8Y132_CQ;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_C5 = CLBLM_R_X5Y132_SLICE_X7Y132_DO6;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_C6 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_D3 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_D4 = CLBLM_L_X8Y141_SLICE_X10Y141_BQ;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_A4 = CLBLM_L_X10Y144_SLICE_X13Y144_AQ;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_A2 = CLBLM_R_X5Y135_SLICE_X7Y135_A5Q;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_A3 = CLBLM_R_X7Y142_SLICE_X8Y142_AQ;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_D5 = CLBLM_R_X13Y140_SLICE_X19Y140_AQ;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_D1 = CLBLM_R_X5Y136_SLICE_X7Y136_DO6;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_D2 = CLBLM_R_X5Y133_SLICE_X7Y133_CO6;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_D3 = 1'b1;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_D4 = CLBLM_R_X7Y133_SLICE_X9Y133_DO6;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_D6 = CLBLM_L_X12Y140_SLICE_X16Y140_CQ;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_D5 = 1'b1;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_D6 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_A6 = CLBLM_L_X12Y144_SLICE_X17Y144_AQ;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_B1 = CLBLM_R_X7Y143_SLICE_X8Y143_DO6;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_B2 = CLBLM_R_X7Y142_SLICE_X9Y142_DO6;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_B3 = CLBLM_L_X8Y141_SLICE_X11Y141_BQ;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_A1 = CLBLL_L_X4Y133_SLICE_X4Y133_AQ;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_A2 = CLBLM_R_X5Y132_SLICE_X7Y132_DO6;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_A1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_A2 = CLBLM_R_X3Y143_SLICE_X2Y143_AO6;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_A5 = CLBLM_R_X5Y132_SLICE_X7Y132_AQ;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_A6 = CLBLM_R_X7Y132_SLICE_X8Y132_CQ;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_A3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_A4 = CLBLM_R_X3Y138_SLICE_X2Y138_AO5;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_A5 = LIOB33_X0Y61_IOB_X0Y61_I;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_A6 = LIOB33_X0Y71_IOB_X0Y71_I;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_B2 = 1'b1;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_B3 = 1'b1;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_B4 = 1'b1;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_B5 = 1'b1;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_B6 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_B1 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_B2 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_B3 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_B4 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_B5 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_B6 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_C1 = 1'b1;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_C5 = 1'b1;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_C6 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_C2 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_C3 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_C4 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_C5 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_C6 = 1'b1;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_C3 = 1'b1;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_C4 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_D1 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_D2 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_D3 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_D4 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_D5 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_D6 = 1'b1;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_D1 = 1'b1;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_D2 = 1'b1;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_D3 = 1'b1;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_D4 = 1'b1;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_D5 = 1'b1;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_D6 = 1'b1;
  assign LIOB33_X0Y157_IOB_X0Y157_O = RIOB33_X105Y115_IOB_X1Y115_I;
  assign LIOB33_X0Y157_IOB_X0Y158_O = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_A1 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_A2 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_A3 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_A4 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_A5 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_A6 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_B1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_B2 = CLBLM_R_X3Y143_SLICE_X2Y143_AO6;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_B3 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_B4 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_B5 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_B6 = 1'b1;
  assign LIOI3_X0Y165_OLOGIC_X0Y166_T1 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_C1 = CLBLL_L_X2Y141_SLICE_X1Y141_AO6;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_C2 = LIOB33_X0Y53_IOB_X0Y54_I;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_C3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_C4 = CLBLM_R_X3Y143_SLICE_X2Y143_AO6;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_C5 = LIOB33_X0Y69_IOB_X0Y70_I;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_C6 = CLBLL_L_X2Y141_SLICE_X1Y141_BO6;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_B5 = CLBLM_R_X13Y144_SLICE_X18Y144_AQ;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_D1 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_D2 = CLBLL_L_X2Y141_SLICE_X0Y141_AO6;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_D3 = LIOB33_X0Y55_IOB_X0Y55_I;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_D4 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_B6 = CLBLM_L_X12Y143_SLICE_X17Y143_BQ;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_D5 = CLBLL_L_X2Y141_SLICE_X1Y141_BO5;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_D6 = CLBLM_L_X10Y140_SLICE_X13Y140_C5Q;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_C4 = CLBLM_L_X12Y142_SLICE_X16Y142_AQ;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_C5 = CLBLM_R_X13Y140_SLICE_X18Y140_BQ;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_C6 = CLBLM_L_X12Y142_SLICE_X16Y142_BQ;
  assign RIOI3_X105Y133_ILOGIC_X1Y134_D = RIOB33_X105Y133_IOB_X1Y134_I;
  assign RIOI3_X105Y133_ILOGIC_X1Y133_D = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_A1 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_A2 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_A3 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_A4 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_A5 = 1'b1;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_A6 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_B1 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_B2 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_B3 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_B4 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_B5 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_B6 = 1'b1;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_D5 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_A1 = CLBLM_L_X10Y140_SLICE_X13Y140_C5Q;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_A2 = CLBLM_R_X7Y143_SLICE_X9Y143_BQ;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_A4 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_A5 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_A6 = CLBLM_L_X10Y144_SLICE_X12Y144_AO5;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_C1 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_C2 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_B1 = CLBLM_R_X3Y137_SLICE_X3Y137_CQ;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_B2 = CLBLM_L_X8Y142_SLICE_X11Y142_CQ;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_B4 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_B5 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_B6 = CLBLM_L_X10Y144_SLICE_X12Y144_AO5;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_D1 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_D2 = 1'b1;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_A1 = CLBLM_R_X5Y135_SLICE_X7Y135_A5Q;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_A2 = CLBLM_R_X5Y135_SLICE_X6Y135_D5Q;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_A3 = CLBLM_R_X3Y137_SLICE_X3Y137_BQ;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_A4 = CLBLM_R_X5Y136_SLICE_X6Y136_DQ;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_A5 = CLBLM_R_X5Y133_SLICE_X6Y133_DO6;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_A6 = CLBLM_R_X5Y134_SLICE_X7Y134_AO6;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_C1 = CLBLM_L_X8Y143_SLICE_X10Y143_DO5;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_C2 = CLBLM_R_X7Y143_SLICE_X9Y143_CQ;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_C3 = CLBLM_R_X7Y135_SLICE_X8Y135_AQ;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_B1 = CLBLM_R_X5Y137_SLICE_X7Y137_B5Q;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_B2 = CLBLM_R_X5Y135_SLICE_X6Y135_DQ;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_B3 = CLBLM_R_X3Y137_SLICE_X3Y137_BQ;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_B4 = CLBLM_R_X5Y135_SLICE_X6Y135_D5Q;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_B5 = CLBLM_R_X5Y136_SLICE_X6Y136_DQ;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_B6 = CLBLM_L_X8Y140_SLICE_X11Y140_A5Q;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_D1 = 1'b1;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_C1 = CLBLM_R_X5Y137_SLICE_X7Y137_C5Q;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_C2 = CLBLL_L_X4Y137_SLICE_X4Y137_A5Q;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_C3 = 1'b1;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_C4 = CLBLM_R_X5Y135_SLICE_X7Y135_A5Q;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_C5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_C6 = CLBLM_R_X5Y133_SLICE_X7Y133_BO6;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_D3 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_D4 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_A1 = CLBLM_L_X8Y143_SLICE_X10Y143_DO6;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_A2 = CLBLM_L_X12Y144_SLICE_X17Y144_AQ;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_A3 = CLBLM_R_X7Y143_SLICE_X8Y143_AQ;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_A5 = CLBLM_R_X7Y143_SLICE_X9Y143_AQ;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_A6 = 1'b1;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_D1 = CLBLM_R_X5Y136_SLICE_X7Y136_DO6;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_D2 = CLBLM_R_X5Y135_SLICE_X7Y135_A5Q;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_D3 = CLBLM_R_X5Y133_SLICE_X6Y133_BO6;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_D4 = 1'b1;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_D5 = 1'b1;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_D6 = CLBLM_R_X7Y133_SLICE_X9Y133_DO6;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_B3 = CLBLM_L_X10Y142_SLICE_X12Y142_BQ;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_B4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_B5 = CLBLM_R_X7Y143_SLICE_X8Y143_A5Q;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_B6 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_B1 = CLBLM_R_X7Y133_SLICE_X8Y133_DO6;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_A1 = CLBLM_R_X5Y135_SLICE_X6Y135_DQ;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_A2 = CLBLM_R_X5Y136_SLICE_X6Y136_DQ;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_A3 = CLBLM_R_X5Y137_SLICE_X7Y137_C5Q;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_A4 = CLBLM_R_X5Y135_SLICE_X6Y135_D5Q;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_A5 = CLBLM_R_X3Y137_SLICE_X3Y137_BQ;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_A6 = 1'b1;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_C1 = CLBLM_L_X10Y144_SLICE_X12Y144_AO6;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_C2 = CLBLM_L_X10Y143_SLICE_X12Y143_CQ;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_B1 = CLBLM_L_X8Y140_SLICE_X11Y140_A5Q;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_B2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_B3 = CLBLM_R_X5Y137_SLICE_X7Y137_B5Q;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_B4 = CLBLM_R_X5Y135_SLICE_X6Y135_D5Q;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_B5 = CLBLM_R_X5Y133_SLICE_X6Y133_AO6;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_B6 = CLBLL_L_X4Y137_SLICE_X4Y137_A5Q;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_C3 = CLBLM_L_X10Y143_SLICE_X13Y143_BO6;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_D1 = CLBLM_R_X3Y143_SLICE_X2Y143_AO5;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_C1 = CLBLL_L_X4Y141_SLICE_X4Y141_DO6;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_C2 = CLBLM_R_X3Y136_SLICE_X3Y136_CQ;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_C3 = CLBLM_L_X12Y135_SLICE_X17Y135_CQ;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_C4 = CLBLM_R_X3Y140_SLICE_X2Y140_DO6;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_C5 = CLBLM_R_X5Y142_SLICE_X6Y142_CO6;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_C6 = CLBLM_R_X5Y134_SLICE_X6Y134_CO5;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_D2 = CLBLM_R_X7Y143_SLICE_X8Y143_AQ;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_D3 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_D4 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_D5 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_D6 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_D1 = CLBLM_R_X5Y137_SLICE_X7Y137_C5Q;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_D2 = 1'b1;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_D3 = CLBLM_R_X5Y135_SLICE_X6Y135_DQ;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_D4 = 1'b1;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_D5 = 1'b1;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_D6 = 1'b1;
  assign LIOI3_X0Y165_OLOGIC_X0Y165_D1 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_D3 = CLBLM_L_X10Y144_SLICE_X13Y144_DO6;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_D4 = CLBLM_L_X10Y145_SLICE_X12Y145_BO6;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_D6 = CLBLM_R_X11Y144_SLICE_X15Y144_BQ;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_C6 = 1'b1;
  assign LIOI3_X0Y161_OLOGIC_X0Y162_D1 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign LIOI3_X0Y161_OLOGIC_X0Y162_T1 = 1'b1;
  assign LIOI3_X0Y101_OLOGIC_X0Y102_D1 = CLBLM_R_X3Y133_SLICE_X2Y133_AO5;
  assign LIOI3_X0Y161_OLOGIC_X0Y161_D1 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_T1 = 1'b1;
  assign LIOI3_X0Y101_OLOGIC_X0Y102_T1 = 1'b1;
  assign LIOI3_X0Y161_OLOGIC_X0Y161_T1 = 1'b1;
  assign LIOI3_X0Y101_OLOGIC_X0Y101_D1 = CLBLM_R_X3Y133_SLICE_X2Y133_AO6;
  assign LIOI3_X0Y101_OLOGIC_X0Y101_T1 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_A1 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_A2 = CLBLM_L_X10Y144_SLICE_X12Y144_AO5;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_A3 = CLBLM_R_X7Y131_SLICE_X9Y131_BQ;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_A4 = CLBLM_R_X7Y143_SLICE_X9Y143_AQ;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_A5 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_B1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_B2 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_B3 = CLBLM_R_X11Y136_SLICE_X14Y136_DQ;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_B6 = CLBLM_R_X7Y144_SLICE_X8Y144_CQ;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_A1 = CLBLM_R_X5Y137_SLICE_X7Y137_B5Q;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_A2 = CLBLM_L_X8Y140_SLICE_X11Y140_A5Q;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_A3 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_A5 = CLBLL_L_X4Y137_SLICE_X4Y137_A5Q;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_A6 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_C1 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_C2 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_C3 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_B1 = CLBLM_R_X5Y136_SLICE_X6Y136_BQ;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_B2 = CLBLM_R_X5Y134_SLICE_X7Y134_BQ;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_B4 = CLBLM_R_X7Y135_SLICE_X8Y135_DO6;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_B5 = CLBLM_L_X8Y135_SLICE_X11Y135_AQ;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_B6 = CLBLM_R_X5Y135_SLICE_X7Y135_CO6;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_D1 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_C1 = CLBLM_R_X5Y137_SLICE_X7Y137_C5Q;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_C2 = CLBLM_R_X5Y134_SLICE_X7Y134_CQ;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_C3 = CLBLM_R_X7Y139_SLICE_X8Y139_A5Q;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_C5 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_C6 = CLBLL_L_X4Y133_SLICE_X5Y133_BO6;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_D3 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_D4 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_A1 = CLBLM_R_X7Y144_SLICE_X8Y144_AQ;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_A2 = CLBLM_R_X7Y144_SLICE_X8Y144_BQ;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_A3 = CLBLM_L_X8Y144_SLICE_X11Y144_BO6;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_A4 = CLBLM_R_X7Y143_SLICE_X9Y143_BQ;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_D1 = CLBLM_L_X8Y140_SLICE_X11Y140_A5Q;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_D2 = CLBLM_R_X3Y139_SLICE_X3Y139_BO6;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_D3 = CLBLM_R_X5Y135_SLICE_X7Y135_A5Q;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_D4 = CLBLM_R_X5Y134_SLICE_X7Y134_AO5;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_D5 = CLBLM_R_X5Y133_SLICE_X6Y133_AO5;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_D6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_A6 = CLBLM_L_X8Y140_SLICE_X10Y140_CQ;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_B1 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_B2 = CLBLM_R_X7Y144_SLICE_X8Y144_BQ;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_B3 = CLBLM_L_X8Y143_SLICE_X10Y143_BQ;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_B4 = CLBLM_R_X7Y143_SLICE_X9Y143_BQ;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_A1 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_A2 = CLBLM_L_X10Y145_SLICE_X12Y145_AQ;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_A3 = CLBLM_R_X5Y134_SLICE_X6Y134_AQ;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_A4 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_A6 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_C1 = CLBLM_R_X11Y136_SLICE_X14Y136_DQ;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_C2 = CLBLM_R_X7Y144_SLICE_X8Y144_CQ;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_AX = CLBLM_R_X5Y134_SLICE_X6Y134_BO6;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_C3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_B1 = CLBLM_R_X5Y134_SLICE_X6Y134_DO6;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_B2 = CLBLM_R_X5Y137_SLICE_X7Y137_C5Q;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_B3 = CLBLM_L_X12Y134_SLICE_X17Y134_AO6;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_B5 = CLBLM_R_X5Y134_SLICE_X6Y134_A5Q;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_B6 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_D1 = CLBLM_R_X3Y143_SLICE_X2Y143_AO5;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_D2 = CLBLM_R_X7Y144_SLICE_X8Y144_CQ;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_C2 = CLBLM_R_X5Y136_SLICE_X6Y136_CQ;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_C3 = CLBLM_R_X7Y134_SLICE_X8Y134_CQ;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_C4 = CLBLM_L_X10Y145_SLICE_X12Y145_AQ;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_C5 = CLBLM_L_X12Y134_SLICE_X17Y134_AQ;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_C6 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_D3 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_D4 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_D5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_D6 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_D2 = CLBLM_R_X7Y134_SLICE_X8Y134_CQ;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_D3 = CLBLM_L_X12Y134_SLICE_X17Y134_AQ;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_D4 = CLBLM_L_X10Y145_SLICE_X12Y145_AQ;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_D5 = CLBLM_R_X5Y136_SLICE_X6Y136_CQ;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_D6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X37Y138_SLICE_X57Y138_B5 = 1'b1;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X37Y138_SLICE_X57Y138_B6 = 1'b1;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_A4 = CLBLM_R_X11Y134_SLICE_X14Y134_AQ;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_A5 = CLBLM_L_X8Y136_SLICE_X10Y136_CQ;
  assign RIOI3_X105Y145_ILOGIC_X1Y146_D = RIOB33_X105Y145_IOB_X1Y146_I;
  assign RIOI3_X105Y145_ILOGIC_X1Y145_D = RIOB33_X105Y145_IOB_X1Y145_I;
  assign CLBLM_R_X37Y138_SLICE_X57Y138_C3 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y64_D = LIOB33_X0Y63_IOB_X0Y64_I;
  assign CLBLM_R_X37Y138_SLICE_X57Y138_C5 = 1'b1;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_B1 = RIOB33_X105Y125_IOB_X1Y126_I;
  assign LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y63_D = LIOB33_X0Y63_IOB_X0Y63_I;
  assign CLBLM_R_X37Y138_SLICE_X57Y138_C6 = 1'b1;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_D4 = CLBLM_R_X11Y139_SLICE_X15Y139_CQ;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_D5 = 1'b1;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_D6 = CLBLM_L_X10Y139_SLICE_X13Y139_AQ;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_C4 = CLBLL_L_X4Y134_SLICE_X5Y134_CQ;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_C5 = CLBLM_R_X7Y143_SLICE_X8Y143_CQ;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_C6 = CLBLL_L_X4Y143_SLICE_X4Y143_AO5;
  assign CLBLM_R_X37Y138_SLICE_X57Y138_D2 = 1'b1;
  assign CLBLM_R_X37Y138_SLICE_X57Y138_D3 = 1'b1;
  assign CLBLM_R_X37Y138_SLICE_X57Y138_D4 = 1'b1;
  assign CLBLM_R_X37Y138_SLICE_X57Y138_D5 = 1'b1;
  assign CLBLM_R_X37Y138_SLICE_X57Y138_D6 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_D1 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_D2 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_D5 = CLBLL_L_X4Y143_SLICE_X5Y143_BO5;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_D6 = CLBLL_L_X4Y138_SLICE_X4Y138_BQ;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_D1 = CLBLL_L_X4Y134_SLICE_X4Y134_AQ;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_D5 = CLBLM_L_X8Y138_SLICE_X10Y138_AQ;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_A1 = CLBLM_R_X5Y135_SLICE_X7Y135_BO5;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_A2 = CLBLM_R_X7Y135_SLICE_X8Y135_DO6;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_A3 = CLBLM_R_X5Y135_SLICE_X7Y135_AQ;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_A4 = 1'b1;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_A6 = CLBLM_R_X7Y139_SLICE_X9Y139_AQ;
  assign LIOB33_X0Y163_IOB_X0Y163_O = RIOB33_X105Y109_IOB_X1Y110_I;
  assign LIOB33_X0Y163_IOB_X0Y164_O = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_AX = CLBLM_R_X5Y135_SLICE_X7Y135_BO6;
  assign CLBLM_R_X37Y138_SLICE_X56Y138_B2 = 1'b1;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_B1 = CLBLM_L_X8Y134_SLICE_X11Y134_DQ;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_B2 = CLBLM_R_X7Y135_SLICE_X8Y135_BQ;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_B4 = CLBLM_R_X7Y134_SLICE_X8Y134_BQ;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_B5 = CLBLM_R_X5Y137_SLICE_X7Y137_AQ;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_B6 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_D4 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_D5 = CLBLM_L_X8Y138_SLICE_X10Y138_BQ;
  assign CLBLM_R_X37Y138_SLICE_X56Y138_B3 = 1'b1;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_C1 = CLBLM_R_X5Y137_SLICE_X7Y137_AQ;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_C2 = CLBLM_R_X7Y135_SLICE_X8Y135_BQ;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_C3 = 1'b1;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_C4 = CLBLM_R_X7Y134_SLICE_X8Y134_BQ;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_C5 = CLBLM_R_X5Y135_SLICE_X7Y135_AQ;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_C6 = 1'b1;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_A2 = CLBLM_R_X11Y135_SLICE_X14Y135_BQ;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_D6 = 1'b1;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_A3 = CLBLM_L_X8Y135_SLICE_X10Y135_AQ;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_D1 = CLBLM_R_X5Y137_SLICE_X7Y137_AQ;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_D2 = CLBLM_R_X7Y135_SLICE_X8Y135_BQ;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_D3 = CLBLM_R_X5Y134_SLICE_X7Y134_BQ;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_D4 = CLBLM_R_X5Y136_SLICE_X6Y136_BQ;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_D5 = CLBLM_R_X5Y135_SLICE_X7Y135_AQ;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_D6 = CLBLM_R_X7Y134_SLICE_X8Y134_BQ;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_A4 = CLBLM_L_X10Y137_SLICE_X13Y137_CO6;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_A5 = CLBLM_L_X8Y138_SLICE_X10Y138_AQ;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_A1 = CLBLM_R_X5Y135_SLICE_X6Y135_AQ;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_A2 = CLBLM_L_X12Y136_SLICE_X17Y136_AQ;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_A3 = CLBLM_R_X5Y134_SLICE_X6Y134_CO6;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_A4 = CLBLM_R_X5Y134_SLICE_X6Y134_BO5;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_A5 = CLBLM_R_X5Y135_SLICE_X6Y135_BQ;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_B5 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_B1 = 1'b1;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_B2 = CLBLM_R_X5Y135_SLICE_X6Y135_BQ;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_B3 = CLBLM_R_X5Y134_SLICE_X6Y134_CO6;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_B4 = CLBLM_R_X5Y134_SLICE_X6Y134_BO5;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_B5 = CLBLM_R_X7Y132_SLICE_X8Y132_BQ;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_B6 = 1'b1;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_C2 = CLBLM_R_X5Y135_SLICE_X6Y135_CQ;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_C3 = CLBLM_R_X5Y135_SLICE_X6Y135_AQ;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_C4 = CLBLM_L_X8Y138_SLICE_X10Y138_AQ;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_C5 = CLBLM_R_X7Y135_SLICE_X9Y135_DO6;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_C6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_B1 = 1'b1;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_B2 = CLBLM_L_X8Y135_SLICE_X10Y135_BQ;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_B3 = CLBLM_L_X8Y135_SLICE_X10Y135_AQ;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_D1 = CLBLM_R_X5Y135_SLICE_X7Y135_AQ;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_D2 = CLBLM_R_X5Y136_SLICE_X6Y136_BQ;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_D3 = CLBLM_R_X5Y136_SLICE_X6Y136_D5Q;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_D4 = CLBLM_R_X5Y139_SLICE_X6Y139_BQ;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_D6 = 1'b1;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_B5 = 1'b1;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_C4 = CLBLM_L_X8Y143_SLICE_X10Y143_BQ;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_C5 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_C6 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_D6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_C4 = CLBLM_L_X8Y135_SLICE_X11Y135_CQ;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_C5 = CLBLM_R_X11Y136_SLICE_X14Y136_DQ;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_C4 = CLBLM_R_X3Y143_SLICE_X3Y143_AO5;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_D1 = CLBLM_L_X12Y139_SLICE_X17Y139_DO5;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_C5 = CLBLL_L_X4Y143_SLICE_X5Y143_BO5;
  assign RIOI3_X105Y183_OLOGIC_X1Y183_D1 = CLBLM_R_X11Y141_SLICE_X14Y141_CO5;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_C6 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_D1 = CLBLM_R_X5Y141_SLICE_X6Y141_BQ;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_T1 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_D2 = CLBLL_L_X4Y139_SLICE_X5Y139_DO6;
  assign RIOI3_X105Y183_OLOGIC_X1Y183_T1 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_D3 = CLBLL_L_X4Y140_SLICE_X5Y140_AO6;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_D4 = CLBLL_L_X4Y141_SLICE_X5Y141_CO6;
  assign LIOB33_X0Y165_IOB_X0Y166_O = RIOB33_X105Y113_IOB_X1Y113_I;
  assign LIOB33_X0Y165_IOB_X0Y165_O = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_D5 = CLBLM_R_X3Y142_SLICE_X2Y142_AO6;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_A1 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_A2 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_A3 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_A4 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_A5 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_A6 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_B1 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_B2 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_B3 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_B4 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_B5 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_B6 = 1'b1;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_A1 = CLBLM_R_X7Y138_SLICE_X8Y138_CQ;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_A2 = CLBLM_R_X5Y135_SLICE_X7Y135_DO6;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_A3 = CLBLM_R_X5Y136_SLICE_X7Y136_AQ;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_A4 = CLBLM_R_X7Y135_SLICE_X8Y135_DO5;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_A5 = CLBLM_R_X5Y137_SLICE_X6Y137_CQ;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_C1 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_C2 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_C3 = 1'b1;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_B1 = CLBLM_R_X3Y137_SLICE_X2Y137_BQ;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_B2 = CLBLM_R_X5Y136_SLICE_X7Y136_BQ;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_B3 = 1'b1;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_B4 = CLBLM_R_X7Y139_SLICE_X9Y139_AQ;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_D1 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_D2 = 1'b1;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_C1 = CLBLM_R_X7Y139_SLICE_X8Y139_AQ;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_C2 = CLBLM_R_X5Y136_SLICE_X7Y136_CQ;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_C3 = CLBLM_R_X7Y134_SLICE_X8Y134_CQ;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_C4 = CLBLM_L_X10Y139_SLICE_X13Y139_B5Q;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_C6 = CLBLM_L_X12Y134_SLICE_X17Y134_AO6;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_D3 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_D4 = 1'b1;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_A1 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_A2 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_A3 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_A4 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_A5 = 1'b1;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_D1 = CLBLM_R_X5Y140_SLICE_X6Y140_AO6;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_D2 = CLBLL_L_X4Y139_SLICE_X4Y139_BO6;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_D3 = CLBLM_R_X3Y137_SLICE_X3Y137_DO6;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_D4 = CLBLM_R_X3Y140_SLICE_X2Y140_DO6;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_D5 = CLBLM_R_X5Y141_SLICE_X7Y141_DO6;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_D6 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_A4 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_A6 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_AX = CLBLM_L_X10Y146_SLICE_X12Y146_AO6;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_B1 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_B2 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_B3 = 1'b1;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_A2 = CLBLM_R_X5Y138_SLICE_X6Y138_CQ;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_A3 = CLBLM_R_X5Y136_SLICE_X6Y136_AQ;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_A4 = CLBLM_L_X8Y143_SLICE_X10Y143_DO5;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_A5 = 1'b1;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_A6 = CLBLL_L_X4Y135_SLICE_X5Y135_CQ;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_C1 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_C2 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_C3 = 1'b1;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_B1 = CLBLM_R_X5Y141_SLICE_X6Y141_CQ;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_B2 = CLBLM_R_X5Y136_SLICE_X6Y136_BQ;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_B3 = CLBLM_R_X5Y135_SLICE_X7Y135_CO6;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_B4 = CLBLM_R_X7Y135_SLICE_X8Y135_DO5;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_B5 = 1'b1;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_D1 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_D2 = 1'b1;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_C1 = CLBLM_R_X5Y135_SLICE_X6Y135_BQ;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_C2 = CLBLM_R_X5Y135_SLICE_X6Y135_AQ;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_C3 = CLBLM_R_X7Y139_SLICE_X9Y139_A5Q;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_C4 = CLBLM_R_X5Y134_SLICE_X6Y134_A5Q;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_C6 = CLBLL_L_X4Y138_SLICE_X5Y138_A5Q;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_D3 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_D4 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_D5 = 1'b1;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_B1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_T1 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_B2 = 1'b1;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_D1 = CLBLL_L_X4Y136_SLICE_X5Y136_BQ;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_D2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_D3 = RIOB33_X105Y127_IOB_X1Y127_I;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_D4 = CLBLM_L_X10Y138_SLICE_X13Y138_CQ;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_D5 = CLBLM_R_X5Y137_SLICE_X6Y137_CQ;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_D6 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_B3 = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_T1 = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_D1 = LIOB33_X0Y57_IOB_X0Y58_I;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_C5 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_C6 = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_T1 = 1'b1;
  assign CLBLM_R_X103Y140_SLICE_X163Y140_A1 = RIOB33_X105Y141_IOB_X1Y141_I;
  assign CLBLM_R_X103Y140_SLICE_X163Y140_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X103Y140_SLICE_X163Y140_A3 = RIOB33_X105Y137_IOB_X1Y138_I;
  assign CLBLM_R_X103Y140_SLICE_X163Y140_A4 = RIOB33_X105Y139_IOB_X1Y139_I;
  assign CLBLM_R_X103Y140_SLICE_X163Y140_A5 = RIOB33_X105Y139_IOB_X1Y140_I;
  assign CLBLM_R_X103Y140_SLICE_X163Y140_A6 = 1'b1;
  assign CLBLM_R_X103Y140_SLICE_X163Y140_B1 = 1'b1;
  assign CLBLM_R_X103Y140_SLICE_X163Y140_B2 = 1'b1;
  assign CLBLM_R_X103Y140_SLICE_X163Y140_B3 = 1'b1;
  assign CLBLM_R_X103Y140_SLICE_X163Y140_B4 = 1'b1;
  assign CLBLM_R_X103Y140_SLICE_X163Y140_B5 = 1'b1;
  assign CLBLM_R_X103Y140_SLICE_X163Y140_B6 = 1'b1;
  assign RIOI3_X105Y147_ILOGIC_X1Y148_D = RIOB33_X105Y147_IOB_X1Y148_I;
  assign RIOI3_X105Y147_ILOGIC_X1Y147_D = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X103Y140_SLICE_X163Y140_C1 = 1'b1;
  assign CLBLM_R_X103Y140_SLICE_X163Y140_C2 = 1'b1;
  assign CLBLM_R_X103Y140_SLICE_X163Y140_C3 = 1'b1;
  assign CLBLM_R_X103Y140_SLICE_X163Y140_C4 = 1'b1;
  assign CLBLM_R_X103Y140_SLICE_X163Y140_C5 = 1'b1;
  assign CLBLM_R_X103Y140_SLICE_X163Y140_C6 = 1'b1;
  assign LIOB33_X0Y167_IOB_X0Y168_O = RIOB33_X105Y123_IOB_X1Y123_I;
  assign LIOB33_X0Y167_IOB_X0Y167_O = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLM_R_X103Y140_SLICE_X163Y140_D1 = 1'b1;
  assign CLBLM_R_X103Y140_SLICE_X163Y140_D2 = 1'b1;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_C4 = 1'b1;
  assign CLBLM_R_X103Y140_SLICE_X163Y140_D3 = 1'b1;
  assign CLBLM_R_X103Y140_SLICE_X163Y140_D4 = 1'b1;
  assign CLBLM_R_X103Y140_SLICE_X163Y140_D5 = 1'b1;
  assign CLBLM_R_X103Y140_SLICE_X163Y140_D6 = 1'b1;
  assign CLBLM_R_X103Y140_SLICE_X162Y140_A1 = 1'b1;
  assign CLBLM_R_X103Y140_SLICE_X162Y140_A2 = 1'b1;
  assign CLBLM_R_X103Y140_SLICE_X162Y140_A3 = 1'b1;
  assign CLBLM_R_X103Y140_SLICE_X162Y140_A4 = 1'b1;
  assign CLBLM_R_X103Y140_SLICE_X162Y140_A5 = 1'b1;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_C4 = CLBLM_L_X12Y143_SLICE_X17Y143_BQ;
  assign CLBLM_R_X103Y140_SLICE_X162Y140_A6 = 1'b1;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_C5 = CLBLM_R_X13Y141_SLICE_X19Y141_CO6;
  assign CLBLM_R_X103Y140_SLICE_X162Y140_B1 = 1'b1;
  assign CLBLM_R_X103Y140_SLICE_X162Y140_B2 = 1'b1;
  assign CLBLM_R_X103Y140_SLICE_X162Y140_B3 = 1'b1;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_C5 = 1'b1;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_C6 = 1'b1;
  assign CLBLM_R_X103Y140_SLICE_X162Y140_B4 = 1'b1;
  assign CLBLM_R_X103Y140_SLICE_X162Y140_B5 = 1'b1;
  assign CLBLM_R_X103Y140_SLICE_X162Y140_B6 = 1'b1;
  assign CLBLM_R_X103Y140_SLICE_X162Y140_C1 = 1'b1;
  assign CLBLM_R_X103Y140_SLICE_X162Y140_C2 = 1'b1;
  assign CLBLM_R_X103Y140_SLICE_X162Y140_C3 = 1'b1;
  assign CLBLM_R_X103Y140_SLICE_X162Y140_C4 = 1'b1;
  assign CLBLM_R_X103Y140_SLICE_X162Y140_C5 = 1'b1;
  assign CLBLM_R_X103Y140_SLICE_X162Y140_C6 = 1'b1;
  assign CLBLM_R_X103Y140_SLICE_X162Y140_D1 = 1'b1;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_C6 = 1'b1;
  assign CLBLM_R_X103Y140_SLICE_X162Y140_D2 = 1'b1;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_A1 = CLBLM_R_X7Y134_SLICE_X8Y134_BQ;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_A3 = CLBLM_R_X5Y137_SLICE_X7Y137_AQ;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_A4 = CLBLM_R_X7Y135_SLICE_X8Y135_DO5;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_A5 = CLBLM_R_X5Y137_SLICE_X6Y137_AQ;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_A6 = CLBLM_R_X7Y135_SLICE_X8Y135_BQ;
  assign CLBLM_R_X103Y140_SLICE_X162Y140_D3 = 1'b1;
  assign CLBLM_R_X103Y140_SLICE_X162Y140_D4 = 1'b1;
  assign CLBLM_R_X103Y140_SLICE_X162Y140_D5 = 1'b1;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_B2 = CLBLM_R_X5Y137_SLICE_X7Y137_BQ;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_B3 = CLBLM_R_X7Y142_SLICE_X8Y142_AQ;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_B4 = CLBLM_R_X5Y136_SLICE_X7Y136_AQ;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_B6 = 1'b1;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_C2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_C3 = CLBLM_L_X8Y139_SLICE_X11Y139_BQ;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_C4 = CLBLM_R_X5Y138_SLICE_X7Y138_BQ;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_C5 = CLBLM_R_X5Y134_SLICE_X7Y134_BQ;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_C6 = 1'b1;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_D2 = CLBLM_L_X12Y140_SLICE_X17Y140_AQ;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_D1 = CLBLM_R_X5Y136_SLICE_X7Y136_AQ;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_D2 = CLBLM_R_X5Y134_SLICE_X7Y134_BQ;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_D3 = CLBLL_L_X4Y137_SLICE_X4Y137_BQ;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_D4 = CLBLM_R_X5Y137_SLICE_X6Y137_CQ;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_D5 = CLBLM_R_X5Y135_SLICE_X7Y135_CO5;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_D6 = CLBLM_R_X5Y136_SLICE_X6Y136_BQ;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_D5 = CLBLM_R_X13Y141_SLICE_X18Y141_CO5;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_A5 = CLBLM_L_X8Y144_SLICE_X11Y144_AQ;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_A1 = CLBLL_L_X4Y137_SLICE_X4Y137_CQ;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_A2 = CLBLM_L_X12Y135_SLICE_X17Y135_AQ;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_A3 = CLBLM_R_X5Y137_SLICE_X6Y137_AQ;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_A4 = CLBLM_R_X5Y137_SLICE_X6Y137_CQ;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_A5 = CLBLM_L_X8Y138_SLICE_X10Y138_BQ;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_A6 = CLBLM_R_X11Y144_SLICE_X14Y144_DO6;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_B1 = CLBLM_R_X7Y143_SLICE_X8Y143_A5Q;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_B3 = CLBLL_L_X4Y136_SLICE_X5Y136_CQ;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_B4 = CLBLM_R_X7Y133_SLICE_X8Y133_CQ;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_B5 = CLBLM_L_X8Y134_SLICE_X10Y134_AQ;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_B6 = CLBLM_R_X3Y138_SLICE_X3Y138_AQ;
  assign RIOI3_X105Y123_ILOGIC_X1Y124_D = RIOB33_X105Y123_IOB_X1Y124_I;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_C1 = CLBLM_R_X7Y143_SLICE_X8Y143_AQ;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_C2 = CLBLM_R_X5Y137_SLICE_X6Y137_CQ;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_C3 = CLBLM_R_X5Y135_SLICE_X7Y135_DO6;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_C4 = CLBLM_R_X7Y135_SLICE_X8Y135_DO5;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_C6 = 1'b1;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_X105Y123_ILOGIC_X1Y123_D = RIOB33_X105Y123_IOB_X1Y123_I;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_B3 = CLBLM_L_X10Y142_SLICE_X12Y142_AQ;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_D1 = CLBLM_R_X5Y135_SLICE_X6Y135_BQ;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_D2 = CLBLM_R_X5Y134_SLICE_X6Y134_DO6;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_D3 = CLBLM_R_X5Y135_SLICE_X6Y135_AQ;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_D4 = CLBLM_R_X5Y134_SLICE_X6Y134_A5Q;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_D5 = CLBLM_L_X12Y134_SLICE_X17Y134_AO6;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_D6 = CLBLL_L_X4Y138_SLICE_X5Y138_A5Q;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_A6 = CLBLM_R_X13Y141_SLICE_X18Y141_AO5;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_B6 = CLBLM_R_X5Y135_SLICE_X7Y135_A5Q;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_D4 = CLBLM_R_X11Y144_SLICE_X14Y144_AQ;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_C4 = CLBLM_L_X12Y143_SLICE_X17Y143_CO5;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_C5 = CLBLM_L_X12Y140_SLICE_X16Y140_BQ;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_C6 = CLBLM_R_X13Y143_SLICE_X18Y143_AO6;
  assign LIOB33_X0Y169_IOB_X0Y169_O = RIOB33_X105Y121_IOB_X1Y122_I;
  assign LIOB33_X0Y169_IOB_X0Y170_O = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_A6 = 1'b1;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_AX = CLBLM_R_X11Y144_SLICE_X14Y144_BO6;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_A1 = 1'b1;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_A2 = CLBLM_R_X7Y144_SLICE_X9Y144_BO6;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_A3 = CLBLM_R_X5Y138_SLICE_X7Y138_AQ;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_A4 = CLBLM_L_X8Y137_SLICE_X10Y137_AQ;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_A6 = CLBLM_R_X7Y134_SLICE_X8Y134_AQ;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_B1 = CLBLM_L_X10Y145_SLICE_X12Y145_BO5;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_B1 = CLBLM_L_X10Y139_SLICE_X13Y139_B5Q;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_B2 = CLBLM_R_X5Y138_SLICE_X7Y138_BQ;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_B4 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_B5 = CLBLM_L_X12Y134_SLICE_X17Y134_AO6;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_B6 = CLBLM_R_X7Y143_SLICE_X8Y143_A5Q;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_B2 = CLBLM_L_X10Y144_SLICE_X12Y144_CO6;
  assign RIOI3_X105Y141_ILOGIC_X1Y141_D = RIOB33_X105Y141_IOB_X1Y141_I;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_C2 = CLBLM_R_X5Y138_SLICE_X7Y138_CQ;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_C3 = CLBLM_L_X12Y138_SLICE_X16Y138_CQ;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_C4 = CLBLL_L_X4Y142_SLICE_X5Y142_DO6;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_C6 = CLBLL_L_X4Y138_SLICE_X5Y138_CO5;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_D1 = CLBLM_R_X5Y137_SLICE_X6Y137_AQ;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_D2 = 1'b1;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_D3 = 1'b1;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_D4 = CLBLM_R_X11Y134_SLICE_X15Y134_AQ;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_D5 = CLBLM_R_X5Y143_SLICE_X6Y143_AO5;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_D6 = CLBLL_L_X4Y143_SLICE_X5Y143_AO5;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_T1 = 1'b1;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_A1 = CLBLM_L_X8Y143_SLICE_X10Y143_DO5;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_A2 = 1'b1;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_A3 = CLBLM_R_X5Y138_SLICE_X6Y138_AQ;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_A4 = CLBLM_L_X10Y137_SLICE_X13Y137_BQ;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_A6 = CLBLM_R_X11Y138_SLICE_X15Y138_CQ;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_B1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_B2 = CLBLL_L_X4Y138_SLICE_X5Y138_A5Q;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_B3 = CLBLM_L_X8Y138_SLICE_X10Y138_AQ;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_B4 = 1'b1;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_B6 = CLBLM_R_X5Y138_SLICE_X6Y138_BQ;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_C1 = CLBLM_L_X8Y142_SLICE_X11Y142_DQ;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_C2 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_C2 = 1'b1;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_C4 = 1'b1;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_C5 = CLBLM_L_X10Y134_SLICE_X13Y134_BQ;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_C6 = CLBLM_R_X5Y138_SLICE_X6Y138_AQ;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_D1 = CLBLM_R_X7Y142_SLICE_X9Y142_CO6;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_D2 = 1'b1;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_D3 = CLBLL_L_X4Y143_SLICE_X4Y143_BO5;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_D4 = 1'b1;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_D5 = CLBLM_R_X7Y137_SLICE_X9Y137_AQ;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_D6 = CLBLM_L_X12Y136_SLICE_X17Y136_AQ;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y167_OLOGIC_X0Y168_D1 = RIOB33_X105Y123_IOB_X1Y123_I;
  assign CLBLM_R_X13Y144_SLICE_X18Y144_C5 = CLBLM_R_X13Y140_SLICE_X18Y140_BQ;
  assign LIOI3_X0Y167_OLOGIC_X0Y168_T1 = 1'b1;
  assign LIOI3_X0Y105_OLOGIC_X0Y106_D1 = CLBLL_L_X4Y138_SLICE_X5Y138_DO6;
  assign CLBLM_R_X103Y170_SLICE_X163Y170_A3 = CLBLM_R_X15Y142_SLICE_X20Y142_AQ;
  assign LIOI3_X0Y167_OLOGIC_X0Y167_D1 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign LIOI3_X0Y105_OLOGIC_X0Y106_T1 = 1'b1;
  assign RIOI3_X105Y151_OLOGIC_X1Y152_D1 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign LIOI3_X0Y167_OLOGIC_X0Y167_T1 = 1'b1;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_D4 = 1'b1;
  assign LIOI3_X0Y105_OLOGIC_X0Y105_D1 = CLBLL_L_X2Y133_SLICE_X0Y133_BO5;
  assign RIOI3_X105Y151_OLOGIC_X1Y152_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_D1 = CLBLM_R_X7Y132_SLICE_X9Y132_DQ;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_C4 = CLBLM_R_X11Y143_SLICE_X14Y143_CO6;
  assign LIOI3_X0Y105_OLOGIC_X0Y105_T1 = 1'b1;
  assign RIOI3_X105Y151_OLOGIC_X1Y151_D1 = LIOB33_X0Y75_IOB_X0Y76_I;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_T1 = 1'b1;
  assign RIOI3_X105Y151_OLOGIC_X1Y151_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_D1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_C5 = CLBLM_L_X10Y145_SLICE_X12Y145_CO6;
  assign LIOB33_X0Y171_IOB_X0Y172_O = CLBLM_R_X103Y140_SLICE_X163Y140_AO6;
  assign LIOB33_X0Y171_IOB_X0Y171_O = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_T1 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_C6 = CLBLM_R_X11Y143_SLICE_X15Y143_BQ;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_A1 = CLBLM_R_X11Y135_SLICE_X14Y135_AQ;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_A2 = 1'b1;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_A3 = CLBLM_R_X5Y139_SLICE_X7Y139_AQ;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_A5 = CLBLM_R_X5Y139_SLICE_X6Y139_AQ;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_A6 = CLBLM_R_X7Y139_SLICE_X8Y139_DO6;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_C4 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_C5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_B1 = CLBLM_R_X5Y139_SLICE_X7Y139_CQ;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_B2 = 1'b1;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_B4 = 1'b1;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_B5 = CLBLM_L_X10Y137_SLICE_X13Y137_BQ;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_C6 = 1'b1;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_C1 = CLBLM_R_X7Y134_SLICE_X9Y134_AQ;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_C2 = CLBLM_R_X5Y139_SLICE_X7Y139_CQ;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_C4 = CLBLL_L_X4Y139_SLICE_X4Y139_BO6;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_C5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_C6 = CLBLL_L_X4Y138_SLICE_X5Y138_CO5;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_D1 = CLBLM_R_X5Y139_SLICE_X6Y139_AQ;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_D2 = CLBLM_R_X5Y139_SLICE_X7Y139_CQ;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_D3 = CLBLM_R_X5Y143_SLICE_X6Y143_AO5;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_D4 = CLBLM_R_X3Y142_SLICE_X3Y142_AO6;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_D5 = 1'b1;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_D6 = 1'b1;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_A1 = CLBLM_L_X8Y143_SLICE_X10Y143_DO6;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_A2 = 1'b1;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_A3 = CLBLM_R_X5Y139_SLICE_X6Y139_AQ;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_A4 = CLBLM_R_X5Y134_SLICE_X6Y134_A5Q;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_A6 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_B1 = CLBLM_L_X8Y142_SLICE_X10Y142_DQ;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_B2 = CLBLM_R_X5Y139_SLICE_X6Y139_BQ;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_B3 = CLBLM_R_X7Y131_SLICE_X9Y131_AQ;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_B4 = CLBLM_L_X12Y134_SLICE_X17Y134_AO6;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_B6 = CLBLM_L_X10Y139_SLICE_X13Y139_B5Q;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_D1 = CLBLM_R_X3Y143_SLICE_X2Y143_AO5;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_D2 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_C1 = CLBLM_L_X8Y137_SLICE_X10Y137_AQ;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_C2 = CLBLM_R_X7Y137_SLICE_X8Y137_BQ;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_C3 = CLBLL_L_X2Y140_SLICE_X1Y140_AO6;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_C4 = CLBLM_R_X3Y143_SLICE_X2Y143_AO5;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_C5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_C6 = CLBLL_L_X2Y141_SLICE_X1Y141_AO6;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_C4 = CLBLM_L_X10Y139_SLICE_X13Y139_CQ;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_D5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_D1 = CLBLL_L_X4Y137_SLICE_X4Y137_AQ;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_D2 = CLBLM_R_X3Y143_SLICE_X2Y143_AO6;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_D3 = CLBLM_R_X5Y134_SLICE_X7Y134_CQ;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_D4 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_D5 = CLBLL_L_X2Y140_SLICE_X1Y140_AO6;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_D6 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_D6 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_C6 = CLBLM_R_X11Y142_SLICE_X14Y142_BQ;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_A4 = CLBLL_L_X4Y133_SLICE_X5Y133_BO6;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_A5 = 1'b1;
  assign LIOB33_X0Y173_IOB_X0Y174_O = CLBLM_R_X11Y153_SLICE_X14Y153_AO6;
  assign LIOB33_X0Y173_IOB_X0Y173_O = CLBLM_R_X103Y140_SLICE_X163Y140_AO5;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_B4 = CLBLM_R_X5Y138_SLICE_X7Y138_CQ;
  assign CLBLM_R_X13Y144_SLICE_X18Y144_D5 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_B5 = CLBLM_R_X3Y142_SLICE_X3Y142_AO6;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_B6 = CLBLL_L_X4Y143_SLICE_X5Y143_AO5;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_C1 = CLBLM_R_X3Y143_SLICE_X2Y143_AO5;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_C2 = CLBLM_R_X7Y138_SLICE_X8Y138_AQ;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_C3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_C4 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_C5 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_C6 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_X105Y173_OLOGIC_X1Y174_T1 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_A1 = CLBLM_R_X5Y136_SLICE_X6Y136_AQ;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_A2 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_A3 = CLBLM_L_X8Y138_SLICE_X10Y138_CQ;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_A4 = CLBLM_L_X8Y143_SLICE_X10Y143_DO5;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_A6 = CLBLM_R_X5Y140_SLICE_X7Y140_AQ;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_D1 = CLBLM_R_X3Y142_SLICE_X3Y142_AO6;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_B1 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_B2 = CLBLM_R_X5Y141_SLICE_X6Y141_AQ;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_B3 = CLBLM_R_X11Y138_SLICE_X15Y138_CQ;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_B4 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_D2 = CLBLM_R_X7Y142_SLICE_X9Y142_CO6;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_D3 = CLBLM_R_X7Y140_SLICE_X8Y140_AQ;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_C1 = CLBLM_R_X5Y135_SLICE_X6Y135_AQ;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_C2 = CLBLM_L_X8Y140_SLICE_X10Y140_CQ;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_C3 = CLBLM_R_X5Y143_SLICE_X6Y143_BO5;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_C4 = CLBLM_R_X5Y143_SLICE_X6Y143_AO6;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_C5 = CLBLM_R_X3Y142_SLICE_X2Y142_AO5;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_C6 = CLBLM_L_X10Y144_SLICE_X12Y144_AQ;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_D4 = CLBLM_R_X7Y142_SLICE_X8Y142_CO6;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_D5 = CLBLM_R_X7Y144_SLICE_X8Y144_DO6;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_D6 = CLBLM_L_X12Y140_SLICE_X16Y140_AQ;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_D1 = CLBLM_R_X5Y141_SLICE_X7Y141_AQ;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_D2 = CLBLL_L_X4Y137_SLICE_X5Y137_CO6;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_D3 = CLBLM_R_X5Y143_SLICE_X6Y143_AO5;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_D4 = CLBLM_L_X8Y142_SLICE_X10Y142_BQ;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_D5 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_D6 = CLBLM_R_X7Y142_SLICE_X9Y142_CO5;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_A1 = CLBLM_R_X5Y140_SLICE_X6Y140_DO6;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_A2 = CLBLM_R_X5Y138_SLICE_X6Y138_DO6;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_A3 = CLBLM_R_X5Y140_SLICE_X7Y140_CO6;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_A4 = CLBLM_R_X3Y142_SLICE_X2Y142_CO6;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_A5 = CLBLM_R_X3Y139_SLICE_X2Y139_CO6;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_A6 = CLBLM_R_X7Y140_SLICE_X9Y140_DO6;
  assign RIOI3_X105Y173_OLOGIC_X1Y173_D1 = CLBLM_R_X11Y144_SLICE_X14Y144_BO5;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_B1 = CLBLM_R_X5Y141_SLICE_X6Y141_CQ;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_B2 = CLBLM_R_X3Y143_SLICE_X2Y143_BO6;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_B3 = CLBLM_R_X5Y139_SLICE_X6Y139_DO6;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_B4 = CLBLM_R_X7Y141_SLICE_X9Y141_CO6;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_B5 = CLBLM_R_X3Y140_SLICE_X3Y140_CO6;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_B6 = CLBLM_R_X5Y143_SLICE_X6Y143_AO6;
  assign LIOB33_X0Y109_IOB_X0Y109_O = CLBLL_L_X2Y127_SLICE_X0Y127_AO6;
  assign LIOB33_X0Y109_IOB_X0Y110_O = CLBLL_L_X2Y127_SLICE_X0Y127_AO5;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_C1 = CLBLM_L_X8Y141_SLICE_X11Y141_AQ;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_C2 = CLBLM_R_X7Y133_SLICE_X8Y133_CQ;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_C3 = CLBLM_R_X3Y141_SLICE_X2Y141_AO5;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_C4 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_C5 = CLBLM_R_X3Y142_SLICE_X2Y142_AO5;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_C6 = CLBLM_R_X5Y143_SLICE_X6Y143_BO6;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_D1 = CLBLM_L_X8Y140_SLICE_X11Y140_BQ;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_D2 = CLBLL_L_X4Y143_SLICE_X5Y143_AO6;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_D3 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_D4 = CLBLM_R_X7Y143_SLICE_X8Y143_A5Q;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_D5 = CLBLM_R_X5Y141_SLICE_X6Y141_DO6;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_D6 = CLBLM_R_X3Y141_SLICE_X2Y141_AO5;
  assign RIOI3_X105Y173_OLOGIC_X1Y173_T1 = 1'b1;
  assign LIOB33_X0Y175_IOB_X0Y176_O = RIOB33_X105Y127_IOB_X1Y128_I;
  assign LIOB33_X0Y175_IOB_X0Y175_O = RIOB33_X105Y127_IOB_X1Y127_I;
  assign LIOI3_X0Y171_OLOGIC_X0Y172_D1 = CLBLM_R_X103Y140_SLICE_X163Y140_AO6;
  assign RIOI3_SING_X105Y100_ILOGIC_X1Y100_D = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_D1 = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign LIOI3_X0Y171_OLOGIC_X0Y172_T1 = 1'b1;
  assign LIOI3_X0Y109_OLOGIC_X0Y110_D1 = CLBLL_L_X2Y127_SLICE_X0Y127_AO5;
  assign LIOI3_X0Y171_OLOGIC_X0Y171_D1 = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_C4 = 1'b1;
  assign LIOI3_X0Y109_OLOGIC_X0Y110_T1 = 1'b1;
  assign RIOI3_X105Y153_OLOGIC_X1Y154_D1 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign LIOI3_X0Y171_OLOGIC_X0Y171_T1 = 1'b1;
  assign LIOI3_X0Y109_OLOGIC_X0Y109_D1 = CLBLL_L_X2Y127_SLICE_X0Y127_AO6;
  assign RIOI3_X105Y153_OLOGIC_X1Y154_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_D1 = CLBLM_R_X3Y136_SLICE_X3Y136_DQ;
  assign LIOI3_X0Y109_OLOGIC_X0Y109_T1 = 1'b1;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_C5 = 1'b1;
  assign RIOI3_X105Y153_OLOGIC_X1Y153_D1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_T1 = 1'b1;
  assign RIOI3_X105Y153_OLOGIC_X1Y153_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_D1 = CLBLM_R_X3Y137_SLICE_X2Y137_BQ;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_B1 = 1'b1;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_C6 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_B2 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_B3 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_T1 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_A1 = CLBLM_L_X8Y143_SLICE_X10Y143_DO6;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_A2 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_A3 = CLBLM_R_X5Y141_SLICE_X7Y141_AQ;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_A4 = CLBLM_R_X11Y139_SLICE_X15Y139_DQ;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_A5 = CLBLM_R_X5Y137_SLICE_X7Y137_AQ;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_B4 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_B5 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_B1 = CLBLM_L_X8Y140_SLICE_X11Y140_A5Q;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_B2 = CLBLM_R_X5Y141_SLICE_X7Y141_BQ;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_B4 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_B5 = CLBLM_R_X7Y135_SLICE_X9Y135_BQ;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_B6 = CLBLL_L_X4Y133_SLICE_X5Y133_BO6;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_C1 = CLBLM_R_X7Y135_SLICE_X9Y135_BQ;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_C2 = CLBLM_R_X7Y140_SLICE_X9Y140_CQ;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_C3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_C4 = CLBLM_R_X3Y143_SLICE_X3Y143_AO6;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_C5 = CLBLM_R_X3Y143_SLICE_X2Y143_AO5;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_C6 = CLBLL_L_X2Y141_SLICE_X1Y141_AO6;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_D1 = CLBLM_R_X5Y143_SLICE_X7Y143_CO6;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_D2 = CLBLM_R_X7Y142_SLICE_X8Y142_DO6;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_D3 = CLBLM_R_X5Y143_SLICE_X6Y143_DO6;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_D4 = CLBLL_L_X2Y141_SLICE_X1Y141_DO6;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_D5 = CLBLM_R_X5Y138_SLICE_X7Y138_DO6;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_D6 = CLBLM_R_X3Y142_SLICE_X2Y142_CO6;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_A1 = CLBLL_L_X4Y137_SLICE_X4Y137_CQ;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_A2 = CLBLM_L_X12Y135_SLICE_X17Y135_AQ;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_A3 = CLBLM_R_X5Y141_SLICE_X6Y141_AQ;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_A4 = CLBLM_R_X7Y137_SLICE_X8Y137_CQ;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_A5 = CLBLL_L_X4Y135_SLICE_X4Y135_BQ;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_AX = CLBLM_L_X8Y141_SLICE_X11Y141_DO6;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_B1 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_B2 = CLBLL_L_X4Y138_SLICE_X5Y138_BQ;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_B4 = CLBLM_L_X8Y143_SLICE_X10Y143_DO5;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_B5 = CLBLM_R_X5Y141_SLICE_X7Y141_AQ;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_B6 = CLBLM_R_X5Y141_SLICE_X6Y141_BQ;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_C1 = CLBLM_L_X8Y143_SLICE_X10Y143_DO5;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_C2 = CLBLM_R_X5Y141_SLICE_X6Y141_CQ;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_C3 = CLBLM_R_X5Y141_SLICE_X6Y141_BQ;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_C5 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_C6 = CLBLM_R_X7Y135_SLICE_X8Y135_CQ;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_D1 = CLBLL_L_X2Y140_SLICE_X1Y140_AO6;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_D2 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_D3 = CLBLL_L_X4Y143_SLICE_X5Y143_BO5;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_D4 = CLBLM_L_X8Y142_SLICE_X10Y142_CQ;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_D5 = CLBLM_R_X3Y143_SLICE_X3Y143_AO5;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_D6 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign LIOB33_X0Y177_IOB_X0Y178_O = RIOB33_X105Y129_IOB_X1Y130_I;
  assign LIOB33_X0Y177_IOB_X0Y177_O = RIOB33_X105Y129_IOB_X1Y129_I;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_T1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_B4 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_B6 = 1'b1;
  assign RIOI3_SING_X105Y149_ILOGIC_X1Y149_D = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_C4 = CLBLM_L_X12Y143_SLICE_X17Y143_BQ;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_C1 = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_T1 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_C5 = CLBLM_R_X13Y144_SLICE_X18Y144_AQ;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_C2 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_C6 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_C3 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_C4 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_C5 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_A1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_A2 = CLBLM_L_X8Y140_SLICE_X10Y140_BQ;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_A3 = CLBLM_R_X3Y143_SLICE_X2Y143_AO5;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_A4 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_A5 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_A6 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_C6 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_B1 = CLBLL_L_X4Y143_SLICE_X5Y143_BO5;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_B2 = CLBLM_R_X7Y143_SLICE_X9Y143_CQ;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_B3 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_B4 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_B5 = CLBLM_R_X7Y134_SLICE_X9Y134_BQ;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_B6 = CLBLM_R_X3Y143_SLICE_X3Y143_AO6;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_C1 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_C2 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_C3 = CLBLM_R_X5Y140_SLICE_X7Y140_AQ;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_C4 = CLBLM_R_X3Y143_SLICE_X3Y143_AO5;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_C5 = CLBLL_L_X4Y143_SLICE_X5Y143_BO5;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_C6 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_D1 = CLBLM_R_X7Y134_SLICE_X9Y134_BQ;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_D2 = CLBLM_R_X5Y143_SLICE_X6Y143_AO6;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_D3 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_D4 = CLBLM_R_X5Y142_SLICE_X7Y142_CO6;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_D2 = CLBLM_R_X13Y140_SLICE_X18Y140_BQ;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_D5 = CLBLM_R_X5Y143_SLICE_X6Y143_BO5;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_D6 = CLBLM_R_X7Y143_SLICE_X9Y143_CQ;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_A1 = CLBLM_R_X5Y142_SLICE_X7Y142_CO6;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_A2 = CLBLM_R_X5Y142_SLICE_X7Y142_BO6;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_A3 = CLBLM_R_X5Y142_SLICE_X7Y142_AO6;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_A4 = CLBLM_R_X5Y142_SLICE_X6Y142_BO6;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_A5 = CLBLM_R_X5Y141_SLICE_X6Y141_AQ;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_A6 = CLBLM_R_X3Y142_SLICE_X3Y142_AO6;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_D5 = CLBLM_R_X13Y144_SLICE_X18Y144_AQ;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_D1 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_B1 = LIOB33_X0Y67_IOB_X0Y68_I;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_B2 = CLBLM_R_X3Y143_SLICE_X2Y143_AO6;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_B3 = CLBLL_L_X4Y138_SLICE_X5Y138_DO5;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_B4 = CLBLM_R_X3Y143_SLICE_X3Y143_AO6;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_B5 = CLBLM_R_X5Y141_SLICE_X7Y141_BQ;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_B6 = CLBLM_R_X3Y143_SLICE_X3Y143_AO5;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_D2 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_D3 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_C1 = CLBLM_R_X5Y143_SLICE_X6Y143_AO5;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_C2 = CLBLM_R_X3Y141_SLICE_X3Y141_DO6;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_C3 = CLBLM_R_X5Y142_SLICE_X7Y142_DO6;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_C4 = CLBLM_R_X3Y143_SLICE_X3Y143_DO6;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_C5 = CLBLM_R_X5Y142_SLICE_X6Y142_DO6;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_C6 = CLBLM_L_X8Y140_SLICE_X10Y140_BQ;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_D4 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_D5 = 1'b1;
  assign LIOB33_X0Y179_IOB_X0Y179_O = RIOB33_X105Y131_IOB_X1Y131_I;
  assign LIOB33_X0Y179_IOB_X0Y180_O = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_D6 = 1'b1;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_D6 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_D1 = CLBLM_R_X5Y141_SLICE_X7Y141_BQ;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_D2 = CLBLL_L_X4Y141_SLICE_X5Y141_BO6;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_D3 = CLBLM_R_X5Y141_SLICE_X6Y141_AQ;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_D4 = CLBLM_R_X3Y142_SLICE_X3Y142_AO6;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_D5 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_D6 = CLBLL_L_X4Y143_SLICE_X4Y143_AO6;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I0 = LIOB33_X0Y77_IOB_X0Y78_I;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_A4 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I1 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_A5 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_A6 = CLBLM_L_X12Y142_SLICE_X16Y142_A5Q;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_B6 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_C6 = CLBLM_L_X10Y144_SLICE_X13Y144_AQ;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_D3 = 1'b1;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_D4 = 1'b1;
  assign RIOI3_SING_X105Y150_OLOGIC_X1Y150_D1 = LIOB33_X0Y75_IOB_X0Y75_I;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_C6 = CLBLM_L_X8Y139_SLICE_X10Y139_BQ;
  assign RIOI3_SING_X105Y150_OLOGIC_X1Y150_T1 = 1'b1;
  assign LIOB33_X0Y181_IOB_X0Y182_O = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_A5 = CLBLM_R_X11Y144_SLICE_X14Y144_AQ;
  assign LIOB33_X0Y181_IOB_X0Y181_O = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_D2 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_D5 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_A1 = CLBLL_L_X4Y143_SLICE_X5Y143_BO5;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_A2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_A3 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_A4 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_A5 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_A6 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign RIOB33_X105Y163_IOB_X1Y164_O = CLBLM_L_X12Y139_SLICE_X17Y139_DO5;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_B1 = CLBLL_L_X4Y134_SLICE_X5Y134_AQ;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_B2 = CLBLL_L_X4Y143_SLICE_X4Y143_AO6;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_B3 = CLBLM_R_X7Y142_SLICE_X8Y142_AQ;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_B4 = CLBLL_L_X4Y143_SLICE_X4Y143_AO5;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_B5 = CLBLM_R_X5Y143_SLICE_X7Y143_AO6;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_B6 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_A2 = CLBLL_L_X4Y134_SLICE_X4Y134_BQ;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_A3 = CLBLM_R_X3Y133_SLICE_X3Y133_AQ;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_A4 = CLBLM_R_X3Y137_SLICE_X3Y137_AQ;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_A5 = CLBLL_L_X4Y132_SLICE_X5Y132_AQ;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_A6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_C1 = CLBLM_R_X5Y143_SLICE_X7Y143_AO6;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_C2 = CLBLL_L_X4Y143_SLICE_X4Y143_AO6;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_C3 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_B1 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_B2 = 1'b1;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_C3 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_B3 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_B4 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_B5 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_B6 = 1'b1;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_C4 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_C1 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_C2 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_C3 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_C4 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_C5 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_C6 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_D3 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_D4 = CLBLM_R_X3Y143_SLICE_X3Y143_AO5;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_A1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_A2 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_A3 = CLBLM_R_X3Y143_SLICE_X2Y143_AO5;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_A4 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_A5 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_D1 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_D2 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_D3 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_D4 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_D5 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_D6 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_A6 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_B1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_B2 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_B3 = CLBLL_L_X4Y143_SLICE_X5Y143_BO6;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_B4 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_A1 = CLBLM_R_X5Y141_SLICE_X7Y141_DO6;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_A2 = CLBLL_L_X4Y142_SLICE_X5Y142_DO6;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_A3 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_A4 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_A5 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_A6 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_C1 = CLBLM_L_X10Y141_SLICE_X13Y141_CQ;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_C2 = CLBLL_L_X2Y141_SLICE_X1Y141_AO5;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_C3 = CLBLL_L_X4Y143_SLICE_X5Y143_BO5;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_B1 = CLBLL_L_X4Y135_SLICE_X5Y135_C5Q;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_B2 = CLBLL_L_X4Y133_SLICE_X4Y133_BO5;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_B3 = CLBLL_L_X4Y139_SLICE_X4Y139_BO6;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_B4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_B5 = CLBLM_R_X3Y133_SLICE_X2Y133_CO6;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_B6 = CLBLM_R_X3Y140_SLICE_X2Y140_DO6;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_D1 = CLBLM_R_X5Y135_SLICE_X6Y135_BQ;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_D2 = CLBLM_R_X5Y139_SLICE_X6Y139_CO6;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_D3 = CLBLM_R_X5Y143_SLICE_X7Y143_DO6;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_C1 = CLBLL_L_X4Y142_SLICE_X5Y142_DO6;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_C2 = CLBLL_L_X4Y135_SLICE_X4Y135_DO5;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_C3 = LIOB33_X0Y51_IOB_X0Y51_I;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_C4 = LIOB33_X0Y53_IOB_X0Y53_I;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_C5 = CLBLM_R_X5Y141_SLICE_X7Y141_DO6;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_C6 = CLBLM_R_X5Y140_SLICE_X6Y140_AO6;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_D6 = CLBLL_L_X4Y143_SLICE_X5Y143_DO6;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_D4 = CLBLM_R_X5Y143_SLICE_X6Y143_CO6;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_D5 = CLBLM_R_X5Y143_SLICE_X6Y143_BO5;
  assign RIOI3_X105Y155_OLOGIC_X1Y155_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_D1 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_D1 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_D2 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_D3 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_D4 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_D5 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_D6 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_T1 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X162Y170_B6 = 1'b1;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_C1 = CLBLM_R_X11Y140_SLICE_X14Y140_AQ;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_C6 = CLBLM_L_X12Y143_SLICE_X17Y143_CO5;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE0 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE1 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE0 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE1 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S0 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S1 = 1'b1;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_D2 = CLBLM_L_X12Y137_SLICE_X17Y137_BO5;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_D5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_D6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOI3_X0Y51_ILOGIC_X0Y52_D = LIOB33_X0Y51_IOB_X0Y52_I;
  assign LIOI3_X0Y51_ILOGIC_X0Y51_D = LIOB33_X0Y51_IOB_X0Y51_I;
  assign RIOI3_SING_X105Y199_OLOGIC_X1Y199_D1 = CLBLM_R_X13Y144_SLICE_X19Y144_AQ;
  assign RIOB33_X105Y151_IOB_X1Y152_O = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign RIOB33_X105Y151_IOB_X1Y151_O = LIOB33_X0Y75_IOB_X0Y76_I;
  assign RIOI3_SING_X105Y199_OLOGIC_X1Y199_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y58_D = LIOB33_X0Y57_IOB_X0Y58_I;
  assign LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y57_D = LIOB33_X0Y57_IOB_X0Y57_I;
  assign LIOB33_X0Y183_IOB_X0Y184_O = RIOB33_X105Y135_IOB_X1Y136_I;
  assign LIOB33_X0Y183_IOB_X0Y183_O = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_C4 = CLBLM_L_X12Y143_SLICE_X16Y143_BQ;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_C5 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_B2 = CLBLM_L_X10Y135_SLICE_X13Y135_CO6;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_B4 = CLBLM_L_X8Y138_SLICE_X10Y138_AQ;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_B5 = CLBLM_R_X11Y141_SLICE_X14Y141_BQ;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_B6 = CLBLM_R_X11Y143_SLICE_X15Y143_BQ;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_C1 = CLBLM_R_X11Y141_SLICE_X14Y141_BQ;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_D2 = 1'b1;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_C2 = CLBLM_R_X7Y133_SLICE_X9Y133_CQ;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_C3 = CLBLM_R_X11Y138_SLICE_X14Y138_DQ;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_C4 = CLBLM_R_X11Y139_SLICE_X14Y139_CQ;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_D5 = 1'b1;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_C5 = CLBLM_L_X8Y133_SLICE_X11Y133_AQ;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_C5 = CLBLM_R_X11Y142_SLICE_X14Y142_DO6;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_D6 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_C6 = 1'b1;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_C6 = CLBLM_L_X10Y145_SLICE_X12Y145_CO6;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_D1 = 1'b1;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_D2 = 1'b1;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_D3 = CLBLM_L_X12Y144_SLICE_X17Y144_AQ;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_D4 = 1'b1;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_D5 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_D6 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_AX = CLBLM_R_X7Y143_SLICE_X8Y143_BO6;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOB33_X0Y111_IOB_X0Y112_O = CLBLM_L_X12Y133_SLICE_X16Y133_C5Q;
  assign LIOB33_X0Y111_IOB_X0Y111_O = 1'b0;
  assign RIOB33_X105Y153_IOB_X1Y154_O = RIOB33_X105Y101_IOB_X1Y102_I;
  assign RIOB33_X105Y153_IOB_X1Y153_O = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_C2 = CLBLM_R_X7Y143_SLICE_X8Y143_CQ;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_C3 = CLBLM_R_X5Y135_SLICE_X6Y135_DQ;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_C4 = CLBLM_L_X12Y141_SLICE_X16Y141_AQ;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_C5 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_C6 = CLBLL_L_X4Y133_SLICE_X5Y133_BO6;
  assign LIOB33_X0Y185_IOB_X0Y186_O = RIOB33_X105Y143_IOB_X1Y143_I;
  assign LIOB33_X0Y185_IOB_X0Y185_O = RIOB33_X105Y137_IOB_X1Y137_I;
  assign LIOB33_X0Y159_IOB_X0Y160_O = RIOB33_X105Y107_IOB_X1Y107_I;
  assign LIOB33_X0Y159_IOB_X0Y159_O = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_A1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_A2 = CLBLL_L_X4Y134_SLICE_X4Y134_BQ;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_A3 = CLBLM_R_X3Y135_SLICE_X3Y135_AQ;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_A4 = CLBLM_R_X7Y142_SLICE_X9Y142_AQ;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_A5 = CLBLM_R_X3Y135_SLICE_X3Y135_CO6;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_B1 = CLBLL_L_X4Y133_SLICE_X5Y133_BO6;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_B2 = CLBLM_R_X3Y135_SLICE_X3Y135_BQ;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_B3 = CLBLM_R_X3Y133_SLICE_X3Y133_AQ;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_B4 = 1'b1;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_B5 = CLBLM_R_X5Y135_SLICE_X6Y135_D5Q;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_C1 = CLBLM_R_X3Y137_SLICE_X3Y137_AQ;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_C2 = CLBLM_R_X3Y136_SLICE_X3Y136_AQ;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_C3 = 1'b1;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_C4 = 1'b1;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_C5 = CLBLM_R_X3Y133_SLICE_X3Y133_AQ;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_C6 = 1'b1;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_D1 = 1'b1;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_D2 = 1'b1;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_D3 = 1'b1;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_D4 = 1'b1;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_D5 = 1'b1;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_D6 = 1'b1;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_A1 = 1'b1;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_A2 = 1'b1;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_A3 = 1'b1;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_A4 = 1'b1;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_A5 = 1'b1;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_A6 = 1'b1;
  assign RIOI3_X105Y189_OLOGIC_X1Y189_D1 = CLBLM_L_X10Y143_SLICE_X13Y143_BQ;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_B1 = 1'b1;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_B2 = 1'b1;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_B3 = 1'b1;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_B4 = 1'b1;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_B5 = 1'b1;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_B6 = 1'b1;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_C1 = 1'b1;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_C2 = 1'b1;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_C3 = 1'b1;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_C4 = 1'b1;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_C5 = 1'b1;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_C6 = 1'b1;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_D1 = 1'b1;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_D2 = 1'b1;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_D3 = 1'b1;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_D4 = 1'b1;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_D5 = 1'b1;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_D6 = 1'b1;
  assign LIOI3_X0Y175_OLOGIC_X0Y176_D1 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y106_D = RIOB33_X105Y105_IOB_X1Y106_I;
  assign LIOI3_X0Y175_OLOGIC_X0Y176_T1 = 1'b1;
  assign LIOI3_X0Y115_OLOGIC_X0Y116_D1 = CLBLM_L_X8Y135_SLICE_X11Y135_BQ;
  assign LIOI3_X0Y175_OLOGIC_X0Y175_D1 = RIOB33_X105Y127_IOB_X1Y127_I;
  assign LIOI3_X0Y115_OLOGIC_X0Y116_T1 = 1'b1;
  assign RIOI3_X105Y159_OLOGIC_X1Y160_D1 = CLBLM_L_X12Y138_SLICE_X17Y138_DO5;
  assign LIOI3_X0Y175_OLOGIC_X0Y175_T1 = 1'b1;
  assign LIOI3_X0Y115_OLOGIC_X0Y115_D1 = CLBLM_L_X12Y133_SLICE_X16Y133_CQ;
  assign RIOI3_X105Y159_OLOGIC_X1Y160_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_D1 = RIOB33_X105Y145_IOB_X1Y145_I;
  assign LIOI3_X0Y115_OLOGIC_X0Y115_T1 = 1'b1;
  assign RIOI3_X105Y159_OLOGIC_X1Y159_D1 = CLBLM_L_X12Y138_SLICE_X17Y138_DO6;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_T1 = 1'b1;
  assign RIOI3_X105Y159_OLOGIC_X1Y159_T1 = 1'b1;
  assign RIOB33_X105Y155_IOB_X1Y156_O = RIOB33_X105Y103_IOB_X1Y104_I;
  assign RIOB33_X105Y155_IOB_X1Y155_O = RIOB33_X105Y103_IOB_X1Y103_I;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_D1 = RIOB33_X105Y143_IOB_X1Y144_I;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_T1 = 1'b1;
  assign RIOI3_X105Y105_ILOGIC_X1Y105_D = RIOB33_X105Y105_IOB_X1Y105_I;
  assign LIOB33_X0Y187_IOB_X0Y188_O = RIOB33_X105Y145_IOB_X1Y145_I;
  assign LIOB33_X0Y187_IOB_X0Y187_O = RIOB33_X105Y143_IOB_X1Y144_I;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_A2 = CLBLM_R_X3Y133_SLICE_X3Y133_AQ;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_A3 = CLBLM_R_X3Y136_SLICE_X3Y136_AQ;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_A4 = CLBLM_R_X3Y139_SLICE_X3Y139_AQ;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_A5 = CLBLM_R_X3Y137_SLICE_X3Y137_AQ;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_A6 = CLBLM_R_X3Y137_SLICE_X3Y137_AO5;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_B1 = CLBLM_R_X3Y137_SLICE_X3Y137_BO5;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_B2 = CLBLM_R_X3Y136_SLICE_X3Y136_BQ;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_B3 = CLBLM_R_X5Y135_SLICE_X6Y135_D5Q;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_B5 = CLBLM_R_X3Y136_SLICE_X2Y136_AQ;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_B6 = CLBLM_R_X3Y137_SLICE_X3Y137_AO5;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_C1 = CLBLM_R_X3Y136_SLICE_X2Y136_AQ;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_C2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_C3 = CLBLM_R_X3Y136_SLICE_X3Y136_BQ;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_C4 = CLBLM_R_X7Y137_SLICE_X8Y137_CQ;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_C5 = CLBLM_R_X3Y137_SLICE_X3Y137_BO5;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_C6 = CLBLL_L_X4Y134_SLICE_X4Y134_BQ;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_D1 = CLBLL_L_X4Y134_SLICE_X4Y134_BQ;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_D2 = CLBLM_L_X8Y135_SLICE_X10Y135_A5Q;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_D3 = CLBLM_R_X3Y136_SLICE_X2Y136_BO6;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_D4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_D5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_D6 = CLBLM_R_X3Y136_SLICE_X3Y136_DQ;
  assign RIOI3_X105Y189_OLOGIC_X1Y189_T1 = 1'b1;
  assign LIOI3_X0Y53_ILOGIC_X0Y54_D = LIOB33_X0Y53_IOB_X0Y54_I;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_A1 = CLBLM_R_X3Y137_SLICE_X3Y137_BO5;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_A2 = CLBLL_L_X4Y134_SLICE_X4Y134_BQ;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_A3 = CLBLM_R_X3Y136_SLICE_X2Y136_AQ;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_A5 = CLBLL_L_X4Y135_SLICE_X5Y135_C5Q;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOI3_X0Y53_ILOGIC_X0Y53_D = LIOB33_X0Y53_IOB_X0Y53_I;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_B1 = CLBLM_R_X3Y137_SLICE_X2Y137_BQ;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_B2 = CLBLM_R_X3Y135_SLICE_X3Y135_AQ;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_B3 = CLBLM_R_X3Y137_SLICE_X3Y137_AQ;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_B4 = CLBLM_R_X3Y133_SLICE_X3Y133_AQ;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_B5 = CLBLM_R_X3Y136_SLICE_X3Y136_AQ;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_B6 = 1'b1;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_C1 = CLBLM_R_X3Y136_SLICE_X3Y136_AQ;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_C2 = CLBLM_R_X3Y135_SLICE_X3Y135_AQ;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_C3 = CLBLM_R_X3Y137_SLICE_X2Y137_BQ;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_C4 = CLBLM_R_X3Y133_SLICE_X3Y133_AQ;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_C5 = CLBLM_R_X3Y136_SLICE_X3Y136_DQ;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_C6 = CLBLM_R_X3Y137_SLICE_X3Y137_AQ;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_C4 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y70_D = LIOB33_X0Y69_IOB_X0Y70_I;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y69_D = LIOB33_X0Y69_IOB_X0Y69_I;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_C5 = 1'b1;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_D1 = 1'b1;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_D2 = 1'b1;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_D3 = 1'b1;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_D4 = 1'b1;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_D5 = 1'b1;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_D6 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_C6 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_D3 = 1'b1;
  assign RIOB33_X105Y157_IOB_X1Y158_O = CLBLM_R_X37Y138_SLICE_X56Y138_AO6;
  assign RIOB33_X105Y157_IOB_X1Y157_O = RIOB33_X105Y125_IOB_X1Y126_I;
  assign LIOB33_X0Y189_IOB_X0Y190_O = RIOB33_X105Y147_IOB_X1Y147_I;
  assign LIOB33_X0Y189_IOB_X0Y189_O = RIOB33_X105Y145_IOB_X1Y146_I;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_D1 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign LIOI3_X0Y111_OLOGIC_X0Y112_D1 = CLBLM_L_X12Y133_SLICE_X16Y133_C5Q;
  assign LIOB33_X0Y161_IOB_X0Y162_O = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_C3 = 1'b1;
  assign LIOB33_X0Y161_IOB_X0Y161_O = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_C4 = 1'b1;
  assign CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_I = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_C5 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_T1 = 1'b1;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_C6 = 1'b1;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_A2 = CLBLM_L_X8Y142_SLICE_X11Y142_BQ;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_A3 = CLBLM_R_X3Y137_SLICE_X3Y137_AQ;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_A4 = CLBLL_L_X4Y134_SLICE_X4Y134_BQ;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_A6 = 1'b1;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_B1 = CLBLL_L_X4Y137_SLICE_X4Y137_BQ;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_B2 = CLBLM_R_X3Y136_SLICE_X3Y136_DQ;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_B3 = CLBLM_R_X3Y136_SLICE_X2Y136_BO6;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_B5 = CLBLM_R_X3Y137_SLICE_X2Y137_AQ;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_B6 = 1'b1;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_C2 = CLBLM_R_X3Y137_SLICE_X3Y137_CQ;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_C3 = CLBLM_R_X3Y137_SLICE_X3Y137_BQ;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_C4 = CLBLL_L_X4Y133_SLICE_X5Y133_BO6;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_C5 = 1'b1;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_C6 = CLBLM_L_X8Y140_SLICE_X10Y140_A5Q;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_D2 = 1'b1;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_D1 = CLBLL_L_X4Y142_SLICE_X5Y142_DO6;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_D2 = CLBLM_R_X5Y142_SLICE_X6Y142_CO6;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_D3 = CLBLL_L_X4Y141_SLICE_X4Y141_DO6;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_D4 = CLBLM_R_X3Y139_SLICE_X2Y139_AO5;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_D5 = CLBLL_L_X4Y142_SLICE_X4Y142_BO6;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_D6 = CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  assign RIOI3_X105Y185_OLOGIC_X1Y186_D1 = CLBLM_R_X13Y139_SLICE_X19Y139_AQ;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_A1 = CLBLM_L_X10Y143_SLICE_X12Y143_CQ;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_D6 = 1'b1;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_A3 = CLBLM_R_X3Y137_SLICE_X2Y137_AQ;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_A4 = CLBLL_L_X4Y134_SLICE_X4Y134_BQ;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_A6 = CLBLM_R_X3Y136_SLICE_X2Y136_CO6;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_B1 = CLBLM_R_X3Y136_SLICE_X2Y136_BO5;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_B2 = CLBLM_R_X7Y138_SLICE_X8Y138_AQ;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_B3 = CLBLM_R_X3Y137_SLICE_X2Y137_BQ;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_B4 = CLBLL_L_X4Y134_SLICE_X4Y134_BQ;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_C1 = 1'b1;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_C2 = 1'b1;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_C3 = 1'b1;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_C4 = 1'b1;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_C5 = 1'b1;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_C6 = 1'b1;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_D1 = 1'b1;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_D2 = 1'b1;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_B4 = 1'b1;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_D3 = 1'b1;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_D4 = 1'b1;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_D5 = 1'b1;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_D6 = 1'b1;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_B5 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_A2 = CLBLM_L_X12Y141_SLICE_X17Y141_AQ;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_A1 = CLBLM_L_X12Y144_SLICE_X16Y144_AO6;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_A3 = CLBLM_L_X10Y132_SLICE_X13Y132_AO6;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_A4 = CLBLM_L_X12Y132_SLICE_X17Y132_BO6;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_B6 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_A6 = CLBLM_L_X12Y133_SLICE_X16Y133_DO5;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_B1 = CLBLM_L_X12Y136_SLICE_X16Y136_CQ;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_B2 = CLBLM_R_X5Y132_SLICE_X7Y132_DO6;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_B3 = CLBLM_L_X12Y132_SLICE_X17Y132_AQ;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_B4 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_B5 = CLBLM_R_X11Y132_SLICE_X15Y132_AO5;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_B6 = CLBLM_L_X12Y133_SLICE_X16Y133_DO5;
  assign RIOI3_X105Y185_OLOGIC_X1Y186_T1 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_C1 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_C2 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_C3 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_C4 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_C5 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_C6 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_D1 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_D2 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_D3 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_D4 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_D5 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_D6 = 1'b1;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_C3 = 1'b1;
  assign RIOB33_X105Y159_IOB_X1Y159_O = CLBLM_L_X12Y138_SLICE_X17Y138_DO6;
  assign RIOB33_X105Y159_IOB_X1Y160_O = CLBLM_L_X12Y138_SLICE_X17Y138_DO5;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_C4 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_A1 = CLBLM_L_X12Y144_SLICE_X16Y144_AO6;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_A2 = CLBLM_L_X12Y136_SLICE_X16Y136_CQ;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_A3 = CLBLM_L_X12Y132_SLICE_X16Y132_AQ;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_A4 = CLBLM_L_X12Y132_SLICE_X16Y132_DO6;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_A5 = CLBLM_L_X10Y132_SLICE_X13Y132_AO6;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_C5 = 1'b1;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_C6 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_B2 = CLBLM_L_X12Y132_SLICE_X16Y132_BQ;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_B3 = CLBLM_R_X11Y133_SLICE_X14Y133_AQ;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_B4 = CLBLM_R_X5Y134_SLICE_X7Y134_DO6;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_B5 = CLBLM_R_X11Y138_SLICE_X14Y138_CQ;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_B6 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_C1 = CLBLM_R_X11Y132_SLICE_X15Y132_BO6;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_C2 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_C3 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_C5 = CLBLM_L_X12Y136_SLICE_X17Y136_DQ;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_C6 = CLBLM_R_X7Y131_SLICE_X9Y131_AQ;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_D1 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_D2 = CLBLM_L_X12Y136_SLICE_X16Y136_CQ;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_D3 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_D4 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_D5 = CLBLM_R_X11Y132_SLICE_X15Y132_AO5;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_D6 = CLBLM_R_X5Y134_SLICE_X7Y134_DO6;
  assign LIOB33_X0Y191_IOB_X0Y191_O = RIOB33_X105Y147_IOB_X1Y148_I;
  assign LIOB33_X0Y191_IOB_X0Y192_O = LIOB33_X0Y51_IOB_X0Y52_I;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_D3 = 1'b1;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_C3 = 1'b1;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_C4 = 1'b1;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_D5 = 1'b1;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_C5 = 1'b1;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_D6 = 1'b1;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_C6 = 1'b1;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_CE = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOI3_X0Y177_OLOGIC_X0Y178_D1 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign LIOI3_X0Y177_OLOGIC_X0Y178_T1 = 1'b1;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_D1 = CLBLL_L_X4Y135_SLICE_X5Y135_DQ;
  assign LIOI3_X0Y177_OLOGIC_X0Y177_D1 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_T1 = 1'b1;
  assign RIOI3_X105Y161_OLOGIC_X1Y162_D1 = CLBLM_R_X11Y141_SLICE_X14Y141_CO5;
  assign LIOI3_X0Y177_OLOGIC_X0Y177_T1 = 1'b1;
  assign LIOI3_X0Y117_OLOGIC_X0Y117_D1 = CLBLM_R_X5Y136_SLICE_X6Y136_D5Q;
  assign RIOI3_X105Y161_OLOGIC_X1Y162_T1 = 1'b1;
  assign LIOI3_X0Y117_OLOGIC_X0Y117_T1 = 1'b1;
  assign RIOI3_X105Y161_OLOGIC_X1Y161_D1 = CLBLM_R_X11Y141_SLICE_X14Y141_CO6;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_D4 = 1'b1;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_D5 = 1'b1;
  assign RIOI3_X105Y161_OLOGIC_X1Y161_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_D1 = CLBLM_L_X12Y139_SLICE_X17Y139_DO6;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_A1 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_A3 = CLBLM_R_X3Y138_SLICE_X3Y138_AQ;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_A4 = CLBLM_R_X7Y133_SLICE_X8Y133_DO6;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_A5 = CLBLL_L_X4Y137_SLICE_X4Y137_D5Q;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_A6 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_B1 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_B2 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_B3 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_B4 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_B5 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_B6 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_C1 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_C2 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_C3 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_C4 = 1'b1;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_B5 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_C5 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_C6 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_B6 = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_T1 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_D1 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_D2 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_D3 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_D4 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_D5 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_D6 = 1'b1;
  assign CLBLM_R_X37Y138_SLICE_X57Y138_A5 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_A1 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_A2 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_A3 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_A4 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_A5 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_A6 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_B1 = LIOB33_X0Y57_IOB_X0Y57_I;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_B2 = CLBLM_R_X3Y135_SLICE_X3Y135_BQ;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_B3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_B4 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_B5 = CLBLM_R_X3Y138_SLICE_X2Y138_AO6;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_B6 = CLBLM_R_X3Y143_SLICE_X2Y143_AO6;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_C1 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_C2 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_C3 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_C4 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_C5 = 1'b1;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_C4 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_C6 = 1'b1;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_C5 = 1'b1;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_C6 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_D1 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_D2 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_D3 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_D4 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_D5 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_D6 = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_D1 = LIOB33_X0Y71_IOB_X0Y71_I;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_A2 = CLBLM_R_X13Y137_SLICE_X18Y137_AQ;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_A3 = CLBLM_L_X12Y133_SLICE_X17Y133_AQ;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_A5 = CLBLM_L_X10Y135_SLICE_X12Y135_DO6;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_A6 = CLBLM_R_X13Y135_SLICE_X18Y135_BQ;
  assign RIOB33_X105Y161_IOB_X1Y161_O = CLBLM_R_X11Y141_SLICE_X14Y141_CO6;
  assign RIOB33_X105Y161_IOB_X1Y162_O = CLBLM_R_X11Y141_SLICE_X14Y141_CO5;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_B1 = CLBLM_R_X11Y134_SLICE_X14Y134_AQ;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_B2 = CLBLM_L_X12Y133_SLICE_X17Y133_BQ;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_B4 = CLBLM_R_X13Y134_SLICE_X19Y134_DQ;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_B5 = CLBLM_L_X10Y135_SLICE_X12Y135_DO6;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_C1 = 1'b1;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_C2 = 1'b1;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_C3 = 1'b1;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_C4 = 1'b1;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_C5 = 1'b1;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_C6 = 1'b1;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_D1 = 1'b1;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_D2 = 1'b1;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_D3 = 1'b1;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_D4 = 1'b1;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_D5 = 1'b1;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_D6 = 1'b1;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_A1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_A2 = CLBLM_L_X10Y135_SLICE_X12Y135_DO6;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_A3 = CLBLM_L_X12Y133_SLICE_X16Y133_AQ;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_A4 = CLBLM_L_X12Y133_SLICE_X17Y133_BQ;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_A6 = CLBLM_R_X11Y140_SLICE_X14Y140_BQ;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_C4 = CLBLM_L_X10Y144_SLICE_X12Y144_AO6;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_C5 = 1'b1;
  assign LIOB33_X0Y193_IOB_X0Y193_O = LIOB33_X0Y55_IOB_X0Y56_I;
  assign LIOB33_X0Y193_IOB_X0Y194_O = LIOB33_X0Y59_IOB_X0Y60_I;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_B1 = CLBLM_R_X13Y133_SLICE_X18Y133_AQ;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_B2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_B3 = CLBLM_L_X10Y135_SLICE_X12Y135_DO6;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_B5 = CLBLM_L_X12Y133_SLICE_X16Y133_BQ;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_B6 = CLBLM_L_X8Y133_SLICE_X11Y133_CQ;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOI3_X0Y55_ILOGIC_X0Y56_D = LIOB33_X0Y55_IOB_X0Y56_I;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_C1 = CLBLM_R_X11Y131_SLICE_X14Y131_BQ;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_C2 = CLBLM_L_X12Y133_SLICE_X16Y133_AQ;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_C4 = CLBLM_R_X11Y136_SLICE_X15Y136_B5Q;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_C5 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_C6 = 1'b1;
  assign CLBLM_R_X37Y138_SLICE_X57Y138_A6 = 1'b1;
  assign LIOI3_X0Y55_ILOGIC_X0Y55_D = LIOB33_X0Y55_IOB_X0Y55_I;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_X105Y101_ILOGIC_X1Y102_D = RIOB33_X105Y101_IOB_X1Y102_I;
  assign RIOI3_X105Y101_ILOGIC_X1Y101_D = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_D1 = CLBLM_R_X7Y132_SLICE_X9Y132_BQ;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_D2 = CLBLM_L_X12Y137_SLICE_X16Y137_AQ;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_D3 = CLBLM_R_X13Y138_SLICE_X18Y138_BO6;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_D4 = CLBLL_L_X4Y142_SLICE_X4Y142_BO6;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_D5 = 1'b1;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_D6 = 1'b1;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_D2 = CLBLM_R_X11Y135_SLICE_X14Y135_DQ;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_D5 = CLBLM_R_X11Y144_SLICE_X14Y144_DO6;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_D6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_A4 = CLBLM_L_X12Y136_SLICE_X17Y136_A5Q;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_A5 = 1'b1;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_A1 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_A2 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_A3 = CLBLM_R_X3Y139_SLICE_X3Y139_AQ;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_A5 = CLBLM_R_X5Y136_SLICE_X6Y136_DQ;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_A6 = CLBLL_L_X4Y133_SLICE_X5Y133_BO6;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_C4 = 1'b1;
  assign RIOI3_X105Y125_ILOGIC_X1Y126_D = RIOB33_X105Y125_IOB_X1Y126_I;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_C5 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_B1 = CLBLM_R_X3Y141_SLICE_X3Y141_CO6;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_B2 = CLBLM_R_X3Y140_SLICE_X3Y140_BO6;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_B3 = CLBLM_R_X5Y140_SLICE_X6Y140_AO6;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_B4 = CLBLL_L_X4Y139_SLICE_X4Y139_BO6;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_B5 = CLBLL_L_X4Y142_SLICE_X5Y142_DO6;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_B6 = CLBLM_R_X5Y141_SLICE_X7Y141_DO6;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_C6 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_C1 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_C2 = CLBLM_R_X3Y139_SLICE_X2Y139_AO5;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_C3 = CLBLL_L_X4Y137_SLICE_X4Y137_D5Q;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_C4 = CLBLL_L_X2Y140_SLICE_X1Y140_AO5;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_C5 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_C6 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_B4 = CLBLL_L_X4Y134_SLICE_X5Y134_CQ;
  assign RIOI3_X105Y125_ILOGIC_X1Y125_D = RIOB33_X105Y125_IOB_X1Y125_I;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_B5 = CLBLM_L_X12Y143_SLICE_X17Y143_CO5;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_D1 = CLBLM_R_X3Y143_SLICE_X2Y143_AO6;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_D2 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_D3 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_D4 = CLBLM_R_X3Y139_SLICE_X3Y139_AQ;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_D5 = CLBLL_L_X2Y140_SLICE_X1Y140_AO6;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_D6 = CLBLM_L_X8Y140_SLICE_X10Y140_A5Q;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_A1 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_A2 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_A3 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_A4 = CLBLM_L_X8Y140_SLICE_X10Y140_A5Q;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_A5 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_A6 = 1'b1;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_C6 = CLBLM_L_X10Y134_SLICE_X13Y134_AQ;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_B1 = CLBLL_L_X2Y140_SLICE_X1Y140_AO6;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_B2 = CLBLM_R_X3Y143_SLICE_X3Y143_AO5;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_B3 = CLBLM_R_X3Y143_SLICE_X2Y143_AO6;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_B4 = LIOB33_X0Y65_IOB_X0Y65_I;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_B5 = CLBLM_R_X3Y139_SLICE_X2Y139_AO6;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_B6 = CLBLM_R_X3Y139_SLICE_X3Y139_AQ;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_D2 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_C1 = CLBLM_R_X3Y138_SLICE_X2Y138_BO6;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_C2 = CLBLM_R_X3Y139_SLICE_X3Y139_CO6;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_C3 = CLBLM_R_X3Y142_SLICE_X2Y142_AO6;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_C4 = CLBLL_L_X4Y138_SLICE_X4Y138_CO6;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_C5 = CLBLM_R_X3Y139_SLICE_X2Y139_DO6;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_C6 = CLBLM_R_X5Y138_SLICE_X6Y138_AQ;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_C3 = CLBLM_L_X10Y144_SLICE_X13Y144_DO6;
  assign RIOB33_X105Y163_IOB_X1Y163_O = CLBLM_L_X12Y139_SLICE_X17Y139_DO6;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_C4 = CLBLM_R_X11Y143_SLICE_X15Y143_CO6;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_D5 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_D1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_D2 = CLBLM_R_X3Y143_SLICE_X3Y143_AO5;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_D3 = CLBLM_R_X3Y143_SLICE_X3Y143_AO6;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_D4 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_D5 = CLBLL_L_X4Y133_SLICE_X5Y133_AQ;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_D6 = CLBLM_R_X3Y143_SLICE_X2Y143_AO6;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_D6 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_A1 = CLBLM_R_X13Y134_SLICE_X18Y134_DO6;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_A2 = CLBLM_L_X12Y134_SLICE_X16Y134_BO6;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_A3 = CLBLM_L_X12Y138_SLICE_X17Y138_BO5;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_A4 = CLBLM_L_X10Y135_SLICE_X12Y135_DO6;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_A5 = CLBLM_L_X12Y133_SLICE_X16Y133_DO6;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_A6 = CLBLM_L_X12Y134_SLICE_X17Y134_CO6;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_AX = CLBLM_R_X13Y134_SLICE_X18Y134_AO6;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_B1 = CLBLM_R_X13Y134_SLICE_X19Y134_AQ;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_B2 = CLBLM_R_X11Y134_SLICE_X14Y134_CQ;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_B3 = CLBLM_L_X12Y133_SLICE_X16Y133_AQ;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_B4 = CLBLM_L_X12Y135_SLICE_X16Y135_BQ;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_B5 = CLBLM_R_X13Y135_SLICE_X18Y135_AQ;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_B6 = CLBLM_L_X12Y133_SLICE_X17Y133_BQ;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_D2 = CLBLM_R_X7Y134_SLICE_X8Y134_DO6;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_C1 = 1'b1;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_D3 = CLBLM_L_X8Y140_SLICE_X11Y140_AQ;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_C2 = CLBLM_R_X11Y134_SLICE_X14Y134_BQ;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_C3 = CLBLM_L_X8Y134_SLICE_X11Y134_AQ;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_C4 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_C5 = CLBLM_L_X12Y135_SLICE_X17Y135_DO6;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_D4 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_C6 = CLBLM_L_X12Y134_SLICE_X17Y134_DO6;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X37Y138_SLICE_X57Y138_A1 = 1'b1;
  assign CLBLM_R_X37Y138_SLICE_X57Y138_A2 = 1'b1;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_D5 = CLBLM_L_X8Y143_SLICE_X10Y143_DO6;
  assign CLBLM_R_X37Y138_SLICE_X57Y138_A3 = 1'b1;
  assign CLBLM_R_X37Y138_SLICE_X57Y138_A4 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_D1 = 1'b1;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_D6 = CLBLM_L_X10Y136_SLICE_X12Y136_CO5;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_D2 = CLBLM_L_X12Y139_SLICE_X17Y139_CQ;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_D3 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_D4 = CLBLM_R_X11Y134_SLICE_X15Y134_BQ;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_D6 = CLBLM_L_X12Y135_SLICE_X16Y135_BQ;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_D5 = CLBLM_R_X7Y133_SLICE_X9Y133_AQ;
  assign CLBLM_R_X37Y138_SLICE_X57Y138_B1 = 1'b1;
  assign CLBLM_R_X37Y138_SLICE_X57Y138_B2 = 1'b1;
  assign CLBLM_R_X37Y138_SLICE_X57Y138_B3 = 1'b1;
  assign CLBLM_R_X37Y138_SLICE_X57Y138_B4 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_A1 = CLBLM_L_X12Y135_SLICE_X17Y135_CQ;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_A2 = CLBLM_R_X11Y134_SLICE_X15Y134_DO6;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_A3 = CLBLM_L_X12Y135_SLICE_X16Y135_AQ;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_A4 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_A5 = CLBLM_R_X13Y134_SLICE_X19Y134_DQ;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_A6 = CLBLM_L_X12Y134_SLICE_X16Y134_CO6;
  assign CLBLM_R_X37Y138_SLICE_X57Y138_C1 = 1'b1;
  assign CLBLM_R_X37Y138_SLICE_X57Y138_C2 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_AX = CLBLM_L_X12Y133_SLICE_X16Y133_CQ;
  assign CLBLM_R_X37Y138_SLICE_X57Y138_C4 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_B1 = CLBLM_L_X12Y134_SLICE_X16Y134_DO6;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_B2 = CLBLM_R_X11Y134_SLICE_X14Y134_CQ;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_B3 = CLBLM_L_X12Y135_SLICE_X16Y135_AQ;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_B4 = CLBLM_R_X13Y134_SLICE_X19Y134_DQ;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_B5 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_B6 = CLBLM_L_X12Y135_SLICE_X16Y135_CQ;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_D3 = CLBLM_L_X10Y143_SLICE_X12Y143_CQ;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_D4 = CLBLM_R_X11Y142_SLICE_X15Y142_CQ;
  assign CLBLM_R_X37Y138_SLICE_X57Y138_D1 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_C1 = CLBLM_R_X7Y132_SLICE_X9Y132_BQ;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_C2 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_C3 = CLBLM_R_X13Y134_SLICE_X19Y134_CQ;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_C4 = CLBLM_R_X11Y134_SLICE_X15Y134_BQ;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_C5 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_C6 = CLBLM_R_X11Y135_SLICE_X14Y135_BQ;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_CE = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X37Y138_SLICE_X56Y138_A1 = RIOB33_X105Y119_IOB_X1Y119_I;
  assign CLBLM_R_X37Y138_SLICE_X56Y138_A2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X37Y138_SLICE_X56Y138_A3 = 1'b1;
  assign CLBLM_R_X37Y138_SLICE_X56Y138_A4 = 1'b1;
  assign CLBLM_R_X37Y138_SLICE_X56Y138_A5 = 1'b1;
  assign CLBLM_R_X37Y138_SLICE_X56Y138_A6 = CLBLM_L_X8Y138_SLICE_X10Y138_DQ;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_D1 = CLBLM_R_X13Y133_SLICE_X18Y133_AQ;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_A3 = CLBLM_L_X10Y136_SLICE_X12Y136_AQ;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_D2 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_D3 = CLBLM_R_X13Y134_SLICE_X19Y134_CQ;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_D4 = CLBLM_R_X13Y134_SLICE_X19Y134_AQ;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_D5 = 1'b1;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_D6 = CLBLM_R_X11Y135_SLICE_X14Y135_BQ;
  assign CLBLM_R_X37Y138_SLICE_X56Y138_B1 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_SR = CLBLM_L_X12Y144_SLICE_X16Y144_AO6;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_A5 = CLBLM_L_X8Y138_SLICE_X10Y138_AQ;
  assign CLBLM_R_X37Y138_SLICE_X56Y138_B5 = 1'b1;
  assign CLBLM_R_X37Y138_SLICE_X56Y138_B6 = 1'b1;
  assign CLBLM_R_X37Y138_SLICE_X56Y138_C1 = 1'b1;
  assign CLBLM_R_X37Y138_SLICE_X56Y138_C2 = 1'b1;
  assign CLBLM_R_X37Y138_SLICE_X56Y138_C3 = 1'b1;
  assign CLBLM_R_X37Y138_SLICE_X56Y138_C4 = 1'b1;
  assign CLBLM_R_X37Y138_SLICE_X56Y138_C5 = 1'b1;
  assign CLBLM_R_X37Y138_SLICE_X56Y138_C6 = 1'b1;
  assign LIOI3_X0Y111_OLOGIC_X0Y112_T1 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_B5 = CLBLM_L_X8Y144_SLICE_X11Y144_BO6;
  assign CLBLM_R_X37Y138_SLICE_X56Y138_D1 = 1'b1;
  assign CLBLM_R_X37Y138_SLICE_X56Y138_D2 = 1'b1;
  assign CLBLM_R_X37Y138_SLICE_X56Y138_D3 = 1'b1;
  assign CLBLM_R_X37Y138_SLICE_X56Y138_D4 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X37Y138_SLICE_X56Y138_D5 = 1'b1;
  assign CLBLM_R_X37Y138_SLICE_X56Y138_D6 = 1'b1;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_B1 = CLBLM_L_X10Y136_SLICE_X12Y136_DO6;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_B2 = CLBLM_L_X10Y136_SLICE_X12Y136_BQ;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_B3 = CLBLM_L_X10Y136_SLICE_X12Y136_AQ;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_B4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_B5 = CLBLM_L_X8Y138_SLICE_X10Y138_AQ;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_C5 = CLBLM_R_X7Y140_SLICE_X8Y140_AQ;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_D1 = 1'b0;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_C6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_A1 = CLBLM_R_X3Y139_SLICE_X2Y139_BO6;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_A2 = CLBLM_L_X10Y134_SLICE_X12Y134_BQ;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_A3 = CLBLM_R_X3Y140_SLICE_X2Y140_AO6;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_A4 = CLBLL_L_X4Y143_SLICE_X4Y143_BO5;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_A5 = CLBLM_R_X11Y140_SLICE_X15Y140_C5Q;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_A6 = CLBLM_R_X7Y142_SLICE_X9Y142_CO6;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_T1 = 1'b1;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_B1 = CLBLM_R_X3Y141_SLICE_X3Y141_BO6;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_B2 = CLBLM_R_X3Y142_SLICE_X2Y142_DO6;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_B3 = CLBLM_R_X5Y142_SLICE_X6Y142_AO6;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_B4 = CLBLM_R_X5Y140_SLICE_X7Y140_DO6;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_B5 = CLBLM_R_X3Y140_SLICE_X3Y140_AO6;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_B6 = CLBLL_L_X4Y140_SLICE_X5Y140_BO6;
  assign CLBLM_R_X103Y170_SLICE_X162Y170_B4 = 1'b1;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_C1 = CLBLL_L_X2Y140_SLICE_X1Y140_AO5;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_C2 = CLBLM_R_X3Y143_SLICE_X2Y143_AO6;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_C3 = CLBLM_R_X3Y143_SLICE_X3Y143_AO6;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_C4 = CLBLL_L_X4Y143_SLICE_X5Y143_BO5;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_C5 = CLBLL_L_X4Y134_SLICE_X5Y134_BQ;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_C6 = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_D1 = CLBLL_L_X4Y143_SLICE_X4Y143_BO5;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_D2 = 1'b1;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_D3 = CLBLM_L_X10Y134_SLICE_X12Y134_BQ;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_D4 = CLBLM_R_X7Y142_SLICE_X9Y142_CO6;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_D5 = 1'b1;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_D6 = CLBLM_R_X11Y140_SLICE_X15Y140_C5Q;
  assign LIOI3_X0Y179_OLOGIC_X0Y180_D1 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign RIOB33_X105Y165_IOB_X1Y165_O = RIOB33_X105Y125_IOB_X1Y125_I;
  assign RIOB33_X105Y165_IOB_X1Y166_O = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_A1 = CLBLM_R_X3Y143_SLICE_X3Y143_AO6;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_A2 = CLBLM_R_X5Y136_SLICE_X6Y136_AQ;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_A3 = CLBLL_L_X4Y136_SLICE_X4Y136_BQ;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_A4 = CLBLL_L_X2Y141_SLICE_X1Y141_AO6;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_A5 = CLBLM_R_X3Y143_SLICE_X2Y143_AO5;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_A6 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_D1 = CLBLL_L_X4Y133_SLICE_X5Y133_A5Q;
  assign LIOI3_X0Y179_OLOGIC_X0Y180_T1 = 1'b1;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_B1 = LIOB33_X0Y65_IOB_X0Y65_I;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_B2 = CLBLM_R_X5Y143_SLICE_X6Y143_AO6;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_B3 = CLBLM_R_X3Y141_SLICE_X2Y141_AO6;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_B4 = CLBLM_R_X3Y139_SLICE_X3Y139_DO6;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_B5 = CLBLL_L_X4Y136_SLICE_X4Y136_BQ;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_B6 = CLBLM_R_X3Y140_SLICE_X2Y140_CO6;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_T1 = 1'b1;
  assign LIOI3_X0Y179_OLOGIC_X0Y179_D1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign RIOI3_X105Y165_OLOGIC_X1Y166_D1 = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_C1 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_C2 = CLBLM_R_X5Y136_SLICE_X6Y136_AQ;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_C3 = CLBLM_R_X3Y143_SLICE_X2Y143_AO5;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_C4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_C5 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_C6 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_D1 = CLBLM_L_X8Y135_SLICE_X11Y135_B5Q;
  assign LIOI3_X0Y179_OLOGIC_X0Y179_T1 = 1'b1;
  assign RIOI3_X105Y165_OLOGIC_X1Y166_T1 = 1'b1;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_D1 = 1'b1;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_D2 = CLBLM_R_X3Y142_SLICE_X2Y142_DO6;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_D3 = CLBLM_R_X3Y140_SLICE_X3Y140_DO6;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_D4 = CLBLL_L_X4Y140_SLICE_X5Y140_BO6;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_D5 = CLBLM_R_X5Y140_SLICE_X7Y140_DO6;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_D6 = CLBLM_R_X3Y140_SLICE_X2Y140_BO6;
  assign LIOB33_X0Y197_IOB_X0Y197_O = LIOB33_X0Y71_IOB_X0Y72_I;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_A1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_A3 = CLBLM_L_X12Y135_SLICE_X17Y135_AQ;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_A4 = CLBLM_L_X12Y135_SLICE_X16Y135_BQ;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_A5 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_A6 = CLBLM_L_X8Y138_SLICE_X10Y138_AQ;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_AX = CLBLM_L_X12Y135_SLICE_X17Y135_BO6;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_B1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_B2 = CLBLM_L_X8Y138_SLICE_X10Y138_AQ;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_B3 = CLBLM_L_X12Y135_SLICE_X17Y135_CQ;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_B5 = CLBLM_R_X11Y135_SLICE_X15Y135_CO6;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_B6 = 1'b1;
  assign RIOI3_X105Y165_OLOGIC_X1Y165_T1 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_C1 = CLBLM_L_X12Y134_SLICE_X16Y134_AO6;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_C2 = CLBLM_L_X12Y133_SLICE_X16Y133_DO5;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_C3 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_C4 = CLBLM_L_X12Y137_SLICE_X17Y137_CQ;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_C6 = CLBLM_L_X8Y138_SLICE_X10Y138_AQ;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_D1 = CLBLM_L_X12Y133_SLICE_X16Y133_BQ;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_D2 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_D3 = CLBLM_R_X13Y136_SLICE_X18Y136_AQ;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_D4 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_D5 = CLBLM_L_X8Y132_SLICE_X11Y132_BQ;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_D6 = CLBLM_R_X11Y139_SLICE_X14Y139_AQ;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_A1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_A3 = CLBLM_L_X12Y135_SLICE_X16Y135_AQ;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_A4 = CLBLM_L_X8Y138_SLICE_X10Y138_AQ;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_A5 = CLBLL_L_X4Y135_SLICE_X5Y135_AQ;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_A6 = CLBLM_L_X12Y142_SLICE_X16Y142_CQ;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_B1 = CLBLM_R_X13Y136_SLICE_X18Y136_AQ;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_B2 = CLBLM_L_X12Y135_SLICE_X16Y135_BQ;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_B5 = CLBLM_L_X10Y135_SLICE_X12Y135_DO6;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_B6 = CLBLM_L_X8Y136_SLICE_X10Y136_AQ;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_C1 = CLBLM_L_X10Y135_SLICE_X12Y135_DO6;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_C2 = CLBLM_L_X12Y135_SLICE_X16Y135_CQ;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_C3 = CLBLM_R_X11Y140_SLICE_X15Y140_CQ;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_C4 = CLBLM_L_X12Y139_SLICE_X17Y139_CQ;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_C5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_D1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_D2 = CLBLM_L_X12Y135_SLICE_X16Y135_AQ;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_D3 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_D4 = CLBLM_L_X8Y135_SLICE_X11Y135_A5Q;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_D5 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_D6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOB33_SING_X0Y100_IOB_X0Y100_O = CLBLL_L_X2Y133_SLICE_X0Y133_BO6;
  assign LIOI3_X0Y173_OLOGIC_X0Y174_D1 = CLBLM_R_X11Y153_SLICE_X14Y153_AO6;
  assign LIOI3_X0Y59_ILOGIC_X0Y60_D = LIOB33_X0Y59_IOB_X0Y60_I;
  assign LIOI3_X0Y59_ILOGIC_X0Y59_D = LIOB33_X0Y59_IOB_X0Y59_I;
  assign LIOB33_X0Y79_IOB_X0Y80_O = CLBLL_L_X2Y133_SLICE_X0Y133_AO6;
  assign RIOI3_X105Y103_ILOGIC_X1Y104_D = RIOB33_X105Y103_IOB_X1Y104_I;
  assign RIOI3_X105Y103_ILOGIC_X1Y103_D = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_A1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_A2 = CLBLL_L_X4Y143_SLICE_X5Y143_BO6;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_A3 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_A4 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_A5 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_A6 = 1'b1;
  assign LIOI3_X0Y173_OLOGIC_X0Y174_T1 = 1'b1;
  assign RIOB33_X105Y167_IOB_X1Y167_O = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign RIOB33_X105Y167_IOB_X1Y168_O = CLBLM_R_X11Y153_SLICE_X14Y153_AO6;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_B1 = CLBLM_R_X3Y143_SLICE_X3Y143_BO6;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_B2 = CLBLM_R_X3Y141_SLICE_X2Y141_BO6;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_B3 = CLBLM_R_X3Y142_SLICE_X2Y142_AO5;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_B4 = CLBLM_R_X3Y143_SLICE_X3Y143_CO6;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_B5 = CLBLM_R_X3Y141_SLICE_X3Y141_AO6;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_B6 = CLBLM_R_X5Y143_SLICE_X6Y143_BO5;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_C1 = CLBLL_L_X4Y142_SLICE_X5Y142_AO6;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_C2 = CLBLL_L_X4Y141_SLICE_X4Y141_BO6;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_C3 = CLBLM_R_X3Y142_SLICE_X3Y142_CO6;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_C4 = CLBLM_R_X3Y142_SLICE_X3Y142_DO6;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_C5 = CLBLL_L_X4Y140_SLICE_X4Y140_AO6;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_C6 = CLBLM_R_X7Y141_SLICE_X9Y141_DO6;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_D1 = CLBLM_R_X3Y143_SLICE_X2Y143_AO6;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_D2 = CLBLM_R_X3Y142_SLICE_X2Y142_AO5;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_D3 = CLBLM_R_X3Y139_SLICE_X2Y139_AO5;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_D4 = CLBLL_L_X2Y141_SLICE_X1Y141_BO6;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_D5 = CLBLM_R_X3Y143_SLICE_X3Y143_BO6;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_D6 = CLBLL_L_X2Y141_SLICE_X1Y141_AO6;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_A1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_A2 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_A3 = CLBLM_R_X3Y143_SLICE_X2Y143_AO6;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_A4 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_A5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_A6 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_B1 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_B2 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_B3 = CLBLM_R_X3Y139_SLICE_X2Y139_AO5;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_B4 = CLBLL_L_X2Y141_SLICE_X1Y141_AO6;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_B5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_B6 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign LIOI3_X0Y173_OLOGIC_X0Y173_D1 = CLBLM_R_X103Y140_SLICE_X163Y140_AO5;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_C1 = CLBLM_R_X3Y143_SLICE_X2Y143_AO6;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_C2 = CLBLL_L_X2Y141_SLICE_X1Y141_BO6;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_C3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_C4 = CLBLM_R_X3Y139_SLICE_X2Y139_AO5;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_C5 = CLBLM_R_X3Y143_SLICE_X2Y143_AO5;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_C6 = CLBLL_L_X2Y141_SLICE_X1Y141_AO6;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_D1 = CLBLM_R_X3Y141_SLICE_X2Y141_AO6;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_D2 = CLBLM_R_X5Y141_SLICE_X6Y141_A5Q;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_D3 = CLBLL_L_X2Y141_SLICE_X1Y141_CO6;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_D4 = LIOB33_X0Y59_IOB_X0Y59_I;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_D5 = CLBLM_R_X3Y139_SLICE_X2Y139_AO5;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_D6 = CLBLM_R_X3Y141_SLICE_X2Y141_BO6;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_A1 = CLBLM_L_X8Y143_SLICE_X10Y143_DO6;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_A2 = 1'b1;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_A3 = CLBLM_L_X12Y136_SLICE_X17Y136_AQ;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_A5 = CLBLM_R_X11Y138_SLICE_X14Y138_CQ;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_A6 = CLBLM_R_X13Y137_SLICE_X19Y137_CQ;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_AX = CLBLM_L_X12Y136_SLICE_X17Y136_BO6;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_B1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_B3 = CLBLM_L_X12Y137_SLICE_X17Y137_CQ;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_B4 = CLBLM_R_X11Y136_SLICE_X15Y136_AQ;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_B5 = CLBLM_R_X3Y136_SLICE_X3Y136_CQ;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_B6 = 1'b1;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_C2 = CLBLM_L_X12Y136_SLICE_X17Y136_CQ;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_C3 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_C4 = CLBLM_L_X8Y138_SLICE_X10Y138_AQ;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_C5 = CLBLM_R_X11Y136_SLICE_X15Y136_CO6;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_C6 = CLBLM_R_X13Y143_SLICE_X18Y143_BQ;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y173_OLOGIC_X0Y173_T1 = 1'b1;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_D1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_D2 = CLBLM_R_X11Y136_SLICE_X15Y136_B5Q;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_D3 = CLBLM_L_X12Y136_SLICE_X17Y136_DQ;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_D4 = CLBLM_L_X8Y138_SLICE_X10Y138_AQ;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_D5 = CLBLM_R_X11Y136_SLICE_X15Y136_CO6;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_D6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_A1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_A2 = CLBLM_R_X7Y139_SLICE_X8Y139_BQ;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_A3 = CLBLM_R_X13Y135_SLICE_X18Y135_BQ;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_A5 = 1'b1;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_A6 = 1'b1;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_B1 = CLBLM_R_X7Y136_SLICE_X8Y136_CQ;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_B2 = CLBLM_L_X12Y132_SLICE_X16Y132_BQ;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_B4 = CLBLM_L_X12Y138_SLICE_X17Y138_BQ;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_B5 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_B6 = 1'b1;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_C1 = CLBLM_L_X12Y132_SLICE_X16Y132_AQ;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_C2 = CLBLM_L_X12Y138_SLICE_X17Y138_A5Q;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_C3 = CLBLM_L_X10Y130_SLICE_X12Y130_AQ;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_C5 = CLBLM_R_X13Y140_SLICE_X18Y140_CQ;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_C6 = 1'b1;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_D1 = CLBLM_R_X5Y132_SLICE_X7Y132_DO6;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_D2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_D3 = CLBLM_L_X12Y136_SLICE_X16Y136_DQ;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_D4 = CLBLM_L_X12Y132_SLICE_X16Y132_BQ;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_D5 = 1'b1;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_D6 = CLBLM_L_X12Y138_SLICE_X17Y138_BQ;
  assign RIOI3_X105Y191_OLOGIC_X1Y192_T1 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_A1 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_A2 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_A3 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_A4 = CLBLM_R_X3Y133_SLICE_X2Y133_BO6;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_A5 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_A6 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_B1 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_B2 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_B3 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_B4 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_B5 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_B6 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_C1 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_C2 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_C3 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_C4 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_C5 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_C6 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_D1 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_D2 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_D3 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_D4 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_D5 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_D6 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_C3 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_C4 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_C5 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_C6 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_A1 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_A2 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_A3 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_A4 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_A5 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_A6 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_B1 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_B2 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_B3 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_B4 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_B5 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_B6 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_C1 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_C2 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_C3 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_C4 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_C5 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_C6 = 1'b1;
  assign RIOB33_X105Y169_IOB_X1Y169_O = CLBLM_R_X103Y169_SLICE_X163Y169_AO6;
  assign RIOB33_X105Y169_IOB_X1Y170_O = CLBLM_R_X103Y170_SLICE_X163Y170_AO6;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_D1 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_D2 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_D3 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_D4 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_D5 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_D6 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_A1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_A2 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_A3 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_A4 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_A5 = CLBLL_L_X4Y143_SLICE_X5Y143_BO6;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_A6 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_D3 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_D4 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_B1 = CLBLL_L_X4Y143_SLICE_X5Y143_AO5;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_B2 = CLBLM_R_X3Y143_SLICE_X3Y143_BO6;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_B3 = CLBLM_R_X3Y141_SLICE_X3Y141_AO6;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_B4 = CLBLM_R_X3Y142_SLICE_X2Y142_AO5;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_B5 = CLBLL_L_X4Y143_SLICE_X5Y143_AO6;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_B6 = CLBLM_R_X3Y143_SLICE_X3Y143_CO6;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_D5 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_D6 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_C1 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_C2 = CLBLM_R_X3Y143_SLICE_X3Y143_CO6;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_C3 = CLBLM_R_X5Y143_SLICE_X6Y143_BO5;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_C4 = CLBLM_R_X3Y142_SLICE_X3Y142_AO5;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_C5 = CLBLM_R_X3Y143_SLICE_X3Y143_BO6;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_C6 = CLBLM_R_X3Y142_SLICE_X2Y142_AO5;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_D1 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_D2 = CLBLM_R_X3Y143_SLICE_X3Y143_CO6;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_D3 = CLBLM_R_X3Y141_SLICE_X2Y141_BO6;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_D4 = CLBLM_R_X3Y142_SLICE_X3Y142_AO5;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_D5 = CLBLM_R_X3Y143_SLICE_X3Y143_BO6;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_D6 = CLBLM_R_X3Y142_SLICE_X2Y142_AO5;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_A1 = CLBLM_R_X3Y143_SLICE_X2Y143_AO5;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_A2 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_A3 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_A4 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_A5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_A6 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_A1 = CLBLM_R_X11Y139_SLICE_X14Y139_B5Q;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_B1 = CLBLL_L_X4Y143_SLICE_X5Y143_BO5;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_B2 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_B3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_B4 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_B5 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_B6 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_A2 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_A3 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_C1 = CLBLM_R_X3Y141_SLICE_X2Y141_BO6;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_C2 = CLBLM_R_X3Y142_SLICE_X3Y142_AO5;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_C3 = CLBLM_R_X3Y143_SLICE_X3Y143_BO6;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_C4 = CLBLM_R_X3Y141_SLICE_X2Y141_CO6;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_C5 = CLBLL_L_X4Y143_SLICE_X4Y143_BO6;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_C6 = CLBLM_R_X3Y142_SLICE_X2Y142_BO6;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_A4 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_A5 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_A6 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_D1 = CLBLM_R_X3Y142_SLICE_X2Y142_AO5;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_D2 = CLBLM_R_X3Y142_SLICE_X3Y142_AO5;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_D3 = CLBLM_R_X3Y143_SLICE_X3Y143_BO6;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_D4 = CLBLM_R_X3Y143_SLICE_X3Y143_CO6;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_D5 = CLBLM_R_X3Y141_SLICE_X2Y141_BO6;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_D6 = CLBLL_L_X4Y143_SLICE_X4Y143_BO6;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_A1 = CLBLM_L_X8Y138_SLICE_X10Y138_AQ;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_A2 = CLBLM_R_X11Y136_SLICE_X15Y136_AQ;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_A3 = CLBLM_L_X12Y137_SLICE_X17Y137_AQ;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_A5 = CLBLM_R_X7Y136_SLICE_X8Y136_DO6;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_A6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_AX = CLBLM_L_X12Y137_SLICE_X17Y137_BO6;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_B1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_B3 = CLBLM_L_X12Y135_SLICE_X16Y135_CQ;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_B4 = CLBLM_R_X5Y137_SLICE_X7Y137_CQ;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_B5 = CLBLM_R_X13Y137_SLICE_X19Y137_AQ;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_B6 = 1'b1;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_C1 = CLBLM_L_X8Y138_SLICE_X10Y138_AQ;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_C2 = CLBLM_L_X12Y137_SLICE_X17Y137_CQ;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_C3 = CLBLM_R_X11Y139_SLICE_X15Y139_CQ;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_C4 = CLBLM_L_X8Y137_SLICE_X11Y137_CO6;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_C5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_B1 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_B2 = 1'b1;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_B3 = 1'b1;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_D1 = 1'b1;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_D2 = CLBLM_R_X13Y136_SLICE_X18Y136_CQ;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_D3 = CLBLM_R_X13Y137_SLICE_X18Y137_AQ;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_D4 = CLBLM_L_X12Y139_SLICE_X16Y139_CQ;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_D5 = 1'b1;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_D6 = CLBLM_L_X10Y136_SLICE_X13Y136_AO6;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_B4 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_B5 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_B6 = 1'b1;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_A1 = CLBLM_L_X12Y137_SLICE_X16Y137_CQ;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_A2 = CLBLM_L_X8Y138_SLICE_X10Y138_AQ;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_A3 = CLBLM_L_X12Y137_SLICE_X16Y137_AQ;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_A5 = CLBLM_R_X11Y139_SLICE_X14Y139_B5Q;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_A6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_AX = CLBLM_L_X12Y137_SLICE_X16Y137_BO6;
  assign LIOI3_X0Y183_OLOGIC_X0Y184_D1 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_B1 = CLBLM_R_X13Y143_SLICE_X18Y143_AO6;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_B3 = CLBLM_R_X11Y139_SLICE_X15Y139_BQ;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_B4 = CLBLM_L_X8Y135_SLICE_X10Y135_BQ;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_B5 = CLBLM_L_X12Y137_SLICE_X16Y137_A5Q;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_B6 = 1'b1;
  assign LIOI3_X0Y183_OLOGIC_X0Y184_T1 = 1'b1;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_C1 = CLBLM_L_X12Y132_SLICE_X16Y132_AQ;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_C2 = CLBLM_L_X8Y138_SLICE_X10Y138_AQ;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_C3 = CLBLM_L_X12Y137_SLICE_X16Y137_DQ;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_C4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_C5 = CLBLM_L_X12Y137_SLICE_X16Y137_CQ;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_C1 = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_D1 = CLBLL_L_X4Y135_SLICE_X5Y135_D5Q;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_C2 = 1'b1;
  assign LIOI3_X0Y183_OLOGIC_X0Y183_D1 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_T1 = 1'b1;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_D1 = CLBLL_L_X4Y136_SLICE_X4Y136_D5Q;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_D2 = CLBLM_L_X8Y138_SLICE_X10Y138_AQ;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_D3 = CLBLM_L_X12Y137_SLICE_X16Y137_DQ;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_D4 = CLBLM_R_X11Y137_SLICE_X14Y137_DO6;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_D6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_C3 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_C4 = 1'b1;
  assign LIOI3_X0Y183_OLOGIC_X0Y183_T1 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_C5 = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_D1 = CLBLM_R_X7Y132_SLICE_X9Y132_D5Q;
  assign RIOI3_X105Y167_OLOGIC_X1Y168_T1 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_C6 = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_T1 = 1'b1;
  assign RIOI3_X105Y167_OLOGIC_X1Y167_D1 = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_D1 = CLBLL_L_X2Y133_SLICE_X0Y133_CO5;
  assign RIOI3_X105Y167_OLOGIC_X1Y167_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_D1 = CLBLL_L_X2Y108_SLICE_X0Y108_AO6;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_D1 = CLBLM_R_X3Y136_SLICE_X3Y136_AQ;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_D1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_T1 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_D2 = 1'b1;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_B5 = CLBLL_L_X4Y134_SLICE_X5Y134_BQ;
  assign RIOB33_X105Y171_IOB_X1Y172_O = CLBLM_R_X103Y170_SLICE_X163Y170_AO5;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_D3 = 1'b1;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_B6 = CLBLM_L_X8Y134_SLICE_X11Y134_CQ;
  assign RIOB33_X105Y171_IOB_X1Y171_O = CLBLM_L_X10Y146_SLICE_X12Y146_AO5;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_D4 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_D5 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_D6 = 1'b1;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_C2 = CLBLL_L_X4Y134_SLICE_X5Y134_CQ;
  assign CLBLM_R_X13Y141_SLICE_X19Y141_C4 = CLBLM_R_X13Y142_SLICE_X19Y142_CO6;
  assign LIOB33_SING_X0Y149_IOB_X0Y149_O = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X13Y141_SLICE_X19Y141_C5 = CLBLM_R_X13Y142_SLICE_X19Y142_DO6;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_T1 = 1'b1;
  assign CLBLM_R_X13Y141_SLICE_X19Y141_C6 = 1'b1;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_A1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_A2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_A3 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_A4 = 1'b1;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_A5 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_A6 = 1'b1;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_B1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_B2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_B3 = CLBLM_R_X3Y143_SLICE_X2Y143_AO6;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_B4 = CLBLM_R_X3Y143_SLICE_X2Y143_AO5;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_B5 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_B6 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_C1 = CLBLM_R_X3Y143_SLICE_X2Y143_AO6;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_C2 = CLBLM_R_X3Y139_SLICE_X2Y139_AO5;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_C3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_C4 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_C5 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_C6 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_D3 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_D4 = 1'b1;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_D1 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_D2 = CLBLL_L_X4Y143_SLICE_X5Y143_BO6;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_D3 = CLBLM_R_X3Y141_SLICE_X2Y141_BO6;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_D4 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_D5 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_D6 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_D5 = 1'b1;
  assign CLBLM_R_X13Y141_SLICE_X19Y141_D2 = CLBLM_R_X13Y144_SLICE_X18Y144_CO6;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_D6 = 1'b1;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_A1 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_A2 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_A3 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_A4 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_A5 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_A6 = 1'b1;
  assign LIOI3_SING_X0Y50_ILOGIC_X0Y50_D = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_B1 = LIOB33_X0Y57_IOB_X0Y58_I;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_B2 = CLBLL_L_X4Y143_SLICE_X5Y143_CO5;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_B3 = CLBLM_R_X3Y143_SLICE_X2Y143_AO6;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_B4 = LIOB33_X0Y63_IOB_X0Y63_I;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_B5 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_B6 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X13Y141_SLICE_X19Y141_D5 = CLBLM_R_X13Y142_SLICE_X19Y142_DO6;
  assign CLBLM_R_X13Y141_SLICE_X19Y141_D6 = CLBLM_R_X13Y141_SLICE_X19Y141_AQ;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_C1 = 1'b1;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_C2 = 1'b1;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_C3 = 1'b1;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_C4 = 1'b1;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_C5 = 1'b1;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_C6 = 1'b1;
  assign LIOI3_X0Y61_ILOGIC_X0Y62_D = LIOB33_X0Y61_IOB_X0Y62_I;
  assign LIOI3_X0Y61_ILOGIC_X0Y61_D = LIOB33_X0Y61_IOB_X0Y61_I;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_D1 = 1'b1;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_D2 = 1'b1;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_D4 = 1'b1;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_D5 = 1'b1;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_D6 = 1'b1;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_D3 = 1'b1;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_A1 = CLBLM_L_X12Y138_SLICE_X17Y138_AQ;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_A3 = CLBLM_L_X10Y145_SLICE_X12Y145_AQ;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_A4 = CLBLM_L_X10Y139_SLICE_X13Y139_AQ;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_A5 = CLBLM_L_X12Y138_SLICE_X17Y138_CO5;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_A4 = 1'b1;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_AX = CLBLM_L_X12Y139_SLICE_X16Y139_BO6;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_B1 = CLBLM_L_X10Y135_SLICE_X12Y135_DO6;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_B2 = CLBLM_R_X13Y138_SLICE_X18Y138_AQ;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_B3 = CLBLM_L_X12Y138_SLICE_X17Y138_AQ;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_B4 = CLBLM_L_X12Y138_SLICE_X16Y138_BQ;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_B5 = CLBLM_L_X12Y138_SLICE_X16Y138_CQ;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_B6 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_A5 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_A6 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_A1 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_A2 = 1'b1;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_C1 = CLBLM_R_X13Y138_SLICE_X18Y138_AQ;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_C2 = CLBLM_L_X10Y135_SLICE_X12Y135_DO6;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_C3 = CLBLM_L_X12Y138_SLICE_X16Y138_BQ;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_C4 = CLBLM_L_X12Y138_SLICE_X16Y138_CQ;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_C5 = CLBLM_L_X12Y138_SLICE_X17Y138_AQ;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_C6 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_A3 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_A5 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_A6 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_A4 = RIOB33_X105Y123_IOB_X1Y124_I;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_B1 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_B2 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_B3 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_B4 = 1'b1;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_D1 = CLBLM_L_X10Y136_SLICE_X12Y136_BQ;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_D2 = CLBLM_L_X12Y137_SLICE_X17Y137_AQ;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_D3 = CLBLM_L_X12Y137_SLICE_X16Y137_DQ;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_D4 = CLBLM_L_X12Y136_SLICE_X17Y136_DQ;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_D5 = CLBLM_R_X11Y138_SLICE_X14Y138_DQ;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_D6 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_B5 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_B6 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_C1 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_C2 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_C3 = 1'b1;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_A1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_A3 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_A4 = CLBLM_R_X13Y139_SLICE_X18Y139_BO6;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_A5 = CLBLM_L_X12Y138_SLICE_X17Y138_A5Q;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_A6 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_D1 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_D2 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_D4 = 1'b1;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_B1 = CLBLM_L_X12Y138_SLICE_X16Y138_BQ;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_B2 = CLBLM_L_X12Y138_SLICE_X17Y138_BO6;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_B3 = CLBLM_L_X12Y137_SLICE_X16Y137_CQ;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_B5 = CLBLM_L_X10Y145_SLICE_X12Y145_AQ;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_D5 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_D6 = 1'b1;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_C4 = CLBLM_L_X10Y143_SLICE_X13Y143_DO6;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_C1 = CLBLM_L_X10Y145_SLICE_X12Y145_AQ;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_C2 = CLBLM_L_X12Y138_SLICE_X17Y138_CO6;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_C5 = CLBLM_L_X12Y139_SLICE_X16Y139_A5Q;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_C6 = CLBLM_L_X12Y138_SLICE_X16Y138_CQ;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_C6 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_B6 = 1'b1;
  assign RIOI3_X105Y191_OLOGIC_X1Y191_T1 = 1'b1;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_D1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_D2 = CLBLM_L_X12Y137_SLICE_X17Y137_A5Q;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_D3 = CLBLM_R_X11Y138_SLICE_X14Y138_CQ;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_D4 = CLBLM_R_X11Y137_SLICE_X14Y137_BO5;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_D5 = 1'b1;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_D6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_A1 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_A2 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_A3 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_A4 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_A5 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_A6 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_B1 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_B2 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_B3 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_B4 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_B5 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_B6 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_C1 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_C1 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_C2 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_C3 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_C4 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_C5 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_C6 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_C2 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_C3 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_C4 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_D1 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_D2 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_D3 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_D4 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_D5 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_D6 = 1'b1;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_D2 = CLBLM_R_X11Y143_SLICE_X14Y143_CO6;
  assign CLBLM_R_X15Y142_SLICE_X21Y142_A1 = 1'b1;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_D3 = CLBLM_L_X10Y144_SLICE_X13Y144_DO6;
  assign CLBLM_R_X15Y142_SLICE_X21Y142_A2 = 1'b1;
  assign CLBLM_R_X15Y142_SLICE_X21Y142_A3 = 1'b1;
  assign CLBLM_R_X15Y142_SLICE_X21Y142_A4 = 1'b1;
  assign CLBLM_R_X15Y142_SLICE_X21Y142_A5 = 1'b1;
  assign CLBLM_R_X13Y141_SLICE_X18Y141_C4 = CLBLM_R_X13Y140_SLICE_X18Y140_BQ;
  assign CLBLM_R_X15Y142_SLICE_X21Y142_A6 = 1'b1;
  assign CLBLM_R_X15Y142_SLICE_X21Y142_B1 = 1'b1;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_D5 = CLBLM_L_X10Y145_SLICE_X12Y145_CO6;
  assign CLBLM_R_X13Y141_SLICE_X18Y141_C5 = CLBLM_L_X12Y143_SLICE_X17Y143_BQ;
  assign CLBLM_R_X15Y142_SLICE_X21Y142_B2 = 1'b1;
  assign CLBLM_R_X15Y142_SLICE_X21Y142_B3 = 1'b1;
  assign CLBLM_R_X15Y142_SLICE_X21Y142_B4 = 1'b1;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_D6 = CLBLM_R_X11Y143_SLICE_X15Y143_BQ;
  assign CLBLM_R_X13Y141_SLICE_X18Y141_C6 = 1'b1;
  assign CLBLM_R_X15Y142_SLICE_X21Y142_B5 = 1'b1;
  assign CLBLM_R_X15Y142_SLICE_X21Y142_B6 = 1'b1;
  assign CLBLM_R_X15Y142_SLICE_X21Y142_C1 = 1'b1;
  assign CLBLM_R_X15Y142_SLICE_X21Y142_C2 = 1'b1;
  assign CLBLM_R_X15Y142_SLICE_X21Y142_C3 = 1'b1;
  assign CLBLM_R_X15Y142_SLICE_X21Y142_C4 = 1'b1;
  assign CLBLM_R_X15Y142_SLICE_X21Y142_C5 = 1'b1;
  assign CLBLM_R_X15Y142_SLICE_X21Y142_C6 = 1'b1;
  assign CLBLM_R_X15Y142_SLICE_X21Y142_D1 = 1'b1;
  assign CLBLM_R_X15Y142_SLICE_X21Y142_D2 = 1'b1;
  assign CLBLM_R_X15Y142_SLICE_X21Y142_D3 = 1'b1;
  assign CLBLM_R_X15Y142_SLICE_X21Y142_D4 = 1'b1;
  assign CLBLM_R_X15Y142_SLICE_X21Y142_D5 = 1'b1;
  assign CLBLM_R_X15Y142_SLICE_X21Y142_D6 = 1'b1;
  assign CLBLM_R_X15Y142_SLICE_X20Y142_A1 = 1'b1;
  assign CLBLM_R_X15Y142_SLICE_X20Y142_A2 = CLBLM_R_X7Y131_SLICE_X9Y131_AQ;
  assign CLBLM_R_X15Y142_SLICE_X20Y142_A3 = CLBLM_R_X15Y142_SLICE_X20Y142_AQ;
  assign CLBLM_R_X15Y142_SLICE_X20Y142_A4 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X15Y142_SLICE_X20Y142_A5 = CLBLM_R_X13Y142_SLICE_X19Y142_AQ;
  assign CLBLM_R_X15Y142_SLICE_X20Y142_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_D1 = 1'b1;
  assign CLBLM_R_X15Y142_SLICE_X20Y142_B1 = 1'b1;
  assign CLBLM_R_X15Y142_SLICE_X20Y142_B2 = 1'b1;
  assign CLBLM_R_X15Y142_SLICE_X20Y142_B3 = 1'b1;
  assign CLBLM_R_X15Y142_SLICE_X20Y142_B4 = 1'b1;
  assign CLBLM_R_X15Y142_SLICE_X20Y142_B5 = 1'b1;
  assign CLBLM_R_X15Y142_SLICE_X20Y142_B6 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_D2 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_D3 = 1'b1;
  assign CLBLM_R_X15Y142_SLICE_X20Y142_C1 = 1'b1;
  assign CLBLM_R_X15Y142_SLICE_X20Y142_C2 = 1'b1;
  assign CLBLM_R_X15Y142_SLICE_X20Y142_C3 = 1'b1;
  assign CLBLM_R_X15Y142_SLICE_X20Y142_C4 = 1'b1;
  assign CLBLM_R_X15Y142_SLICE_X20Y142_C5 = 1'b1;
  assign CLBLM_R_X15Y142_SLICE_X20Y142_C6 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_D4 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_D5 = 1'b1;
  assign CLBLM_R_X15Y142_SLICE_X20Y142_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_D6 = 1'b1;
  assign CLBLM_R_X15Y142_SLICE_X20Y142_D1 = 1'b1;
  assign CLBLM_R_X15Y142_SLICE_X20Y142_D2 = 1'b1;
  assign CLBLM_R_X15Y142_SLICE_X20Y142_D3 = 1'b1;
  assign CLBLM_R_X15Y142_SLICE_X20Y142_D4 = 1'b1;
  assign CLBLM_R_X15Y142_SLICE_X20Y142_D5 = 1'b1;
  assign CLBLM_R_X15Y142_SLICE_X20Y142_D6 = 1'b1;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_B5 = CLBLM_R_X11Y144_SLICE_X14Y144_AQ;
  assign LIOI3_X0Y197_OLOGIC_X0Y197_D1 = LIOB33_X0Y71_IOB_X0Y72_I;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_B6 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_C5 = CLBLM_R_X11Y138_SLICE_X15Y138_B5Q;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_C6 = CLBLM_L_X8Y137_SLICE_X10Y137_BO6;
  assign LIOI3_X0Y75_ILOGIC_X0Y76_D = LIOB33_X0Y75_IOB_X0Y76_I;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_C4 = CLBLM_R_X11Y144_SLICE_X14Y144_CO6;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_A2 = CLBLM_R_X13Y139_SLICE_X18Y139_AQ;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_A3 = CLBLM_L_X12Y139_SLICE_X17Y139_AQ;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_A4 = CLBLM_L_X8Y138_SLICE_X10Y138_AQ;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_A5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_A6 = CLBLM_L_X10Y135_SLICE_X12Y135_CO6;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_C5 = CLBLM_L_X10Y143_SLICE_X12Y143_CQ;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_C6 = 1'b1;
  assign LIOI3_X0Y197_OLOGIC_X0Y197_T1 = 1'b1;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_B1 = CLBLM_L_X8Y141_SLICE_X10Y141_DQ;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_B4 = CLBLM_L_X12Y140_SLICE_X16Y140_CQ;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_B5 = CLBLM_L_X10Y145_SLICE_X12Y145_AQ;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_B6 = 1'b1;
  assign LIOI3_X0Y75_ILOGIC_X0Y75_D = LIOB33_X0Y75_IOB_X0Y75_I;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_C1 = CLBLM_L_X10Y144_SLICE_X13Y144_AQ;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_D1 = CLBLM_R_X11Y137_SLICE_X14Y137_AQ;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_C2 = CLBLM_L_X12Y139_SLICE_X17Y139_CQ;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_C4 = CLBLM_L_X12Y133_SLICE_X16Y133_BQ;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_D2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_C6 = CLBLM_L_X10Y135_SLICE_X12Y135_DO6;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_D3 = CLBLM_L_X10Y137_SLICE_X13Y137_BQ;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_D1 = CLBLM_R_X11Y138_SLICE_X14Y138_DQ;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_D2 = CLBLM_L_X12Y135_SLICE_X17Y135_A5Q;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_D3 = CLBLL_L_X4Y138_SLICE_X5Y138_B5Q;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_D4 = CLBLM_L_X8Y136_SLICE_X10Y136_BQ;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_D5 = CLBLM_L_X12Y139_SLICE_X17Y139_AQ;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_D6 = 1'b1;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_A1 = 1'b1;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_A2 = CLBLM_L_X12Y134_SLICE_X17Y134_AQ;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_A3 = 1'b1;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_A5 = CLBLM_R_X11Y139_SLICE_X15Y139_BQ;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_A6 = CLBLM_R_X13Y141_SLICE_X18Y141_AO6;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_AX = CLBLM_L_X12Y139_SLICE_X17Y139_BO6;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_B1 = CLBLM_R_X7Y139_SLICE_X8Y139_A5Q;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_B2 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_B3 = CLBLM_L_X12Y139_SLICE_X16Y139_CQ;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_B5 = CLBLM_R_X11Y137_SLICE_X15Y137_AQ;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_B6 = 1'b1;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_D2 = CLBLM_R_X11Y143_SLICE_X15Y143_CO6;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_C2 = 1'b1;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_C3 = 1'b1;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_C4 = CLBLM_L_X12Y140_SLICE_X17Y140_AQ;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_C5 = CLBLM_R_X7Y139_SLICE_X8Y139_A5Q;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_D3 = CLBLM_R_X11Y142_SLICE_X14Y142_AQ;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_D5 = CLBLM_L_X10Y145_SLICE_X12Y145_CO6;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_A1 = CLBLM_L_X8Y137_SLICE_X11Y137_DO6;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_D1 = CLBLM_L_X8Y136_SLICE_X10Y136_DQ;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_D3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_D2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_D4 = CLBLM_L_X12Y139_SLICE_X17Y139_CQ;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_D5 = CLBLM_R_X7Y139_SLICE_X8Y139_BQ;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_D6 = 1'b1;
  assign LIOB33_X0Y123_IOB_X0Y124_O = CLBLL_L_X4Y135_SLICE_X5Y135_D5Q;
  assign RIOB33_X105Y175_IOB_X1Y175_O = CLBLM_L_X12Y146_SLICE_X16Y146_AO6;
  assign RIOB33_X105Y175_IOB_X1Y176_O = CLBLM_R_X103Y173_SLICE_X163Y173_AO5;
  assign LIOB33_X0Y123_IOB_X0Y123_O = CLBLM_R_X7Y132_SLICE_X9Y132_D5Q;
  assign CLBLM_R_X13Y133_SLICE_X19Y133_A1 = 1'b1;
  assign CLBLM_R_X13Y133_SLICE_X19Y133_A2 = 1'b1;
  assign CLBLM_R_X13Y133_SLICE_X19Y133_A3 = 1'b1;
  assign CLBLM_R_X13Y133_SLICE_X19Y133_A4 = 1'b1;
  assign CLBLM_R_X13Y133_SLICE_X19Y133_A5 = 1'b1;
  assign CLBLM_R_X13Y133_SLICE_X19Y133_A6 = 1'b1;
  assign CLBLM_R_X13Y133_SLICE_X19Y133_B1 = 1'b1;
  assign CLBLM_R_X13Y133_SLICE_X19Y133_B2 = 1'b1;
  assign CLBLM_R_X13Y133_SLICE_X19Y133_B3 = 1'b1;
  assign CLBLM_R_X13Y133_SLICE_X19Y133_B4 = 1'b1;
  assign CLBLM_R_X13Y133_SLICE_X19Y133_B5 = 1'b1;
  assign CLBLM_R_X13Y133_SLICE_X19Y133_B6 = 1'b1;
  assign CLBLM_R_X13Y133_SLICE_X19Y133_C1 = 1'b1;
  assign CLBLM_R_X13Y133_SLICE_X19Y133_C2 = 1'b1;
  assign CLBLM_R_X13Y133_SLICE_X19Y133_C3 = 1'b1;
  assign CLBLM_R_X13Y133_SLICE_X19Y133_C4 = 1'b1;
  assign CLBLM_R_X13Y133_SLICE_X19Y133_C5 = 1'b1;
  assign CLBLM_R_X13Y133_SLICE_X19Y133_C6 = 1'b1;
  assign LIOI3_X0Y185_OLOGIC_X0Y186_D1 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_R_X13Y133_SLICE_X19Y133_D1 = 1'b1;
  assign CLBLM_R_X13Y133_SLICE_X19Y133_D2 = 1'b1;
  assign CLBLM_R_X13Y133_SLICE_X19Y133_D3 = 1'b1;
  assign CLBLM_R_X13Y133_SLICE_X19Y133_D4 = 1'b1;
  assign CLBLM_R_X13Y133_SLICE_X19Y133_D5 = 1'b1;
  assign CLBLM_R_X13Y133_SLICE_X19Y133_D6 = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_D1 = CLBLM_R_X3Y136_SLICE_X3Y136_CQ;
  assign LIOI3_X0Y185_OLOGIC_X0Y186_T1 = 1'b1;
  assign CLBLM_R_X13Y133_SLICE_X18Y133_A1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X13Y133_SLICE_X18Y133_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y133_SLICE_X18Y133_A3 = CLBLM_R_X13Y133_SLICE_X18Y133_AQ;
  assign CLBLM_R_X13Y133_SLICE_X18Y133_A4 = CLBLM_L_X10Y142_SLICE_X13Y142_CQ;
  assign CLBLM_R_X13Y133_SLICE_X18Y133_A5 = CLBLM_L_X10Y135_SLICE_X12Y135_DO6;
  assign CLBLM_R_X13Y133_SLICE_X18Y133_A6 = CLBLM_R_X11Y134_SLICE_X14Y134_BQ;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_T1 = 1'b1;
  assign LIOI3_X0Y185_OLOGIC_X0Y185_D1 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign RIOI3_X105Y171_OLOGIC_X1Y172_D1 = CLBLM_R_X103Y170_SLICE_X163Y170_AO5;
  assign CLBLM_R_X13Y133_SLICE_X18Y133_B1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X13Y133_SLICE_X18Y133_B2 = CLBLM_R_X13Y133_SLICE_X18Y133_BQ;
  assign CLBLM_R_X13Y133_SLICE_X18Y133_B3 = CLBLM_R_X11Y131_SLICE_X14Y131_BQ;
  assign CLBLM_R_X13Y133_SLICE_X18Y133_B4 = CLBLM_L_X12Y133_SLICE_X17Y133_AQ;
  assign CLBLM_R_X13Y133_SLICE_X18Y133_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y133_SLICE_X18Y133_B6 = CLBLM_L_X8Y138_SLICE_X10Y138_AQ;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_D1 = CLBLM_R_X11Y138_SLICE_X15Y138_D5Q;
  assign LIOI3_X0Y185_OLOGIC_X0Y185_T1 = 1'b1;
  assign RIOI3_X105Y171_OLOGIC_X1Y172_T1 = 1'b1;
  assign CLBLM_R_X13Y133_SLICE_X18Y133_C1 = 1'b1;
  assign CLBLM_R_X13Y133_SLICE_X18Y133_C2 = 1'b1;
  assign CLBLM_R_X13Y133_SLICE_X18Y133_C3 = 1'b1;
  assign CLBLM_R_X13Y133_SLICE_X18Y133_C4 = 1'b1;
  assign CLBLM_R_X13Y133_SLICE_X18Y133_C5 = 1'b1;
  assign CLBLM_R_X13Y133_SLICE_X18Y133_C6 = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_T1 = 1'b1;
  assign CLBLM_R_X13Y133_SLICE_X18Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_X105Y171_OLOGIC_X1Y171_D1 = CLBLM_L_X10Y146_SLICE_X12Y146_AO5;
  assign CLBLM_R_X13Y133_SLICE_X18Y133_D1 = 1'b1;
  assign CLBLM_R_X13Y133_SLICE_X18Y133_D2 = 1'b1;
  assign CLBLM_R_X13Y133_SLICE_X18Y133_D3 = 1'b1;
  assign CLBLM_R_X13Y133_SLICE_X18Y133_D4 = 1'b1;
  assign CLBLM_R_X13Y133_SLICE_X18Y133_D5 = 1'b1;
  assign CLBLM_R_X13Y133_SLICE_X18Y133_D6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_D1 = CLBLM_L_X12Y136_SLICE_X16Y136_BQ;
  assign RIOI3_X105Y171_OLOGIC_X1Y171_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_D1 = CLBLM_L_X10Y135_SLICE_X13Y135_BQ;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_T1 = 1'b1;
  assign LIOB33_SING_X0Y150_IOB_X0Y150_O = LIOB33_X0Y63_IOB_X0Y63_I;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_A1 = CLBLM_L_X12Y140_SLICE_X17Y140_DO6;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_A2 = CLBLM_L_X8Y134_SLICE_X11Y134_BQ;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_A3 = 1'b1;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_A5 = CLBLM_L_X12Y143_SLICE_X17Y143_DO6;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_A6 = CLBLM_R_X13Y141_SLICE_X18Y141_AO5;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_B1 = CLBLM_L_X12Y142_SLICE_X16Y142_CQ;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_B3 = CLBLM_R_X13Y143_SLICE_X18Y143_AO6;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_B4 = CLBLM_L_X12Y143_SLICE_X17Y143_CO5;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_B5 = CLBLM_L_X8Y141_SLICE_X11Y141_CQ;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_B6 = CLBLM_L_X12Y140_SLICE_X17Y140_BQ;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_A1 = CLBLL_L_X4Y135_SLICE_X5Y135_CQ;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_A2 = CLBLM_R_X11Y131_SLICE_X15Y131_BQ;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_A3 = CLBLM_L_X8Y131_SLICE_X11Y131_BQ;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_A4 = CLBLM_L_X10Y131_SLICE_X12Y131_BQ;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_A5 = CLBLM_L_X10Y130_SLICE_X12Y130_AQ;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_A6 = 1'b1;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_C1 = CLBLM_R_X13Y143_SLICE_X18Y143_AO6;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_C2 = CLBLM_L_X12Y140_SLICE_X17Y140_CQ;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_C3 = CLBLM_L_X12Y136_SLICE_X16Y136_AQ;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_B1 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_B2 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_B3 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_B4 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_B5 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_B6 = 1'b1;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_D4 = CLBLM_L_X12Y140_SLICE_X17Y140_BQ;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_C1 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_C2 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_C3 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_C4 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_C5 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_C6 = 1'b1;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_D5 = CLBLM_L_X12Y140_SLICE_X17Y140_AQ;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_D6 = 1'b1;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_A1 = CLBLM_L_X8Y143_SLICE_X10Y143_DO6;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_A2 = CLBLM_L_X12Y138_SLICE_X16Y138_DQ;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_A3 = CLBLM_L_X12Y140_SLICE_X16Y140_AQ;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_A5 = CLBLM_R_X13Y135_SLICE_X18Y135_AQ;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_A6 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_D1 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_D2 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_D3 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_D4 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_D5 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_D6 = 1'b1;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_B1 = CLBLM_L_X12Y143_SLICE_X16Y143_CQ;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_B2 = CLBLM_L_X12Y140_SLICE_X16Y140_BQ;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_B3 = CLBLM_R_X13Y143_SLICE_X18Y143_AO6;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_B4 = CLBLM_R_X5Y138_SLICE_X7Y138_AQ;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_A1 = CLBLM_L_X10Y130_SLICE_X12Y130_BO5;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_A2 = CLBLM_L_X12Y132_SLICE_X17Y132_AQ;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_A3 = CLBLM_L_X10Y130_SLICE_X12Y130_AQ;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_A6 = CLBLM_R_X11Y140_SLICE_X15Y140_CQ;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_C1 = CLBLM_L_X8Y140_SLICE_X10Y140_AQ;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_C2 = 1'b1;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_C3 = CLBLM_L_X12Y141_SLICE_X16Y141_BQ;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_B1 = CLBLL_L_X4Y135_SLICE_X5Y135_CQ;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_B2 = CLBLM_L_X10Y131_SLICE_X12Y131_BQ;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_B3 = CLBLM_L_X10Y130_SLICE_X12Y130_AQ;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_B4 = CLBLM_R_X11Y131_SLICE_X15Y131_BQ;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_B5 = CLBLM_R_X5Y132_SLICE_X7Y132_DO6;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_B6 = 1'b1;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_D1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_D2 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_C1 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_C2 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_C3 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_C4 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_C5 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_C6 = 1'b1;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_D3 = CLBLM_L_X12Y139_SLICE_X16Y139_BO5;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_D4 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_D5 = CLBLM_L_X12Y139_SLICE_X16Y139_AQ;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_D6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOI3_X0Y65_ILOGIC_X0Y65_D = LIOB33_X0Y65_IOB_X0Y65_I;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_D1 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_D2 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_D3 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_D4 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_D5 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_D6 = 1'b1;
  assign RIOI3_X105Y109_ILOGIC_X1Y110_D = RIOB33_X105Y109_IOB_X1Y110_I;
  assign RIOI3_X105Y109_ILOGIC_X1Y109_D = RIOB33_X105Y109_IOB_X1Y109_I;
  assign RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y138_D = RIOB33_X105Y137_IOB_X1Y138_I;
  assign RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y137_D = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_A2 = CLBLM_R_X13Y134_SLICE_X19Y134_BQ;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_A3 = CLBLM_R_X13Y134_SLICE_X19Y134_AQ;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_A4 = CLBLM_L_X10Y135_SLICE_X12Y135_DO6;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_A6 = CLBLM_R_X13Y134_SLICE_X18Y134_CO6;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_B2 = CLBLM_R_X13Y134_SLICE_X19Y134_BQ;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_B3 = CLBLM_L_X12Y136_SLICE_X16Y136_B5Q;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_B4 = 1'b1;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_B5 = CLBLM_R_X7Y131_SLICE_X9Y131_AQ;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_B6 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_C1 = CLBLM_L_X8Y134_SLICE_X10Y134_AQ;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_C2 = CLBLM_R_X13Y134_SLICE_X19Y134_CQ;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_C4 = CLBLM_L_X12Y140_SLICE_X16Y140_BQ;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_C5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_C6 = CLBLM_L_X8Y138_SLICE_X10Y138_AQ;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_D1 = CLBLM_R_X13Y139_SLICE_X19Y139_AQ;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_D2 = CLBLM_R_X13Y133_SLICE_X18Y133_BQ;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_D3 = CLBLM_R_X13Y134_SLICE_X19Y134_DQ;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_D4 = CLBLM_L_X8Y138_SLICE_X10Y138_AQ;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_D5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_D6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_A2 = CLBLM_L_X12Y139_SLICE_X17Y139_CQ;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_A3 = CLBLM_R_X13Y133_SLICE_X18Y133_AQ;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_A4 = CLBLM_L_X12Y134_SLICE_X17Y134_AO6;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_A5 = CLBLM_L_X12Y133_SLICE_X16Y133_BQ;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_A6 = 1'b1;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_B1 = CLBLM_R_X13Y135_SLICE_X18Y135_BQ;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_B2 = CLBLM_L_X12Y139_SLICE_X17Y139_CQ;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_B3 = CLBLM_L_X12Y134_SLICE_X17Y134_BO6;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_B4 = CLBLM_L_X12Y133_SLICE_X16Y133_BQ;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_B5 = CLBLM_R_X13Y133_SLICE_X18Y133_AQ;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_B6 = CLBLM_R_X13Y135_SLICE_X18Y135_CO6;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_C1 = CLBLM_L_X12Y133_SLICE_X17Y133_AQ;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_C2 = CLBLM_R_X13Y135_SLICE_X18Y135_BQ;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_C3 = CLBLM_L_X12Y133_SLICE_X16Y133_DO6;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_C4 = CLBLM_L_X12Y138_SLICE_X17Y138_BO5;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_C5 = 1'b1;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_C6 = CLBLM_R_X13Y134_SLICE_X18Y134_BO6;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_D1 = CLBLM_L_X12Y134_SLICE_X17Y134_BO6;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_D2 = CLBLM_R_X13Y135_SLICE_X18Y135_CO6;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_D3 = CLBLM_R_X13Y135_SLICE_X18Y135_BQ;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_D4 = CLBLM_R_X13Y134_SLICE_X18Y134_AO5;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_D5 = 1'b1;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_D6 = CLBLM_L_X12Y133_SLICE_X17Y133_AQ;
  assign LIOB33_X0Y139_IOB_X0Y140_O = CLBLM_R_X3Y136_SLICE_X2Y136_AQ;
  assign LIOB33_X0Y139_IOB_X0Y139_O = CLBLM_R_X3Y137_SLICE_X2Y137_AQ;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_AX = CLBLM_L_X10Y133_SLICE_X12Y133_BQ;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_A1 = CLBLM_R_X13Y140_SLICE_X18Y140_BQ;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_A3 = CLBLM_R_X13Y140_SLICE_X19Y140_AQ;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_A4 = CLBLM_L_X12Y142_SLICE_X16Y142_BQ;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_A5 = CLBLM_R_X13Y144_SLICE_X18Y144_AQ;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_A6 = CLBLM_L_X12Y143_SLICE_X17Y143_BQ;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_B1 = CLBLM_L_X12Y142_SLICE_X17Y142_AQ;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_B2 = CLBLM_L_X12Y142_SLICE_X16Y142_BQ;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_B3 = 1'b1;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_B4 = CLBLM_R_X13Y140_SLICE_X18Y140_BQ;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_B5 = CLBLM_R_X13Y144_SLICE_X18Y144_AQ;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_B6 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_A1 = CLBLM_R_X5Y133_SLICE_X7Y133_DO6;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_A3 = CLBLM_L_X10Y131_SLICE_X13Y131_AQ;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_A4 = CLBLM_R_X11Y132_SLICE_X14Y132_AQ;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_A5 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_A6 = CLBLM_R_X11Y133_SLICE_X15Y133_CQ;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_C1 = CLBLM_L_X12Y143_SLICE_X17Y143_AQ;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_C2 = CLBLM_R_X13Y140_SLICE_X18Y140_CQ;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_C3 = CLBLM_R_X13Y141_SLICE_X18Y141_CO6;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_B1 = CLBLM_L_X10Y131_SLICE_X13Y131_CQ;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_B2 = CLBLM_L_X10Y131_SLICE_X13Y131_BQ;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_B3 = CLBLM_L_X10Y131_SLICE_X13Y131_AQ;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_B5 = CLBLM_R_X5Y132_SLICE_X7Y132_DO6;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_B6 = 1'b1;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_D1 = CLBLM_R_X13Y144_SLICE_X18Y144_AQ;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_C1 = CLBLM_L_X10Y133_SLICE_X13Y133_AQ;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_C2 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_C3 = CLBLM_L_X8Y131_SLICE_X11Y131_AQ;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_C4 = CLBLM_R_X5Y132_SLICE_X7Y132_DO6;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_C5 = CLBLM_L_X10Y131_SLICE_X13Y131_CQ;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_D3 = CLBLM_R_X13Y140_SLICE_X18Y140_BQ;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_D4 = CLBLM_L_X12Y142_SLICE_X16Y142_BQ;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_A1 = CLBLM_L_X12Y141_SLICE_X16Y141_DO6;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_A2 = CLBLM_L_X12Y143_SLICE_X17Y143_DO6;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_A4 = CLBLM_R_X13Y141_SLICE_X18Y141_AO5;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_A5 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_D1 = CLBLM_R_X11Y131_SLICE_X14Y131_AO6;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_D2 = CLBLM_R_X3Y139_SLICE_X3Y139_BO6;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_D3 = CLBLM_R_X5Y133_SLICE_X7Y133_CO6;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_D4 = CLBLM_L_X8Y135_SLICE_X11Y135_AQ;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_D5 = CLBLM_L_X12Y136_SLICE_X16Y136_B5Q;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_D6 = CLBLM_L_X10Y131_SLICE_X12Y131_AO6;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_A6 = CLBLM_L_X8Y141_SLICE_X10Y141_DQ;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_B1 = CLBLM_R_X13Y140_SLICE_X18Y140_BQ;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_B2 = CLBLM_L_X12Y142_SLICE_X16Y142_BQ;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_B3 = CLBLM_L_X12Y139_SLICE_X16Y139_AQ;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_A1 = CLBLM_R_X11Y131_SLICE_X15Y131_BQ;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_A2 = CLBLM_L_X10Y131_SLICE_X12Y131_BQ;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_A3 = CLBLM_L_X10Y133_SLICE_X13Y133_AQ;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_A4 = CLBLL_L_X4Y135_SLICE_X5Y135_CQ;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_A5 = CLBLM_L_X10Y130_SLICE_X12Y130_AQ;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_A6 = 1'b1;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_C1 = CLBLM_R_X13Y144_SLICE_X18Y144_AQ;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_C2 = CLBLM_L_X12Y140_SLICE_X17Y140_AQ;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_C3 = CLBLM_L_X12Y142_SLICE_X17Y142_AQ;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_B2 = CLBLM_L_X10Y131_SLICE_X12Y131_BQ;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_B4 = CLBLM_R_X11Y140_SLICE_X15Y140_CQ;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_B5 = CLBLM_L_X10Y130_SLICE_X12Y130_BO6;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_B6 = CLBLM_L_X8Y131_SLICE_X10Y131_A5Q;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_D1 = CLBLM_R_X11Y140_SLICE_X14Y140_AQ;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_D2 = CLBLM_R_X13Y141_SLICE_X18Y141_BO5;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_C1 = CLBLM_L_X10Y130_SLICE_X12Y130_AQ;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_C2 = CLBLL_L_X4Y135_SLICE_X5Y135_CQ;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_C3 = CLBLM_L_X10Y131_SLICE_X12Y131_BQ;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_C4 = CLBLM_L_X8Y131_SLICE_X10Y131_A5Q;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_C5 = CLBLM_R_X11Y131_SLICE_X15Y131_BQ;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_C6 = 1'b1;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_D3 = CLBLM_R_X13Y144_SLICE_X18Y144_CO6;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_D4 = CLBLM_L_X12Y141_SLICE_X16Y141_CO6;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_D6 = CLBLM_L_X12Y141_SLICE_X16Y141_AQ;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_D1 = CLBLM_L_X10Y133_SLICE_X13Y133_AQ;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_D2 = CLBLM_L_X8Y135_SLICE_X11Y135_AQ;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_D3 = CLBLM_R_X5Y132_SLICE_X7Y132_DO6;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_D4 = CLBLM_L_X10Y131_SLICE_X12Y131_CO6;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_D5 = CLBLM_L_X10Y131_SLICE_X12Y131_AO5;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_D6 = CLBLM_L_X8Y133_SLICE_X11Y133_CQ;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_B2 = 1'b1;
  assign CLBLM_R_X13Y135_SLICE_X19Y135_A1 = 1'b1;
  assign CLBLM_R_X13Y135_SLICE_X19Y135_A2 = 1'b1;
  assign CLBLM_R_X13Y135_SLICE_X19Y135_A3 = 1'b1;
  assign CLBLM_R_X13Y135_SLICE_X19Y135_A4 = 1'b1;
  assign CLBLM_R_X13Y135_SLICE_X19Y135_A5 = 1'b1;
  assign CLBLM_R_X13Y135_SLICE_X19Y135_A6 = 1'b1;
  assign CLBLM_R_X13Y135_SLICE_X19Y135_B1 = 1'b1;
  assign CLBLM_R_X13Y135_SLICE_X19Y135_B2 = 1'b1;
  assign CLBLM_R_X13Y135_SLICE_X19Y135_B3 = 1'b1;
  assign CLBLM_R_X13Y135_SLICE_X19Y135_B4 = 1'b1;
  assign CLBLM_R_X13Y135_SLICE_X19Y135_B5 = 1'b1;
  assign CLBLM_R_X13Y135_SLICE_X19Y135_B6 = 1'b1;
  assign CLBLM_R_X13Y135_SLICE_X19Y135_C1 = 1'b1;
  assign CLBLM_R_X13Y135_SLICE_X19Y135_C2 = 1'b1;
  assign CLBLM_R_X13Y135_SLICE_X19Y135_C3 = 1'b1;
  assign CLBLM_R_X13Y135_SLICE_X19Y135_C4 = 1'b1;
  assign CLBLM_R_X13Y135_SLICE_X19Y135_C5 = 1'b1;
  assign CLBLM_R_X13Y135_SLICE_X19Y135_C6 = 1'b1;
  assign CLBLM_R_X13Y135_SLICE_X19Y135_D1 = 1'b1;
  assign CLBLM_R_X13Y135_SLICE_X19Y135_D2 = 1'b1;
  assign CLBLM_R_X13Y135_SLICE_X19Y135_D3 = 1'b1;
  assign CLBLM_R_X13Y135_SLICE_X19Y135_D4 = 1'b1;
  assign CLBLM_R_X13Y135_SLICE_X19Y135_D5 = 1'b1;
  assign CLBLM_R_X13Y135_SLICE_X19Y135_D6 = 1'b1;
  assign CLBLM_R_X13Y135_SLICE_X18Y135_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y135_SLICE_X18Y135_A2 = CLBLM_L_X8Y136_SLICE_X11Y136_BQ;
  assign CLBLM_R_X13Y135_SLICE_X18Y135_A3 = CLBLM_R_X13Y135_SLICE_X18Y135_AQ;
  assign CLBLM_R_X13Y135_SLICE_X18Y135_A4 = CLBLM_L_X10Y135_SLICE_X12Y135_DO6;
  assign CLBLM_R_X13Y135_SLICE_X18Y135_A5 = CLBLM_L_X12Y133_SLICE_X16Y133_AQ;
  assign CLBLM_R_X13Y135_SLICE_X18Y135_A6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X13Y135_SLICE_X18Y135_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y135_SLICE_X18Y135_B2 = CLBLM_R_X13Y135_SLICE_X18Y135_BQ;
  assign CLBLM_R_X13Y135_SLICE_X18Y135_B3 = CLBLM_R_X13Y135_SLICE_X18Y135_AQ;
  assign CLBLM_R_X13Y135_SLICE_X18Y135_B4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X13Y135_SLICE_X18Y135_B5 = CLBLM_R_X11Y134_SLICE_X15Y134_AQ;
  assign CLBLM_R_X13Y135_SLICE_X18Y135_B6 = CLBLM_L_X10Y135_SLICE_X12Y135_DO6;
  assign CLBLM_R_X13Y135_SLICE_X18Y135_C1 = CLBLM_R_X11Y134_SLICE_X14Y134_AQ;
  assign CLBLM_R_X13Y135_SLICE_X18Y135_C2 = 1'b1;
  assign CLBLM_R_X13Y135_SLICE_X18Y135_C3 = 1'b1;
  assign CLBLM_R_X13Y135_SLICE_X18Y135_C4 = CLBLM_R_X11Y134_SLICE_X14Y134_BQ;
  assign CLBLM_R_X13Y135_SLICE_X18Y135_C5 = CLBLM_L_X12Y135_SLICE_X16Y135_CQ;
  assign CLBLM_R_X13Y135_SLICE_X18Y135_C6 = CLBLM_R_X13Y136_SLICE_X18Y136_AQ;
  assign CLBLM_R_X13Y135_SLICE_X18Y135_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y135_SLICE_X18Y135_D1 = 1'b1;
  assign CLBLM_R_X13Y135_SLICE_X18Y135_D2 = 1'b1;
  assign CLBLM_R_X13Y135_SLICE_X18Y135_D3 = 1'b1;
  assign CLBLM_R_X13Y135_SLICE_X18Y135_D4 = 1'b1;
  assign CLBLM_R_X13Y135_SLICE_X18Y135_D5 = 1'b1;
  assign CLBLM_R_X13Y135_SLICE_X18Y135_D6 = 1'b1;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_C5 = CLBLM_R_X11Y142_SLICE_X15Y142_CQ;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_D1 = 1'b1;
  assign LIOI3_X0Y189_OLOGIC_X0Y190_D1 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign LIOI3_X0Y189_OLOGIC_X0Y190_T1 = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_D1 = CLBLL_L_X4Y134_SLICE_X5Y134_A5Q;
  assign LIOI3_X0Y189_OLOGIC_X0Y189_D1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_T1 = 1'b1;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_A1 = CLBLM_L_X12Y143_SLICE_X17Y143_DO6;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_A3 = CLBLM_R_X11Y141_SLICE_X15Y141_AQ;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_A4 = CLBLM_L_X12Y142_SLICE_X17Y142_DO6;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_A5 = 1'b1;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_A6 = CLBLM_R_X13Y141_SLICE_X18Y141_AO5;
  assign LIOI3_X0Y189_OLOGIC_X0Y189_T1 = 1'b1;
  assign RIOI3_X105Y173_OLOGIC_X1Y174_D1 = CLBLM_R_X103Y173_SLICE_X163Y173_AO6;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_B1 = CLBLM_L_X12Y143_SLICE_X17Y143_DO6;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_B2 = CLBLM_L_X12Y142_SLICE_X17Y142_BQ;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_B4 = CLBLM_L_X10Y141_SLICE_X13Y141_BQ;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_B5 = CLBLM_R_X13Y142_SLICE_X18Y142_BO6;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_B6 = CLBLM_R_X13Y141_SLICE_X18Y141_AO5;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_A1 = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_D1 = CLBLM_R_X5Y137_SLICE_X6Y137_BQ;
  assign RIOB33_X105Y181_IOB_X1Y181_O = CLBLM_L_X12Y138_SLICE_X17Y138_DO5;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_A1 = CLBLM_L_X10Y131_SLICE_X13Y131_DO6;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_A2 = CLBLM_R_X11Y131_SLICE_X14Y131_CO6;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_A3 = CLBLM_L_X10Y132_SLICE_X12Y132_CO6;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_A4 = CLBLM_L_X10Y132_SLICE_X13Y132_BO6;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_A5 = CLBLM_L_X8Y132_SLICE_X10Y132_CO6;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_A6 = CLBLM_L_X10Y132_SLICE_X13Y132_CO6;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_C1 = CLBLM_L_X12Y143_SLICE_X17Y143_AQ;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_C2 = CLBLM_R_X13Y144_SLICE_X18Y144_AQ;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_C3 = CLBLM_R_X13Y140_SLICE_X19Y140_AQ;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_B1 = CLBLM_L_X10Y137_SLICE_X12Y137_B5Q;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_B2 = CLBLM_L_X10Y133_SLICE_X12Y133_DO5;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_B3 = CLBLM_L_X10Y130_SLICE_X13Y130_AO6;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_B4 = CLBLM_R_X3Y139_SLICE_X3Y139_BO6;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_B5 = CLBLM_R_X5Y133_SLICE_X7Y133_CO6;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_B6 = CLBLM_L_X10Y141_SLICE_X12Y141_CQ;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_D1 = CLBLM_L_X12Y140_SLICE_X17Y140_CQ;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_C1 = CLBLM_R_X5Y133_SLICE_X7Y133_CO6;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_C2 = CLBLM_L_X10Y137_SLICE_X12Y137_CQ;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_C3 = CLBLM_L_X10Y134_SLICE_X13Y134_B5Q;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_C4 = CLBLM_R_X5Y136_SLICE_X7Y136_DO6;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_C5 = CLBLM_R_X7Y133_SLICE_X9Y133_DO6;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_C6 = CLBLM_R_X11Y132_SLICE_X15Y132_AO6;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_D3 = CLBLM_L_X12Y142_SLICE_X17Y142_AQ;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_D4 = CLBLM_R_X13Y141_SLICE_X18Y141_BO5;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_A1 = CLBLM_L_X12Y142_SLICE_X16Y142_DO6;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_D6 = CLBLM_R_X13Y144_SLICE_X18Y144_CO6;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_A2 = CLBLM_R_X11Y144_SLICE_X15Y144_BQ;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_A3 = CLBLM_L_X12Y142_SLICE_X16Y142_AQ;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_A4 = CLBLM_L_X12Y143_SLICE_X17Y143_DO6;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_D1 = CLBLM_R_X11Y134_SLICE_X15Y134_CQ;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_D2 = CLBLM_L_X10Y141_SLICE_X12Y141_CQ;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_D3 = CLBLM_L_X10Y132_SLICE_X12Y132_DO6;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_D4 = CLBLM_R_X11Y133_SLICE_X15Y133_CQ;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_D5 = CLBLM_L_X10Y134_SLICE_X13Y134_B5Q;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_D6 = 1'b1;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_AX = CLBLM_L_X12Y139_SLICE_X16Y139_DO6;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_B4 = CLBLM_R_X13Y141_SLICE_X19Y141_CO6;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_B5 = CLBLM_R_X13Y140_SLICE_X18Y140_BQ;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_B2 = CLBLM_L_X12Y142_SLICE_X16Y142_BQ;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_B3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_A1 = CLBLM_L_X8Y134_SLICE_X11Y134_BQ;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_A2 = CLBLM_L_X12Y136_SLICE_X16Y136_CQ;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_A3 = CLBLM_L_X10Y132_SLICE_X13Y132_DO6;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_A4 = CLBLM_L_X10Y132_SLICE_X12Y132_BO6;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_A5 = CLBLM_L_X8Y131_SLICE_X11Y131_DO6;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_A6 = CLBLM_L_X12Y136_SLICE_X16Y136_B5Q;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_C1 = CLBLM_L_X10Y142_SLICE_X12Y142_AQ;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_C2 = CLBLM_L_X12Y142_SLICE_X16Y142_CQ;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_B1 = CLBLM_L_X10Y133_SLICE_X12Y133_CQ;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_B2 = CLBLM_L_X12Y136_SLICE_X16Y136_CQ;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_B3 = CLBLM_L_X10Y133_SLICE_X12Y133_BQ;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_B4 = CLBLM_L_X8Y132_SLICE_X11Y132_DO6;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_B5 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_B6 = CLBLM_R_X5Y132_SLICE_X7Y132_BO5;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_D1 = CLBLM_L_X12Y142_SLICE_X17Y142_AQ;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_D2 = CLBLM_R_X13Y141_SLICE_X18Y141_BO5;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_C1 = CLBLM_L_X10Y131_SLICE_X12Y131_CO5;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_C2 = CLBLM_R_X5Y133_SLICE_X7Y133_CO6;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_C3 = CLBLM_R_X5Y136_SLICE_X7Y136_DO6;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_C4 = CLBLM_R_X11Y146_SLICE_X14Y146_AQ;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_C5 = CLBLM_R_X7Y133_SLICE_X9Y133_DO6;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_C6 = 1'b1;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_D3 = CLBLM_R_X13Y141_SLICE_X18Y141_CO5;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_D4 = CLBLM_L_X12Y140_SLICE_X17Y140_AQ;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_D5 = CLBLM_R_X11Y140_SLICE_X14Y140_BQ;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_D6 = CLBLM_R_X13Y144_SLICE_X18Y144_CO6;
  assign CLBLM_R_X103Y170_SLICE_X163Y170_A5 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_R_X103Y170_SLICE_X163Y170_A6 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_D1 = CLBLM_L_X10Y133_SLICE_X12Y133_AQ;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_D2 = CLBLM_L_X10Y134_SLICE_X12Y134_AQ;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_D3 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_D4 = CLBLM_R_X7Y134_SLICE_X8Y134_C5Q;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_D5 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_D6 = CLBLM_R_X13Y137_SLICE_X18Y137_A5Q;
  assign CLBLM_R_X103Y170_SLICE_X163Y170_B4 = 1'b1;
  assign CLBLM_R_X13Y136_SLICE_X19Y136_A1 = 1'b1;
  assign CLBLM_R_X13Y136_SLICE_X19Y136_A2 = 1'b1;
  assign CLBLM_R_X13Y136_SLICE_X19Y136_A3 = 1'b1;
  assign CLBLM_R_X13Y136_SLICE_X19Y136_A4 = 1'b1;
  assign CLBLM_R_X13Y136_SLICE_X19Y136_A5 = 1'b1;
  assign CLBLM_R_X13Y136_SLICE_X19Y136_A6 = 1'b1;
  assign CLBLM_R_X13Y136_SLICE_X19Y136_B1 = 1'b1;
  assign CLBLM_R_X13Y136_SLICE_X19Y136_B2 = 1'b1;
  assign CLBLM_R_X13Y136_SLICE_X19Y136_B3 = 1'b1;
  assign CLBLM_R_X13Y136_SLICE_X19Y136_B4 = 1'b1;
  assign CLBLM_R_X13Y136_SLICE_X19Y136_B5 = 1'b1;
  assign CLBLM_R_X13Y136_SLICE_X19Y136_B6 = 1'b1;
  assign CLBLM_R_X13Y136_SLICE_X19Y136_C1 = 1'b1;
  assign CLBLM_R_X13Y136_SLICE_X19Y136_C2 = 1'b1;
  assign CLBLM_R_X13Y136_SLICE_X19Y136_C3 = 1'b1;
  assign CLBLM_R_X13Y136_SLICE_X19Y136_C4 = 1'b1;
  assign CLBLM_R_X13Y136_SLICE_X19Y136_C5 = 1'b1;
  assign CLBLM_R_X13Y136_SLICE_X19Y136_C6 = 1'b1;
  assign CLBLM_R_X13Y136_SLICE_X19Y136_D1 = 1'b1;
  assign CLBLM_R_X13Y136_SLICE_X19Y136_D2 = 1'b1;
  assign CLBLM_R_X13Y136_SLICE_X19Y136_D3 = 1'b1;
  assign CLBLM_R_X13Y136_SLICE_X19Y136_D4 = 1'b1;
  assign CLBLM_R_X13Y136_SLICE_X19Y136_D5 = 1'b1;
  assign CLBLM_R_X13Y136_SLICE_X19Y136_D6 = 1'b1;
  assign CLBLM_R_X13Y136_SLICE_X18Y136_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y136_SLICE_X18Y136_A2 = CLBLM_L_X10Y135_SLICE_X12Y135_DO6;
  assign CLBLM_R_X13Y136_SLICE_X18Y136_A3 = CLBLM_R_X13Y136_SLICE_X18Y136_AQ;
  assign CLBLM_R_X13Y136_SLICE_X18Y136_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X13Y136_SLICE_X18Y136_A5 = CLBLM_L_X12Y135_SLICE_X16Y135_CQ;
  assign CLBLM_R_X13Y136_SLICE_X18Y136_A6 = CLBLM_R_X13Y140_SLICE_X19Y140_BQ;
  assign CLBLM_R_X13Y136_SLICE_X18Y136_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y136_SLICE_X18Y136_B2 = CLBLM_R_X13Y136_SLICE_X18Y136_BQ;
  assign CLBLM_R_X13Y136_SLICE_X18Y136_B3 = CLBLM_R_X13Y137_SLICE_X19Y137_CQ;
  assign CLBLM_R_X13Y136_SLICE_X18Y136_B4 = CLBLM_R_X13Y137_SLICE_X18Y137_BO5;
  assign CLBLM_R_X13Y136_SLICE_X18Y136_B5 = CLBLM_R_X13Y133_SLICE_X18Y133_BQ;
  assign CLBLM_R_X13Y136_SLICE_X18Y136_B6 = CLBLM_R_X13Y143_SLICE_X18Y143_AO6;
  assign CLBLM_R_X13Y142_SLICE_X19Y142_C4 = CLBLM_L_X12Y142_SLICE_X17Y142_BQ;
  assign LIOI3_X0Y67_ILOGIC_X0Y68_D = LIOB33_X0Y67_IOB_X0Y68_I;
  assign LIOI3_X0Y67_ILOGIC_X0Y67_D = LIOB33_X0Y67_IOB_X0Y67_I;
  assign CLBLM_R_X13Y142_SLICE_X19Y142_C5 = CLBLM_R_X13Y140_SLICE_X18Y140_AQ;
  assign CLBLM_R_X13Y136_SLICE_X18Y136_C1 = 1'b1;
  assign CLBLM_R_X13Y136_SLICE_X18Y136_C2 = CLBLM_R_X13Y137_SLICE_X18Y137_A5Q;
  assign CLBLM_R_X13Y136_SLICE_X18Y136_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y136_SLICE_X18Y136_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X13Y136_SLICE_X18Y136_C5 = 1'b1;
  assign CLBLM_R_X13Y136_SLICE_X18Y136_C6 = CLBLM_R_X11Y135_SLICE_X15Y135_BQ;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_D4 = 1'b1;
  assign CLBLM_R_X13Y142_SLICE_X19Y142_C6 = CLBLM_R_X13Y142_SLICE_X19Y142_AQ;
  assign RIOI3_X105Y111_ILOGIC_X1Y112_D = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X13Y136_SLICE_X18Y136_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_X105Y111_ILOGIC_X1Y111_D = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_D6 = 1'b1;
  assign CLBLM_R_X13Y136_SLICE_X18Y136_D1 = 1'b1;
  assign CLBLM_R_X13Y136_SLICE_X18Y136_D2 = 1'b1;
  assign CLBLM_R_X13Y136_SLICE_X18Y136_D3 = 1'b1;
  assign CLBLM_R_X13Y136_SLICE_X18Y136_D4 = 1'b1;
  assign CLBLM_R_X13Y136_SLICE_X18Y136_D5 = 1'b1;
  assign CLBLM_R_X13Y136_SLICE_X18Y136_D6 = 1'b1;
  assign CLBLM_R_X13Y142_SLICE_X19Y142_D2 = CLBLM_L_X12Y142_SLICE_X17Y142_BQ;
  assign CLBLM_R_X13Y142_SLICE_X19Y142_D5 = CLBLM_L_X12Y141_SLICE_X16Y141_AQ;
  assign RIOB33_X105Y183_IOB_X1Y184_O = CLBLM_L_X12Y139_SLICE_X17Y139_DO6;
  assign CLBLM_R_X13Y142_SLICE_X19Y142_D6 = CLBLM_R_X13Y142_SLICE_X19Y142_AQ;
  assign RIOB33_X105Y183_IOB_X1Y183_O = CLBLM_R_X11Y141_SLICE_X14Y141_CO5;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_A2 = CLBLM_R_X13Y144_SLICE_X18Y144_BO6;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_A3 = CLBLM_L_X12Y143_SLICE_X17Y143_AQ;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_A4 = CLBLM_L_X12Y142_SLICE_X17Y142_CO6;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_A5 = CLBLM_L_X8Y137_SLICE_X11Y137_AQ;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_A6 = CLBLM_R_X13Y141_SLICE_X18Y141_AO5;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_B1 = CLBLM_R_X7Y141_SLICE_X9Y141_BQ;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_B2 = CLBLM_L_X12Y143_SLICE_X17Y143_BQ;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_B3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_B5 = CLBLM_L_X12Y142_SLICE_X17Y142_CO6;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_B6 = CLBLM_L_X12Y143_SLICE_X17Y143_CO6;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_A1 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_A3 = CLBLM_L_X10Y133_SLICE_X13Y133_AQ;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_A4 = CLBLM_R_X5Y132_SLICE_X7Y132_DO6;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_A5 = CLBLM_L_X8Y137_SLICE_X11Y137_BQ;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_A6 = CLBLM_L_X10Y134_SLICE_X13Y134_A5Q;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_C1 = CLBLM_R_X13Y141_SLICE_X19Y141_CO5;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_C2 = CLBLM_R_X13Y140_SLICE_X19Y140_AQ;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_C3 = CLBLM_R_X13Y137_SLICE_X18Y137_CO5;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_B1 = CLBLM_L_X10Y133_SLICE_X13Y133_DO6;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_B3 = CLBLM_R_X7Y131_SLICE_X9Y131_AQ;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_B4 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_B5 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_B6 = CLBLM_L_X10Y134_SLICE_X13Y134_BQ;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_D1 = CLBLM_R_X13Y141_SLICE_X19Y141_CO5;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_C1 = CLBLM_L_X10Y131_SLICE_X13Y131_BQ;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_C2 = CLBLM_L_X10Y137_SLICE_X12Y137_CQ;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_C3 = CLBLM_L_X10Y131_SLICE_X13Y131_CQ;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_C4 = CLBLM_L_X8Y137_SLICE_X11Y137_BQ;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_C5 = CLBLM_L_X10Y133_SLICE_X13Y133_AQ;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_C6 = CLBLM_R_X11Y132_SLICE_X14Y132_AQ;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_D3 = CLBLM_L_X12Y142_SLICE_X16Y142_BQ;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_D4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_D6 = CLBLM_R_X13Y144_SLICE_X18Y144_BO6;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_A1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_A3 = CLBLM_R_X13Y139_SLICE_X18Y139_BO6;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_D1 = CLBLM_L_X10Y137_SLICE_X12Y137_CQ;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_D2 = CLBLM_R_X11Y132_SLICE_X15Y132_AO6;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_D3 = CLBLM_L_X10Y133_SLICE_X13Y133_BQ;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_D4 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_D5 = CLBLM_L_X10Y134_SLICE_X13Y134_B5Q;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_D6 = CLBLM_R_X5Y132_SLICE_X7Y132_DO6;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_B1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_B2 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_B3 = CLBLM_R_X13Y139_SLICE_X18Y139_BO6;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_B5 = CLBLM_L_X12Y141_SLICE_X16Y141_BQ;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_A1 = CLBLM_L_X8Y134_SLICE_X11Y134_BQ;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_A2 = CLBLL_L_X4Y134_SLICE_X4Y134_AQ;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_A3 = CLBLM_L_X10Y133_SLICE_X12Y133_AQ;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_C2 = CLBLM_L_X12Y143_SLICE_X16Y143_CQ;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_C3 = CLBLM_L_X12Y143_SLICE_X17Y143_CO5;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_C4 = CLBLM_R_X11Y142_SLICE_X14Y142_BQ;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_A5 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_A6 = CLBLM_R_X5Y133_SLICE_X7Y133_DO6;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_C1 = CLBLM_R_X13Y143_SLICE_X18Y143_AO6;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_B1 = CLBLM_L_X8Y131_SLICE_X11Y131_AQ;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_B2 = CLBLM_L_X10Y133_SLICE_X12Y133_BQ;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_B4 = CLBLM_L_X10Y134_SLICE_X12Y134_BQ;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_B5 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_B6 = CLBLM_R_X5Y133_SLICE_X7Y133_DO6;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_D1 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_C1 = CLBLM_L_X10Y133_SLICE_X12Y133_BQ;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_C2 = CLBLM_L_X10Y133_SLICE_X12Y133_CQ;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_C4 = CLBLM_R_X5Y132_SLICE_X7Y132_DO6;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_C5 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_C6 = CLBLM_R_X11Y133_SLICE_X15Y133_CQ;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_D3 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_D4 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_D6 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_D1 = CLBLM_R_X11Y131_SLICE_X15Y131_BQ;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_D2 = CLBLM_L_X8Y137_SLICE_X11Y137_BQ;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_D3 = CLBLL_L_X4Y135_SLICE_X5Y135_CQ;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_D4 = CLBLM_L_X10Y131_SLICE_X12Y131_BQ;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_D5 = CLBLM_L_X10Y130_SLICE_X12Y130_AQ;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_D6 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X162Y170_C3 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_D2 = 1'b1;
  assign LIOI3_X0Y65_ILOGIC_X0Y66_D = LIOB33_X0Y65_IOB_X0Y66_I;
  assign CLBLM_R_X13Y137_SLICE_X19Y137_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y137_SLICE_X19Y137_A2 = CLBLM_R_X15Y142_SLICE_X20Y142_AQ;
  assign CLBLM_R_X13Y137_SLICE_X19Y137_A3 = CLBLM_R_X13Y137_SLICE_X19Y137_AQ;
  assign CLBLM_R_X13Y137_SLICE_X19Y137_A4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X13Y137_SLICE_X19Y137_A5 = CLBLM_L_X10Y136_SLICE_X13Y136_BO6;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_D5 = CLBLM_L_X10Y145_SLICE_X12Y145_CO6;
  assign CLBLM_R_X13Y137_SLICE_X19Y137_A6 = CLBLM_L_X8Y138_SLICE_X10Y138_AQ;
  assign CLBLM_R_X13Y142_SLICE_X18Y142_C4 = CLBLM_L_X12Y140_SLICE_X17Y140_AQ;
  assign CLBLM_R_X13Y142_SLICE_X18Y142_C5 = CLBLM_L_X12Y142_SLICE_X17Y142_AQ;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_D6 = 1'b1;
  assign CLBLM_R_X13Y137_SLICE_X19Y137_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y137_SLICE_X19Y137_B2 = CLBLM_L_X12Y134_SLICE_X16Y134_AQ;
  assign CLBLM_R_X13Y137_SLICE_X19Y137_B3 = CLBLM_R_X13Y137_SLICE_X18Y137_CO5;
  assign CLBLM_R_X13Y137_SLICE_X19Y137_B4 = CLBLM_R_X13Y143_SLICE_X18Y143_AO6;
  assign CLBLM_R_X13Y137_SLICE_X19Y137_B5 = CLBLM_L_X12Y137_SLICE_X16Y137_BO5;
  assign CLBLM_R_X13Y137_SLICE_X19Y137_B6 = CLBLM_R_X13Y137_SLICE_X19Y137_BQ;
  assign CLBLM_R_X13Y142_SLICE_X18Y142_C6 = CLBLM_L_X12Y142_SLICE_X16Y142_AQ;
  assign CLBLM_R_X13Y137_SLICE_X19Y137_C1 = 1'b1;
  assign CLBLM_R_X13Y137_SLICE_X19Y137_C2 = CLBLM_R_X13Y137_SLICE_X18Y137_CO6;
  assign CLBLM_R_X13Y137_SLICE_X19Y137_C3 = CLBLM_R_X13Y143_SLICE_X18Y143_AO6;
  assign CLBLM_R_X13Y137_SLICE_X19Y137_C4 = CLBLM_R_X5Y136_SLICE_X7Y136_CQ;
  assign CLBLM_R_X13Y137_SLICE_X19Y137_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y137_SLICE_X19Y137_C6 = CLBLM_R_X13Y137_SLICE_X19Y137_CQ;
  assign CLBLM_R_X13Y137_SLICE_X19Y137_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y137_SLICE_X19Y137_D1 = 1'b1;
  assign CLBLM_R_X13Y137_SLICE_X19Y137_D2 = 1'b1;
  assign CLBLM_R_X13Y137_SLICE_X19Y137_D3 = 1'b1;
  assign CLBLM_R_X13Y137_SLICE_X19Y137_D4 = 1'b1;
  assign CLBLM_R_X13Y137_SLICE_X19Y137_D5 = 1'b1;
  assign CLBLM_R_X13Y137_SLICE_X19Y137_D6 = 1'b1;
  assign CLBLM_R_X13Y137_SLICE_X18Y137_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y137_SLICE_X18Y137_A2 = CLBLM_R_X11Y135_SLICE_X15Y135_BQ;
  assign CLBLM_R_X13Y137_SLICE_X18Y137_A3 = CLBLM_R_X13Y137_SLICE_X18Y137_AQ;
  assign CLBLM_R_X13Y137_SLICE_X18Y137_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X13Y137_SLICE_X18Y137_A5 = CLBLM_R_X11Y138_SLICE_X15Y138_B5Q;
  assign CLBLM_R_X13Y137_SLICE_X18Y137_A6 = CLBLM_L_X12Y137_SLICE_X17Y137_DO6;
  assign CLBLM_R_X13Y137_SLICE_X18Y137_AX = CLBLM_R_X13Y137_SLICE_X18Y137_BO6;
  assign CLBLM_R_X13Y137_SLICE_X18Y137_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y137_SLICE_X18Y137_B2 = CLBLM_L_X12Y137_SLICE_X17Y137_A5Q;
  assign CLBLM_R_X13Y137_SLICE_X18Y137_B3 = CLBLM_L_X12Y137_SLICE_X16Y137_A5Q;
  assign CLBLM_R_X13Y137_SLICE_X18Y137_B4 = CLBLM_R_X13Y137_SLICE_X19Y137_BQ;
  assign CLBLM_R_X13Y137_SLICE_X18Y137_B5 = CLBLM_R_X11Y139_SLICE_X15Y139_BQ;
  assign CLBLM_R_X13Y137_SLICE_X18Y137_B6 = 1'b1;
  assign CLBLM_R_X13Y137_SLICE_X18Y137_C1 = CLBLM_R_X13Y136_SLICE_X18Y136_BQ;
  assign CLBLM_R_X13Y137_SLICE_X18Y137_C2 = CLBLM_R_X13Y137_SLICE_X19Y137_BQ;
  assign CLBLM_R_X13Y137_SLICE_X18Y137_C3 = CLBLM_R_X11Y139_SLICE_X15Y139_BQ;
  assign CLBLM_R_X13Y137_SLICE_X18Y137_C4 = CLBLM_R_X13Y137_SLICE_X19Y137_CQ;
  assign CLBLM_R_X13Y137_SLICE_X18Y137_C5 = CLBLM_L_X12Y137_SLICE_X16Y137_A5Q;
  assign CLBLM_R_X13Y137_SLICE_X18Y137_C6 = 1'b1;
  assign CLBLM_R_X13Y137_SLICE_X18Y137_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_X105Y189_OLOGIC_X1Y190_D1 = CLBLM_R_X15Y142_SLICE_X20Y142_AQ;
  assign CLBLM_R_X13Y137_SLICE_X18Y137_D1 = 1'b1;
  assign CLBLM_R_X13Y137_SLICE_X18Y137_D2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X13Y137_SLICE_X18Y137_D3 = CLBLM_R_X13Y137_SLICE_X18Y137_AQ;
  assign CLBLM_R_X13Y137_SLICE_X18Y137_D4 = CLBLM_L_X12Y137_SLICE_X17Y137_DO6;
  assign CLBLM_R_X13Y137_SLICE_X18Y137_D5 = 1'b1;
  assign CLBLM_R_X13Y137_SLICE_X18Y137_D6 = CLBLM_R_X11Y135_SLICE_X15Y135_BQ;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_C4 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_C5 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_C6 = 1'b1;
  assign RIOB33_X105Y185_IOB_X1Y186_O = CLBLM_R_X13Y139_SLICE_X19Y139_AQ;
  assign RIOB33_X105Y185_IOB_X1Y185_O = CLBLM_L_X12Y139_SLICE_X17Y139_DO5;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_B6 = 1'b1;
  assign RIOI3_X105Y189_OLOGIC_X1Y190_T1 = 1'b1;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_A1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_A2 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_A3 = CLBLM_R_X13Y143_SLICE_X18Y143_AQ;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_A5 = CLBLM_L_X8Y140_SLICE_X11Y140_AQ;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_A6 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_C4 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_B1 = 1'b1;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_B2 = 1'b1;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_B3 = 1'b1;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_B4 = 1'b1;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_B5 = 1'b1;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_B6 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_D5 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_D6 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_C5 = CLBLM_R_X11Y144_SLICE_X15Y144_BQ;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_A1 = CLBLM_L_X10Y134_SLICE_X13Y134_DO6;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_A3 = CLBLM_L_X10Y134_SLICE_X13Y134_AQ;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_A4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_A5 = CLBLM_L_X8Y138_SLICE_X10Y138_AQ;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_A6 = CLBLM_R_X11Y134_SLICE_X15Y134_CQ;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_C1 = 1'b1;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_C2 = 1'b1;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_AX = CLBLM_L_X10Y140_SLICE_X13Y140_AO6;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_B1 = CLBLM_L_X10Y137_SLICE_X13Y137_DO6;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_B2 = CLBLM_L_X10Y134_SLICE_X13Y134_A5Q;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_B3 = CLBLM_L_X10Y133_SLICE_X13Y133_BQ;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_B4 = CLBLM_L_X10Y137_SLICE_X13Y137_AQ;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_B6 = 1'b1;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_D1 = 1'b1;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_D4 = 1'b1;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_C2 = CLBLM_L_X10Y135_SLICE_X12Y135_AQ;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_C3 = CLBLM_R_X5Y140_SLICE_X7Y140_BQ;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_C4 = CLBLM_R_X11Y134_SLICE_X15Y134_BQ;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_C5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_C6 = 1'b1;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_D3 = 1'b1;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_D5 = 1'b1;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_A1 = 1'b1;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_A2 = 1'b1;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_A3 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_A6 = CLBLM_R_X7Y131_SLICE_X9Y131_AQ;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_A5 = 1'b1;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_D1 = CLBLL_L_X4Y139_SLICE_X4Y139_BO6;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_AX = CLBLM_L_X10Y141_SLICE_X12Y141_C5Q;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_D2 = CLBLM_R_X13Y138_SLICE_X18Y138_BO6;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_D3 = 1'b1;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_D4 = CLBLL_L_X4Y142_SLICE_X5Y142_DO6;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_D5 = CLBLM_L_X8Y135_SLICE_X10Y135_CO6;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_D6 = CLBLM_R_X5Y136_SLICE_X7Y136_DO6;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_B1 = 1'b1;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_B2 = 1'b1;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_B3 = 1'b1;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_B4 = 1'b1;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_B5 = 1'b1;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_B6 = 1'b1;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_A1 = 1'b1;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_A2 = CLBLM_L_X10Y140_SLICE_X12Y140_AQ;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_A3 = CLBLM_L_X10Y134_SLICE_X12Y134_AQ;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_A5 = CLBLM_L_X10Y133_SLICE_X12Y133_AQ;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_A6 = CLBLM_R_X5Y133_SLICE_X7Y133_DO6;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_C1 = 1'b1;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_C2 = 1'b1;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_B1 = CLBLM_L_X8Y143_SLICE_X10Y143_DO6;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_B2 = CLBLM_L_X10Y134_SLICE_X12Y134_BQ;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_B3 = 1'b1;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_B5 = CLBLM_L_X10Y140_SLICE_X12Y140_A5Q;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_B6 = CLBLM_R_X11Y134_SLICE_X14Y134_CQ;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_D1 = 1'b1;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_C1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_C2 = CLBLM_L_X10Y134_SLICE_X12Y134_CQ;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_C3 = CLBLM_L_X10Y134_SLICE_X12Y134_DQ;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_C4 = CLBLM_L_X8Y138_SLICE_X10Y138_AQ;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_C5 = 1'b1;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_D2 = 1'b1;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_D3 = 1'b1;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_D6 = 1'b1;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_SR = CLBLM_L_X12Y144_SLICE_X16Y144_AO6;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_D1 = CLBLL_L_X52Y126_SLICE_X78Y126_AO6;
  assign LIOI3_X0Y191_OLOGIC_X0Y192_T1 = 1'b1;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_D1 = 1'b1;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_D2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_D3 = CLBLM_L_X10Y134_SLICE_X12Y134_DQ;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_D4 = CLBLM_L_X10Y134_SLICE_X13Y134_B5Q;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_D5 = 1'b1;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_D6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_T1 = 1'b1;
  assign LIOI3_X0Y191_OLOGIC_X0Y191_D1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign RIOI3_X105Y175_OLOGIC_X1Y176_D1 = CLBLM_R_X103Y173_SLICE_X163Y173_AO5;
  assign LIOI3_X0Y191_OLOGIC_X0Y191_T1 = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_D1 = CLBLM_R_X5Y136_SLICE_X6Y136_CQ;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_B4 = 1'b1;
  assign RIOI3_X105Y175_OLOGIC_X1Y176_T1 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_B5 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_B6 = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_T1 = 1'b1;
  assign RIOI3_X105Y175_OLOGIC_X1Y175_D1 = CLBLM_L_X12Y146_SLICE_X16Y146_AO6;
  assign CLBLM_R_X13Y138_SLICE_X19Y138_A1 = 1'b1;
  assign CLBLM_R_X13Y138_SLICE_X19Y138_A2 = 1'b1;
  assign CLBLM_R_X13Y138_SLICE_X19Y138_A3 = 1'b1;
  assign CLBLM_R_X13Y138_SLICE_X19Y138_A4 = 1'b1;
  assign CLBLM_R_X13Y138_SLICE_X19Y138_A5 = 1'b1;
  assign CLBLM_R_X13Y138_SLICE_X19Y138_A6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_D1 = LIOB33_X0Y57_IOB_X0Y57_I;
  assign RIOI3_X105Y175_OLOGIC_X1Y175_T1 = 1'b1;
  assign CLBLM_R_X13Y138_SLICE_X19Y138_B1 = 1'b1;
  assign CLBLM_R_X13Y138_SLICE_X19Y138_B2 = 1'b1;
  assign CLBLM_R_X13Y138_SLICE_X19Y138_B3 = 1'b1;
  assign CLBLM_R_X13Y138_SLICE_X19Y138_B4 = 1'b1;
  assign CLBLM_R_X13Y138_SLICE_X19Y138_B5 = 1'b1;
  assign CLBLM_R_X13Y138_SLICE_X19Y138_B6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_D1 = CLBLM_R_X11Y144_SLICE_X15Y144_AQ;
  assign CLBLM_R_X13Y138_SLICE_X19Y138_C1 = 1'b1;
  assign CLBLM_R_X13Y138_SLICE_X19Y138_C2 = 1'b1;
  assign CLBLM_R_X13Y138_SLICE_X19Y138_C3 = 1'b1;
  assign CLBLM_R_X13Y138_SLICE_X19Y138_C4 = 1'b1;
  assign CLBLM_R_X13Y138_SLICE_X19Y138_C5 = 1'b1;
  assign CLBLM_R_X13Y138_SLICE_X19Y138_C6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_D1 = LIOB33_X0Y55_IOB_X0Y55_I;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_T1 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_C4 = 1'b1;
  assign CLBLM_R_X13Y138_SLICE_X19Y138_D1 = 1'b1;
  assign CLBLM_R_X13Y138_SLICE_X19Y138_D2 = 1'b1;
  assign CLBLM_R_X13Y138_SLICE_X19Y138_D3 = 1'b1;
  assign CLBLM_R_X13Y138_SLICE_X19Y138_D4 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_C5 = 1'b1;
  assign CLBLM_R_X13Y138_SLICE_X19Y138_D6 = 1'b1;
  assign CLBLM_R_X13Y138_SLICE_X19Y138_D5 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_T1 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_C6 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_D1 = CLBLM_L_X12Y134_SLICE_X16Y134_AQ;
  assign CLBLM_R_X13Y138_SLICE_X18Y138_A1 = CLBLM_L_X12Y139_SLICE_X17Y139_BO5;
  assign CLBLM_R_X13Y138_SLICE_X18Y138_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y138_SLICE_X18Y138_A3 = CLBLM_R_X13Y138_SLICE_X18Y138_AQ;
  assign CLBLM_R_X13Y138_SLICE_X18Y138_A4 = CLBLM_L_X10Y135_SLICE_X12Y135_DO6;
  assign CLBLM_R_X13Y138_SLICE_X18Y138_A5 = CLBLM_R_X13Y140_SLICE_X18Y140_CQ;
  assign CLBLM_R_X13Y138_SLICE_X18Y138_A6 = CLBLM_L_X12Y138_SLICE_X17Y138_BO5;
  assign LIOB33_X0Y101_IOB_X0Y101_O = CLBLM_R_X3Y133_SLICE_X2Y133_AO6;
  assign LIOB33_X0Y101_IOB_X0Y102_O = CLBLM_R_X3Y133_SLICE_X2Y133_AO5;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_T1 = 1'b1;
  assign CLBLM_R_X13Y138_SLICE_X18Y138_B1 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X13Y138_SLICE_X18Y138_B2 = CLBLM_R_X13Y139_SLICE_X18Y139_BO6;
  assign CLBLM_R_X13Y138_SLICE_X18Y138_B3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X13Y138_SLICE_X18Y138_B4 = 1'b1;
  assign CLBLM_R_X13Y138_SLICE_X18Y138_B5 = 1'b1;
  assign CLBLM_R_X13Y138_SLICE_X18Y138_B6 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X13Y138_SLICE_X18Y138_C1 = 1'b1;
  assign CLBLM_R_X13Y138_SLICE_X18Y138_C2 = 1'b1;
  assign CLBLM_R_X13Y138_SLICE_X18Y138_C3 = 1'b1;
  assign CLBLM_R_X13Y138_SLICE_X18Y138_C4 = 1'b1;
  assign CLBLM_R_X13Y138_SLICE_X18Y138_C5 = 1'b1;
  assign CLBLM_R_X13Y138_SLICE_X18Y138_C6 = 1'b1;
  assign CLBLM_R_X13Y138_SLICE_X18Y138_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y138_SLICE_X18Y138_D1 = 1'b1;
  assign CLBLM_R_X13Y138_SLICE_X18Y138_D2 = 1'b1;
  assign CLBLM_R_X13Y138_SLICE_X18Y138_D3 = 1'b1;
  assign CLBLM_R_X13Y138_SLICE_X18Y138_D4 = 1'b1;
  assign CLBLM_R_X13Y138_SLICE_X18Y138_D5 = 1'b1;
  assign CLBLM_R_X13Y138_SLICE_X18Y138_D6 = 1'b1;
  assign RIOB33_X105Y187_IOB_X1Y187_O = CLBLM_L_X12Y134_SLICE_X16Y134_AQ;
  assign RIOB33_X105Y187_IOB_X1Y188_O = CLBLM_R_X11Y144_SLICE_X15Y144_AQ;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_D1 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_D6 = 1'b1;
  assign LIOI3_X0Y71_ILOGIC_X0Y72_D = LIOB33_X0Y71_IOB_X0Y72_I;
  assign LIOI3_X0Y71_ILOGIC_X0Y71_D = LIOB33_X0Y71_IOB_X0Y71_I;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_T1 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_A1 = CLBLM_L_X10Y135_SLICE_X13Y135_B5Q;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_A3 = CLBLM_R_X11Y135_SLICE_X14Y135_DQ;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_A4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_A5 = CLBLM_L_X10Y133_SLICE_X13Y133_AQ;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_A6 = 1'b1;
  assign RIOI3_X105Y115_ILOGIC_X1Y116_D = RIOB33_X105Y115_IOB_X1Y116_I;
  assign RIOI3_X105Y115_ILOGIC_X1Y115_D = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_B2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_B3 = CLBLM_R_X11Y134_SLICE_X14Y134_DQ;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_B4 = CLBLM_R_X11Y138_SLICE_X14Y138_BQ;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_B5 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_B6 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_C1 = CLBLM_R_X11Y135_SLICE_X15Y135_CO5;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_C2 = CLBLL_L_X4Y142_SLICE_X5Y142_DO6;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_C3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_C4 = CLBLM_L_X10Y138_SLICE_X13Y138_CQ;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_C5 = CLBLM_L_X10Y135_SLICE_X13Y135_B5Q;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_C6 = CLBLM_L_X8Y137_SLICE_X11Y137_CO5;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_D1 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_D2 = CLBLM_L_X8Y133_SLICE_X11Y133_BQ;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_D3 = CLBLM_L_X12Y135_SLICE_X16Y135_DQ;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_D4 = CLBLM_R_X11Y134_SLICE_X14Y134_DQ;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_D5 = CLBLM_L_X10Y135_SLICE_X13Y135_B5Q;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_D6 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_A1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_A3 = CLBLM_L_X10Y135_SLICE_X12Y135_AQ;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_A4 = CLBLM_L_X8Y138_SLICE_X10Y138_AQ;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_A5 = CLBLM_R_X7Y132_SLICE_X8Y132_AQ;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_A6 = CLBLM_L_X10Y135_SLICE_X12Y135_CO6;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_D1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_B1 = CLBLM_L_X12Y135_SLICE_X16Y135_DQ;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_B2 = CLBLM_R_X11Y139_SLICE_X15Y139_A5Q;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_B3 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_B4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_B6 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_C1 = CLBLL_L_X4Y134_SLICE_X4Y134_AQ;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_C2 = CLBLM_L_X10Y137_SLICE_X12Y137_AQ;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_C3 = CLBLM_L_X8Y135_SLICE_X11Y135_DO6;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_C4 = CLBLM_R_X5Y140_SLICE_X7Y140_BQ;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_C5 = CLBLM_L_X8Y135_SLICE_X10Y135_CO6;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_C6 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_D1 = CLBLM_R_X5Y134_SLICE_X6Y134_AQ;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_D2 = CLBLM_R_X11Y135_SLICE_X14Y135_AQ;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_D3 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_D4 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_D5 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_D6 = CLBLM_L_X8Y138_SLICE_X10Y138_AQ;
  assign LIOB33_X0Y141_IOB_X0Y142_O = LIOB33_X0Y53_IOB_X0Y54_I;
  assign LIOB33_X0Y141_IOB_X0Y141_O = CLBLM_R_X3Y136_SLICE_X3Y136_BQ;
  assign CLBLM_R_X13Y139_SLICE_X19Y139_A1 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X13Y139_SLICE_X19Y139_A2 = CLBLM_L_X8Y139_SLICE_X11Y139_AQ;
  assign CLBLM_R_X13Y139_SLICE_X19Y139_A3 = CLBLM_R_X13Y139_SLICE_X19Y139_AQ;
  assign CLBLM_R_X13Y139_SLICE_X19Y139_A4 = 1'b1;
  assign CLBLM_R_X13Y139_SLICE_X19Y139_A5 = CLBLM_R_X7Y131_SLICE_X9Y131_AQ;
  assign CLBLM_R_X13Y139_SLICE_X19Y139_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y139_SLICE_X19Y139_B1 = 1'b1;
  assign CLBLM_R_X13Y139_SLICE_X19Y139_B2 = 1'b1;
  assign CLBLM_R_X13Y139_SLICE_X19Y139_B3 = 1'b1;
  assign CLBLM_R_X13Y139_SLICE_X19Y139_B4 = 1'b1;
  assign CLBLM_R_X13Y139_SLICE_X19Y139_B5 = 1'b1;
  assign CLBLM_R_X13Y139_SLICE_X19Y139_B6 = 1'b1;
  assign LIOB33_X0Y103_IOB_X0Y104_O = CLBLL_L_X2Y133_SLICE_X0Y133_CO6;
  assign LIOB33_X0Y103_IOB_X0Y103_O = CLBLL_L_X2Y133_SLICE_X0Y133_AO5;
  assign CLBLM_R_X13Y139_SLICE_X19Y139_C1 = 1'b1;
  assign CLBLM_R_X13Y139_SLICE_X19Y139_C2 = 1'b1;
  assign CLBLM_R_X13Y139_SLICE_X19Y139_C3 = 1'b1;
  assign CLBLM_R_X13Y139_SLICE_X19Y139_C4 = 1'b1;
  assign CLBLM_R_X13Y139_SLICE_X19Y139_C5 = 1'b1;
  assign CLBLM_R_X13Y139_SLICE_X19Y139_C6 = 1'b1;
  assign CLBLM_R_X13Y139_SLICE_X19Y139_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y139_SLICE_X19Y139_D1 = 1'b1;
  assign CLBLM_R_X13Y139_SLICE_X19Y139_D2 = 1'b1;
  assign CLBLM_R_X13Y139_SLICE_X19Y139_D3 = 1'b1;
  assign CLBLM_R_X13Y139_SLICE_X19Y139_D4 = 1'b1;
  assign CLBLM_R_X13Y139_SLICE_X19Y139_D5 = 1'b1;
  assign CLBLM_R_X13Y139_SLICE_X19Y139_D6 = 1'b1;
  assign CLBLM_R_X13Y139_SLICE_X18Y139_A1 = CLBLM_R_X13Y143_SLICE_X18Y143_AO6;
  assign CLBLM_R_X13Y139_SLICE_X18Y139_A2 = CLBLM_R_X13Y137_SLICE_X18Y137_CO5;
  assign CLBLM_R_X13Y139_SLICE_X18Y139_A3 = CLBLM_R_X13Y139_SLICE_X18Y139_AQ;
  assign CLBLM_R_X13Y139_SLICE_X18Y139_A4 = CLBLM_R_X13Y141_SLICE_X18Y141_BO6;
  assign CLBLM_R_X13Y139_SLICE_X18Y139_A5 = CLBLM_R_X7Y132_SLICE_X9Y132_AQ;
  assign CLBLM_R_X13Y139_SLICE_X18Y139_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign RIOB33_X105Y189_IOB_X1Y190_O = CLBLM_R_X15Y142_SLICE_X20Y142_AQ;
  assign RIOB33_X105Y189_IOB_X1Y189_O = CLBLM_L_X10Y143_SLICE_X13Y143_BQ;
  assign CLBLM_R_X13Y139_SLICE_X18Y139_B1 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLM_R_X13Y139_SLICE_X18Y139_B2 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X13Y139_SLICE_X18Y139_B3 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLM_R_X13Y139_SLICE_X18Y139_B4 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X13Y139_SLICE_X18Y139_B5 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X13Y139_SLICE_X18Y139_B6 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X13Y139_SLICE_X18Y139_C1 = 1'b1;
  assign CLBLM_R_X13Y139_SLICE_X18Y139_C2 = 1'b1;
  assign CLBLM_R_X13Y139_SLICE_X18Y139_C3 = 1'b1;
  assign CLBLM_R_X13Y139_SLICE_X18Y139_C4 = 1'b1;
  assign CLBLM_R_X13Y139_SLICE_X18Y139_C5 = 1'b1;
  assign CLBLM_R_X13Y139_SLICE_X18Y139_C6 = 1'b1;
  assign CLBLM_R_X13Y139_SLICE_X18Y139_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y139_SLICE_X18Y139_D1 = 1'b1;
  assign CLBLM_R_X13Y139_SLICE_X18Y139_D2 = 1'b1;
  assign CLBLM_R_X13Y139_SLICE_X18Y139_D3 = 1'b1;
  assign CLBLM_R_X13Y139_SLICE_X18Y139_D4 = 1'b1;
  assign CLBLM_R_X13Y139_SLICE_X18Y139_D5 = 1'b1;
  assign CLBLM_R_X13Y139_SLICE_X18Y139_D6 = 1'b1;
  assign CLBLM_R_X13Y143_SLICE_X19Y143_C4 = 1'b1;
  assign CLBLM_R_X13Y143_SLICE_X19Y143_C5 = 1'b1;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_A1 = 1'b1;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_A2 = 1'b1;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_A3 = 1'b1;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_A4 = 1'b1;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_A5 = 1'b1;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_A6 = 1'b1;
  assign CLBLM_R_X13Y143_SLICE_X19Y143_C6 = 1'b1;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_B1 = 1'b1;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_B2 = 1'b1;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_B3 = 1'b1;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_B4 = 1'b1;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_B5 = 1'b1;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_B6 = 1'b1;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_C1 = 1'b1;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_C2 = 1'b1;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_C3 = 1'b1;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_C4 = 1'b1;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_C5 = 1'b1;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_C6 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_A1 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_A2 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_A3 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_A4 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_A5 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_A6 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_B1 = 1'b1;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_D1 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_B3 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_B4 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_B5 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_B6 = 1'b1;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_D2 = 1'b1;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_D3 = 1'b1;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_D4 = 1'b1;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_D5 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_C1 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_C2 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_C3 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_C4 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_C5 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_C6 = 1'b1;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_A1 = CLBLM_R_X7Y139_SLICE_X8Y139_A5Q;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_A2 = CLBLM_R_X11Y137_SLICE_X15Y137_BO6;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_A3 = CLBLM_L_X10Y135_SLICE_X13Y135_DO6;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_A4 = CLBLM_R_X11Y136_SLICE_X15Y136_BQ;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_A5 = CLBLM_L_X10Y141_SLICE_X13Y141_BQ;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_A6 = CLBLM_R_X7Y139_SLICE_X9Y139_A5Q;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_B1 = CLBLL_L_X4Y141_SLICE_X4Y141_DO6;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_B2 = CLBLM_L_X12Y135_SLICE_X17Y135_BO5;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_D2 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_D3 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_D4 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_D5 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_D6 = 1'b1;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_B3 = CLBLL_L_X4Y134_SLICE_X4Y134_AQ;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_B4 = CLBLM_L_X8Y136_SLICE_X11Y136_DO5;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_B6 = CLBLM_L_X10Y134_SLICE_X12Y134_CQ;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_C1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_C2 = CLBLM_L_X10Y136_SLICE_X12Y136_CO5;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_C3 = CLBLL_L_X4Y141_SLICE_X4Y141_DO6;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_C4 = CLBLM_R_X13Y137_SLICE_X18Y137_AQ;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_C5 = CLBLM_R_X13Y138_SLICE_X18Y138_BO6;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_A2 = 1'b1;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_A3 = CLBLM_L_X10Y131_SLICE_X13Y131_AQ;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_A4 = CLBLM_R_X5Y136_SLICE_X6Y136_DQ;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_A5 = CLBLM_R_X5Y133_SLICE_X7Y133_DO6;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_A6 = CLBLL_L_X4Y132_SLICE_X5Y132_AQ;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_D1 = CLBLM_R_X13Y135_SLICE_X18Y135_BQ;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_B1 = 1'b1;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_B2 = 1'b1;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_B3 = 1'b1;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_B4 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_B6 = 1'b1;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_B5 = 1'b1;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_B6 = 1'b1;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_C1 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_C1 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_C2 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_C3 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_C4 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_C5 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_C6 = 1'b1;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_C2 = 1'b1;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_A1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_A2 = CLBLM_L_X10Y134_SLICE_X13Y134_AQ;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_C5 = 1'b1;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_C6 = 1'b1;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_A6 = 1'b1;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_AX = CLBLM_R_X11Y136_SLICE_X14Y136_CO6;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_D1 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_D2 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_D3 = 1'b1;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_D1 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_D5 = 1'b1;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_D2 = 1'b1;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_D3 = 1'b1;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_D4 = 1'b1;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_D5 = 1'b1;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_D6 = 1'b1;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_C1 = CLBLM_L_X10Y134_SLICE_X13Y134_AQ;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_C2 = CLBLL_L_X4Y136_SLICE_X4Y136_CQ;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_C3 = CLBLM_R_X5Y138_SLICE_X6Y138_BQ;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_C6 = 1'b1;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_C4 = CLBLM_R_X11Y136_SLICE_X14Y136_BQ;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_C5 = CLBLM_L_X10Y136_SLICE_X12Y136_AQ;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_D1 = CLBLL_L_X4Y134_SLICE_X4Y134_AQ;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_D2 = CLBLM_L_X8Y138_SLICE_X11Y138_CO6;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_D3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_D4 = CLBLM_L_X10Y134_SLICE_X12Y134_CQ;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_D5 = 1'b1;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_D6 = CLBLL_L_X4Y142_SLICE_X4Y142_BO6;
  assign LIOB33_X0Y105_IOB_X0Y106_O = CLBLL_L_X4Y138_SLICE_X5Y138_DO6;
  assign LIOB33_X0Y105_IOB_X0Y105_O = CLBLL_L_X2Y133_SLICE_X0Y133_BO5;
  assign CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_CE = 1'b1;
  assign CLBLM_R_X13Y140_SLICE_X19Y140_A1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X13Y140_SLICE_X19Y140_A2 = CLBLM_R_X13Y143_SLICE_X18Y143_AO5;
  assign CLBLM_R_X13Y140_SLICE_X19Y140_A3 = CLBLM_R_X13Y140_SLICE_X19Y140_AQ;
  assign CLBLM_R_X13Y140_SLICE_X19Y140_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y140_SLICE_X19Y140_A5 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_R_X13Y140_SLICE_X19Y140_A6 = CLBLM_R_X13Y140_SLICE_X19Y140_CO6;
  assign CLBLM_R_X13Y140_SLICE_X19Y140_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y140_SLICE_X19Y140_B2 = CLBLM_L_X12Y143_SLICE_X17Y143_DO6;
  assign CLBLM_R_X13Y140_SLICE_X19Y140_B3 = 1'b1;
  assign CLBLM_R_X13Y140_SLICE_X19Y140_B4 = CLBLM_R_X13Y141_SLICE_X18Y141_AO5;
  assign CLBLM_R_X13Y140_SLICE_X19Y140_B5 = CLBLM_R_X7Y133_SLICE_X9Y133_BQ;
  assign CLBLM_R_X13Y140_SLICE_X19Y140_B6 = CLBLM_R_X13Y140_SLICE_X18Y140_DO6;
  assign CLBLM_R_X13Y140_SLICE_X19Y140_C1 = 1'b1;
  assign CLBLM_R_X13Y140_SLICE_X19Y140_C2 = CLBLM_L_X12Y143_SLICE_X17Y143_CO5;
  assign CLBLM_R_X13Y140_SLICE_X19Y140_C3 = CLBLM_L_X12Y142_SLICE_X16Y142_CQ;
  assign CLBLM_R_X13Y140_SLICE_X19Y140_C4 = 1'b1;
  assign CLBLM_R_X13Y140_SLICE_X19Y140_C5 = 1'b1;
  assign CLBLM_R_X13Y140_SLICE_X19Y140_C6 = 1'b1;
  assign RIOB33_X105Y191_IOB_X1Y191_O = CLBLM_L_X10Y143_SLICE_X13Y143_AQ;
  assign RIOB33_X105Y191_IOB_X1Y192_O = CLBLM_R_X13Y134_SLICE_X19Y134_BQ;
  assign CLBLM_R_X13Y140_SLICE_X19Y140_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y140_SLICE_X19Y140_D1 = 1'b1;
  assign CLBLM_R_X13Y140_SLICE_X19Y140_D2 = 1'b1;
  assign CLBLM_R_X13Y140_SLICE_X19Y140_D3 = 1'b1;
  assign CLBLM_R_X13Y140_SLICE_X19Y140_D4 = 1'b1;
  assign CLBLM_R_X13Y140_SLICE_X19Y140_D5 = 1'b1;
  assign CLBLM_R_X13Y140_SLICE_X19Y140_D6 = 1'b1;
  assign CLBLM_R_X13Y140_SLICE_X18Y140_A1 = CLBLM_R_X13Y140_SLICE_X18Y140_AQ;
  assign CLBLM_R_X13Y140_SLICE_X18Y140_A2 = CLBLM_R_X13Y141_SLICE_X18Y141_AO5;
  assign CLBLM_R_X13Y140_SLICE_X18Y140_A3 = CLBLM_R_X13Y142_SLICE_X18Y142_AO6;
  assign CLBLM_R_X13Y140_SLICE_X18Y140_A4 = CLBLM_L_X12Y143_SLICE_X17Y143_DO6;
  assign CLBLM_R_X13Y140_SLICE_X18Y140_A5 = CLBLM_L_X8Y141_SLICE_X11Y141_AQ;
  assign CLBLM_R_X13Y140_SLICE_X18Y140_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOI3_X0Y195_OLOGIC_X0Y196_D1 = LIOB33_X0Y69_IOB_X0Y69_I;
  assign CLBLM_R_X13Y140_SLICE_X18Y140_B1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X13Y140_SLICE_X18Y140_B2 = CLBLM_R_X13Y140_SLICE_X18Y140_BQ;
  assign CLBLM_R_X13Y140_SLICE_X18Y140_B3 = CLBLM_R_X13Y138_SLICE_X18Y138_AQ;
  assign CLBLM_R_X13Y140_SLICE_X18Y140_B4 = CLBLM_R_X13Y141_SLICE_X18Y141_DO6;
  assign CLBLM_R_X13Y140_SLICE_X18Y140_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y140_SLICE_X18Y140_B6 = CLBLM_R_X13Y143_SLICE_X18Y143_AO6;
  assign LIOI3_X0Y195_OLOGIC_X0Y196_T1 = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_D1 = CLBLM_R_X3Y133_SLICE_X3Y133_AQ;
  assign CLBLM_R_X13Y140_SLICE_X18Y140_C1 = CLBLM_R_X13Y141_SLICE_X19Y141_AQ;
  assign CLBLM_R_X13Y140_SLICE_X18Y140_C2 = CLBLM_R_X13Y143_SLICE_X18Y143_AO6;
  assign CLBLM_R_X13Y140_SLICE_X18Y140_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y140_SLICE_X18Y140_C4 = CLBLM_L_X12Y141_SLICE_X17Y141_CO6;
  assign CLBLM_R_X13Y140_SLICE_X18Y140_C5 = 1'b1;
  assign CLBLM_R_X13Y140_SLICE_X18Y140_C6 = CLBLM_R_X5Y137_SLICE_X7Y137_DO6;
  assign LIOI3_X0Y195_OLOGIC_X0Y195_D1 = LIOB33_X0Y63_IOB_X0Y64_I;
  assign CLBLM_R_X13Y140_SLICE_X18Y140_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_T1 = 1'b1;
  assign RIOI3_X105Y177_OLOGIC_X1Y178_D1 = CLBLM_R_X103Y177_SLICE_X163Y177_AO5;
  assign CLBLM_R_X13Y140_SLICE_X18Y140_D1 = 1'b1;
  assign CLBLM_R_X13Y140_SLICE_X18Y140_D2 = CLBLM_R_X13Y144_SLICE_X18Y144_CO6;
  assign CLBLM_R_X13Y140_SLICE_X18Y140_D3 = CLBLM_R_X11Y142_SLICE_X14Y142_BQ;
  assign CLBLM_R_X13Y140_SLICE_X18Y140_D4 = CLBLM_R_X13Y143_SLICE_X18Y143_BO6;
  assign CLBLM_R_X13Y140_SLICE_X18Y140_D5 = CLBLM_R_X13Y141_SLICE_X18Y141_BO5;
  assign CLBLM_R_X13Y140_SLICE_X18Y140_D6 = CLBLM_R_X13Y140_SLICE_X19Y140_BQ;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_D1 = CLBLM_R_X3Y137_SLICE_X3Y137_AQ;
  assign LIOI3_X0Y195_OLOGIC_X0Y195_T1 = 1'b1;
  assign RIOI3_X105Y177_OLOGIC_X1Y178_T1 = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_T1 = 1'b1;
  assign RIOI3_X105Y177_OLOGIC_X1Y177_D1 = CLBLM_R_X103Y177_SLICE_X163Y177_AO6;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_D1 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign RIOI3_X105Y177_OLOGIC_X1Y177_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_T1 = 1'b1;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_A3 = CLBLL_L_X4Y133_SLICE_X4Y133_AQ;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_A4 = CLBLM_R_X3Y135_SLICE_X3Y135_BQ;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_A5 = CLBLM_R_X5Y132_SLICE_X7Y132_CO5;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_A6 = CLBLM_R_X11Y138_SLICE_X15Y138_BQ;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_D1 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_B1 = CLBLL_L_X4Y134_SLICE_X5Y134_A5Q;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_B2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_B3 = CLBLL_L_X4Y135_SLICE_X5Y135_C5Q;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_B4 = CLBLM_R_X11Y138_SLICE_X15Y138_BQ;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_B5 = CLBLL_L_X4Y134_SLICE_X4Y134_B5Q;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_B6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_T1 = 1'b1;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_C2 = CLBLL_L_X4Y139_SLICE_X4Y139_BO6;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_C3 = CLBLL_L_X4Y142_SLICE_X4Y142_BO6;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_C4 = CLBLL_L_X4Y136_SLICE_X4Y136_AO5;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_C5 = CLBLM_L_X12Y134_SLICE_X17Y134_AQ;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_C6 = CLBLM_R_X5Y133_SLICE_X6Y133_CO6;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_D1 = 1'b1;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_D2 = 1'b1;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_D3 = 1'b1;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_D4 = 1'b1;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_D5 = 1'b1;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_D6 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_A2 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_A3 = CLBLM_L_X8Y139_SLICE_X10Y139_BQ;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_A5 = CLBLM_L_X12Y137_SLICE_X16Y137_AQ;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_A6 = CLBLM_L_X10Y138_SLICE_X12Y138_CO6;
  assign LIOI3_X0Y103_OLOGIC_X0Y104_D1 = CLBLL_L_X2Y133_SLICE_X0Y133_CO6;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_B2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_B3 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_B4 = CLBLM_R_X11Y137_SLICE_X14Y137_CO6;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_B5 = CLBLM_R_X11Y137_SLICE_X14Y137_AQ;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_B6 = CLBLM_L_X8Y135_SLICE_X11Y135_A5Q;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_C1 = CLBLM_L_X10Y141_SLICE_X13Y141_BQ;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_C2 = CLBLM_L_X10Y139_SLICE_X13Y139_AQ;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_A1 = CLBLL_L_X4Y133_SLICE_X5Y133_DO6;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_A2 = CLBLM_R_X11Y133_SLICE_X15Y133_BQ;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_A3 = CLBLL_L_X4Y133_SLICE_X5Y133_AQ;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_A5 = CLBLL_L_X4Y133_SLICE_X4Y133_BO6;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_A6 = CLBLL_L_X4Y134_SLICE_X5Y134_CQ;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_C3 = CLBLM_R_X11Y139_SLICE_X15Y139_CQ;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_AX = CLBLL_L_X4Y136_SLICE_X5Y136_DO6;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_C4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_B1 = CLBLM_R_X5Y132_SLICE_X7Y132_DO6;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_B2 = CLBLL_L_X4Y133_SLICE_X4Y133_BO5;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_B4 = CLBLM_L_X10Y132_SLICE_X12Y132_AO6;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_B5 = CLBLL_L_X4Y135_SLICE_X5Y135_C5Q;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_B6 = CLBLM_R_X5Y132_SLICE_X7Y132_BO5;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_D4 = CLBLL_L_X4Y138_SLICE_X5Y138_BQ;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_D5 = 1'b1;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_C1 = CLBLM_L_X10Y132_SLICE_X12Y132_AO6;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_C2 = CLBLL_L_X4Y134_SLICE_X5Y134_CQ;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_C3 = CLBLL_L_X4Y134_SLICE_X5Y134_AQ;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_C4 = CLBLM_R_X5Y132_SLICE_X7Y132_BO5;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_C5 = CLBLL_L_X4Y133_SLICE_X5Y133_AQ;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_C6 = CLBLM_R_X5Y132_SLICE_X7Y132_DO6;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_D6 = CLBLM_L_X10Y134_SLICE_X13Y134_BQ;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_A3 = CLBLM_L_X10Y137_SLICE_X12Y137_AQ;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_A4 = CLBLM_R_X11Y142_SLICE_X15Y142_BQ;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_A5 = CLBLM_L_X8Y138_SLICE_X10Y138_AQ;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_A2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_D1 = CLBLM_L_X10Y132_SLICE_X12Y132_AO6;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_D2 = CLBLL_L_X4Y134_SLICE_X5Y134_AQ;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_B1 = CLBLM_L_X10Y136_SLICE_X12Y136_A5Q;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_B2 = CLBLL_L_X4Y137_SLICE_X5Y137_BQ;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_B3 = CLBLM_L_X10Y143_SLICE_X12Y143_AQ;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_B5 = CLBLM_L_X12Y136_SLICE_X17Y136_A5Q;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_B6 = 1'b1;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_D3 = 1'b1;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_D4 = CLBLM_R_X5Y132_SLICE_X7Y132_BO5;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_D5 = 1'b1;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_D6 = CLBLM_R_X5Y132_SLICE_X7Y132_DO6;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_C2 = CLBLM_L_X10Y137_SLICE_X12Y137_CQ;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_C3 = CLBLM_L_X8Y140_SLICE_X11Y140_BQ;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_C5 = CLBLM_R_X11Y133_SLICE_X15Y133_AQ;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_C6 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_C1 = CLBLM_R_X5Y132_SLICE_X7Y132_DO6;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOB33_X0Y107_IOB_X0Y108_O = CLBLL_L_X2Y133_SLICE_X0Y133_CO5;
  assign LIOB33_X0Y107_IOB_X0Y107_O = CLBLL_L_X2Y108_SLICE_X0Y108_AO6;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_D1 = CLBLM_R_X7Y132_SLICE_X8Y132_BQ;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_D2 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_D3 = CLBLM_R_X11Y138_SLICE_X15Y138_B5Q;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_D4 = CLBLM_R_X11Y133_SLICE_X14Y133_CQ;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_D5 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_D6 = CLBLM_L_X8Y135_SLICE_X10Y135_BQ;
  assign LIOI3_X0Y73_ILOGIC_X0Y74_D = LIOB33_X0Y73_IOB_X0Y74_I;
  assign LIOI3_X0Y73_ILOGIC_X0Y73_D = LIOB33_X0Y73_IOB_X0Y73_I;
  assign RIOI3_X105Y117_ILOGIC_X1Y118_D = RIOB33_X105Y117_IOB_X1Y118_I;
  assign RIOI3_X105Y117_ILOGIC_X1Y117_D = RIOB33_X105Y117_IOB_X1Y117_I;
  assign RIOB33_X105Y193_IOB_X1Y194_O = CLBLM_R_X13Y144_SLICE_X19Y144_AQ;
  assign RIOB33_X105Y193_IOB_X1Y193_O = CLBLM_L_X12Y144_SLICE_X16Y144_AQ;
  assign CLBLM_R_X13Y141_SLICE_X19Y141_A1 = CLBLM_R_X13Y141_SLICE_X19Y141_DO6;
  assign CLBLM_R_X13Y141_SLICE_X19Y141_A2 = CLBLM_R_X13Y144_SLICE_X18Y144_AQ;
  assign CLBLM_R_X13Y141_SLICE_X19Y141_A3 = CLBLM_R_X13Y141_SLICE_X18Y141_AO5;
  assign CLBLM_R_X13Y141_SLICE_X19Y141_A4 = 1'b1;
  assign CLBLM_R_X13Y141_SLICE_X19Y141_A5 = CLBLM_L_X12Y143_SLICE_X17Y143_DO6;
  assign CLBLM_R_X13Y141_SLICE_X19Y141_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y141_SLICE_X19Y141_B1 = 1'b1;
  assign CLBLM_R_X13Y141_SLICE_X19Y141_B2 = CLBLM_R_X13Y141_SLICE_X19Y141_BQ;
  assign CLBLM_R_X13Y141_SLICE_X19Y141_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X13Y141_SLICE_X19Y141_B4 = CLBLM_L_X12Y142_SLICE_X17Y142_BQ;
  assign CLBLM_R_X13Y141_SLICE_X19Y141_B5 = 1'b1;
  assign CLBLM_R_X13Y141_SLICE_X19Y141_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOB33_X0Y119_IOB_X0Y120_O = CLBLM_L_X12Y136_SLICE_X16Y136_BQ;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_A1 = CLBLM_L_X10Y131_SLICE_X12Y131_BQ;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_A2 = CLBLM_R_X11Y131_SLICE_X15Y131_BQ;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_A3 = CLBLM_L_X10Y130_SLICE_X12Y130_AQ;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_A4 = CLBLM_L_X10Y131_SLICE_X13Y131_CQ;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_A5 = CLBLL_L_X4Y135_SLICE_X5Y135_CQ;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_A6 = 1'b1;
  assign CLBLM_R_X13Y141_SLICE_X19Y141_C1 = 1'b1;
  assign CLBLM_R_X13Y141_SLICE_X19Y141_C2 = CLBLM_R_X13Y141_SLICE_X19Y141_AQ;
  assign CLBLM_R_X13Y141_SLICE_X19Y141_C3 = CLBLM_R_X13Y141_SLICE_X18Y141_BO5;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_B1 = CLBLM_R_X11Y131_SLICE_X15Y131_DO6;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_B2 = CLBLM_R_X11Y131_SLICE_X15Y131_BQ;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_B3 = CLBLM_R_X13Y140_SLICE_X18Y140_AQ;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_B5 = CLBLM_R_X11Y140_SLICE_X15Y140_CQ;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X13Y141_SLICE_X19Y141_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y141_SLICE_X19Y141_D1 = CLBLM_L_X12Y142_SLICE_X16Y142_CQ;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_C1 = CLBLL_L_X4Y135_SLICE_X5Y135_CQ;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_C2 = CLBLM_R_X11Y133_SLICE_X15Y133_AQ;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_C3 = CLBLM_R_X11Y131_SLICE_X15Y131_BQ;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_C4 = CLBLM_L_X10Y131_SLICE_X12Y131_BQ;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_C5 = CLBLM_L_X10Y130_SLICE_X12Y130_AQ;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_C6 = 1'b1;
  assign CLBLM_R_X13Y141_SLICE_X19Y141_D3 = CLBLM_R_X13Y141_SLICE_X18Y141_BO5;
  assign CLBLM_R_X13Y141_SLICE_X19Y141_D4 = CLBLM_R_X13Y142_SLICE_X19Y142_CO6;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y141_SLICE_X18Y141_A1 = CLBLM_L_X12Y143_SLICE_X17Y143_BQ;
  assign CLBLM_R_X13Y141_SLICE_X18Y141_A2 = CLBLM_L_X12Y142_SLICE_X16Y142_BQ;
  assign CLBLM_R_X13Y141_SLICE_X18Y141_A3 = CLBLM_R_X13Y141_SLICE_X19Y141_CO5;
  assign CLBLM_R_X13Y141_SLICE_X18Y141_A4 = CLBLM_R_X13Y144_SLICE_X18Y144_AQ;
  assign CLBLM_R_X13Y141_SLICE_X18Y141_A5 = CLBLM_R_X13Y140_SLICE_X18Y140_BQ;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_D1 = CLBLL_L_X4Y135_SLICE_X5Y135_CQ;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_D2 = CLBLM_L_X10Y131_SLICE_X12Y131_BQ;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_D3 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_D4 = CLBLM_R_X11Y131_SLICE_X15Y131_BQ;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_D5 = CLBLM_L_X10Y130_SLICE_X12Y130_AQ;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_D6 = CLBLM_R_X5Y132_SLICE_X7Y132_DO6;
  assign CLBLM_R_X13Y141_SLICE_X18Y141_A6 = 1'b1;
  assign CLBLM_R_X13Y141_SLICE_X18Y141_B1 = CLBLM_L_X12Y142_SLICE_X17Y142_CO5;
  assign CLBLM_R_X13Y141_SLICE_X18Y141_B2 = CLBLM_L_X12Y142_SLICE_X16Y142_BQ;
  assign CLBLM_R_X13Y141_SLICE_X18Y141_B3 = CLBLM_R_X13Y139_SLICE_X18Y139_AQ;
  assign CLBLM_R_X13Y141_SLICE_X18Y141_B4 = CLBLM_R_X13Y140_SLICE_X18Y140_BQ;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_A1 = CLBLL_L_X4Y135_SLICE_X5Y135_CQ;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_A2 = CLBLM_R_X7Y131_SLICE_X9Y131_BQ;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_A3 = CLBLM_L_X10Y130_SLICE_X12Y130_AQ;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_A4 = CLBLM_R_X11Y131_SLICE_X15Y131_BQ;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_A5 = CLBLM_L_X10Y131_SLICE_X12Y131_BQ;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_A6 = 1'b1;
  assign CLBLM_R_X13Y141_SLICE_X18Y141_C1 = CLBLM_R_X13Y139_SLICE_X18Y139_AQ;
  assign CLBLM_R_X13Y141_SLICE_X18Y141_C2 = CLBLM_R_X13Y144_SLICE_X18Y144_AQ;
  assign CLBLM_R_X13Y141_SLICE_X18Y141_C3 = CLBLM_L_X12Y142_SLICE_X16Y142_BQ;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_B1 = CLBLM_R_X11Y131_SLICE_X14Y131_DO6;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_B3 = CLBLM_R_X7Y141_SLICE_X9Y141_AQ;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_B4 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_B5 = CLBLM_R_X7Y131_SLICE_X9Y131_AQ;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_B6 = 1'b1;
  assign CLBLM_R_X13Y141_SLICE_X18Y141_D1 = CLBLM_L_X12Y143_SLICE_X17Y143_AQ;
  assign CLBLM_R_X13Y141_SLICE_X18Y141_D2 = CLBLM_R_X13Y140_SLICE_X18Y140_BQ;
  assign CLBLM_R_X13Y141_SLICE_X18Y141_D3 = CLBLM_L_X12Y142_SLICE_X17Y142_CO5;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_C1 = CLBLM_R_X11Y131_SLICE_X15Y131_AO6;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_C2 = CLBLM_R_X11Y131_SLICE_X15Y131_CO6;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_C3 = CLBLM_R_X5Y133_SLICE_X7Y133_CO6;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_C4 = CLBLM_L_X10Y137_SLICE_X12Y137_BQ;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_C5 = CLBLM_R_X3Y139_SLICE_X3Y139_BO6;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_C6 = CLBLM_R_X13Y137_SLICE_X18Y137_A5Q;
  assign CLBLM_R_X13Y141_SLICE_X18Y141_D4 = CLBLM_R_X13Y141_SLICE_X19Y141_CO5;
  assign CLBLM_R_X13Y141_SLICE_X18Y141_D5 = CLBLM_L_X12Y142_SLICE_X16Y142_BQ;
  assign CLBLM_R_X13Y141_SLICE_X18Y141_D6 = CLBLM_R_X13Y144_SLICE_X18Y144_AQ;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_SING_X0Y100_OLOGIC_X0Y100_D1 = CLBLL_L_X2Y133_SLICE_X0Y133_BO6;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_D1 = CLBLM_R_X5Y132_SLICE_X7Y132_DO6;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_D2 = CLBLM_R_X11Y146_SLICE_X14Y146_AQ;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_D3 = CLBLM_L_X8Y131_SLICE_X10Y131_A5Q;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_D4 = CLBLM_R_X11Y131_SLICE_X14Y131_AO5;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_D5 = CLBLM_R_X11Y131_SLICE_X14Y131_BQ;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_D6 = CLBLM_L_X10Y130_SLICE_X13Y130_AO5;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_A2 = CLBLM_L_X8Y138_SLICE_X10Y138_AQ;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_A3 = CLBLL_L_X4Y134_SLICE_X4Y134_AQ;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_A4 = CLBLM_R_X11Y135_SLICE_X14Y135_AQ;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_A5 = CLBLM_R_X3Y137_SLICE_X3Y137_AQ;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_A6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X13Y143_SLICE_X19Y143_D2 = 1'b1;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_B2 = CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_B3 = 1'b1;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_B4 = CLBLM_R_X11Y135_SLICE_X14Y135_AQ;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_B5 = CLBLL_L_X4Y134_SLICE_X5Y134_A5Q;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_B6 = 1'b1;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_C1 = 1'b1;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_C2 = 1'b1;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_C3 = 1'b1;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_C4 = 1'b1;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_C5 = 1'b1;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_C6 = 1'b1;
  assign CLBLM_R_X13Y143_SLICE_X19Y143_D5 = 1'b1;
  assign CLBLM_R_X13Y143_SLICE_X19Y143_D6 = 1'b1;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_D1 = 1'b1;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_D2 = 1'b1;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_D3 = 1'b1;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_D4 = 1'b1;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_D5 = 1'b1;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_D6 = 1'b1;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_A1 = CLBLM_L_X10Y139_SLICE_X13Y139_DO6;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_A2 = CLBLM_L_X12Y135_SLICE_X17Y135_BO5;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_A3 = CLBLM_L_X10Y138_SLICE_X13Y138_AQ;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_A4 = CLBLM_L_X10Y136_SLICE_X13Y136_CO6;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_A6 = CLBLM_L_X10Y140_SLICE_X13Y140_BQ;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_B1 = CLBLM_R_X11Y140_SLICE_X15Y140_DQ;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_B2 = CLBLM_L_X10Y138_SLICE_X13Y138_BQ;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_B3 = 1'b1;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_B4 = CLBLM_R_X7Y136_SLICE_X9Y136_CQ;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_B5 = CLBLM_L_X8Y143_SLICE_X10Y143_DO6;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_A2 = CLBLL_L_X4Y134_SLICE_X5Y134_BQ;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_A3 = CLBLL_L_X4Y133_SLICE_X4Y133_BO6;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_C1 = CLBLM_L_X8Y138_SLICE_X10Y138_AQ;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_C2 = CLBLM_L_X10Y138_SLICE_X13Y138_CQ;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_C3 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_C4 = CLBLM_R_X13Y136_SLICE_X18Y136_BQ;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_C5 = CLBLM_L_X10Y138_SLICE_X13Y138_DO6;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_A4 = CLBLM_R_X5Y132_SLICE_X6Y132_AO6;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_A5 = 1'b1;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_A6 = CLBLL_L_X4Y134_SLICE_X5Y134_AQ;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_AX = CLBLL_L_X4Y134_SLICE_X5Y134_DO5;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_B1 = CLBLL_L_X4Y134_SLICE_X5Y134_DO6;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_B3 = CLBLL_L_X4Y133_SLICE_X4Y133_BO6;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_B4 = CLBLL_L_X4Y133_SLICE_X5Y133_CO6;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_D1 = CLBLM_R_X7Y136_SLICE_X9Y136_CQ;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_D2 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_D3 = CLBLM_R_X11Y139_SLICE_X14Y139_DO6;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_D4 = CLBLM_L_X10Y135_SLICE_X12Y135_BQ;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_D5 = CLBLM_R_X5Y136_SLICE_X7Y136_BQ;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_D6 = CLBLM_L_X10Y139_SLICE_X12Y139_BQ;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_C1 = CLBLM_R_X5Y132_SLICE_X6Y132_AO6;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_C4 = CLBLM_R_X7Y133_SLICE_X8Y133_CQ;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_C6 = CLBLL_L_X4Y133_SLICE_X4Y133_BO6;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_C5 = CLBLL_L_X4Y134_SLICE_X5Y134_AQ;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_A1 = CLBLM_R_X11Y135_SLICE_X14Y135_AQ;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_A3 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_A4 = 1'b1;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_A2 = CLBLM_R_X11Y133_SLICE_X14Y133_BQ;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_D1 = CLBLL_L_X4Y134_SLICE_X5Y134_BQ;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_A5 = CLBLM_R_X7Y138_SLICE_X9Y138_CO6;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_D2 = CLBLL_L_X4Y134_SLICE_X5Y134_CQ;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_D3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_D4 = CLBLL_L_X4Y134_SLICE_X5Y134_AQ;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_D6 = 1'b1;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_AX = CLBLM_R_X11Y137_SLICE_X14Y137_BO6;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_D5 = CLBLL_L_X4Y133_SLICE_X5Y133_AQ;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_B1 = CLBLM_R_X5Y136_SLICE_X7Y136_BQ;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_B2 = CLBLM_R_X7Y136_SLICE_X9Y136_CQ;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_B3 = CLBLM_L_X10Y139_SLICE_X13Y139_AQ;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_B4 = CLBLM_L_X10Y139_SLICE_X13Y139_BQ;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_B5 = CLBLM_R_X11Y139_SLICE_X15Y139_CQ;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_B6 = 1'b1;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_C1 = CLBLM_L_X10Y139_SLICE_X13Y139_AQ;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_C2 = CLBLM_R_X11Y139_SLICE_X15Y139_CQ;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_C3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_C4 = CLBLM_R_X11Y136_SLICE_X15Y136_BQ;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_C5 = CLBLM_L_X10Y138_SLICE_X12Y138_DO6;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_C6 = CLBLM_L_X8Y138_SLICE_X11Y138_BQ;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_C6 = 1'b1;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_C4 = 1'b1;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_D1 = CLBLM_R_X7Y136_SLICE_X9Y136_CQ;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_D2 = 1'b1;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_D3 = CLBLM_R_X5Y136_SLICE_X7Y136_BQ;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_D4 = 1'b1;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_D5 = 1'b1;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_D6 = 1'b1;
  assign CLBLM_R_X13Y143_SLICE_X18Y143_B5 = CLBLM_R_X13Y141_SLICE_X18Y141_CO5;
  assign CLBLM_R_X13Y143_SLICE_X18Y143_B6 = CLBLM_L_X12Y140_SLICE_X17Y140_AQ;
  assign RIOB33_X105Y195_IOB_X1Y195_O = CLBLM_R_X13Y143_SLICE_X18Y143_BQ;
  assign RIOB33_X105Y195_IOB_X1Y196_O = CLBLM_R_X13Y143_SLICE_X18Y143_AQ;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_C5 = 1'b1;
  assign CLBLM_R_X13Y142_SLICE_X19Y142_A1 = CLBLM_L_X12Y143_SLICE_X17Y143_DO6;
  assign CLBLM_R_X13Y142_SLICE_X19Y142_A2 = CLBLM_R_X13Y141_SLICE_X18Y141_AO5;
  assign CLBLM_R_X13Y142_SLICE_X19Y142_A3 = CLBLM_L_X12Y137_SLICE_X17Y137_AQ;
  assign CLBLM_R_X13Y142_SLICE_X19Y142_A4 = CLBLM_R_X13Y142_SLICE_X19Y142_BO6;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_D3 = 1'b1;
  assign CLBLM_R_X13Y142_SLICE_X19Y142_A5 = 1'b1;
  assign CLBLM_R_X13Y142_SLICE_X19Y142_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y142_SLICE_X19Y142_B1 = CLBLM_R_X13Y141_SLICE_X18Y141_BO5;
  assign CLBLM_R_X13Y142_SLICE_X19Y142_B2 = CLBLM_R_X13Y143_SLICE_X19Y143_BO6;
  assign CLBLM_R_X13Y142_SLICE_X19Y142_B3 = CLBLM_L_X12Y140_SLICE_X16Y140_BQ;
  assign CLBLM_R_X13Y142_SLICE_X19Y142_B4 = CLBLM_R_X13Y142_SLICE_X19Y142_AQ;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_D5 = 1'b1;
  assign CLBLM_R_X13Y142_SLICE_X19Y142_B5 = CLBLM_R_X13Y144_SLICE_X18Y144_CO6;
  assign CLBLM_R_X13Y142_SLICE_X19Y142_B6 = CLBLM_R_X13Y143_SLICE_X19Y143_AO6;
  assign CLBLM_R_X13Y143_SLICE_X18Y143_C4 = CLBLM_L_X12Y140_SLICE_X17Y140_AQ;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_D6 = 1'b1;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_A1 = CLBLL_L_X4Y135_SLICE_X5Y135_CQ;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_A2 = CLBLM_L_X10Y131_SLICE_X12Y131_BQ;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_A3 = CLBLM_L_X10Y130_SLICE_X12Y130_AQ;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_A4 = CLBLM_R_X11Y131_SLICE_X15Y131_BQ;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_A5 = CLBLM_R_X11Y132_SLICE_X15Y132_CO6;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_A6 = 1'b1;
  assign CLBLM_R_X13Y142_SLICE_X19Y142_C1 = CLBLM_R_X13Y140_SLICE_X19Y140_BQ;
  assign CLBLM_R_X13Y142_SLICE_X19Y142_C2 = CLBLM_L_X12Y141_SLICE_X16Y141_AQ;
  assign CLBLM_R_X13Y142_SLICE_X19Y142_C3 = CLBLM_R_X13Y143_SLICE_X18Y143_DO6;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_B1 = CLBLM_L_X12Y132_SLICE_X16Y132_CQ;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_B2 = CLBLM_R_X11Y131_SLICE_X15Y131_BQ;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_B3 = CLBLM_R_X5Y132_SLICE_X7Y132_DO6;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_B4 = CLBLM_R_X7Y131_SLICE_X9Y131_BQ;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_B5 = CLBLM_R_X11Y131_SLICE_X15Y131_AO5;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_B6 = CLBLM_L_X12Y136_SLICE_X16Y136_B5Q;
  assign CLBLM_R_X13Y142_SLICE_X19Y142_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y142_SLICE_X19Y142_D1 = CLBLM_R_X13Y143_SLICE_X18Y143_CO6;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_C1 = CLBLM_L_X12Y132_SLICE_X16Y132_BQ;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_C2 = CLBLM_R_X11Y132_SLICE_X14Y132_CO6;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_C3 = CLBLM_L_X12Y136_SLICE_X16Y136_DQ;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_C4 = CLBLM_L_X10Y133_SLICE_X13Y133_CO6;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_C5 = 1'b1;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_C6 = 1'b1;
  assign CLBLM_R_X13Y142_SLICE_X19Y142_D3 = CLBLM_R_X13Y140_SLICE_X19Y140_BQ;
  assign CLBLM_R_X13Y142_SLICE_X19Y142_D4 = CLBLM_R_X13Y140_SLICE_X18Y140_AQ;
  assign CLBLM_R_X13Y142_SLICE_X18Y142_A1 = CLBLM_R_X13Y143_SLICE_X18Y143_DO6;
  assign CLBLM_R_X13Y142_SLICE_X18Y142_A2 = CLBLM_R_X11Y141_SLICE_X15Y141_CQ;
  assign CLBLM_R_X13Y142_SLICE_X18Y142_A3 = CLBLM_L_X12Y141_SLICE_X16Y141_AQ;
  assign CLBLM_R_X13Y142_SLICE_X18Y142_A4 = CLBLM_R_X13Y144_SLICE_X18Y144_CO6;
  assign CLBLM_R_X13Y142_SLICE_X18Y142_A5 = CLBLM_R_X13Y143_SLICE_X18Y143_CO6;
  assign CLBLM_R_X13Y142_SLICE_X18Y142_A6 = CLBLM_R_X13Y141_SLICE_X18Y141_BO5;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_D1 = 1'b1;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_D2 = CLBLM_R_X11Y133_SLICE_X15Y133_CQ;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_D3 = CLBLM_R_X11Y134_SLICE_X15Y134_CQ;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_D4 = 1'b1;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_D5 = CLBLM_L_X8Y134_SLICE_X11Y134_BQ;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_D6 = CLBLM_L_X10Y134_SLICE_X12Y134_AQ;
  assign CLBLM_R_X13Y142_SLICE_X18Y142_B2 = CLBLM_R_X13Y140_SLICE_X19Y140_BQ;
  assign CLBLM_R_X13Y142_SLICE_X18Y142_B3 = CLBLM_R_X13Y144_SLICE_X18Y144_CO6;
  assign CLBLM_R_X13Y142_SLICE_X18Y142_B4 = CLBLM_R_X13Y141_SLICE_X18Y141_BO5;
  assign CLBLM_R_X13Y142_SLICE_X18Y142_B5 = CLBLM_L_X12Y143_SLICE_X16Y143_CQ;
  assign CLBLM_R_X13Y142_SLICE_X18Y142_B6 = CLBLM_R_X13Y142_SLICE_X18Y142_CO6;
  assign CLBLM_R_X13Y142_SLICE_X18Y142_B1 = CLBLM_R_X13Y142_SLICE_X18Y142_DO6;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_A1 = 1'b1;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_A2 = CLBLM_L_X10Y131_SLICE_X13Y131_BQ;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_A3 = CLBLM_R_X11Y132_SLICE_X14Y132_AQ;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_A4 = CLBLM_R_X11Y134_SLICE_X14Y134_BQ;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_A5 = CLBLM_R_X5Y132_SLICE_X7Y132_DO6;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y142_SLICE_X18Y142_C1 = CLBLM_R_X13Y141_SLICE_X18Y141_CO5;
  assign CLBLM_R_X13Y142_SLICE_X18Y142_C2 = CLBLM_R_X13Y140_SLICE_X18Y140_AQ;
  assign CLBLM_R_X13Y142_SLICE_X18Y142_C3 = CLBLM_L_X12Y141_SLICE_X16Y141_AQ;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_B1 = CLBLM_R_X11Y132_SLICE_X14Y132_DO6;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_B2 = CLBLM_R_X11Y133_SLICE_X14Y133_CQ;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_B3 = CLBLM_R_X7Y131_SLICE_X9Y131_AQ;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_B4 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_B5 = 1'b1;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y142_SLICE_X18Y142_D1 = CLBLM_R_X13Y141_SLICE_X18Y141_CO5;
  assign CLBLM_R_X13Y142_SLICE_X18Y142_D2 = CLBLM_R_X13Y140_SLICE_X18Y140_AQ;
  assign CLBLM_R_X13Y142_SLICE_X18Y142_D3 = CLBLM_L_X12Y141_SLICE_X16Y141_AQ;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_C1 = CLBLM_R_X11Y133_SLICE_X15Y133_AQ;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_C2 = CLBLM_R_X11Y133_SLICE_X14Y133_BQ;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_C3 = CLBLM_L_X8Y131_SLICE_X10Y131_BO5;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_C4 = CLBLM_R_X11Y133_SLICE_X14Y133_AQ;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_C5 = CLBLM_R_X7Y131_SLICE_X9Y131_BQ;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_C6 = CLBLM_R_X11Y133_SLICE_X15Y133_BQ;
  assign CLBLM_R_X13Y142_SLICE_X18Y142_D4 = CLBLM_L_X12Y140_SLICE_X17Y140_AQ;
  assign CLBLM_R_X13Y142_SLICE_X18Y142_D5 = CLBLM_L_X12Y142_SLICE_X17Y142_AQ;
  assign CLBLM_R_X13Y142_SLICE_X18Y142_D6 = CLBLM_L_X12Y142_SLICE_X16Y142_AQ;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_B4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y143_SLICE_X18Y143_D5 = CLBLM_R_X13Y144_SLICE_X18Y144_AQ;
  assign CLBLM_R_X103Y140_SLICE_X162Y140_D6 = 1'b1;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_D1 = CLBLM_R_X5Y132_SLICE_X7Y132_DO6;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_D2 = 1'b1;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_D3 = CLBLM_R_X11Y132_SLICE_X14Y132_BQ;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_D4 = 1'b1;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_D5 = CLBLM_L_X10Y130_SLICE_X13Y130_AO6;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_D6 = CLBLM_L_X10Y137_SLICE_X12Y137_B5Q;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_B1 = CLBLM_L_X10Y143_SLICE_X13Y143_DO6;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_A1 = 1'b1;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_A2 = CLBLM_R_X7Y137_SLICE_X9Y137_BQ;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_A3 = CLBLL_L_X4Y135_SLICE_X4Y135_AQ;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_A5 = CLBLM_L_X12Y133_SLICE_X16Y133_C5Q;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_A6 = CLBLM_R_X7Y144_SLICE_X9Y144_BO6;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_C1 = 1'b1;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_B5 = 1'b1;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_AX = CLBLL_L_X4Y135_SLICE_X4Y135_DO6;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_C2 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_B1 = CLBLL_L_X4Y135_SLICE_X5Y135_DQ;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_B2 = CLBLL_L_X4Y135_SLICE_X4Y135_BQ;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_B4 = 1'b1;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_B5 = CLBLM_L_X10Y134_SLICE_X13Y134_BQ;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_B6 = CLBLM_R_X7Y144_SLICE_X9Y144_BO6;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_B6 = 1'b1;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_C1 = 1'b1;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_C2 = CLBLL_L_X4Y135_SLICE_X4Y135_CQ;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_C3 = CLBLM_R_X3Y135_SLICE_X3Y135_AQ;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_C4 = CLBLM_R_X7Y135_SLICE_X9Y135_A5Q;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_C6 = CLBLM_R_X7Y144_SLICE_X9Y144_BO6;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_D1 = CLBLM_R_X3Y136_SLICE_X2Y136_AQ;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_D1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_D2 = CLBLM_R_X5Y137_SLICE_X6Y137_BQ;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_D3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_D4 = CLBLL_L_X4Y135_SLICE_X4Y135_A5Q;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_D5 = CLBLM_R_X5Y138_SLICE_X7Y138_CQ;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_D6 = 1'b1;
  assign LIOI3_X0Y197_OLOGIC_X0Y198_D1 = LIOB33_X0Y73_IOB_X0Y73_I;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y197_OLOGIC_X0Y198_T1 = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_D1 = CLBLM_R_X3Y135_SLICE_X3Y135_AQ;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_C4 = 1'b1;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_A1 = 1'b1;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_A2 = CLBLM_R_X7Y139_SLICE_X9Y139_AQ;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_A3 = CLBLM_L_X10Y139_SLICE_X13Y139_AQ;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_A4 = CLBLM_L_X10Y139_SLICE_X12Y139_BQ;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_C5 = 1'b1;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_C6 = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_T1 = 1'b1;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_B1 = CLBLM_R_X7Y136_SLICE_X8Y136_AQ;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_A1 = CLBLM_L_X8Y138_SLICE_X10Y138_AQ;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_A2 = CLBLM_L_X8Y134_SLICE_X11Y134_DQ;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_A3 = CLBLL_L_X4Y135_SLICE_X5Y135_AQ;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_B6 = 1'b1;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_A5 = CLBLL_L_X4Y135_SLICE_X4Y135_AQ;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_A6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_B2 = CLBLM_L_X10Y139_SLICE_X13Y139_BQ;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_B3 = CLBLM_R_X11Y144_SLICE_X15Y144_AQ;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_C3 = CLBLM_L_X8Y142_SLICE_X11Y142_AQ;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_C4 = CLBLM_R_X11Y135_SLICE_X15Y135_DO6;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_C6 = CLBLM_R_X7Y131_SLICE_X9Y131_AQ;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_B1 = 1'b1;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_B4 = CLBLL_L_X4Y135_SLICE_X5Y135_D5Q;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_B5 = CLBLM_R_X7Y137_SLICE_X9Y137_BQ;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_B6 = CLBLM_R_X7Y135_SLICE_X9Y135_DO6;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_C1 = CLBLM_R_X7Y137_SLICE_X9Y137_BQ;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_C2 = CLBLM_L_X8Y134_SLICE_X10Y134_DO6;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_C4 = CLBLL_L_X4Y135_SLICE_X4Y135_CQ;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_C5 = CLBLM_R_X5Y132_SLICE_X6Y132_AO6;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_C6 = 1'b1;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_D6 = CLBLM_R_X13Y141_SLICE_X19Y141_BQ;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_D1 = CLBLM_L_X8Y137_SLICE_X10Y137_BO6;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_D2 = CLBLM_L_X10Y140_SLICE_X13Y140_CQ;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_D3 = CLBLM_L_X10Y139_SLICE_X12Y139_DO6;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_D4 = CLBLM_R_X11Y139_SLICE_X14Y139_DO6;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_D5 = CLBLM_L_X12Y135_SLICE_X17Y135_AQ;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_D1 = CLBLM_R_X7Y135_SLICE_X8Y135_AQ;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_D2 = CLBLM_R_X7Y136_SLICE_X8Y136_BQ;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_D3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_A2 = CLBLM_L_X10Y140_SLICE_X12Y140_BQ;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_A3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_A4 = CLBLM_R_X13Y139_SLICE_X18Y139_BO6;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_A5 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_D4 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_D5 = 1'b1;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_D6 = 1'b1;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_B1 = 1'b1;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_B2 = CLBLM_L_X10Y139_SLICE_X12Y139_BQ;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_B5 = 1'b1;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_B6 = CLBLM_L_X8Y136_SLICE_X11Y136_CQ;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_D1 = RIOB33_X105Y121_IOB_X1Y122_I;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_C1 = CLBLM_R_X11Y139_SLICE_X14Y139_BQ;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_C2 = CLBLM_R_X5Y137_SLICE_X7Y137_BQ;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_C3 = CLBLM_L_X10Y139_SLICE_X12Y139_BQ;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_C4 = CLBLM_L_X8Y138_SLICE_X11Y138_BQ;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_C5 = CLBLM_L_X10Y134_SLICE_X12Y134_DQ;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_C6 = CLBLM_L_X8Y144_SLICE_X11Y144_AQ;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_T1 = 1'b1;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_B4 = CLBLM_L_X12Y135_SLICE_X17Y135_AQ;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_A1 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_D1 = CLBLM_L_X10Y140_SLICE_X12Y140_BQ;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_D2 = CLBLM_R_X13Y141_SLICE_X19Y141_BQ;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_D4 = CLBLM_L_X10Y139_SLICE_X12Y139_CO6;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_D5 = CLBLM_L_X8Y141_SLICE_X10Y141_CQ;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_D6 = CLBLM_L_X10Y139_SLICE_X13Y139_BQ;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_D3 = CLBLM_L_X10Y137_SLICE_X12Y137_DO6;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_D1 = CLBLM_R_X7Y131_SLICE_X9Y131_AQ;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_C1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_C2 = CLBLM_L_X8Y141_SLICE_X11Y141_CQ;
  assign CLBLM_R_X13Y143_SLICE_X19Y143_A1 = CLBLM_L_X12Y141_SLICE_X16Y141_AQ;
  assign CLBLM_R_X13Y143_SLICE_X19Y143_A2 = CLBLM_R_X13Y140_SLICE_X18Y140_AQ;
  assign CLBLM_R_X13Y143_SLICE_X19Y143_A3 = CLBLM_R_X13Y140_SLICE_X19Y140_BQ;
  assign CLBLM_R_X13Y143_SLICE_X19Y143_A4 = CLBLM_R_X13Y143_SLICE_X18Y143_CO6;
  assign CLBLM_R_X13Y143_SLICE_X19Y143_A5 = CLBLM_L_X12Y142_SLICE_X17Y142_BQ;
  assign CLBLM_R_X13Y143_SLICE_X19Y143_A6 = 1'b1;
  assign CLBLM_R_X13Y143_SLICE_X19Y143_B1 = CLBLM_L_X12Y141_SLICE_X16Y141_AQ;
  assign CLBLM_R_X13Y143_SLICE_X19Y143_B2 = CLBLM_R_X13Y140_SLICE_X18Y140_AQ;
  assign CLBLM_R_X13Y143_SLICE_X19Y143_B3 = CLBLM_R_X13Y140_SLICE_X19Y140_BQ;
  assign CLBLM_R_X13Y143_SLICE_X19Y143_B4 = CLBLM_R_X13Y143_SLICE_X18Y143_DO6;
  assign CLBLM_R_X13Y143_SLICE_X19Y143_B5 = CLBLM_L_X12Y142_SLICE_X17Y142_BQ;
  assign CLBLM_R_X13Y143_SLICE_X19Y143_B6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_T1 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_A2 = CLBLM_R_X11Y133_SLICE_X15Y133_BQ;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_A3 = CLBLM_R_X11Y133_SLICE_X15Y133_AQ;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_A4 = CLBLM_R_X5Y133_SLICE_X7Y133_DO6;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_A5 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_A6 = CLBLM_L_X10Y140_SLICE_X12Y140_A5Q;
  assign CLBLM_R_X13Y143_SLICE_X19Y143_C1 = 1'b1;
  assign CLBLM_R_X13Y143_SLICE_X19Y143_C2 = 1'b1;
  assign CLBLM_R_X13Y143_SLICE_X19Y143_C3 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_B2 = CLBLM_R_X11Y133_SLICE_X15Y133_BQ;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_B3 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_B4 = CLBLM_R_X5Y134_SLICE_X7Y134_DO6;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_B5 = CLBLM_R_X7Y131_SLICE_X9Y131_BQ;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_B6 = CLBLM_L_X12Y136_SLICE_X17Y136_CQ;
  assign CLBLM_R_X13Y143_SLICE_X19Y143_D1 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_C2 = CLBLM_R_X11Y133_SLICE_X15Y133_CQ;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_C3 = CLBLM_R_X11Y134_SLICE_X15Y134_CQ;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_C4 = CLBLM_R_X11Y140_SLICE_X15Y140_BQ;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_C5 = CLBLM_R_X5Y132_SLICE_X7Y132_DO6;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_C6 = 1'b1;
  assign CLBLM_R_X13Y143_SLICE_X19Y143_D3 = 1'b1;
  assign CLBLM_R_X13Y143_SLICE_X19Y143_D4 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y143_SLICE_X18Y143_A1 = CLBLM_R_X13Y137_SLICE_X18Y137_CO5;
  assign CLBLM_R_X13Y143_SLICE_X18Y143_A2 = CLBLM_R_X13Y140_SLICE_X18Y140_BQ;
  assign CLBLM_R_X13Y143_SLICE_X18Y143_A3 = CLBLM_L_X12Y142_SLICE_X16Y142_BQ;
  assign CLBLM_R_X13Y143_SLICE_X18Y143_A4 = CLBLM_R_X13Y144_SLICE_X18Y144_AQ;
  assign CLBLM_R_X13Y143_SLICE_X18Y143_A5 = CLBLM_L_X12Y143_SLICE_X17Y143_BQ;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_D1 = CLBLM_R_X7Y131_SLICE_X9Y131_AQ;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_D2 = CLBLM_L_X12Y133_SLICE_X17Y133_BQ;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_D3 = CLBLM_R_X11Y133_SLICE_X14Y133_DO6;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_D4 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_D6 = 1'b1;
  assign CLBLM_R_X13Y143_SLICE_X18Y143_A6 = 1'b1;
  assign CLBLM_R_X13Y143_SLICE_X18Y143_AX = CLBLM_R_X13Y140_SLICE_X18Y140_BQ;
  assign CLBLM_R_X13Y143_SLICE_X18Y143_B1 = CLBLM_L_X12Y141_SLICE_X16Y141_AQ;
  assign CLBLM_R_X13Y143_SLICE_X18Y143_B2 = CLBLM_L_X12Y142_SLICE_X16Y142_AQ;
  assign CLBLM_R_X13Y143_SLICE_X18Y143_B3 = CLBLM_L_X12Y142_SLICE_X17Y142_AQ;
  assign CLBLM_R_X13Y143_SLICE_X18Y143_B4 = CLBLM_R_X13Y140_SLICE_X18Y140_AQ;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_A1 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_A2 = CLBLM_R_X11Y133_SLICE_X14Y133_BQ;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_A3 = CLBLM_R_X11Y133_SLICE_X14Y133_AQ;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_A4 = CLBLM_R_X5Y134_SLICE_X7Y134_DO6;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_A5 = CLBLM_L_X10Y142_SLICE_X13Y142_AQ;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y143_SLICE_X18Y143_BX = CLBLM_L_X12Y143_SLICE_X16Y143_CQ;
  assign CLBLM_R_X13Y143_SLICE_X18Y143_C1 = CLBLM_L_X12Y142_SLICE_X17Y142_AQ;
  assign CLBLM_R_X13Y143_SLICE_X18Y143_C2 = CLBLM_R_X13Y140_SLICE_X18Y140_BQ;
  assign CLBLM_R_X13Y143_SLICE_X18Y143_C3 = CLBLM_L_X12Y142_SLICE_X16Y142_BQ;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_B1 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_B2 = CLBLM_R_X11Y133_SLICE_X14Y133_BQ;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_B4 = CLBLM_R_X5Y134_SLICE_X7Y134_DO6;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_B5 = CLBLM_R_X11Y132_SLICE_X14Y132_AQ;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_B6 = CLBLM_R_X11Y140_SLICE_X14Y140_AQ;
  assign CLBLM_R_X13Y143_SLICE_X18Y143_CE = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y143_SLICE_X18Y143_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y143_SLICE_X18Y143_D1 = CLBLM_L_X12Y142_SLICE_X17Y142_AQ;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_C1 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_C2 = CLBLM_R_X11Y133_SLICE_X14Y133_CQ;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_C5 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_C6 = CLBLM_R_X7Y134_SLICE_X8Y134_AQ;
  assign CLBLM_R_X13Y143_SLICE_X18Y143_D2 = CLBLM_R_X13Y140_SLICE_X18Y140_BQ;
  assign CLBLM_R_X13Y143_SLICE_X18Y143_D3 = CLBLM_L_X12Y142_SLICE_X16Y142_BQ;
  assign CLBLM_R_X13Y143_SLICE_X18Y143_D4 = CLBLM_L_X12Y140_SLICE_X17Y140_AQ;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y143_SLICE_X18Y143_D6 = CLBLM_L_X12Y142_SLICE_X16Y142_AQ;
  assign CLBLM_R_X13Y143_SLICE_X18Y143_SR = CLBLM_L_X12Y144_SLICE_X16Y144_AO6;
  assign RIOI3_X105Y121_ILOGIC_X1Y122_D = RIOB33_X105Y121_IOB_X1Y122_I;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_D1 = CLBLM_R_X11Y131_SLICE_X15Y131_BQ;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_D2 = CLBLM_L_X10Y131_SLICE_X13Y131_CQ;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_D3 = CLBLM_R_X5Y132_SLICE_X7Y132_DO6;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_D4 = CLBLM_L_X10Y137_SLICE_X12Y137_BQ;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_D5 = CLBLM_R_X11Y133_SLICE_X15Y133_DQ;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_D6 = CLBLM_L_X10Y133_SLICE_X12Y133_DO6;
  assign RIOI3_X105Y121_ILOGIC_X1Y121_D = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_A1 = CLBLL_L_X4Y137_SLICE_X4Y137_CQ;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_A2 = CLBLL_L_X4Y136_SLICE_X4Y136_BQ;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_A3 = CLBLM_L_X12Y135_SLICE_X17Y135_AQ;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_A6 = 1'b1;
  assign CLBLM_R_X13Y143_SLICE_X18Y143_C5 = CLBLM_L_X12Y142_SLICE_X16Y142_AQ;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_B2 = CLBLL_L_X4Y136_SLICE_X4Y136_BQ;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_B3 = CLBLM_R_X7Y144_SLICE_X9Y144_BO6;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_B4 = 1'b1;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_B5 = CLBLM_R_X7Y132_SLICE_X8Y132_CQ;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_B6 = CLBLL_L_X4Y136_SLICE_X4Y136_DQ;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_T1 = 1'b1;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_C1 = 1'b1;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_C2 = CLBLL_L_X4Y136_SLICE_X4Y136_CQ;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_C3 = CLBLL_L_X4Y137_SLICE_X4Y137_DQ;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_C4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_C5 = CLBLM_L_X8Y138_SLICE_X10Y138_AQ;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y143_SLICE_X18Y143_C6 = CLBLM_R_X13Y144_SLICE_X18Y144_AQ;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_D1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_D2 = CLBLM_R_X5Y141_SLICE_X6Y141_A5Q;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_D3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_D4 = CLBLM_R_X7Y135_SLICE_X9Y135_A5Q;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_D5 = CLBLL_L_X4Y136_SLICE_X4Y136_AQ;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_D6 = 1'b1;
  assign LIOB33_X0Y113_IOB_X0Y114_O = CLBLM_R_X7Y132_SLICE_X9Y132_DQ;
  assign LIOB33_X0Y113_IOB_X0Y113_O = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_A1 = CLBLM_L_X10Y135_SLICE_X12Y135_BQ;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_A2 = CLBLM_L_X10Y140_SLICE_X12Y140_CQ;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_A3 = CLBLM_R_X3Y138_SLICE_X3Y138_AQ;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_A5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_A6 = 1'b1;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_A1 = CLBLM_R_X11Y138_SLICE_X14Y138_BQ;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_A2 = CLBLM_R_X5Y135_SLICE_X6Y135_CQ;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_A3 = CLBLL_L_X4Y136_SLICE_X5Y136_AQ;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_A4 = CLBLM_L_X12Y135_SLICE_X17Y135_AQ;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_A6 = CLBLL_L_X4Y137_SLICE_X4Y137_CQ;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_B1 = CLBLM_L_X12Y138_SLICE_X16Y138_DQ;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_AX = CLBLL_L_X4Y137_SLICE_X5Y137_AO6;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_B2 = CLBLL_L_X4Y136_SLICE_X5Y136_BQ;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_B3 = CLBLL_L_X4Y133_SLICE_X4Y133_AQ;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_B4 = CLBLM_R_X7Y139_SLICE_X8Y139_AQ;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_B5 = CLBLM_L_X12Y135_SLICE_X17Y135_AQ;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_B6 = CLBLL_L_X4Y137_SLICE_X4Y137_CQ;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_B4 = 1'b1;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_C1 = CLBLL_L_X4Y135_SLICE_X5Y135_AQ;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_C2 = CLBLL_L_X4Y136_SLICE_X5Y136_CQ;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_C4 = CLBLM_R_X7Y133_SLICE_X8Y133_DO6;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_C5 = 1'b1;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_C6 = 1'b1;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_C5 = CLBLM_R_X5Y141_SLICE_X7Y141_DO6;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_D1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_D2 = CLBLM_R_X7Y133_SLICE_X9Y133_CQ;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_D3 = CLBLM_R_X11Y141_SLICE_X15Y141_DQ;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_D1 = CLBLM_R_X5Y136_SLICE_X7Y136_AQ;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_D2 = CLBLM_R_X5Y137_SLICE_X6Y137_CQ;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_D3 = RIOB33_X105Y127_IOB_X1Y127_I;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_D4 = CLBLM_R_X5Y135_SLICE_X7Y135_DO6;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_D6 = 1'b1;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_D4 = 1'b1;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_A1 = CLBLM_L_X12Y140_SLICE_X16Y140_DQ;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_A2 = CLBLM_L_X8Y143_SLICE_X10Y143_DO6;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_A3 = CLBLM_L_X10Y140_SLICE_X12Y140_AQ;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_A5 = 1'b1;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_A6 = CLBLM_L_X10Y141_SLICE_X12Y141_CQ;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_AX = CLBLM_L_X10Y141_SLICE_X12Y141_BO6;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_B2 = CLBLM_L_X10Y140_SLICE_X12Y140_BQ;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_B3 = CLBLM_L_X10Y140_SLICE_X12Y140_CQ;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_B5 = CLBLM_L_X8Y140_SLICE_X11Y140_AQ;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_B6 = 1'b1;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_C1 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_C2 = CLBLM_L_X10Y140_SLICE_X12Y140_CQ;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_C3 = CLBLM_L_X10Y136_SLICE_X12Y136_DO6;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_C4 = CLBLM_L_X8Y138_SLICE_X10Y138_AQ;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_C5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOB33_X105Y173_IOB_X1Y174_O = CLBLM_R_X103Y173_SLICE_X163Y173_AO6;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_D1 = CLBLM_L_X10Y140_SLICE_X12Y140_A5Q;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_D2 = CLBLM_R_X11Y140_SLICE_X14Y140_DO6;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_D3 = CLBLM_R_X11Y141_SLICE_X15Y141_DQ;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_D4 = CLBLM_R_X11Y140_SLICE_X15Y140_BQ;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_D5 = CLBLM_L_X10Y140_SLICE_X12Y140_BO5;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_D6 = CLBLM_L_X10Y140_SLICE_X13Y140_BQ;
  assign RIOB33_X105Y173_IOB_X1Y173_O = CLBLM_R_X11Y144_SLICE_X14Y144_BO5;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_A1 = CLBLM_L_X12Y134_SLICE_X16Y134_AQ;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_A2 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_A3 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_A4 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_A5 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_A6 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_B1 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_B2 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_B3 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_B4 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_B5 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_B6 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_C1 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_C2 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_C3 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_C4 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_C5 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_C6 = 1'b1;
  assign CLBLM_R_X13Y144_SLICE_X19Y144_A1 = CLBLM_L_X10Y145_SLICE_X13Y145_AQ;
  assign CLBLM_R_X13Y144_SLICE_X19Y144_A2 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X13Y144_SLICE_X19Y144_A3 = CLBLM_R_X13Y144_SLICE_X19Y144_AQ;
  assign CLBLM_R_X13Y144_SLICE_X19Y144_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y144_SLICE_X19Y144_A5 = 1'b1;
  assign CLBLM_R_X13Y144_SLICE_X19Y144_A6 = CLBLM_R_X7Y131_SLICE_X9Y131_AQ;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_D1 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_D2 = 1'b1;
  assign CLBLM_R_X13Y144_SLICE_X19Y144_B1 = 1'b1;
  assign CLBLM_R_X13Y144_SLICE_X19Y144_B2 = 1'b1;
  assign CLBLM_R_X13Y144_SLICE_X19Y144_B3 = 1'b1;
  assign CLBLM_R_X13Y144_SLICE_X19Y144_B4 = 1'b1;
  assign CLBLM_R_X13Y144_SLICE_X19Y144_B5 = 1'b1;
  assign CLBLM_R_X13Y144_SLICE_X19Y144_B6 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_A1 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_A2 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_A3 = 1'b1;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_A1 = 1'b1;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_A2 = CLBLM_L_X8Y133_SLICE_X11Y133_BQ;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_A3 = CLBLM_R_X11Y134_SLICE_X15Y134_AQ;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_A5 = CLBLM_L_X8Y143_SLICE_X10Y143_DO6;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_A6 = CLBLM_L_X8Y140_SLICE_X11Y140_AQ;
  assign CLBLM_R_X13Y144_SLICE_X19Y144_C1 = 1'b1;
  assign CLBLM_R_X13Y144_SLICE_X19Y144_C2 = 1'b1;
  assign CLBLM_R_X13Y144_SLICE_X19Y144_C3 = 1'b1;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_B1 = CLBLM_L_X8Y134_SLICE_X11Y134_CQ;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_B2 = CLBLM_R_X11Y134_SLICE_X15Y134_BQ;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_B3 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_B4 = CLBLM_L_X8Y138_SLICE_X10Y138_AQ;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_B5 = CLBLM_R_X11Y139_SLICE_X15Y139_BQ;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y144_SLICE_X19Y144_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y144_SLICE_X19Y144_D1 = 1'b1;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_C1 = CLBLM_R_X5Y133_SLICE_X7Y133_DO6;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_C2 = CLBLM_R_X11Y134_SLICE_X15Y134_CQ;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_C3 = CLBLM_L_X12Y138_SLICE_X17Y138_AQ;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_C4 = 1'b1;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_C5 = CLBLM_L_X10Y134_SLICE_X12Y134_AQ;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y144_SLICE_X19Y144_D3 = 1'b1;
  assign CLBLM_R_X13Y144_SLICE_X19Y144_D4 = 1'b1;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y144_SLICE_X18Y144_A1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X13Y144_SLICE_X18Y144_A2 = CLBLM_R_X13Y144_SLICE_X18Y144_BO5;
  assign CLBLM_R_X13Y144_SLICE_X18Y144_A3 = CLBLM_R_X13Y144_SLICE_X18Y144_AQ;
  assign CLBLM_R_X13Y144_SLICE_X18Y144_A4 = CLBLM_R_X13Y141_SLICE_X19Y141_CO5;
  assign CLBLM_R_X13Y144_SLICE_X18Y144_A5 = CLBLM_L_X12Y143_SLICE_X16Y143_AQ;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_D1 = CLBLM_L_X8Y132_SLICE_X11Y132_BQ;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_D2 = CLBLM_R_X11Y139_SLICE_X14Y139_AQ;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_D3 = 1'b1;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_D4 = CLBLM_L_X8Y134_SLICE_X11Y134_AQ;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_D5 = 1'b1;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_D6 = CLBLM_R_X7Y133_SLICE_X9Y133_AQ;
  assign CLBLM_R_X13Y144_SLICE_X18Y144_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y144_SLICE_X18Y144_B1 = CLBLM_R_X13Y140_SLICE_X18Y140_BQ;
  assign CLBLM_R_X13Y144_SLICE_X18Y144_B2 = CLBLM_L_X12Y143_SLICE_X17Y143_BQ;
  assign CLBLM_R_X13Y144_SLICE_X18Y144_B3 = CLBLM_R_X13Y144_SLICE_X18Y144_AQ;
  assign CLBLM_R_X13Y144_SLICE_X18Y144_B4 = CLBLM_R_X13Y140_SLICE_X19Y140_AQ;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_A1 = CLBLM_L_X10Y135_SLICE_X12Y135_DO6;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_A3 = CLBLM_R_X11Y134_SLICE_X14Y134_AQ;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_A4 = CLBLM_L_X12Y135_SLICE_X16Y135_BQ;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_A5 = CLBLM_R_X5Y136_SLICE_X7Y136_BQ;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_A6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X13Y141_SLICE_X18Y141_B5 = CLBLM_R_X13Y137_SLICE_X18Y137_CO5;
  assign CLBLM_R_X13Y144_SLICE_X18Y144_C1 = CLBLM_L_X12Y142_SLICE_X16Y142_BQ;
  assign CLBLM_R_X13Y144_SLICE_X18Y144_C2 = CLBLM_L_X12Y143_SLICE_X17Y143_BQ;
  assign CLBLM_R_X13Y144_SLICE_X18Y144_C3 = CLBLM_R_X13Y144_SLICE_X18Y144_AQ;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_B1 = CLBLM_L_X10Y135_SLICE_X12Y135_DO6;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_B2 = CLBLM_R_X11Y134_SLICE_X14Y134_BQ;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_B3 = CLBLM_R_X11Y134_SLICE_X14Y134_CQ;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_B5 = CLBLL_L_X4Y138_SLICE_X5Y138_BQ;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X13Y144_SLICE_X18Y144_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y144_SLICE_X18Y144_D1 = 1'b1;
  assign CLBLM_R_X13Y144_SLICE_X18Y144_D2 = 1'b1;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_C2 = CLBLM_R_X11Y134_SLICE_X14Y134_CQ;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_C3 = CLBLM_L_X10Y135_SLICE_X12Y135_DO6;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_C4 = CLBLM_R_X13Y134_SLICE_X19Y134_AQ;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_C5 = CLBLM_L_X10Y138_SLICE_X13Y138_AQ;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y144_SLICE_X18Y144_D3 = 1'b1;
  assign CLBLM_R_X13Y141_SLICE_X18Y141_B6 = 1'b1;
  assign CLBLM_R_X13Y144_SLICE_X18Y144_D4 = 1'b1;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y144_SLICE_X18Y144_D6 = 1'b1;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_D1 = CLBLM_R_X11Y136_SLICE_X15Y136_AQ;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_D2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_D3 = 1'b1;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_D4 = CLBLM_L_X10Y131_SLICE_X12Y131_BQ;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_D5 = 1'b1;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_D6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_A1 = CLBLM_R_X7Y135_SLICE_X8Y135_BQ;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_A2 = CLBLL_L_X4Y134_SLICE_X4Y134_BQ;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_A4 = CLBLL_L_X4Y139_SLICE_X4Y139_BO6;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_A5 = 1'b1;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_A6 = 1'b1;
  assign LIOI3_X0Y77_ILOGIC_X0Y78_D = LIOB33_X0Y77_IOB_X0Y78_I;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_B1 = CLBLM_R_X5Y139_SLICE_X7Y139_AQ;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_B2 = CLBLL_L_X4Y137_SLICE_X4Y137_BQ;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_B3 = CLBLM_R_X7Y135_SLICE_X8Y135_DO5;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_B4 = 1'b1;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_B5 = CLBLL_L_X4Y136_SLICE_X5Y136_DO5;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOI3_X0Y103_OLOGIC_X0Y103_D1 = CLBLL_L_X2Y133_SLICE_X0Y133_AO5;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_C1 = CLBLL_L_X4Y136_SLICE_X4Y136_D5Q;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_C2 = 1'b1;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_C3 = 1'b1;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_C4 = CLBLM_L_X12Y135_SLICE_X17Y135_AQ;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_C6 = CLBLL_L_X4Y138_SLICE_X5Y138_AQ;
  assign LIOB33_X0Y115_IOB_X0Y116_O = CLBLM_L_X8Y135_SLICE_X11Y135_BQ;
  assign LIOB33_X0Y115_IOB_X0Y115_O = CLBLM_L_X12Y133_SLICE_X16Y133_CQ;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y77_ILOGIC_X0Y77_D = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_D1 = CLBLM_R_X5Y140_SLICE_X6Y140_AO6;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_D2 = CLBLM_L_X10Y134_SLICE_X12Y134_CQ;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_D3 = CLBLL_L_X4Y136_SLICE_X4Y136_AQ;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_D4 = CLBLL_L_X4Y142_SLICE_X4Y142_BO6;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_D6 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_A1 = CLBLM_R_X11Y142_SLICE_X15Y142_CQ;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_A1 = CLBLM_L_X8Y137_SLICE_X10Y137_CO6;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_A3 = CLBLM_L_X8Y138_SLICE_X10Y138_AQ;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_A4 = CLBLM_R_X3Y136_SLICE_X3Y136_BQ;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_A5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_A6 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_A2 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_A3 = CLBLL_L_X4Y134_SLICE_X5Y134_AQ;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_B1 = 1'b1;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_B1 = 1'b1;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_B2 = CLBLL_L_X4Y137_SLICE_X5Y137_BQ;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_B3 = CLBLM_R_X3Y136_SLICE_X2Y136_AQ;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_B4 = 1'b1;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_B5 = CLBLM_R_X7Y138_SLICE_X9Y138_AQ;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_A1 = CLBLM_R_X7Y132_SLICE_X9Y132_DQ;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_C2 = CLBLL_L_X4Y144_SLICE_X4Y144_AO6;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_C3 = CLBLM_L_X8Y136_SLICE_X10Y136_AQ;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_C4 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_C5 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_C6 = CLBLL_L_X4Y136_SLICE_X5Y136_BQ;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_A3 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_A4 = CLBLM_R_X5Y133_SLICE_X7Y133_DO6;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_A5 = CLBLM_L_X8Y132_SLICE_X11Y132_AQ;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_A6 = CLBLM_L_X8Y131_SLICE_X11Y131_AQ;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_B5 = CLBLM_R_X11Y132_SLICE_X15Y132_CO6;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_B2 = CLBLM_L_X8Y131_SLICE_X11Y131_BQ;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_D1 = CLBLM_R_X5Y140_SLICE_X6Y140_AO6;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_D2 = CLBLL_L_X4Y138_SLICE_X5Y138_B5Q;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_B3 = 1'b1;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_D4 = CLBLM_L_X10Y134_SLICE_X12Y134_CQ;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_B4 = CLBLM_R_X7Y134_SLICE_X8Y134_BQ;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_D6 = CLBLL_L_X4Y134_SLICE_X4Y134_AQ;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_C3 = CLBLM_L_X8Y131_SLICE_X10Y131_AQ;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_C4 = CLBLM_L_X8Y133_SLICE_X10Y133_CQ;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_C1 = CLBLM_L_X8Y132_SLICE_X11Y132_AQ;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_C2 = CLBLM_L_X8Y132_SLICE_X10Y132_AQ;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_C5 = CLBLM_L_X8Y131_SLICE_X11Y131_AQ;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_C6 = CLBLM_L_X10Y131_SLICE_X13Y131_AQ;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_SR = CLBLM_R_X7Y144_SLICE_X9Y144_BO6;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_A1 = CLBLM_L_X10Y141_SLICE_X12Y141_DO6;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_D1 = CLBLM_L_X8Y132_SLICE_X10Y132_AQ;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_D2 = CLBLM_L_X8Y131_SLICE_X10Y131_CO6;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_D3 = CLBLM_L_X10Y137_SLICE_X12Y137_B5Q;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_D4 = CLBLM_L_X8Y133_SLICE_X10Y133_CQ;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_D5 = CLBLM_R_X11Y146_SLICE_X14Y146_AQ;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_D6 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_A6 = CLBLM_L_X10Y140_SLICE_X12Y140_DO6;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_B2 = CLBLM_R_X11Y141_SLICE_X14Y141_AQ;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_B4 = CLBLM_R_X7Y135_SLICE_X9Y135_AQ;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_A1 = CLBLM_R_X5Y133_SLICE_X7Y133_DO6;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_A2 = CLBLM_L_X10Y137_SLICE_X12Y137_BQ;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_A3 = CLBLM_L_X8Y131_SLICE_X10Y131_AQ;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_A5 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_A6 = CLBLL_L_X4Y132_SLICE_X5Y132_AQ;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_C2 = CLBLM_R_X11Y135_SLICE_X14Y135_AQ;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_AX = CLBLM_L_X8Y131_SLICE_X10Y131_BO6;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_C3 = CLBLM_L_X10Y145_SLICE_X13Y145_CO6;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_B1 = CLBLM_L_X8Y131_SLICE_X11Y131_BQ;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_B3 = CLBLM_R_X5Y132_SLICE_X7Y132_DO6;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_B4 = CLBLM_L_X8Y135_SLICE_X11Y135_BQ;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_B5 = CLBLM_L_X8Y131_SLICE_X10Y131_A5Q;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_B6 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_D1 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_D2 = CLBLM_L_X12Y144_SLICE_X17Y144_AQ;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_C1 = CLBLM_L_X10Y131_SLICE_X13Y131_AQ;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_C2 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_C3 = CLBLM_L_X10Y137_SLICE_X12Y137_BQ;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_C4 = CLBLM_L_X8Y135_SLICE_X11Y135_AQ;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_C5 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_C6 = CLBLL_L_X4Y132_SLICE_X5Y132_AQ;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_D3 = CLBLM_R_X11Y141_SLICE_X15Y141_AQ;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_D4 = CLBLM_R_X11Y139_SLICE_X15Y139_DQ;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_D5 = CLBLM_L_X10Y141_SLICE_X12Y141_BO5;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_D6 = CLBLM_L_X8Y140_SLICE_X11Y140_CO5;
  assign CLBLM_R_X103Y170_SLICE_X163Y170_A1 = CLBLM_R_X11Y144_SLICE_X15Y144_AQ;
  assign CLBLM_R_X103Y170_SLICE_X163Y170_A2 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X163Y170_A4 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_D1 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_D2 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_D3 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_D4 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_D5 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_D6 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X163Y170_B1 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X163Y170_B2 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X163Y170_B3 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X163Y170_B5 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X163Y170_B6 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X163Y170_C1 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X163Y170_C2 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X163Y170_C3 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X163Y170_C4 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X163Y170_C5 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X163Y170_C6 = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_T1 = 1'b1;
  assign RIOI3_X105Y183_OLOGIC_X1Y184_D1 = CLBLM_L_X12Y139_SLICE_X17Y139_DO6;
  assign CLBLM_R_X103Y170_SLICE_X163Y170_D1 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X163Y170_D2 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X163Y170_D3 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X163Y170_D4 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X163Y170_D5 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X163Y170_D6 = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_D1 = CLBLM_R_X3Y137_SLICE_X2Y137_AQ;
  assign RIOI3_X105Y183_OLOGIC_X1Y184_T1 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X162Y170_A1 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X162Y170_A2 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X162Y170_A3 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X162Y170_A4 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X162Y170_A5 = 1'b1;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_A1 = CLBLM_R_X11Y136_SLICE_X14Y136_DQ;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_A3 = CLBLM_R_X11Y135_SLICE_X15Y135_AQ;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_A4 = CLBLM_L_X8Y135_SLICE_X11Y135_CQ;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_A5 = CLBLM_R_X13Y137_SLICE_X19Y137_AQ;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_A6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X103Y170_SLICE_X162Y170_A6 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X162Y170_B1 = 1'b1;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_B2 = CLBLM_L_X8Y133_SLICE_X11Y133_BQ;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_B3 = 1'b1;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_B4 = CLBLM_L_X10Y136_SLICE_X12Y136_BQ;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_B6 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X162Y170_B2 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X162Y170_B3 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X162Y170_B5 = 1'b1;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_C1 = CLBLL_L_X4Y139_SLICE_X4Y139_BO6;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_C2 = CLBLM_L_X10Y134_SLICE_X12Y134_CQ;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_C3 = CLBLM_L_X12Y135_SLICE_X17Y135_A5Q;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_C5 = CLBLL_L_X4Y134_SLICE_X4Y134_AQ;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_C6 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X162Y170_C1 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X162Y170_C2 = 1'b1;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X103Y170_SLICE_X162Y170_C4 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X162Y170_C5 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X162Y170_C6 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X162Y170_D1 = 1'b1;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_D1 = CLBLM_R_X5Y132_SLICE_X7Y132_DO6;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_D2 = CLBLM_R_X11Y131_SLICE_X15Y131_AO5;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_D3 = CLBLM_L_X10Y139_SLICE_X13Y139_CQ;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_D4 = CLBLM_R_X11Y131_SLICE_X15Y131_BQ;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_D5 = CLBLM_R_X11Y133_SLICE_X15Y133_AQ;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_D6 = CLBLM_R_X13Y137_SLICE_X18Y137_A5Q;
  assign CLBLM_R_X103Y170_SLICE_X162Y170_D2 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X162Y170_D3 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X162Y170_D4 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X162Y170_D5 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X162Y170_D6 = 1'b1;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_A1 = CLBLM_R_X11Y135_SLICE_X14Y135_CQ;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_A2 = CLBLM_R_X11Y138_SLICE_X14Y138_D5Q;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_A3 = CLBLM_R_X11Y135_SLICE_X14Y135_AQ;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_A5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_A6 = CLBLM_L_X8Y138_SLICE_X10Y138_AQ;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_T1 = 1'b1;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_B1 = CLBLM_R_X11Y135_SLICE_X14Y135_CQ;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_B2 = CLBLM_R_X11Y135_SLICE_X14Y135_BQ;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_B3 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_B4 = CLBLM_L_X8Y138_SLICE_X10Y138_AQ;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_B5 = CLBLM_L_X10Y144_SLICE_X12Y144_AQ;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_C1 = CLBLM_R_X11Y132_SLICE_X14Y132_BQ;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_C2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_C3 = CLBLM_L_X8Y136_SLICE_X11Y136_AQ;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_C5 = CLBLM_R_X11Y135_SLICE_X14Y135_CQ;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_C6 = CLBLM_L_X8Y138_SLICE_X10Y138_AQ;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_D1 = CLBLM_R_X11Y133_SLICE_X14Y133_AQ;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_D2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_D3 = CLBLM_R_X11Y135_SLICE_X14Y135_DQ;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_D4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_D5 = CLBLM_L_X10Y135_SLICE_X13Y135_CO6;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_D6 = CLBLM_L_X8Y138_SLICE_X10Y138_AQ;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y114_D = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_A1 = 1'b1;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_A3 = CLBLL_L_X4Y138_SLICE_X4Y138_AQ;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_A4 = 1'b1;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_A5 = CLBLL_L_X4Y139_SLICE_X4Y139_AQ;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_A6 = CLBLM_L_X8Y136_SLICE_X11Y136_CQ;
  assign LIOB33_X0Y117_IOB_X0Y117_O = CLBLM_R_X5Y136_SLICE_X6Y136_D5Q;
  assign LIOB33_X0Y117_IOB_X0Y118_O = CLBLL_L_X4Y135_SLICE_X5Y135_DQ;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_B2 = CLBLL_L_X4Y138_SLICE_X4Y138_BQ;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_B3 = CLBLL_L_X4Y138_SLICE_X5Y138_B5Q;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_B4 = 1'b1;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_B5 = 1'b1;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_B6 = CLBLM_R_X5Y139_SLICE_X7Y139_BQ;
  assign LIOI3_X0Y165_OLOGIC_X0Y166_D1 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_C1 = CLBLL_L_X4Y144_SLICE_X4Y144_AO6;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_C2 = CLBLL_L_X4Y139_SLICE_X4Y139_AQ;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_C3 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_C4 = CLBLM_R_X7Y136_SLICE_X8Y136_BQ;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_C5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_C6 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_D = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_D1 = CLBLL_L_X4Y136_SLICE_X5Y136_AQ;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_D2 = 1'b1;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_D3 = CLBLM_L_X10Y138_SLICE_X13Y138_BQ;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_D4 = CLBLL_L_X4Y143_SLICE_X5Y143_AO5;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_D5 = 1'b1;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_D6 = CLBLM_R_X7Y142_SLICE_X9Y142_CO6;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_SR = CLBLM_R_X7Y144_SLICE_X9Y144_BO6;
  assign LIOB33_SING_X0Y199_IOB_X0Y199_O = LIOB33_X0Y73_IOB_X0Y74_I;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_A1 = CLBLM_R_X5Y137_SLICE_X6Y137_DO6;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_A3 = CLBLM_R_X5Y142_SLICE_X6Y142_CO6;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_A4 = CLBLL_L_X4Y138_SLICE_X4Y138_BQ;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_A5 = CLBLM_R_X7Y141_SLICE_X8Y141_AQ;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_A6 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_A2 = CLBLM_L_X10Y142_SLICE_X13Y142_BQ;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_A3 = CLBLM_L_X10Y142_SLICE_X13Y142_AQ;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_B1 = 1'b1;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_B2 = CLBLM_R_X5Y139_SLICE_X7Y139_BQ;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_B3 = CLBLL_L_X4Y136_SLICE_X5Y136_AQ;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_B6 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_A4 = CLBLM_L_X8Y144_SLICE_X11Y144_CO6;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_A5 = CLBLM_L_X10Y135_SLICE_X12Y135_AQ;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_BX = CLBLL_L_X4Y138_SLICE_X5Y138_CO6;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_C1 = CLBLL_L_X4Y135_SLICE_X5Y135_BQ;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_C2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_C3 = CLBLM_L_X8Y138_SLICE_X10Y138_AQ;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_C4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_C5 = CLBLL_L_X4Y137_SLICE_X5Y137_DO6;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_C6 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_A1 = CLBLM_L_X8Y132_SLICE_X11Y132_CQ;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_A2 = CLBLM_R_X5Y133_SLICE_X7Y133_DO6;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_A3 = CLBLM_L_X8Y132_SLICE_X11Y132_AQ;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_A5 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_A6 = CLBLM_L_X8Y133_SLICE_X10Y133_BQ;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_D1 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_D2 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_D3 = CLBLL_L_X4Y141_SLICE_X4Y141_DO6;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_D1 = CLBLM_L_X10Y142_SLICE_X13Y142_BQ;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_D4 = CLBLL_L_X4Y138_SLICE_X5Y138_AQ;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_D5 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_D6 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_D5 = CLBLM_L_X10Y145_SLICE_X12Y145_CO6;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_D6 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_B4 = CLBLM_L_X10Y133_SLICE_X12Y133_AQ;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_B6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_C1 = CLBLM_L_X8Y138_SLICE_X10Y138_AQ;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_C2 = CLBLM_L_X8Y132_SLICE_X11Y132_CQ;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_C3 = CLBLM_L_X8Y133_SLICE_X11Y133_CQ;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_C4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_C5 = CLBLL_L_X4Y136_SLICE_X4Y136_DQ;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_A1 = CLBLM_L_X10Y145_SLICE_X13Y145_BO6;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_A2 = CLBLM_L_X8Y144_SLICE_X11Y144_CO6;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_D1 = CLBLL_L_X4Y132_SLICE_X5Y132_AQ;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_D2 = CLBLM_L_X8Y131_SLICE_X11Y131_CO6;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_D3 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_D4 = CLBLM_L_X8Y133_SLICE_X10Y133_BQ;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_D5 = CLBLM_R_X11Y132_SLICE_X15Y132_DO6;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_D6 = CLBLM_L_X10Y133_SLICE_X12Y133_AQ;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_A6 = CLBLL_L_X4Y136_SLICE_X5Y136_CQ;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_B1 = CLBLM_L_X10Y145_SLICE_X13Y145_BO6;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_B2 = CLBLM_L_X10Y142_SLICE_X12Y142_BQ;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_A1 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_A3 = CLBLM_L_X8Y132_SLICE_X10Y132_AQ;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_A4 = CLBLM_L_X8Y140_SLICE_X10Y140_BQ;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_A5 = CLBLM_R_X5Y134_SLICE_X7Y134_DO6;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_A6 = CLBLM_L_X10Y132_SLICE_X12Y132_BO6;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_C2 = CLBLM_L_X10Y142_SLICE_X12Y142_CQ;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_C3 = CLBLM_L_X10Y145_SLICE_X13Y145_BO6;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_B1 = CLBLM_L_X10Y137_SLICE_X12Y137_AQ;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_B2 = CLBLM_L_X8Y132_SLICE_X10Y132_BQ;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_B3 = CLBLM_L_X12Y132_SLICE_X17Y132_AQ;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_B4 = CLBLM_L_X8Y138_SLICE_X10Y138_AQ;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_B6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_D2 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_C1 = CLBLM_L_X8Y132_SLICE_X10Y132_DO6;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_C2 = CLBLM_R_X5Y133_SLICE_X7Y133_AO6;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_C3 = CLBLM_R_X7Y133_SLICE_X9Y133_DO6;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_C4 = CLBLM_R_X5Y136_SLICE_X7Y136_DO6;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_C5 = CLBLM_R_X5Y133_SLICE_X7Y133_CO6;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_C6 = CLBLM_R_X7Y134_SLICE_X8Y134_C5Q;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_D3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_D4 = CLBLM_R_X7Y135_SLICE_X8Y135_CQ;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_D5 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_D6 = CLBLM_L_X10Y142_SLICE_X13Y142_BQ;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_D1 = CLBLM_R_X11Y133_SLICE_X15Y133_BQ;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_D2 = CLBLM_L_X10Y130_SLICE_X12Y130_AQ;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_D3 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_D4 = CLBLM_L_X10Y131_SLICE_X12Y131_BQ;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_D5 = CLBLL_L_X4Y135_SLICE_X5Y135_CQ;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_D6 = CLBLM_R_X11Y131_SLICE_X15Y131_BQ;
  assign LIOI3_X0Y165_OLOGIC_X0Y165_T1 = 1'b1;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_C1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_A1 = CLBLM_R_X13Y136_SLICE_X18Y136_CQ;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_A3 = CLBLM_L_X10Y139_SLICE_X13Y139_CQ;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_A5 = CLBLM_R_X5Y140_SLICE_X7Y140_BQ;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_A6 = 1'b1;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_B1 = CLBLM_L_X8Y132_SLICE_X10Y132_AQ;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_B2 = CLBLM_R_X11Y136_SLICE_X15Y136_A5Q;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_B4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_B5 = CLBLM_L_X10Y141_SLICE_X13Y141_AQ;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_B6 = 1'b1;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_C1 = CLBLL_L_X4Y134_SLICE_X4Y134_AQ;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_C2 = CLBLM_R_X11Y137_SLICE_X14Y137_CO5;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_C3 = CLBLM_R_X5Y141_SLICE_X7Y141_DO6;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_C4 = CLBLM_L_X10Y134_SLICE_X12Y134_CQ;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_C5 = CLBLM_L_X12Y135_SLICE_X17Y135_BO5;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_C6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_D1 = CLBLM_L_X8Y136_SLICE_X10Y136_CQ;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_D2 = CLBLM_L_X8Y135_SLICE_X11Y135_A5Q;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_D3 = 1'b1;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_D4 = CLBLM_R_X13Y136_SLICE_X18Y136_CQ;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_D5 = 1'b1;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_D6 = CLBLM_R_X11Y135_SLICE_X15Y135_BQ;
  assign RIOI3_X105Y167_OLOGIC_X1Y168_D1 = CLBLM_R_X11Y153_SLICE_X14Y153_AO6;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_A1 = CLBLM_R_X7Y139_SLICE_X9Y139_BO6;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_A3 = CLBLM_R_X11Y136_SLICE_X14Y136_AQ;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_A4 = CLBLM_R_X13Y136_SLICE_X18Y136_AQ;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_A5 = CLBLM_R_X11Y135_SLICE_X14Y135_AQ;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_A6 = 1'b1;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_B1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_B2 = CLBLM_R_X11Y136_SLICE_X14Y136_BQ;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_B4 = CLBLM_R_X11Y138_SLICE_X14Y138_D5Q;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_B5 = CLBLM_L_X8Y138_SLICE_X10Y138_AQ;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_B6 = 1'b1;
  assign CLBLM_R_X13Y144_SLICE_X19Y144_C4 = 1'b1;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_D3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign LIOB33_X0Y119_IOB_X0Y119_O = CLBLM_L_X10Y135_SLICE_X13Y135_BQ;
  assign CLBLM_R_X13Y144_SLICE_X19Y144_C5 = 1'b1;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_C2 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_C3 = CLBLM_L_X10Y141_SLICE_X13Y141_BQ;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_C4 = CLBLM_R_X11Y133_SLICE_X15Y133_DQ;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_C5 = CLBLM_L_X12Y136_SLICE_X17Y136_CQ;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_C6 = 1'b1;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_D5 = 1'b1;
  assign CLBLM_R_X13Y144_SLICE_X19Y144_C6 = 1'b1;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOB33_X105Y197_IOB_X1Y197_O = CLBLM_R_X103Y175_SLICE_X163Y175_AO6;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_D2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_D3 = CLBLM_R_X13Y137_SLICE_X18Y137_AQ;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_D4 = CLBLM_R_X11Y136_SLICE_X14Y136_BQ;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_A1 = CLBLL_L_X4Y138_SLICE_X5Y138_CO5;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_A2 = CLBLM_R_X5Y140_SLICE_X6Y140_AO6;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_A3 = CLBLL_L_X4Y139_SLICE_X4Y139_AQ;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_A6 = CLBLM_L_X10Y142_SLICE_X12Y142_CQ;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_D5 = CLBLM_R_X11Y135_SLICE_X15Y135_AQ;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_D6 = CLBLM_L_X10Y136_SLICE_X13Y136_AO6;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_B1 = CLBLL_L_X4Y138_SLICE_X4Y138_DO6;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_B2 = CLBLM_R_X5Y139_SLICE_X7Y139_DO6;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_B3 = CLBLM_R_X5Y140_SLICE_X6Y140_CO6;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_B4 = CLBLM_R_X3Y142_SLICE_X2Y142_CO6;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_B5 = CLBLM_R_X5Y140_SLICE_X6Y140_BO6;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_B6 = CLBLL_L_X4Y139_SLICE_X4Y139_CO6;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_C1 = CLBLM_L_X8Y137_SLICE_X11Y137_AQ;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_C2 = CLBLL_L_X4Y139_SLICE_X5Y139_CO6;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_C3 = 1'b1;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_C4 = CLBLL_L_X4Y143_SLICE_X5Y143_AO6;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_C5 = CLBLM_R_X3Y142_SLICE_X2Y142_AO6;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_C6 = CLBLL_L_X4Y139_SLICE_X5Y139_BQ;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_D1 = CLBLL_L_X4Y135_SLICE_X4Y135_CQ;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_D2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_D3 = CLBLM_R_X3Y143_SLICE_X2Y143_AO5;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_D4 = CLBLL_L_X2Y141_SLICE_X1Y141_AO5;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_D5 = 1'b1;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_D6 = CLBLM_R_X7Y136_SLICE_X8Y136_CQ;
  assign CLBLM_R_X13Y144_SLICE_X19Y144_D2 = 1'b1;
  assign CLBLM_R_X13Y144_SLICE_X19Y144_D5 = 1'b1;
  assign CLBLM_R_X13Y144_SLICE_X19Y144_D6 = 1'b1;
  assign RIOI3_X105Y141_ILOGIC_X1Y142_D = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_A2 = CLBLL_L_X4Y139_SLICE_X5Y139_BQ;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_A3 = CLBLL_L_X4Y139_SLICE_X5Y139_AQ;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_A4 = CLBLM_L_X8Y143_SLICE_X10Y143_DO5;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_A5 = 1'b1;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_A6 = CLBLM_R_X7Y134_SLICE_X9Y134_AQ;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_A1 = CLBLM_R_X11Y144_SLICE_X14Y144_AQ;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_B1 = CLBLM_L_X10Y139_SLICE_X13Y139_B5Q;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_B2 = CLBLL_L_X4Y139_SLICE_X5Y139_BQ;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_A5 = CLBLM_L_X10Y142_SLICE_X12Y142_CQ;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_A6 = CLBLM_L_X10Y143_SLICE_X12Y143_AQ;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_B4 = CLBLM_R_X11Y138_SLICE_X14Y138_BQ;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_B5 = CLBLM_R_X7Y139_SLICE_X8Y139_AQ;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_B6 = CLBLM_L_X12Y134_SLICE_X17Y134_AO6;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_A2 = CLBLM_R_X11Y144_SLICE_X15Y144_BQ;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_A3 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_B2 = CLBLM_R_X11Y142_SLICE_X15Y142_CQ;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_B3 = CLBLM_L_X10Y142_SLICE_X12Y142_BQ;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_B4 = CLBLM_L_X10Y145_SLICE_X12Y145_CO6;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_B5 = CLBLM_R_X11Y143_SLICE_X14Y143_CO5;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_B6 = CLBLM_L_X10Y144_SLICE_X13Y144_DO6;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_C1 = CLBLM_R_X7Y135_SLICE_X9Y135_AQ;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_BX = CLBLM_R_X7Y135_SLICE_X8Y135_CQ;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_C2 = CLBLL_L_X4Y138_SLICE_X5Y138_A5Q;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_C1 = CLBLM_L_X10Y142_SLICE_X13Y142_AQ;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_C2 = CLBLM_R_X11Y142_SLICE_X15Y142_CQ;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_C3 = CLBLM_L_X10Y145_SLICE_X12Y145_CO6;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_C4 = CLBLM_L_X10Y144_SLICE_X13Y144_DO6;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_C5 = CLBLM_L_X10Y143_SLICE_X13Y143_DO6;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_C6 = CLBLM_R_X11Y143_SLICE_X14Y143_CO5;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_CE = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_A2 = CLBLM_L_X8Y138_SLICE_X10Y138_AQ;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_A3 = CLBLM_L_X8Y133_SLICE_X11Y133_AQ;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_A4 = CLBLM_L_X10Y131_SLICE_X13Y131_BQ;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_D1 = CLBLM_R_X5Y138_SLICE_X7Y138_BQ;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_D1 = CLBLM_L_X10Y143_SLICE_X13Y143_AO6;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_D2 = CLBLM_L_X10Y142_SLICE_X13Y142_CQ;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_D3 = 1'b1;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_D4 = 1'b1;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_D5 = 1'b1;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_D6 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_B4 = CLBLM_R_X13Y137_SLICE_X18Y137_AQ;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_SR = CLBLM_L_X12Y144_SLICE_X16Y144_AO6;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_C1 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_C2 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_C3 = CLBLM_R_X7Y142_SLICE_X9Y142_BQ;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_C4 = CLBLM_L_X10Y131_SLICE_X12Y131_DO6;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_C6 = CLBLM_R_X7Y131_SLICE_X9Y131_AQ;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_A1 = CLBLM_L_X10Y143_SLICE_X12Y143_DO6;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_A2 = 1'b1;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_A3 = CLBLM_L_X10Y144_SLICE_X12Y144_AO6;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_A4 = CLBLM_R_X11Y144_SLICE_X14Y144_DO6;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_A5 = CLBLM_R_X5Y134_SLICE_X6Y134_AQ;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_D1 = CLBLM_R_X5Y132_SLICE_X7Y132_DO6;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_D2 = CLBLM_R_X11Y131_SLICE_X15Y131_BQ;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_D3 = CLBLM_L_X10Y133_SLICE_X12Y133_DO6;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_D4 = CLBLM_L_X10Y141_SLICE_X12Y141_CQ;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_B6 = CLBLM_L_X10Y145_SLICE_X13Y145_BO6;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_D5 = CLBLM_L_X8Y134_SLICE_X11Y134_DQ;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_D6 = CLBLM_L_X8Y137_SLICE_X11Y137_BQ;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_B1 = CLBLL_L_X4Y137_SLICE_X4Y137_BQ;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_B2 = CLBLM_L_X10Y143_SLICE_X12Y143_BQ;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_B3 = CLBLM_L_X10Y145_SLICE_X13Y145_AQ;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_B4 = CLBLM_L_X8Y144_SLICE_X11Y144_CO6;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_A1 = CLBLM_L_X8Y133_SLICE_X10Y133_DO6;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_C5 = CLBLM_R_X11Y144_SLICE_X14Y144_DO6;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_C6 = CLBLM_L_X10Y145_SLICE_X12Y145_AQ;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_A3 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_A4 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_A5 = CLBLM_R_X7Y131_SLICE_X9Y131_AQ;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_A6 = CLBLM_L_X10Y139_SLICE_X13Y139_B5Q;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_B1 = CLBLM_R_X5Y137_SLICE_X7Y137_B5Q;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_B2 = CLBLM_L_X8Y133_SLICE_X10Y133_BQ;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_B3 = CLBLM_L_X8Y131_SLICE_X10Y131_AQ;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_B5 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_B6 = CLBLM_R_X5Y133_SLICE_X7Y133_DO6;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_D1 = CLBLM_L_X10Y143_SLICE_X12Y143_BQ;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_D2 = CLBLM_L_X10Y143_SLICE_X12Y143_AQ;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_C1 = CLBLM_R_X5Y134_SLICE_X7Y134_DO6;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_C2 = CLBLM_L_X8Y133_SLICE_X10Y133_CQ;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_C4 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_C5 = CLBLM_L_X8Y132_SLICE_X10Y132_AQ;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_C6 = CLBLM_L_X8Y133_SLICE_X10Y133_AQ;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_D5 = CLBLM_L_X10Y145_SLICE_X12Y145_CO6;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y144_SLICE_X18Y144_B5 = CLBLM_L_X12Y142_SLICE_X16Y142_BQ;
  assign CLBLM_R_X13Y144_SLICE_X18Y144_B6 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_D1 = CLBLM_R_X5Y132_SLICE_X7Y132_DO6;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_D2 = CLBLM_L_X8Y133_SLICE_X10Y133_AQ;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_D3 = CLBLM_R_X7Y134_SLICE_X8Y134_C5Q;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_D4 = CLBLM_R_X5Y133_SLICE_X7Y133_DO6;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_D5 = CLBLM_L_X8Y132_SLICE_X10Y132_DO6;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_D6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y143_D = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_D1 = 1'b1;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_D2 = 1'b1;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_D3 = 1'b1;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_D4 = 1'b1;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_A1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_A2 = CLBLM_L_X10Y137_SLICE_X12Y137_CQ;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_A3 = CLBLM_R_X11Y137_SLICE_X15Y137_AQ;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_A4 = CLBLM_R_X11Y137_SLICE_X14Y137_DO6;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_A6 = CLBLM_L_X8Y138_SLICE_X10Y138_AQ;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_D5 = 1'b1;
  assign CLBLM_R_X13Y144_SLICE_X18Y144_C4 = CLBLM_R_X13Y140_SLICE_X19Y140_AQ;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_D6 = 1'b1;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_B1 = CLBLM_R_X11Y136_SLICE_X15Y136_DO6;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_B2 = CLBLM_R_X11Y138_SLICE_X15Y138_AQ;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_B3 = CLBLM_R_X5Y137_SLICE_X7Y137_CQ;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_B4 = CLBLM_R_X11Y137_SLICE_X15Y137_DO6;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_B5 = CLBLM_R_X11Y136_SLICE_X15Y136_AQ;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_B6 = CLBLM_R_X11Y137_SLICE_X15Y137_CO6;
  assign CLBLM_R_X13Y144_SLICE_X18Y144_C6 = CLBLM_R_X13Y137_SLICE_X18Y137_CO5;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_C1 = 1'b1;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_C2 = CLBLM_L_X10Y135_SLICE_X12Y135_BQ;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_C3 = 1'b1;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_C4 = CLBLM_R_X5Y140_SLICE_X7Y140_BQ;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_C5 = CLBLM_L_X12Y136_SLICE_X16Y136_AQ;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_C6 = CLBLM_R_X7Y139_SLICE_X8Y139_BQ;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOB33_X0Y121_IOB_X0Y121_O = CLBLM_L_X8Y135_SLICE_X11Y135_B5Q;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_D1 = CLBLM_R_X11Y136_SLICE_X15Y136_A5Q;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_D2 = CLBLM_L_X12Y139_SLICE_X16Y139_CQ;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_D3 = CLBLM_R_X11Y138_SLICE_X15Y138_CQ;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_D4 = CLBLM_L_X8Y139_SLICE_X11Y139_BQ;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_D5 = 1'b1;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_D6 = 1'b1;
  assign LIOB33_X0Y121_IOB_X0Y122_O = CLBLL_L_X4Y133_SLICE_X5Y133_A5Q;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_A1 = CLBLM_L_X12Y137_SLICE_X16Y137_A5Q;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_A4 = 1'b1;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_A5 = CLBLM_R_X11Y137_SLICE_X14Y137_CO5;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_A6 = CLBLM_R_X7Y134_SLICE_X8Y134_AQ;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_B1 = CLBLM_R_X11Y133_SLICE_X15Y133_AQ;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_B3 = CLBLM_R_X7Y136_SLICE_X9Y136_AQ;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_B4 = CLBLM_L_X8Y135_SLICE_X11Y135_A5Q;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_B5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_B6 = 1'b1;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_C1 = CLBLM_R_X11Y138_SLICE_X14Y138_AQ;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_C2 = CLBLM_R_X7Y139_SLICE_X8Y139_A5Q;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_C3 = CLBLM_L_X10Y138_SLICE_X13Y138_AQ;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_C4 = CLBLM_L_X10Y141_SLICE_X13Y141_BQ;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_C5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_C6 = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_D1 = LIOB33_X0Y53_IOB_X0Y54_I;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_B3 = CLBLM_R_X5Y138_SLICE_X6Y138_BQ;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_A1 = CLBLL_L_X4Y139_SLICE_X4Y139_DO6;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_A2 = CLBLL_L_X4Y140_SLICE_X5Y140_DO6;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_A3 = LIOB33_X0Y65_IOB_X0Y66_I;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_A4 = CLBLL_L_X4Y140_SLICE_X4Y140_BO6;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_A5 = CLBLL_L_X4Y140_SLICE_X4Y140_CO6;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_A6 = CLBLM_R_X3Y141_SLICE_X2Y141_AO6;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_D1 = CLBLL_L_X4Y134_SLICE_X4Y134_AQ;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_D2 = CLBLM_L_X10Y134_SLICE_X12Y134_CQ;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_B1 = CLBLL_L_X4Y143_SLICE_X5Y143_BO5;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_B2 = CLBLM_R_X5Y139_SLICE_X6Y139_BQ;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_B3 = CLBLL_L_X2Y140_SLICE_X1Y140_AO6;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_B4 = CLBLL_L_X4Y135_SLICE_X4Y135_BQ;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_B5 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_B6 = CLBLM_R_X3Y141_SLICE_X3Y141_AO5;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_B6 = CLBLM_L_X10Y140_SLICE_X13Y140_AO5;
  assign LIOI3_X0Y79_OLOGIC_X0Y80_T1 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_C1 = CLBLL_L_X2Y140_SLICE_X1Y140_AO6;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_C2 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_C3 = CLBLM_R_X3Y143_SLICE_X2Y143_AO6;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_C4 = CLBLM_L_X8Y139_SLICE_X10Y139_DQ;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_C5 = CLBLM_L_X8Y140_SLICE_X10Y140_AQ;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_C6 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_T1 = 1'b1;
  assign RIOI3_X105Y185_OLOGIC_X1Y185_D1 = CLBLM_L_X12Y139_SLICE_X17Y139_DO5;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_D1 = CLBLL_L_X4Y143_SLICE_X5Y143_AO6;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_D2 = CLBLM_R_X5Y139_SLICE_X6Y139_BQ;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_D3 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_D4 = CLBLM_R_X3Y142_SLICE_X2Y142_AO5;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_D5 = CLBLL_L_X4Y139_SLICE_X4Y139_DO6;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_D6 = CLBLL_L_X4Y135_SLICE_X4Y135_BQ;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_C1 = CLBLM_R_X11Y140_SLICE_X15Y140_DQ;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_B4 = 1'b1;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_C2 = CLBLM_L_X10Y140_SLICE_X13Y140_CQ;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_B5 = 1'b1;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_B6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_D1 = LIOB33_X0Y59_IOB_X0Y60_I;
  assign RIOI3_X105Y185_OLOGIC_X1Y185_T1 = 1'b1;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_D1 = LIOB33_X0Y55_IOB_X0Y56_I;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_C6 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_A1 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_A2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_A3 = CLBLM_R_X3Y138_SLICE_X3Y138_AQ;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_A4 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_A5 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_A6 = CLBLM_R_X3Y143_SLICE_X2Y143_AO6;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_T1 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_B1 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_B2 = CLBLM_R_X5Y136_SLICE_X7Y136_CQ;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_B3 = CLBLL_L_X4Y143_SLICE_X5Y143_AO6;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_B4 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_B5 = CLBLM_R_X5Y143_SLICE_X6Y143_BO6;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_B6 = CLBLL_L_X4Y140_SLICE_X5Y140_CO6;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_A1 = CLBLM_L_X10Y144_SLICE_X13Y144_AQ;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_A3 = CLBLM_L_X10Y144_SLICE_X12Y144_AO6;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_C1 = CLBLL_L_X2Y140_SLICE_X1Y140_AO6;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_C2 = CLBLM_R_X5Y138_SLICE_X7Y138_AQ;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_C3 = CLBLM_R_X3Y143_SLICE_X3Y143_AO5;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_C4 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_C5 = CLBLM_R_X3Y143_SLICE_X2Y143_AO5;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_C6 = CLBLL_L_X4Y135_SLICE_X4Y135_AQ;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_A4 = CLBLM_L_X10Y144_SLICE_X13Y144_BO6;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_B4 = CLBLM_L_X10Y145_SLICE_X12Y145_CO6;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_B5 = CLBLM_R_X11Y144_SLICE_X15Y144_BQ;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_B6 = CLBLM_L_X10Y145_SLICE_X12Y145_BO6;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_B1 = CLBLM_L_X10Y144_SLICE_X13Y144_DO6;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_B2 = CLBLM_L_X10Y143_SLICE_X12Y143_AQ;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_C1 = CLBLM_R_X11Y144_SLICE_X15Y144_BQ;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_C2 = CLBLM_L_X10Y143_SLICE_X12Y143_AQ;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_C3 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_C4 = CLBLM_R_X11Y144_SLICE_X14Y144_AQ;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_C5 = CLBLM_L_X10Y144_SLICE_X13Y144_AQ;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_C6 = CLBLM_L_X10Y142_SLICE_X12Y142_CQ;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_A1 = CLBLM_L_X8Y134_SLICE_X11Y134_AQ;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_D1 = CLBLL_L_X4Y139_SLICE_X5Y139_AQ;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_D2 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_D3 = CLBLM_R_X3Y143_SLICE_X3Y143_AO5;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_D4 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_D5 = CLBLL_L_X4Y143_SLICE_X5Y143_BO5;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_D1 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_D2 = CLBLM_L_X8Y142_SLICE_X10Y142_D5Q;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_D3 = CLBLM_L_X10Y141_SLICE_X12Y141_C5Q;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_D5 = CLBLM_L_X8Y144_SLICE_X11Y144_BO5;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_D6 = CLBLM_L_X10Y142_SLICE_X12Y142_CQ;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_B3 = CLBLM_R_X5Y134_SLICE_X7Y134_DO6;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_B4 = CLBLM_R_X5Y136_SLICE_X6Y136_BQ;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_B6 = CLBLM_L_X8Y133_SLICE_X10Y133_CQ;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_C1 = CLBLM_L_X8Y138_SLICE_X10Y138_AQ;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_C2 = CLBLM_L_X8Y134_SLICE_X11Y134_CQ;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_C4 = CLBLM_R_X5Y137_SLICE_X6Y137_BQ;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_C5 = CLBLM_R_X11Y133_SLICE_X15Y133_DQ;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_C6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_A5 = CLBLM_R_X11Y144_SLICE_X14Y144_AQ;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_A1 = CLBLM_L_X8Y142_SLICE_X10Y142_D5Q;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_A2 = CLBLM_L_X10Y142_SLICE_X12Y142_CQ;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_D5 = CLBLM_L_X10Y134_SLICE_X13Y134_CO5;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_A3 = CLBLM_R_X11Y143_SLICE_X14Y143_DO6;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_A4 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_D1 = CLBLM_R_X7Y131_SLICE_X9Y131_AQ;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_D2 = CLBLM_L_X8Y133_SLICE_X11Y133_DO6;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_B4 = CLBLM_R_X7Y142_SLICE_X9Y142_AQ;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_B5 = CLBLM_R_X11Y143_SLICE_X14Y143_AQ;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_B6 = CLBLM_L_X10Y144_SLICE_X12Y144_AO5;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_D3 = CLBLM_L_X8Y140_SLICE_X11Y140_AQ;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_D4 = 1'b1;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_D5 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_D6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_B3 = CLBLM_L_X10Y141_SLICE_X12Y141_C5Q;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_A1 = CLBLM_R_X11Y135_SLICE_X15Y135_AQ;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_C3 = CLBLM_L_X8Y135_SLICE_X10Y135_CO6;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_C4 = CLBLM_L_X8Y142_SLICE_X10Y142_D5Q;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_C5 = CLBLM_R_X11Y144_SLICE_X14Y144_AQ;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_C6 = CLBLM_L_X10Y142_SLICE_X12Y142_CQ;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_A2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_A3 = CLBLM_L_X8Y134_SLICE_X10Y134_AQ;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_A4 = CLBLM_L_X8Y133_SLICE_X10Y133_AQ;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_A5 = CLBLM_L_X8Y138_SLICE_X10Y138_AQ;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_AX = CLBLM_L_X10Y134_SLICE_X13Y134_CO6;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_B1 = CLBLL_L_X4Y136_SLICE_X4Y136_CQ;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_B2 = CLBLM_R_X7Y133_SLICE_X8Y133_BQ;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_B3 = CLBLM_R_X11Y140_SLICE_X15Y140_CQ;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_D2 = 1'b1;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_B6 = 1'b1;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_D1 = 1'b1;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_D3 = 1'b1;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_C1 = CLBLM_L_X8Y137_SLICE_X11Y137_CO5;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_C2 = CLBLL_L_X4Y139_SLICE_X4Y139_BO6;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_C3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_C4 = CLBLM_R_X7Y134_SLICE_X9Y134_DO6;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_C5 = CLBLM_R_X11Y136_SLICE_X15Y136_BQ;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_C6 = CLBLM_L_X8Y135_SLICE_X10Y135_AQ;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_D5 = 1'b1;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_D6 = 1'b1;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_SR = CLBLM_R_X7Y144_SLICE_X9Y144_BO6;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_A4 = CLBLM_R_X13Y134_SLICE_X19Y134_BQ;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_D1 = CLBLM_R_X5Y132_SLICE_X7Y132_DO6;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_D2 = CLBLM_L_X10Y131_SLICE_X12Y131_BQ;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_D3 = CLBLM_L_X10Y130_SLICE_X12Y130_AQ;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_D4 = CLBLM_R_X11Y131_SLICE_X15Y131_BQ;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_D5 = CLBLL_L_X4Y135_SLICE_X5Y135_CQ;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_D6 = CLBLM_L_X8Y134_SLICE_X10Y134_BO6;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_B1 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_B2 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_B3 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_B5 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_B6 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_C1 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_C2 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_C3 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_C4 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_C5 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_C6 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_D1 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_D2 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_D3 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_B1 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_D4 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_D5 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_D6 = 1'b1;
  assign LIOI3_X0Y79_ILOGIC_X0Y79_D = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_A1 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_A2 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_A3 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_A4 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_A5 = 1'b1;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_A1 = 1'b1;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_A2 = CLBLM_R_X11Y138_SLICE_X15Y138_BQ;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_A3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_A4 = CLBLM_L_X10Y141_SLICE_X13Y141_BQ;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_A6 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_A6 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_B1 = 1'b1;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_B1 = CLBLM_R_X11Y138_SLICE_X15Y138_B5Q;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_B4 = CLBLM_R_X11Y138_SLICE_X15Y138_D5Q;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_B5 = CLBLM_L_X12Y138_SLICE_X16Y138_AQ;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_B6 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_B2 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_B3 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_B5 = 1'b1;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_C1 = CLBLM_R_X5Y137_SLICE_X7Y137_CQ;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_C2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_C3 = 1'b1;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_C4 = CLBLM_L_X12Y135_SLICE_X17Y135_A5Q;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_C5 = 1'b1;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_C6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_C1 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_C2 = 1'b1;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_C4 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_C5 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_C6 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_D1 = 1'b1;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_D1 = CLBLM_L_X8Y136_SLICE_X10Y136_DQ;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_D2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_D3 = CLBLM_R_X11Y142_SLICE_X15Y142_AQ;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_D4 = CLBLM_L_X10Y141_SLICE_X13Y141_A5Q;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_D5 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_D6 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_B3 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_D2 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_D3 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_D4 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_D5 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_D6 = 1'b1;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_A1 = CLBLM_L_X12Y139_SLICE_X17Y139_AQ;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_A3 = CLBLM_R_X11Y138_SLICE_X14Y138_AQ;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_A4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_A5 = CLBLM_L_X10Y138_SLICE_X12Y138_BO6;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_A6 = CLBLM_L_X8Y138_SLICE_X10Y138_AQ;
  assign RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_D = RIOB33_X105Y119_IOB_X1Y119_I;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_B1 = CLBLM_R_X7Y139_SLICE_X9Y139_BO6;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_B2 = CLBLM_R_X11Y138_SLICE_X14Y138_BQ;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_B3 = CLBLM_R_X11Y138_SLICE_X14Y138_AQ;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_B4 = CLBLM_R_X11Y135_SLICE_X14Y135_AQ;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_B5 = CLBLM_R_X11Y136_SLICE_X14Y136_AQ;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_B4 = 1'b1;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_C2 = 1'b1;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_C3 = CLBLM_R_X11Y136_SLICE_X14Y136_DQ;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_C5 = CLBLM_R_X11Y140_SLICE_X15Y140_DQ;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_C6 = CLBLM_L_X10Y135_SLICE_X13Y135_AO5;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_A1 = CLBLM_R_X3Y143_SLICE_X3Y143_AO6;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_A2 = CLBLL_L_X4Y143_SLICE_X5Y143_BO5;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_A3 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_A4 = CLBLM_R_X3Y143_SLICE_X3Y143_AO5;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_A5 = CLBLM_R_X7Y137_SLICE_X8Y137_AQ;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_A6 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_D1 = CLBLM_R_X5Y135_SLICE_X6Y135_BQ;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_D2 = CLBLM_L_X8Y138_SLICE_X10Y138_DQ;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_B1 = CLBLL_L_X4Y143_SLICE_X4Y143_DO6;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_B2 = LIOB33_X0Y67_IOB_X0Y67_I;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_B3 = CLBLL_L_X4Y143_SLICE_X5Y143_AO6;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_B4 = CLBLM_R_X3Y141_SLICE_X2Y141_AO6;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_B5 = CLBLL_L_X4Y141_SLICE_X4Y141_AO6;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_B6 = CLBLM_L_X8Y139_SLICE_X10Y139_CQ;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_D3 = CLBLM_R_X11Y138_SLICE_X14Y138_DQ;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_D4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_D5 = RIOB33_X105Y119_IOB_X1Y119_I;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_C1 = LIOB33_X0Y65_IOB_X0Y66_I;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_C2 = CLBLM_R_X3Y139_SLICE_X2Y139_AO5;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_C3 = CLBLL_L_X4Y143_SLICE_X4Y143_AO5;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_C4 = CLBLM_L_X8Y140_SLICE_X10Y140_AQ;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_C5 = CLBLM_L_X8Y139_SLICE_X10Y139_DQ;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_C6 = CLBLM_R_X3Y141_SLICE_X2Y141_AO6;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_D1 = CLBLL_L_X4Y140_SLICE_X5Y140_DO6;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_D2 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_D3 = CLBLM_R_X7Y141_SLICE_X9Y141_DO6;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_D4 = CLBLL_L_X4Y141_SLICE_X4Y141_CO6;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_D5 = CLBLM_R_X3Y142_SLICE_X3Y142_DO6;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_D6 = CLBLL_L_X4Y140_SLICE_X4Y140_DO6;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_A1 = CLBLM_R_X5Y143_SLICE_X6Y143_AO6;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_A2 = CLBLM_R_X5Y143_SLICE_X6Y143_BO6;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_A3 = CLBLM_R_X7Y137_SLICE_X8Y137_AQ;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_A4 = CLBLL_L_X4Y143_SLICE_X5Y143_AO6;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_A5 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_A6 = CLBLM_L_X8Y139_SLICE_X10Y139_CQ;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_B1 = LIOB33_X0Y67_IOB_X0Y68_I;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_B2 = CLBLM_R_X3Y143_SLICE_X3Y143_AO5;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_B3 = CLBLL_L_X4Y138_SLICE_X5Y138_AQ;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_B4 = CLBLM_R_X3Y143_SLICE_X2Y143_AO6;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_B5 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_B6 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_A1 = CLBLL_L_X4Y133_SLICE_X4Y133_CO6;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_A2 = CLBLM_R_X5Y136_SLICE_X7Y136_DO5;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_A1 = CLBLM_R_X11Y142_SLICE_X15Y142_AQ;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_A2 = CLBLM_L_X8Y144_SLICE_X11Y144_CO6;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_A3 = CLBLM_L_X10Y145_SLICE_X13Y145_AQ;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_A4 = CLBLM_L_X10Y145_SLICE_X13Y145_BO6;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_A6 = CLBLM_R_X7Y144_SLICE_X8Y144_CQ;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_C1 = CLBLL_L_X4Y138_SLICE_X4Y138_AQ;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_C2 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_C3 = CLBLL_L_X2Y140_SLICE_X1Y140_AO6;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_B1 = CLBLM_L_X8Y144_SLICE_X11Y144_BO5;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_B2 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_B3 = CLBLM_R_X11Y144_SLICE_X14Y144_AQ;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_B4 = CLBLM_L_X8Y142_SLICE_X10Y142_D5Q;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_B5 = CLBLM_L_X10Y142_SLICE_X12Y142_CQ;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_B6 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_C3 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_C4 = 1'b1;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_C1 = CLBLM_L_X8Y144_SLICE_X11Y144_CO6;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_C2 = CLBLM_L_X10Y141_SLICE_X12Y141_C5Q;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_C3 = CLBLM_R_X11Y142_SLICE_X15Y142_AQ;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_C4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_C5 = CLBLM_L_X10Y145_SLICE_X13Y145_BO5;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_A3 = CLBLM_L_X8Y135_SLICE_X10Y135_A5Q;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_A6 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_D6 = CLBLM_R_X5Y141_SLICE_X7Y141_CO6;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_B2 = CLBLM_L_X12Y142_SLICE_X16Y142_AQ;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_B3 = CLBLM_R_X3Y136_SLICE_X3Y136_AQ;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_D1 = 1'b1;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_D2 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_D3 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_D4 = 1'b1;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_D5 = 1'b1;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_D6 = 1'b1;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_B5 = 1'b1;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_B6 = 1'b1;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_C1 = CLBLM_L_X10Y136_SLICE_X13Y136_AO6;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_C2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_C3 = 1'b1;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_C5 = CLBLM_L_X8Y135_SLICE_X11Y135_B5Q;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_C6 = CLBLM_R_X13Y137_SLICE_X18Y137_AQ;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_A6 = 1'b1;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_A2 = CLBLM_L_X10Y141_SLICE_X12Y141_C5Q;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_A3 = CLBLM_L_X12Y143_SLICE_X16Y143_BQ;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_A4 = CLBLM_L_X8Y142_SLICE_X10Y142_D5Q;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_B1 = 1'b1;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_B2 = CLBLM_L_X10Y142_SLICE_X12Y142_CQ;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_B3 = CLBLM_R_X11Y144_SLICE_X14Y144_AQ;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_B4 = CLBLM_L_X8Y142_SLICE_X10Y142_D5Q;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_B5 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_B6 = 1'b1;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_D2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_D3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_D4 = CLBLM_L_X10Y134_SLICE_X12Y134_CQ;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_D6 = 1'b1;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_C1 = CLBLM_L_X8Y142_SLICE_X11Y142_DQ;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_C2 = 1'b1;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_C3 = CLBLM_L_X10Y142_SLICE_X12Y142_CQ;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_A6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_C4 = CLBLM_L_X10Y145_SLICE_X12Y145_AO5;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_C5 = CLBLM_L_X8Y144_SLICE_X11Y144_BO5;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_C6 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_AX = CLBLM_L_X10Y135_SLICE_X13Y135_AO6;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_B1 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_B2 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_B3 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_B4 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_B6 = 1'b1;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_D1 = 1'b1;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_D2 = 1'b1;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_D3 = 1'b1;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_D4 = 1'b1;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_D5 = 1'b1;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_D6 = 1'b1;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_C2 = CLBLM_R_X11Y135_SLICE_X15Y135_AQ;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_C5 = 1'b1;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_C6 = 1'b1;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_C1 = CLBLM_R_X3Y140_SLICE_X2Y140_DO6;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_D1 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_D2 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_D3 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_D4 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_D5 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_D6 = 1'b1;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_D1 = CLBLM_L_X8Y135_SLICE_X10Y135_CO5;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_D2 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_D3 = CLBLM_L_X10Y137_SLICE_X12Y137_AQ;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_D4 = CLBLM_R_X11Y132_SLICE_X15Y132_DO6;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_D5 = CLBLM_L_X8Y135_SLICE_X11Y135_DO5;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_D6 = CLBLM_R_X5Y135_SLICE_X6Y135_AQ;
  assign LIOB33_X0Y125_IOB_X0Y126_O = CLBLM_R_X3Y136_SLICE_X3Y136_CQ;
  assign LIOB33_X0Y125_IOB_X0Y125_O = CLBLM_R_X11Y138_SLICE_X15Y138_D5Q;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_A1 = CLBLM_R_X11Y138_SLICE_X15Y138_DQ;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_A2 = CLBLM_L_X12Y140_SLICE_X16Y140_CQ;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_A4 = CLBLM_L_X10Y135_SLICE_X12Y135_BQ;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_A5 = CLBLM_R_X13Y141_SLICE_X18Y141_AO6;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_A6 = 1'b1;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_B1 = 1'b1;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_B3 = CLBLM_R_X11Y139_SLICE_X15Y139_AQ;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_B4 = CLBLM_R_X11Y139_SLICE_X15Y139_DQ;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_B5 = CLBLM_R_X13Y141_SLICE_X18Y141_AO6;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_B6 = 1'b1;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_C2 = CLBLM_R_X11Y139_SLICE_X15Y139_CQ;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_C3 = 1'b1;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_C4 = CLBLM_R_X7Y139_SLICE_X9Y139_AQ;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_C5 = CLBLM_R_X11Y139_SLICE_X15Y139_AQ;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_C6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign RIOI3_X105Y191_OLOGIC_X1Y192_D1 = CLBLM_R_X13Y134_SLICE_X19Y134_BQ;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_D1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_D2 = CLBLM_L_X12Y139_SLICE_X16Y139_DO5;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_D3 = 1'b1;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_D4 = CLBLM_R_X11Y138_SLICE_X15Y138_AQ;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_D5 = CLBLM_R_X11Y140_SLICE_X15Y140_BQ;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_D6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_A1 = CLBLM_R_X11Y140_SLICE_X14Y140_CQ;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_A3 = CLBLM_R_X11Y139_SLICE_X14Y139_AQ;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_A4 = CLBLM_L_X8Y138_SLICE_X10Y138_AQ;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_A5 = CLBLM_R_X7Y136_SLICE_X9Y136_AQ;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_A6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_C5 = 1'b1;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_B2 = CLBLM_R_X11Y139_SLICE_X14Y139_BQ;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_B4 = CLBLM_L_X12Y133_SLICE_X16Y133_BQ;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_B5 = CLBLM_R_X7Y141_SLICE_X8Y141_AQ;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_B6 = 1'b1;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_C2 = CLBLM_R_X11Y139_SLICE_X14Y139_CQ;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_C3 = CLBLM_L_X8Y137_SLICE_X11Y137_CO6;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_C4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_C5 = CLBLM_L_X8Y138_SLICE_X10Y138_AQ;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_A1 = CLBLM_R_X3Y143_SLICE_X3Y143_AO6;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_A2 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_A3 = CLBLL_L_X4Y137_SLICE_X4Y137_DQ;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_A4 = CLBLL_L_X4Y143_SLICE_X5Y143_BO6;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_A5 = CLBLM_R_X7Y141_SLICE_X9Y141_BQ;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_A6 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_C6 = CLBLM_L_X10Y138_SLICE_X13Y138_BQ;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_B1 = CLBLM_R_X5Y143_SLICE_X6Y143_BO5;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_B2 = CLBLL_L_X4Y143_SLICE_X4Y143_CO6;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_B3 = CLBLM_R_X3Y142_SLICE_X3Y142_BO6;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_B4 = CLBLL_L_X4Y142_SLICE_X5Y142_CO6;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_B5 = CLBLL_L_X4Y141_SLICE_X5Y141_AO6;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_B6 = CLBLL_L_X4Y142_SLICE_X4Y142_CO6;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_D1 = 1'b1;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_D2 = 1'b1;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_D3 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_C1 = CLBLM_R_X7Y141_SLICE_X9Y141_BQ;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_C2 = CLBLM_R_X5Y143_SLICE_X6Y143_BO5;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_C3 = CLBLM_R_X3Y142_SLICE_X2Y142_AO6;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_C4 = CLBLL_L_X4Y137_SLICE_X5Y137_BQ;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_C5 = CLBLL_L_X4Y137_SLICE_X4Y137_DQ;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_C6 = CLBLM_R_X3Y139_SLICE_X2Y139_AO5;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_D1 = CLBLM_R_X3Y142_SLICE_X3Y142_BO6;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_D2 = CLBLM_R_X5Y143_SLICE_X6Y143_BO5;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_D3 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_D4 = CLBLL_L_X4Y143_SLICE_X4Y143_CO6;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_D5 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_D6 = CLBLL_L_X4Y141_SLICE_X5Y141_AO6;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_B6 = CLBLM_R_X5Y133_SLICE_X7Y133_DO6;
  assign RIOI3_X105Y191_OLOGIC_X1Y191_D1 = CLBLM_L_X10Y143_SLICE_X13Y143_AQ;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_A1 = CLBLM_R_X3Y142_SLICE_X2Y142_AO6;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_A2 = CLBLL_L_X4Y137_SLICE_X5Y137_BQ;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_A3 = CLBLL_L_X4Y142_SLICE_X4Y142_AO6;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_A4 = CLBLL_L_X4Y142_SLICE_X5Y142_BO6;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_A5 = CLBLM_R_X7Y140_SLICE_X9Y140_AQ;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_A6 = CLBLM_R_X5Y143_SLICE_X6Y143_AO5;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_B1 = CLBLM_L_X8Y132_SLICE_X11Y132_CQ;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_B1 = CLBLM_L_X8Y142_SLICE_X10Y142_AQ;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_B2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_B3 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_B4 = CLBLM_L_X8Y142_SLICE_X11Y142_AQ;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_B2 = CLBLM_L_X8Y132_SLICE_X11Y132_BQ;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_B5 = CLBLL_L_X4Y144_SLICE_X4Y144_AO6;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_B6 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_C1 = CLBLM_L_X8Y142_SLICE_X11Y142_AQ;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_C2 = CLBLM_R_X7Y140_SLICE_X9Y140_AQ;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_C3 = CLBLL_L_X4Y143_SLICE_X5Y143_AO5;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_C4 = CLBLM_R_X5Y143_SLICE_X6Y143_AO5;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_C5 = CLBLM_L_X8Y142_SLICE_X10Y142_AQ;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_C6 = CLBLM_R_X3Y142_SLICE_X3Y142_AO6;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_A1 = 1'b1;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_A2 = 1'b1;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_A3 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_B5 = CLBLM_L_X8Y138_SLICE_X10Y138_AQ;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_A4 = 1'b1;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_A5 = 1'b1;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_A6 = 1'b1;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_B1 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_D1 = CLBLM_R_X3Y142_SLICE_X2Y142_CO6;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_D2 = CLBLL_L_X4Y141_SLICE_X5Y141_DO6;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_D3 = CLBLL_L_X4Y143_SLICE_X5Y143_CO6;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_D4 = CLBLM_R_X3Y141_SLICE_X2Y141_DO6;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_D5 = CLBLM_R_X7Y142_SLICE_X8Y142_BO6;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_D6 = CLBLM_R_X5Y143_SLICE_X7Y143_BO6;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_B2 = 1'b1;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_B3 = 1'b1;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_A1 = CLBLM_R_X7Y138_SLICE_X8Y138_CQ;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_A2 = 1'b1;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_A3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_A5 = CLBLM_L_X8Y132_SLICE_X11Y132_AQ;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_A6 = CLBLM_L_X8Y138_SLICE_X11Y138_CO6;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_C1 = 1'b1;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_C2 = 1'b1;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_B2 = CLBLM_L_X8Y136_SLICE_X11Y136_BQ;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_B3 = CLBLM_L_X8Y138_SLICE_X10Y138_AQ;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_B4 = CLBLM_R_X3Y137_SLICE_X3Y137_BQ;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_B5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_B6 = CLBLM_L_X10Y138_SLICE_X12Y138_CO6;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_D1 = 1'b1;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_D2 = 1'b1;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_C1 = 1'b1;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_C2 = CLBLM_L_X8Y137_SLICE_X11Y137_DO6;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_C3 = CLBLM_L_X8Y134_SLICE_X11Y134_AQ;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_C4 = CLBLM_L_X10Y137_SLICE_X13Y137_AQ;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_C5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_D4 = 1'b1;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_A1 = 1'b1;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_A3 = CLBLM_R_X5Y136_SLICE_X7Y136_DO5;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_A4 = CLBLM_L_X10Y143_SLICE_X13Y143_BQ;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_A5 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_D1 = CLBLM_L_X10Y135_SLICE_X13Y135_B5Q;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_D2 = CLBLM_L_X10Y138_SLICE_X13Y138_CQ;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_D3 = CLBLM_L_X8Y136_SLICE_X11Y136_BQ;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_D4 = CLBLM_R_X5Y137_SLICE_X7Y137_CQ;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_D5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_D6 = 1'b1;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_A6 = 1'b1;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_B1 = 1'b1;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_B2 = 1'b1;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_B3 = 1'b1;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_B4 = 1'b1;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_A1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_A2 = CLBLM_L_X8Y135_SLICE_X10Y135_CO6;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_A3 = CLBLM_L_X8Y136_SLICE_X10Y136_AQ;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_A5 = CLBLM_L_X8Y138_SLICE_X10Y138_AQ;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_A6 = CLBLL_L_X4Y137_SLICE_X4Y137_CQ;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_C1 = 1'b1;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_C2 = 1'b1;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_C3 = 1'b1;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_B1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_B2 = CLBLM_L_X8Y136_SLICE_X10Y136_BQ;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_B3 = CLBLM_L_X8Y138_SLICE_X10Y138_AQ;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_B4 = CLBLM_L_X10Y136_SLICE_X13Y136_BO6;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_B6 = CLBLM_R_X7Y132_SLICE_X9Y132_D5Q;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_D1 = 1'b1;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_D2 = 1'b1;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_D3 = 1'b1;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_C1 = CLBLM_L_X10Y135_SLICE_X13Y135_B5Q;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_C2 = 1'b1;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_C4 = 1'b1;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_C5 = CLBLM_L_X8Y139_SLICE_X10Y139_DQ;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_D4 = 1'b1;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_D5 = 1'b1;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_D6 = 1'b1;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X103Y175_SLICE_X163Y175_A6 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLM_R_X103Y175_SLICE_X163Y175_B1 = 1'b1;
  assign CLBLM_R_X103Y175_SLICE_X163Y175_B2 = 1'b1;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_D1 = CLBLM_L_X8Y138_SLICE_X10Y138_AQ;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_D2 = CLBLM_R_X5Y137_SLICE_X7Y137_CQ;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_D3 = CLBLM_L_X8Y136_SLICE_X10Y136_DQ;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_D4 = CLBLM_R_X7Y134_SLICE_X9Y134_CO6;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_D5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_D6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X103Y175_SLICE_X163Y175_B3 = 1'b1;
  assign CLBLM_R_X103Y175_SLICE_X163Y175_B4 = 1'b1;
  assign CLBLM_R_X103Y175_SLICE_X163Y175_B5 = 1'b1;
  assign CLBLM_R_X103Y175_SLICE_X163Y175_B6 = 1'b1;
  assign CLBLM_R_X103Y175_SLICE_X163Y175_C1 = 1'b1;
  assign CLBLM_R_X103Y175_SLICE_X163Y175_C2 = 1'b1;
  assign CLBLM_R_X103Y175_SLICE_X163Y175_C3 = 1'b1;
  assign CLBLM_R_X103Y175_SLICE_X163Y175_C4 = 1'b1;
  assign CLBLM_R_X103Y175_SLICE_X163Y175_C5 = 1'b1;
  assign CLBLM_R_X103Y175_SLICE_X163Y175_C6 = 1'b1;
  assign CLBLM_R_X103Y175_SLICE_X163Y175_D1 = 1'b1;
  assign CLBLM_R_X103Y175_SLICE_X163Y175_D2 = 1'b1;
  assign CLBLM_R_X103Y175_SLICE_X163Y175_D3 = 1'b1;
  assign CLBLM_R_X103Y175_SLICE_X163Y175_D4 = 1'b1;
  assign CLBLM_R_X103Y175_SLICE_X163Y175_D5 = 1'b1;
  assign CLBLM_R_X103Y175_SLICE_X163Y175_D6 = 1'b1;
  assign CLBLM_R_X103Y175_SLICE_X162Y175_A1 = 1'b1;
  assign CLBLM_R_X103Y175_SLICE_X162Y175_A2 = 1'b1;
  assign CLBLM_R_X103Y175_SLICE_X162Y175_A3 = 1'b1;
  assign CLBLM_R_X103Y175_SLICE_X162Y175_A4 = 1'b1;
  assign CLBLM_R_X103Y175_SLICE_X162Y175_A5 = 1'b1;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_A1 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_A2 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_A3 = CLBLM_R_X11Y136_SLICE_X15Y136_BQ;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_A5 = CLBLM_R_X11Y140_SLICE_X15Y140_C5Q;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_A6 = 1'b1;
  assign CLBLM_R_X103Y175_SLICE_X162Y175_A6 = 1'b1;
  assign CLBLM_R_X103Y175_SLICE_X162Y175_B1 = 1'b1;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_B2 = 1'b1;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_B3 = CLBLM_L_X10Y140_SLICE_X13Y140_DQ;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_B4 = CLBLM_L_X8Y142_SLICE_X11Y142_CQ;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_B6 = CLBLM_R_X11Y140_SLICE_X15Y140_AO5;
  assign CLBLM_R_X103Y175_SLICE_X162Y175_B2 = 1'b1;
  assign CLBLM_R_X103Y175_SLICE_X162Y175_B3 = 1'b1;
  assign CLBLM_R_X103Y175_SLICE_X162Y175_B5 = 1'b1;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_C1 = CLBLM_R_X11Y132_SLICE_X14Y132_BQ;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_C2 = CLBLM_L_X12Y138_SLICE_X16Y138_DQ;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_C3 = CLBLM_R_X11Y143_SLICE_X14Y143_AQ;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_C5 = CLBLM_L_X12Y143_SLICE_X16Y143_AQ;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_C6 = 1'b1;
  assign CLBLM_R_X103Y175_SLICE_X162Y175_C1 = 1'b1;
  assign CLBLM_R_X103Y175_SLICE_X162Y175_C2 = 1'b1;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X103Y175_SLICE_X162Y175_C4 = 1'b1;
  assign CLBLM_R_X103Y175_SLICE_X162Y175_C5 = 1'b1;
  assign CLBLM_R_X103Y175_SLICE_X162Y175_C6 = 1'b1;
  assign CLBLM_R_X103Y175_SLICE_X162Y175_D1 = 1'b1;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_D1 = CLBLM_L_X12Y142_SLICE_X17Y142_AQ;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_D2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_D3 = CLBLM_L_X10Y140_SLICE_X12Y140_A5Q;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_D4 = 1'b1;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_D5 = CLBLM_L_X12Y136_SLICE_X17Y136_BO5;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_D6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X103Y175_SLICE_X162Y175_D2 = 1'b1;
  assign CLBLM_R_X103Y175_SLICE_X162Y175_D3 = 1'b1;
  assign CLBLM_R_X103Y175_SLICE_X162Y175_D4 = 1'b1;
  assign CLBLM_R_X103Y175_SLICE_X162Y175_D5 = 1'b1;
  assign CLBLM_R_X103Y175_SLICE_X162Y175_D6 = 1'b1;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_A1 = CLBLM_R_X13Y143_SLICE_X18Y143_AO6;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_A2 = CLBLM_R_X11Y140_SLICE_X14Y140_BQ;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_A3 = CLBLM_R_X11Y140_SLICE_X14Y140_AQ;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_A4 = CLBLM_L_X12Y143_SLICE_X17Y143_CO5;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_A6 = CLBLM_R_X7Y140_SLICE_X9Y140_CQ;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_B1 = CLBLM_R_X13Y143_SLICE_X18Y143_AO6;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_B2 = CLBLM_R_X11Y140_SLICE_X14Y140_BQ;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_B3 = CLBLM_R_X11Y136_SLICE_X14Y136_AQ;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_B5 = CLBLM_L_X12Y143_SLICE_X17Y143_CO5;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_B6 = CLBLM_L_X12Y140_SLICE_X17Y140_CQ;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_A1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_A2 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_A3 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_A4 = CLBLM_R_X3Y143_SLICE_X2Y143_AO6;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_A5 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_A6 = 1'b1;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_C1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_C2 = CLBLM_R_X11Y140_SLICE_X14Y140_CQ;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_C3 = CLBLM_L_X8Y138_SLICE_X10Y138_AQ;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_B1 = CLBLM_R_X3Y143_SLICE_X2Y143_AO5;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_B2 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_B3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_B4 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_B5 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_B6 = 1'b1;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_D1 = CLBLM_L_X10Y140_SLICE_X13Y140_DQ;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_D2 = 1'b1;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_C1 = CLBLL_L_X4Y143_SLICE_X4Y143_AO6;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_C2 = CLBLM_R_X3Y137_SLICE_X3Y137_CQ;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_C3 = CLBLM_L_X8Y143_SLICE_X10Y143_CQ;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_C4 = CLBLL_L_X4Y143_SLICE_X4Y143_AO5;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_C5 = CLBLM_R_X3Y141_SLICE_X2Y141_AO6;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_C6 = LIOB33_X0Y67_IOB_X0Y67_I;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_D3 = 1'b1;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_D4 = CLBLM_L_X12Y138_SLICE_X16Y138_DQ;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_D5 = CLBLM_R_X11Y140_SLICE_X15Y140_DQ;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_D6 = CLBLM_R_X11Y138_SLICE_X14Y138_CQ;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_D1 = 1'b1;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_D2 = CLBLL_L_X2Y141_SLICE_X1Y141_AO5;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_D3 = CLBLM_L_X8Y143_SLICE_X10Y143_CQ;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_D4 = CLBLM_R_X3Y137_SLICE_X3Y137_CQ;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_D5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_D6 = CLBLM_R_X3Y143_SLICE_X2Y143_AO6;
  assign RIOI3_X105Y127_ILOGIC_X1Y128_D = RIOB33_X105Y127_IOB_X1Y128_I;
  assign RIOI3_X105Y127_ILOGIC_X1Y127_D = RIOB33_X105Y127_IOB_X1Y127_I;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_A1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_A2 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_A3 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_A4 = CLBLL_L_X4Y143_SLICE_X5Y143_BO6;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_A5 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_A6 = 1'b1;
  assign RIOB33_X105Y197_IOB_X1Y198_O = CLBLM_R_X103Y175_SLICE_X163Y175_AO6;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_B1 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_B2 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_B3 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_B4 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_B5 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_B6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y132_D = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_C1 = CLBLM_L_X10Y141_SLICE_X12Y141_AQ;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_C2 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_C3 = CLBLL_L_X4Y143_SLICE_X4Y143_BO6;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_C4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_C5 = CLBLM_R_X11Y141_SLICE_X15Y141_AQ;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_C6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y131_D = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_D1 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_D2 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_D3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_D4 = CLBLL_L_X4Y136_SLICE_X5Y136_CQ;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_D5 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_D6 = CLBLM_R_X3Y143_SLICE_X2Y143_AO6;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_D1 = CLBLM_R_X7Y131_SLICE_X9Y131_AO5;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_A1 = CLBLM_L_X10Y137_SLICE_X12Y137_B5Q;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_A3 = CLBLM_L_X8Y137_SLICE_X11Y137_AQ;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_A4 = CLBLM_L_X8Y143_SLICE_X10Y143_DO5;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_A5 = CLBLM_R_X11Y137_SLICE_X14Y137_AQ;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_A6 = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y156_D1 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_B1 = CLBLM_L_X10Y137_SLICE_X12Y137_CQ;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_B2 = CLBLM_L_X8Y137_SLICE_X11Y137_BQ;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_B3 = CLBLM_R_X5Y132_SLICE_X7Y132_DO6;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_B5 = 1'b1;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_B6 = CLBLM_R_X7Y137_SLICE_X9Y137_AQ;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_C1 = CLBLM_R_X7Y136_SLICE_X9Y136_BO5;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_C2 = CLBLL_L_X4Y134_SLICE_X4Y134_AQ;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_C3 = CLBLM_R_X5Y141_SLICE_X7Y141_DO6;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_C5 = CLBLM_L_X10Y134_SLICE_X12Y134_CQ;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_C6 = 1'b1;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_D1 = CLBLM_L_X10Y139_SLICE_X13Y139_AQ;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_D2 = CLBLM_R_X5Y137_SLICE_X7Y137_BQ;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_D3 = CLBLM_R_X11Y139_SLICE_X15Y139_CQ;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_D4 = CLBLM_L_X8Y137_SLICE_X10Y137_BO6;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_D5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_D6 = CLBLM_R_X7Y139_SLICE_X8Y139_BQ;
  assign LIOB33_X0Y129_IOB_X0Y129_O = CLBLM_R_X5Y136_SLICE_X6Y136_CQ;
  assign LIOB33_X0Y129_IOB_X0Y130_O = CLBLL_L_X52Y126_SLICE_X78Y126_AO6;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_A1 = 1'b1;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_A2 = CLBLM_R_X11Y135_SLICE_X15Y135_BQ;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_A3 = CLBLM_L_X8Y137_SLICE_X10Y137_AQ;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_A4 = CLBLM_R_X7Y144_SLICE_X9Y144_BO6;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_A6 = CLBLM_L_X10Y137_SLICE_X13Y137_AQ;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_B1 = 1'b1;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_B2 = CLBLM_R_X7Y136_SLICE_X9Y136_CQ;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_B3 = CLBLM_L_X10Y139_SLICE_X13Y139_AQ;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_B4 = CLBLM_R_X5Y136_SLICE_X7Y136_BQ;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_B5 = 1'b1;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_B6 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_A1 = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y156_T1 = 1'b1;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_C1 = CLBLM_L_X10Y139_SLICE_X13Y139_AQ;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_C2 = CLBLL_L_X4Y136_SLICE_X5Y136_A5Q;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_C3 = CLBLM_R_X5Y136_SLICE_X7Y136_BQ;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_C4 = CLBLM_R_X7Y136_SLICE_X9Y136_CQ;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_C5 = CLBLM_R_X11Y139_SLICE_X15Y139_CQ;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_C6 = CLBLM_L_X8Y135_SLICE_X10Y135_BQ;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_A2 = CLBLM_R_X13Y144_SLICE_X19Y144_AQ;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_A3 = 1'b1;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_A5 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_D1 = CLBLM_R_X7Y137_SLICE_X8Y137_DO6;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_D2 = CLBLM_L_X10Y136_SLICE_X12Y136_CO6;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_D3 = CLBLM_L_X8Y135_SLICE_X10Y135_DO6;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_D4 = CLBLM_R_X5Y135_SLICE_X7Y135_CO5;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_D5 = CLBLM_L_X8Y137_SLICE_X10Y137_BO5;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_D6 = CLBLM_L_X10Y145_SLICE_X12Y145_CO6;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_A6 = 1'b1;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_A1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_A2 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_A3 = CLBLM_R_X11Y141_SLICE_X15Y141_AQ;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_A4 = CLBLM_L_X10Y131_SLICE_X13Y131_CQ;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_A5 = CLBLM_R_X11Y136_SLICE_X14Y136_DQ;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_B4 = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y155_D1 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_B1 = 1'b1;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_B2 = CLBLM_R_X11Y141_SLICE_X15Y141_BQ;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_B3 = CLBLM_R_X11Y140_SLICE_X15Y140_BQ;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_B4 = CLBLM_R_X11Y141_SLICE_X14Y141_BQ;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_B5 = CLBLM_L_X8Y143_SLICE_X10Y143_DO6;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_A1 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_A3 = CLBLM_R_X7Y131_SLICE_X9Y131_AQ;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_A4 = CLBLM_R_X11Y139_SLICE_X15Y139_A5Q;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_A5 = CLBLM_L_X8Y131_SLICE_X11Y131_BQ;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_A6 = 1'b1;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_C2 = CLBLM_R_X11Y141_SLICE_X15Y141_CQ;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_C3 = CLBLM_R_X13Y143_SLICE_X18Y143_AO6;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_C4 = CLBLM_R_X11Y139_SLICE_X14Y139_CQ;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_B1 = CLBLM_L_X8Y131_SLICE_X10Y131_A5Q;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_B2 = CLBLM_R_X7Y131_SLICE_X9Y131_BQ;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_B4 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_B5 = CLBLM_R_X5Y134_SLICE_X7Y134_DO6;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_B6 = CLBLM_R_X5Y136_SLICE_X6Y136_CQ;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_D1 = CLBLM_L_X10Y140_SLICE_X13Y140_BQ;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_C1 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_C2 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_C3 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_C4 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_C5 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_C6 = 1'b1;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_D3 = 1'b1;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_D4 = CLBLM_R_X11Y143_SLICE_X15Y143_AQ;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_A1 = CLBLM_L_X10Y141_SLICE_X13Y141_AQ;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_A2 = CLBLM_L_X12Y140_SLICE_X16Y140_DQ;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_A3 = CLBLM_R_X11Y141_SLICE_X14Y141_AQ;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_A4 = CLBLM_R_X11Y141_SLICE_X14Y141_DO6;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_D1 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_D2 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_D3 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_D4 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_D5 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_D6 = 1'b1;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_B1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_A1 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_A2 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_A3 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_A4 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_A5 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_A6 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_A1 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_A2 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_A3 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_B1 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_B2 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_B3 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_B4 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_B5 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_B6 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_A5 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_A6 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_C1 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_C2 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_C3 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_C4 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_C5 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_C6 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_B4 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_B5 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_B6 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_C1 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_C2 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_C3 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_C4 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_D1 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_D2 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_D3 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_D4 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_D5 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_D6 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_D1 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_D2 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_D3 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_D4 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_D5 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_D6 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_A1 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_A2 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_A3 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_A4 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_A5 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_A6 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_B1 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_B2 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_B3 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_B4 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_B5 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_B6 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_C1 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_C2 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_C3 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_C4 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_C5 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_C6 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_D1 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_D2 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_D3 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_D4 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_D5 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_D6 = 1'b1;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_A1 = CLBLM_L_X8Y138_SLICE_X11Y138_DO6;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_A3 = CLBLM_L_X8Y139_SLICE_X11Y139_BQ;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_A5 = CLBLM_L_X10Y136_SLICE_X13Y136_CO6;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_A6 = 1'b1;
  assign LIOB33_X0Y131_IOB_X0Y131_O = CLBLM_R_X7Y131_SLICE_X9Y131_AO5;
  assign LIOB33_X0Y131_IOB_X0Y132_O = CLBLM_R_X7Y131_SLICE_X9Y131_AQ;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_B2 = CLBLM_L_X8Y138_SLICE_X11Y138_BQ;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_B3 = CLBLM_L_X8Y138_SLICE_X11Y138_AQ;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_B5 = 1'b1;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_B6 = 1'b1;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_C1 = CLBLM_L_X8Y139_SLICE_X11Y139_AQ;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_C2 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_C3 = CLBLM_L_X10Y137_SLICE_X12Y137_AQ;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_C4 = CLBLM_R_X5Y140_SLICE_X7Y140_BQ;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_C5 = CLBLM_L_X10Y135_SLICE_X12Y135_BQ;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_C6 = 1'b1;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_D1 = 1'b1;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_D2 = CLBLM_L_X10Y142_SLICE_X12Y142_DQ;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_D3 = CLBLM_L_X12Y139_SLICE_X16Y139_A5Q;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_D4 = CLBLM_R_X7Y135_SLICE_X8Y135_CQ;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_D5 = 1'b1;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_D6 = CLBLM_L_X8Y138_SLICE_X11Y138_AQ;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_A1 = CLBLL_L_X4Y138_SLICE_X4Y138_AQ;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_A2 = CLBLM_L_X8Y138_SLICE_X10Y138_DQ;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_A3 = CLBLM_L_X8Y138_SLICE_X10Y138_AQ;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_A5 = RIOB33_X105Y119_IOB_X1Y119_I;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_A6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_B2 = 1'b1;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_B1 = CLBLM_R_X7Y138_SLICE_X9Y138_CO6;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_B2 = CLBLM_L_X8Y138_SLICE_X10Y138_BQ;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_B3 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_B4 = CLBLM_R_X7Y139_SLICE_X8Y139_BQ;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_B6 = CLBLM_R_X11Y135_SLICE_X14Y135_AQ;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_B4 = 1'b1;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_C1 = CLBLM_L_X8Y136_SLICE_X11Y136_AQ;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_C2 = 1'b1;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_C3 = CLBLM_L_X8Y136_SLICE_X11Y136_DO5;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_C5 = CLBLM_L_X8Y142_SLICE_X10Y142_AQ;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_B6 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_A1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_A2 = CLBLM_R_X13Y143_SLICE_X18Y143_BQ;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_A3 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_A4 = CLBLM_R_X13Y139_SLICE_X19Y139_AQ;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_A5 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_A6 = 1'b1;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_D1 = CLBLM_L_X10Y135_SLICE_X13Y135_B5Q;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_D2 = CLBLM_L_X8Y138_SLICE_X10Y138_CQ;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_D3 = RIOB33_X105Y119_IOB_X1Y119_I;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_D4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_D5 = CLBLM_L_X8Y138_SLICE_X10Y138_D5Q;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_D6 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_B6 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_C1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_C2 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_C3 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_C4 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_C5 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_C6 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_D1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_D2 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_D3 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_D4 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_C3 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_D5 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_D6 = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_D1 = LIOB33_X0Y61_IOB_X0Y61_I;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_A1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_A2 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_A3 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_A4 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_A5 = 1'b1;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_A1 = CLBLM_L_X8Y144_SLICE_X11Y144_CO6;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_A3 = CLBLM_R_X11Y142_SLICE_X15Y142_AQ;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_A4 = CLBLM_L_X10Y135_SLICE_X13Y135_BQ;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_A5 = CLBLM_R_X11Y143_SLICE_X15Y143_AQ;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_A6 = CLBLM_L_X10Y145_SLICE_X13Y145_BO6;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_A6 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_B1 = 1'b1;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_B1 = CLBLM_L_X8Y144_SLICE_X11Y144_CO6;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_B2 = CLBLM_R_X11Y142_SLICE_X15Y142_BQ;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_B3 = CLBLM_L_X10Y142_SLICE_X12Y142_BQ;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_B4 = CLBLM_L_X8Y138_SLICE_X10Y138_AQ;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_B6 = CLBLM_L_X10Y145_SLICE_X13Y145_BO6;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_B2 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_B3 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_B5 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_A1 = CLBLM_L_X12Y132_SLICE_X16Y132_CQ;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_A2 = CLBLL_L_X4Y135_SLICE_X4Y135_A5Q;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_A4 = CLBLM_R_X5Y137_SLICE_X6Y137_BQ;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_A6 = LIOB33_X0Y53_IOB_X0Y53_I;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_C1 = CLBLM_R_X11Y137_SLICE_X15Y137_AQ;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_C2 = CLBLM_L_X10Y143_SLICE_X13Y143_CO6;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_C3 = CLBLM_R_X11Y144_SLICE_X14Y144_DO6;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_B1 = CLBLM_R_X5Y135_SLICE_X6Y135_DQ;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_B2 = CLBLM_R_X7Y132_SLICE_X9Y132_BQ;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_B4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_B5 = CLBLM_L_X8Y138_SLICE_X10Y138_AQ;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_B6 = CLBLM_L_X8Y132_SLICE_X10Y132_BQ;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_D1 = CLBLM_R_X11Y144_SLICE_X15Y144_CO6;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_C1 = CLBLL_L_X4Y134_SLICE_X4Y134_B5Q;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_C2 = CLBLM_R_X7Y132_SLICE_X9Y132_CQ;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_C3 = CLBLM_L_X8Y138_SLICE_X10Y138_AQ;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_C4 = CLBLM_L_X12Y132_SLICE_X16Y132_CQ;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_C6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_D3 = CLBLM_R_X11Y142_SLICE_X15Y142_DQ;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_D4 = CLBLM_L_X10Y144_SLICE_X12Y144_AO6;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_A1 = CLBLM_R_X11Y144_SLICE_X14Y144_DO6;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_A2 = CLBLM_L_X10Y144_SLICE_X12Y144_AO6;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_A5 = RIOB33_X105Y143_IOB_X1Y144_I;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_D2 = CLBLM_L_X8Y132_SLICE_X10Y132_BQ;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_D3 = CLBLM_R_X7Y137_SLICE_X8Y137_BQ;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_A6 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_D4 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_D5 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_D6 = 1'b1;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_A6 = CLBLM_R_X11Y142_SLICE_X14Y142_CO6;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_B1 = CLBLM_R_X13Y143_SLICE_X18Y143_AO6;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_B2 = CLBLM_R_X11Y142_SLICE_X14Y142_BQ;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_B3 = CLBLM_R_X11Y141_SLICE_X15Y141_CQ;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_A1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_A2 = CLBLM_R_X5Y132_SLICE_X7Y132_BO6;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_A3 = CLBLM_L_X8Y133_SLICE_X11Y133_AQ;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_A4 = CLBLM_R_X11Y138_SLICE_X15Y138_BQ;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_A6 = 1'b1;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_C1 = CLBLM_R_X11Y142_SLICE_X15Y142_AQ;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_C2 = CLBLM_R_X11Y142_SLICE_X14Y142_AQ;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_B2 = CLBLM_R_X7Y132_SLICE_X8Y132_BQ;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_B3 = CLBLM_R_X7Y134_SLICE_X8Y134_C5Q;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_B4 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_B6 = 1'b1;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_D1 = CLBLM_R_X11Y142_SLICE_X15Y142_DQ;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_D2 = CLBLM_R_X11Y144_SLICE_X14Y144_CO6;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_C2 = CLBLM_R_X7Y132_SLICE_X8Y132_CQ;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_C3 = CLBLM_R_X5Y132_SLICE_X7Y132_BO5;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_C4 = CLBLM_R_X7Y132_SLICE_X8Y132_AO5;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_C5 = CLBLM_R_X7Y144_SLICE_X8Y144_AQ;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_C6 = CLBLM_R_X5Y132_SLICE_X7Y132_DO6;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_D5 = CLBLM_R_X11Y143_SLICE_X15Y143_BQ;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_D6 = CLBLM_L_X10Y142_SLICE_X13Y142_CQ;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_B4 = CLBLM_L_X12Y136_SLICE_X16Y136_AQ;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_B5 = CLBLM_L_X10Y141_SLICE_X12Y141_AQ;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_D1 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_D2 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_D3 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_B6 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_D4 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_D5 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_D6 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_C1 = CLBLM_L_X12Y136_SLICE_X16Y136_DQ;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_C2 = CLBLM_L_X10Y141_SLICE_X13Y141_CQ;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_C3 = CLBLM_L_X10Y139_SLICE_X13Y139_B5Q;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_C4 = CLBLM_L_X12Y134_SLICE_X17Y134_AO6;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_C5 = CLBLM_L_X8Y138_SLICE_X10Y138_BQ;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOB33_X0Y133_IOB_X0Y134_O = CLBLM_R_X3Y133_SLICE_X3Y133_AQ;
  assign LIOB33_X0Y133_IOB_X0Y133_O = CLBLM_R_X3Y137_SLICE_X3Y137_AQ;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_A1 = CLBLM_L_X10Y142_SLICE_X12Y142_DQ;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_A3 = CLBLM_L_X8Y139_SLICE_X11Y139_AQ;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_A4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_A5 = CLBLM_L_X8Y138_SLICE_X10Y138_AQ;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_A6 = CLBLM_L_X8Y139_SLICE_X11Y139_CO6;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_B1 = CLBLM_R_X7Y144_SLICE_X8Y144_BQ;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_B3 = 1'b1;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_B4 = CLBLM_L_X10Y135_SLICE_X12Y135_BQ;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_B6 = 1'b1;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_C1 = CLBLM_L_X10Y139_SLICE_X13Y139_AQ;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_C2 = CLBLM_L_X8Y144_SLICE_X11Y144_AQ;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_C3 = CLBLM_R_X5Y140_SLICE_X7Y140_BQ;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_C4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_C5 = CLBLM_R_X11Y139_SLICE_X15Y139_CQ;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_C6 = CLBLM_L_X10Y138_SLICE_X12Y138_DO6;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_D1 = CLBLM_R_X7Y140_SLICE_X8Y140_DO6;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_D2 = CLBLM_L_X12Y141_SLICE_X17Y141_BO6;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_D3 = CLBLM_R_X13Y137_SLICE_X18Y137_DO6;
  assign RIOI3_X105Y129_ILOGIC_X1Y130_D = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_D1 = CLBLM_L_X10Y139_SLICE_X13Y139_AQ;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_D2 = CLBLM_L_X8Y141_SLICE_X10Y141_CQ;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_D3 = CLBLM_R_X7Y139_SLICE_X8Y139_A5Q;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_D4 = CLBLM_R_X11Y139_SLICE_X15Y139_CQ;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_D5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_D6 = CLBLM_L_X10Y138_SLICE_X12Y138_DO6;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_D4 = CLBLM_R_X11Y143_SLICE_X14Y143_BO6;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_D5 = CLBLL_L_X4Y141_SLICE_X4Y141_DO6;
  assign RIOI3_X105Y129_ILOGIC_X1Y129_D = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_D6 = CLBLM_L_X10Y136_SLICE_X13Y136_DO6;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_A1 = CLBLM_L_X8Y139_SLICE_X10Y139_CQ;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_A2 = 1'b1;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_A3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_A5 = CLBLM_R_X11Y136_SLICE_X14Y136_CO5;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_A6 = CLBLM_R_X11Y139_SLICE_X15Y139_DQ;
  assign LIOB33_X0Y195_IOB_X0Y196_O = LIOB33_X0Y69_IOB_X0Y69_I;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_B1 = 1'b1;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_B2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_B3 = CLBLM_L_X8Y139_SLICE_X11Y139_CO6;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_B4 = CLBLM_R_X11Y141_SLICE_X15Y141_BQ;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_B5 = CLBLL_L_X4Y135_SLICE_X5Y135_BQ;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOB33_X0Y195_IOB_X0Y195_O = LIOB33_X0Y63_IOB_X0Y64_I;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_C1 = CLBLM_L_X8Y138_SLICE_X11Y138_BQ;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_C2 = CLBLM_L_X8Y139_SLICE_X10Y139_CQ;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_C4 = CLBLM_L_X12Y134_SLICE_X17Y134_AO6;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_C5 = CLBLM_L_X10Y139_SLICE_X13Y139_B5Q;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_C6 = CLBLM_R_X5Y139_SLICE_X7Y139_AQ;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y144_D = RIOB33_X105Y143_IOB_X1Y144_I;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_D1 = CLBLL_L_X4Y133_SLICE_X5Y133_BO6;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_D2 = 1'b1;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_D3 = CLBLM_L_X8Y139_SLICE_X10Y139_DQ;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_D4 = CLBLM_L_X12Y140_SLICE_X17Y140_BQ;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_D5 = CLBLM_R_X5Y137_SLICE_X7Y137_B5Q;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_D6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign RIOB33_X105Y177_IOB_X1Y177_O = CLBLM_R_X103Y177_SLICE_X163Y177_AO6;
  assign RIOB33_X105Y177_IOB_X1Y178_O = CLBLM_R_X103Y177_SLICE_X163Y177_AO5;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_A3 = CLBLM_L_X10Y141_SLICE_X12Y141_AQ;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_A5 = CLBLM_L_X8Y131_SLICE_X10Y131_AQ;
  assign LIOI3_X0Y79_OLOGIC_X0Y80_D1 = CLBLL_L_X2Y133_SLICE_X0Y133_AO6;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_A1 = CLBLM_R_X11Y142_SLICE_X15Y142_BQ;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_A3 = CLBLM_R_X11Y143_SLICE_X15Y143_AQ;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_A4 = CLBLM_L_X8Y143_SLICE_X10Y143_CQ;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_A5 = CLBLM_L_X10Y145_SLICE_X13Y145_BO6;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_A6 = CLBLM_L_X8Y144_SLICE_X11Y144_CO6;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_B1 = CLBLM_R_X11Y143_SLICE_X15Y143_DO6;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_B3 = CLBLM_R_X11Y144_SLICE_X14Y144_DO6;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_B4 = CLBLM_L_X10Y144_SLICE_X12Y144_AO6;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_B5 = CLBLM_L_X12Y143_SLICE_X17Y143_AQ;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_B6 = 1'b1;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_A2 = CLBLM_R_X7Y133_SLICE_X9Y133_BQ;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_A3 = CLBLM_R_X7Y133_SLICE_X9Y133_AQ;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_A4 = CLBLM_R_X5Y134_SLICE_X7Y134_CQ;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_A5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_A6 = CLBLM_L_X8Y138_SLICE_X10Y138_AQ;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_C1 = CLBLM_R_X11Y143_SLICE_X15Y143_BQ;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_C2 = CLBLM_R_X11Y142_SLICE_X15Y142_DQ;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_C3 = CLBLM_L_X10Y143_SLICE_X12Y143_CQ;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_B1 = CLBLL_L_X4Y137_SLICE_X4Y137_A5Q;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_B2 = CLBLM_R_X7Y133_SLICE_X9Y133_BQ;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_B4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_B5 = CLBLM_L_X10Y133_SLICE_X13Y133_BQ;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_B5 = CLBLM_L_X12Y140_SLICE_X16Y140_DQ;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_B6 = CLBLM_L_X8Y138_SLICE_X10Y138_AQ;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_D1 = CLBLM_R_X11Y143_SLICE_X15Y143_CO5;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_B6 = 1'b1;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_C1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_C2 = CLBLM_R_X7Y133_SLICE_X9Y133_CQ;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_C3 = CLBLM_R_X7Y134_SLICE_X9Y134_CO6;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_C4 = CLBLM_L_X8Y138_SLICE_X10Y138_AQ;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_C5 = CLBLL_L_X4Y133_SLICE_X5Y133_A5Q;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_D4 = CLBLM_R_X11Y142_SLICE_X15Y142_BQ;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_A1 = CLBLM_R_X11Y143_SLICE_X14Y143_BO5;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_A2 = CLBLM_L_X12Y142_SLICE_X16Y142_BQ;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_A3 = CLBLM_L_X8Y141_SLICE_X11Y141_DO5;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_A4 = CLBLM_L_X10Y144_SLICE_X12Y144_BO6;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_A5 = CLBLM_L_X10Y145_SLICE_X13Y145_BO6;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_D1 = CLBLL_L_X4Y141_SLICE_X4Y141_DO6;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_D2 = CLBLM_R_X3Y140_SLICE_X2Y140_DO6;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_D3 = CLBLL_L_X4Y142_SLICE_X4Y142_BO6;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_D4 = CLBLL_L_X4Y142_SLICE_X5Y142_DO6;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_D5 = CLBLM_R_X5Y142_SLICE_X6Y142_CO6;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_D6 = CLBLL_L_X4Y139_SLICE_X4Y139_BO6;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_B1 = CLBLM_R_X11Y143_SLICE_X14Y143_DO6;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_B2 = 1'b1;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_B3 = CLBLM_L_X10Y142_SLICE_X12Y142_CQ;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_B4 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_A1 = CLBLM_L_X8Y138_SLICE_X10Y138_AQ;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_A2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_A3 = CLBLM_R_X7Y133_SLICE_X8Y133_AQ;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_A4 = CLBLM_R_X7Y134_SLICE_X9Y134_BQ;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_A5 = CLBLM_L_X8Y139_SLICE_X11Y139_DO6;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_C1 = 1'b1;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_C2 = CLBLM_R_X11Y142_SLICE_X15Y142_CQ;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_C3 = CLBLM_L_X10Y142_SLICE_X13Y142_CQ;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_B1 = 1'b1;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_B2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_B3 = CLBLM_R_X7Y135_SLICE_X8Y135_AQ;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_B5 = CLBLM_R_X7Y133_SLICE_X9Y133_AQ;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_B6 = CLBLM_L_X8Y139_SLICE_X11Y139_DO6;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_C4 = CLBLM_L_X10Y138_SLICE_X12Y138_A5Q;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_D1 = CLBLM_R_X11Y143_SLICE_X15Y143_BQ;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_C1 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_C5 = 1'b1;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_C2 = CLBLM_R_X7Y133_SLICE_X8Y133_CQ;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_C3 = CLBLM_R_X11Y131_SLICE_X15Y131_BQ;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_C4 = 1'b1;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_C5 = CLBLM_R_X7Y133_SLICE_X8Y133_DO6;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_C6 = 1'b1;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_D4 = CLBLM_R_X11Y143_SLICE_X14Y143_CO6;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_D6 = CLBLM_R_X11Y142_SLICE_X15Y142_DQ;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_D2 = LIOB33_X0Y53_IOB_X0Y53_I;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_D3 = CLBLM_R_X7Y135_SLICE_X9Y135_B5Q;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_D4 = CLBLL_L_X4Y135_SLICE_X4Y135_A5Q;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_D5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_D6 = CLBLM_R_X5Y137_SLICE_X6Y137_BQ;
  assign LIOB33_X0Y135_IOB_X0Y136_O = CLBLM_R_X3Y135_SLICE_X3Y135_AQ;
  assign LIOB33_X0Y135_IOB_X0Y135_O = CLBLM_R_X3Y136_SLICE_X3Y136_AQ;
  assign RIOI3_X105Y179_OLOGIC_X1Y180_D1 = CLBLM_L_X12Y138_SLICE_X17Y138_DO6;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_A1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_A3 = CLBLM_R_X7Y138_SLICE_X8Y138_BQ;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_A4 = CLBLM_L_X12Y140_SLICE_X16Y140_DQ;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_A5 = CLBLM_R_X7Y134_SLICE_X8Y134_BQ;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_A6 = 1'b1;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_B1 = CLBLM_L_X12Y134_SLICE_X17Y134_AO6;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_B2 = CLBLM_L_X8Y140_SLICE_X11Y140_BQ;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_B3 = CLBLM_L_X10Y139_SLICE_X13Y139_B5Q;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_B5 = CLBLM_R_X11Y136_SLICE_X14Y136_AQ;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_B6 = CLBLM_L_X8Y141_SLICE_X10Y141_CQ;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_C1 = CLBLM_L_X10Y137_SLICE_X13Y137_BQ;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_C2 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_C3 = CLBLM_R_X11Y136_SLICE_X14Y136_DQ;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_C4 = 1'b1;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_C5 = CLBLM_R_X7Y144_SLICE_X8Y144_CQ;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_C6 = 1'b1;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_D1 = CLBLM_L_X8Y140_SLICE_X11Y140_CO5;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_D2 = CLBLM_L_X8Y136_SLICE_X11Y136_CQ;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_D3 = CLBLM_R_X7Y144_SLICE_X8Y144_CQ;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_D4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_D5 = CLBLM_L_X8Y141_SLICE_X10Y141_DQ;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_D6 = CLBLM_L_X10Y142_SLICE_X12Y142_DQ;
  assign RIOI3_X105Y179_OLOGIC_X1Y180_T1 = 1'b1;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_A1 = CLBLL_L_X4Y141_SLICE_X4Y141_DO6;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_A2 = CLBLM_L_X8Y132_SLICE_X11Y132_BQ;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_A3 = CLBLM_L_X10Y143_SLICE_X12Y143_BQ;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_A5 = CLBLM_R_X3Y140_SLICE_X2Y140_DO6;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_A6 = 1'b1;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_B1 = CLBLM_R_X11Y141_SLICE_X15Y141_DQ;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_B2 = CLBLM_L_X8Y140_SLICE_X10Y140_BQ;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_B3 = CLBLM_L_X8Y143_SLICE_X10Y143_DO6;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_B4 = CLBLM_L_X8Y142_SLICE_X10Y142_BQ;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_B5 = 1'b1;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_C2 = CLBLM_L_X8Y140_SLICE_X10Y140_CQ;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_C3 = CLBLM_R_X11Y140_SLICE_X14Y140_CQ;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_C4 = 1'b1;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_C5 = CLBLM_L_X8Y143_SLICE_X10Y143_DO5;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_C6 = CLBLM_L_X10Y142_SLICE_X12Y142_DQ;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_D1 = CLBLM_R_X7Y138_SLICE_X8Y138_BQ;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_D2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_D3 = CLBLM_L_X8Y136_SLICE_X11Y136_DO6;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_D4 = CLBLM_R_X7Y143_SLICE_X9Y143_CQ;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_D5 = 1'b1;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_D6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign RIOI3_X105Y179_OLOGIC_X1Y179_D1 = CLBLM_L_X12Y144_SLICE_X17Y144_AO5;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_A2 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_A3 = CLBLM_R_X11Y144_SLICE_X15Y144_AQ;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_A4 = CLBLM_R_X11Y142_SLICE_X15Y142_DQ;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_A5 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_A6 = CLBLM_R_X7Y131_SLICE_X9Y131_AQ;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_B1 = CLBLM_R_X11Y144_SLICE_X15Y144_DO6;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_B2 = CLBLM_L_X10Y144_SLICE_X12Y144_AO6;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_B4 = CLBLM_R_X11Y144_SLICE_X14Y144_DO6;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_B5 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_B6 = CLBLM_L_X10Y141_SLICE_X13Y141_CQ;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_A1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_A2 = CLBLM_R_X7Y135_SLICE_X9Y135_CO5;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_A3 = 1'b1;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_A5 = CLBLM_R_X7Y138_SLICE_X9Y138_AQ;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_A6 = CLBLM_R_X7Y132_SLICE_X9Y132_CQ;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_C1 = CLBLM_R_X11Y143_SLICE_X15Y143_CO5;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_C2 = CLBLM_L_X10Y144_SLICE_X13Y144_DO6;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_C3 = CLBLM_R_X11Y143_SLICE_X15Y143_AQ;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_B1 = CLBLM_L_X10Y139_SLICE_X13Y139_B5Q;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_B2 = CLBLM_R_X7Y134_SLICE_X9Y134_BQ;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_B3 = CLBLM_R_X13Y134_SLICE_X19Y134_AQ;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_B4 = CLBLM_L_X12Y134_SLICE_X17Y134_AO6;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_B6 = CLBLM_R_X7Y137_SLICE_X8Y137_CQ;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_D1 = CLBLM_L_X10Y144_SLICE_X13Y144_DO6;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_C1 = CLBLM_R_X7Y133_SLICE_X8Y133_AQ;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_C2 = CLBLM_R_X7Y139_SLICE_X8Y139_BQ;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_C3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_C4 = CLBLM_R_X5Y140_SLICE_X6Y140_AO6;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_C5 = CLBLM_R_X7Y134_SLICE_X9Y134_DO6;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_C6 = CLBLM_L_X8Y137_SLICE_X11Y137_CO5;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_D3 = CLBLM_R_X11Y144_SLICE_X15Y144_BQ;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_D4 = CLBLM_L_X10Y145_SLICE_X13Y145_AQ;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_A2 = CLBLM_R_X11Y141_SLICE_X14Y141_AQ;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_A3 = CLBLM_R_X11Y144_SLICE_X14Y144_AQ;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_A4 = CLBLM_R_X11Y145_SLICE_X14Y145_AO6;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_A5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_D2 = CLBLM_L_X8Y138_SLICE_X10Y138_AQ;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_D3 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_D4 = CLBLM_L_X10Y134_SLICE_X12Y134_CQ;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_D5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_D6 = CLBLL_L_X4Y134_SLICE_X4Y134_AQ;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_A6 = CLBLM_R_X11Y143_SLICE_X14Y143_DO6;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_B1 = CLBLM_L_X10Y144_SLICE_X12Y144_AQ;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_B2 = CLBLM_L_X8Y140_SLICE_X10Y140_DQ;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_B3 = CLBLM_L_X10Y143_SLICE_X13Y143_AQ;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_B4 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_A1 = 1'b1;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_A4 = CLBLM_R_X7Y134_SLICE_X8Y134_DO5;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_A5 = CLBLM_R_X7Y135_SLICE_X9Y135_B5Q;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_A6 = CLBLM_R_X7Y134_SLICE_X9Y134_AQ;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_C1 = CLBLM_L_X10Y142_SLICE_X12Y142_CQ;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_C2 = CLBLM_R_X11Y144_SLICE_X14Y144_AQ;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_C3 = CLBLM_L_X10Y143_SLICE_X12Y143_AQ;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_B1 = 1'b1;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_B2 = CLBLM_R_X7Y134_SLICE_X8Y134_BQ;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_B4 = CLBLM_R_X7Y135_SLICE_X8Y135_BQ;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_B5 = CLBLM_R_X7Y135_SLICE_X8Y135_DO6;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_B6 = CLBLM_R_X13Y134_SLICE_X19Y134_CQ;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_D2 = 1'b1;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_C2 = CLBLM_R_X5Y136_SLICE_X6Y136_CQ;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_C3 = CLBLM_L_X8Y134_SLICE_X10Y134_A5Q;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_C4 = 1'b1;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_C5 = CLBLM_R_X7Y137_SLICE_X8Y137_AQ;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_C6 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_D3 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_D4 = CLBLM_R_X11Y145_SLICE_X14Y145_AO5;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_D5 = 1'b1;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_D6 = CLBLM_R_X11Y143_SLICE_X14Y143_DO6;
  assign LIOB33_X0Y137_IOB_X0Y137_O = CLBLM_R_X3Y137_SLICE_X2Y137_BQ;
  assign LIOB33_X0Y137_IOB_X0Y138_O = CLBLM_R_X3Y136_SLICE_X3Y136_DQ;
  assign LIOI3_X0Y151_OLOGIC_X0Y152_D1 = LIOB33_X0Y65_IOB_X0Y66_I;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_D1 = CLBLM_R_X7Y133_SLICE_X8Y133_AQ;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_D2 = CLBLM_L_X10Y134_SLICE_X12Y134_CQ;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_D3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_D4 = CLBLL_L_X4Y134_SLICE_X4Y134_AQ;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_D5 = CLBLM_R_X7Y139_SLICE_X8Y139_BQ;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_D6 = 1'b1;
  assign LIOI3_X0Y151_OLOGIC_X0Y152_T1 = 1'b1;
  assign RIOI3_X105Y195_OLOGIC_X1Y196_D1 = CLBLM_R_X13Y143_SLICE_X18Y143_AQ;
  assign LIOI3_X0Y151_OLOGIC_X0Y151_D1 = LIOB33_X0Y65_IOB_X0Y65_I;
  assign RIOI3_X105Y195_OLOGIC_X1Y196_T1 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_A1 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_A2 = CLBLL_L_X4Y142_SLICE_X4Y142_BO6;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_A3 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_A4 = CLBLM_R_X5Y140_SLICE_X6Y140_AO6;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_A5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_A5 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_A6 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_A6 = CLBLM_L_X8Y134_SLICE_X10Y134_CO6;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_B1 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_B2 = CLBLM_R_X3Y140_SLICE_X2Y140_DO6;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_B3 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_B4 = CLBLM_R_X5Y142_SLICE_X6Y142_CO6;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_B5 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_B6 = 1'b1;
  assign LIOI3_X0Y151_OLOGIC_X0Y151_T1 = 1'b1;
  assign RIOI3_X105Y195_OLOGIC_X1Y195_D1 = CLBLM_R_X13Y143_SLICE_X18Y143_BQ;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_C1 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_C2 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_C3 = CLBLL_L_X4Y139_SLICE_X4Y139_BO6;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_C4 = CLBLM_R_X5Y136_SLICE_X7Y136_DO5;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_C5 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_C6 = 1'b1;
  assign RIOI3_X105Y195_OLOGIC_X1Y195_T1 = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_T1 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_D1 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_D2 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_D3 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_D4 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_B2 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_D5 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_D6 = 1'b1;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_D3 = CLBLL_L_X4Y142_SLICE_X5Y142_DO6;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_B3 = CLBLM_R_X5Y132_SLICE_X7Y132_AQ;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_D4 = CLBLM_R_X11Y137_SLICE_X14Y137_CO6;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_D5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_D6 = CLBLM_L_X12Y135_SLICE_X17Y135_BO5;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_D1 = CLBLM_R_X37Y138_SLICE_X56Y138_AO6;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_B5 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_A2 = CLBLM_L_X8Y141_SLICE_X11Y141_BQ;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_A3 = CLBLM_L_X8Y141_SLICE_X11Y141_AQ;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_A4 = CLBLM_L_X10Y141_SLICE_X13Y141_DO6;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_A5 = CLBLM_R_X7Y138_SLICE_X8Y138_BQ;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_A6 = CLBLM_L_X8Y143_SLICE_X10Y143_DO5;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_T1 = 1'b1;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_A1 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_A2 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_A3 = 1'b1;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_B5 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_B6 = CLBLL_L_X4Y137_SLICE_X4Y137_CQ;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_A4 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_A5 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_A6 = 1'b1;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_B2 = CLBLM_L_X8Y141_SLICE_X11Y141_BQ;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_B3 = CLBLM_R_X13Y141_SLICE_X19Y141_BQ;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_C4 = CLBLM_R_X11Y136_SLICE_X14Y136_DQ;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_C5 = CLBLM_L_X8Y142_SLICE_X11Y142_DQ;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_B1 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_B2 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_B3 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_B4 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_B5 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_B6 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_C1 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_C2 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_C3 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_C4 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_C5 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_C6 = 1'b1;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_D1 = CLBLM_R_X5Y139_SLICE_X7Y139_AQ;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_D2 = CLBLM_R_X11Y139_SLICE_X14Y139_AQ;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_D3 = CLBLL_L_X4Y142_SLICE_X5Y142_DO6;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_D4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_D5 = CLBLM_R_X11Y138_SLICE_X14Y138_DQ;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_D6 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_D1 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_D2 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_D3 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_D4 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_D5 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_D6 = 1'b1;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_A1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_A2 = CLBLM_L_X8Y141_SLICE_X10Y141_BQ;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_A3 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_A5 = CLBLM_L_X8Y138_SLICE_X10Y138_AQ;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_A6 = CLBLM_L_X8Y134_SLICE_X10Y134_CO6;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_B1 = CLBLM_L_X8Y143_SLICE_X10Y143_DO6;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_B2 = CLBLM_L_X8Y141_SLICE_X10Y141_BQ;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_B3 = CLBLM_L_X10Y140_SLICE_X13Y140_BQ;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_B4 = 1'b1;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_B5 = CLBLM_R_X5Y140_SLICE_X7Y140_AQ;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_C1 = 1'b1;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_C2 = CLBLM_L_X8Y141_SLICE_X10Y141_CQ;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_C3 = 1'b1;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_C5 = CLBLM_L_X8Y142_SLICE_X10Y142_CQ;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_D1 = CLBLM_R_X11Y141_SLICE_X15Y141_DQ;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_D2 = CLBLM_L_X10Y142_SLICE_X12Y142_DQ;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_D3 = 1'b1;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_D4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_D5 = 1'b1;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_D6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_A1 = 1'b1;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_A2 = 1'b1;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_A3 = 1'b1;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_A4 = 1'b1;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_A5 = 1'b1;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_A6 = 1'b1;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_B1 = 1'b1;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_B2 = 1'b1;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_B3 = 1'b1;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_B4 = 1'b1;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_B5 = 1'b1;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_B6 = 1'b1;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_A1 = CLBLL_L_X4Y135_SLICE_X5Y135_BQ;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_A2 = CLBLM_L_X8Y133_SLICE_X10Y133_CQ;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_A3 = CLBLM_R_X7Y135_SLICE_X9Y135_AQ;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_A4 = 1'b1;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_A6 = CLBLM_L_X8Y143_SLICE_X10Y143_DO5;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_C1 = 1'b1;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_C2 = 1'b1;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_AX = CLBLM_L_X8Y134_SLICE_X10Y134_BO5;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_C3 = 1'b1;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_B1 = 1'b1;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_B2 = CLBLM_R_X7Y135_SLICE_X9Y135_BQ;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_B4 = CLBLM_L_X8Y135_SLICE_X11Y135_CQ;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_B5 = CLBLM_L_X8Y136_SLICE_X11Y136_AQ;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_B6 = CLBLM_L_X8Y143_SLICE_X10Y143_DO5;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_D1 = 1'b1;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_BX = CLBLM_R_X7Y136_SLICE_X9Y136_BO6;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_D2 = 1'b1;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_C1 = CLBLM_L_X8Y135_SLICE_X10Y135_AQ;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_C2 = CLBLM_R_X11Y136_SLICE_X15Y136_BQ;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_C3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_C4 = CLBLM_R_X5Y135_SLICE_X6Y135_CQ;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_C5 = CLBLM_L_X8Y135_SLICE_X11Y135_A5Q;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_C6 = 1'b1;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_D4 = 1'b1;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_A1 = CLBLM_R_X11Y144_SLICE_X14Y144_AQ;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_A2 = CLBLM_L_X8Y142_SLICE_X10Y142_D5Q;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_A3 = CLBLM_L_X10Y142_SLICE_X12Y142_CQ;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_A4 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_A5 = CLBLM_L_X10Y141_SLICE_X12Y141_C5Q;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_D1 = CLBLM_R_X7Y132_SLICE_X8Y132_BQ;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_D2 = CLBLM_L_X10Y138_SLICE_X12Y138_BO5;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_D3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_D4 = CLBLM_R_X5Y137_SLICE_X7Y137_CQ;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_D5 = CLBLM_R_X5Y136_SLICE_X7Y136_BQ;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_D6 = 1'b1;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_A6 = 1'b1;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_B1 = 1'b1;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_B2 = 1'b1;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_B3 = 1'b1;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_B4 = 1'b1;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_A1 = 1'b1;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_A2 = CLBLM_L_X10Y137_SLICE_X13Y137_CO6;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_A5 = CLBLM_R_X5Y135_SLICE_X7Y135_AQ;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_A6 = CLBLM_L_X8Y136_SLICE_X11Y136_CQ;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_C1 = 1'b1;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_C2 = 1'b1;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_C3 = 1'b1;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_B1 = CLBLM_L_X10Y135_SLICE_X12Y135_B5Q;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_B2 = CLBLM_R_X7Y135_SLICE_X8Y135_BQ;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_B4 = CLBLM_R_X11Y139_SLICE_X15Y139_A5Q;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_B5 = CLBLM_R_X7Y136_SLICE_X8Y136_AQ;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_D1 = 1'b1;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_D2 = 1'b1;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_D3 = 1'b1;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_C2 = 1'b1;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_C3 = CLBLM_L_X10Y135_SLICE_X12Y135_B5Q;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_C5 = CLBLL_L_X4Y136_SLICE_X4Y136_DQ;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_C6 = 1'b1;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_D4 = 1'b1;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_D5 = 1'b1;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_D6 = 1'b1;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_D2 = CLBLM_R_X11Y139_SLICE_X15Y139_A5Q;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_D3 = CLBLM_L_X10Y135_SLICE_X12Y135_B5Q;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_D4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_D5 = 1'b1;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_D6 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_A2 = CLBLM_R_X11Y141_SLICE_X15Y141_CQ;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_A3 = CLBLM_L_X8Y142_SLICE_X11Y142_AQ;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_A4 = CLBLM_R_X5Y139_SLICE_X7Y139_AQ;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_A5 = CLBLM_L_X12Y135_SLICE_X17Y135_AQ;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_A6 = CLBLL_L_X4Y137_SLICE_X4Y137_CQ;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_D = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_B1 = CLBLM_L_X10Y145_SLICE_X13Y145_BO6;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_B2 = CLBLM_L_X8Y142_SLICE_X11Y142_BQ;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_B4 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_B5 = CLBLM_R_X7Y133_SLICE_X8Y133_BQ;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_B6 = CLBLM_L_X8Y143_SLICE_X11Y143_CO6;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_C1 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_C2 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_C3 = CLBLM_L_X10Y144_SLICE_X12Y144_AO5;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_C5 = CLBLM_L_X12Y140_SLICE_X17Y140_CQ;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_C6 = CLBLM_R_X7Y142_SLICE_X9Y142_AQ;
  assign LIOI3_X0Y103_OLOGIC_X0Y104_T1 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_D1 = CLBLM_L_X10Y134_SLICE_X12Y134_AQ;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_D2 = CLBLM_R_X7Y141_SLICE_X8Y141_CO6;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_D3 = CLBLM_R_X7Y139_SLICE_X9Y139_CO6;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_D4 = CLBLM_L_X10Y145_SLICE_X13Y145_BO6;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_D6 = CLBLM_L_X8Y143_SLICE_X11Y143_BO6;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_A2 = CLBLM_R_X11Y142_SLICE_X14Y142_AQ;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_A3 = CLBLM_L_X8Y142_SLICE_X10Y142_AQ;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_A4 = CLBLM_R_X7Y140_SLICE_X9Y140_BQ;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_A5 = CLBLM_L_X12Y135_SLICE_X17Y135_AQ;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_A6 = CLBLL_L_X4Y137_SLICE_X4Y137_CQ;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_B1 = CLBLM_R_X11Y144_SLICE_X14Y144_AQ;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_B2 = CLBLL_L_X4Y135_SLICE_X4Y135_A5Q;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_B3 = CLBLM_L_X10Y142_SLICE_X12Y142_CQ;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_B4 = CLBLM_L_X8Y142_SLICE_X10Y142_D5Q;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_B6 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_C1 = CLBLM_L_X8Y142_SLICE_X10Y142_CQ;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_C2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_C3 = CLBLM_L_X8Y143_SLICE_X10Y143_DO5;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_C4 = CLBLM_L_X8Y139_SLICE_X10Y139_BQ;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_C5 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_C6 = CLBLM_L_X8Y142_SLICE_X10Y142_D5Q;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_D1 = RIOB33_X105Y125_IOB_X1Y126_I;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_C3 = CLBLL_L_X4Y143_SLICE_X5Y143_BO5;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_D1 = CLBLM_L_X8Y143_SLICE_X11Y143_AO6;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_D2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_D3 = CLBLM_R_X7Y140_SLICE_X9Y140_BQ;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_D4 = CLBLM_R_X7Y140_SLICE_X8Y140_DO6;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_C4 = CLBLL_L_X2Y141_SLICE_X1Y141_AO5;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_D5 = CLBLM_R_X5Y141_SLICE_X7Y141_BQ;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_D6 = 1'b1;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_C5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_C6 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_A1 = 1'b1;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_A2 = 1'b1;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_A3 = 1'b1;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_A4 = 1'b1;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_A5 = 1'b1;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_A6 = 1'b1;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_B1 = 1'b1;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_B2 = 1'b1;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_B3 = 1'b1;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_B4 = 1'b1;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_B5 = 1'b1;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_B6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_T1 = 1'b1;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_A1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_A2 = CLBLM_R_X7Y136_SLICE_X8Y136_DO6;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_A3 = CLBLM_R_X7Y136_SLICE_X9Y136_AQ;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_A4 = CLBLM_L_X8Y138_SLICE_X10Y138_AQ;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_A6 = CLBLM_R_X5Y138_SLICE_X6Y138_CQ;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_C1 = 1'b1;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_C2 = 1'b1;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_C3 = 1'b1;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_B1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_D2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_B3 = CLBLM_R_X7Y132_SLICE_X9Y132_AQ;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_B4 = CLBLL_L_X4Y136_SLICE_X5Y136_A5Q;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_B5 = CLBLM_R_X11Y136_SLICE_X15Y136_AQ;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_D3 = CLBLM_R_X5Y134_SLICE_X6Y134_A5Q;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_B6 = 1'b1;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_C1 = CLBLM_R_X7Y138_SLICE_X9Y138_AQ;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_D4 = CLBLL_L_X2Y141_SLICE_X1Y141_AO5;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_C2 = CLBLM_R_X7Y136_SLICE_X9Y136_CQ;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_C3 = CLBLM_R_X7Y139_SLICE_X9Y139_AQ;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_C5 = 1'b1;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_D5 = 1'b1;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_C6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_A1 = 1'b1;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_A2 = 1'b1;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_D6 = CLBLL_L_X4Y143_SLICE_X5Y143_BO6;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_A3 = 1'b1;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_A4 = 1'b1;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_D1 = CLBLM_L_X8Y138_SLICE_X11Y138_AQ;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_D2 = CLBLM_R_X7Y135_SLICE_X8Y135_AQ;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_D3 = 1'b1;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_D4 = CLBLM_R_X7Y135_SLICE_X8Y135_CQ;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_D5 = 1'b1;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_D6 = CLBLM_R_X7Y135_SLICE_X9Y135_A5Q;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_A5 = 1'b1;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_A6 = 1'b1;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_AX = CLBLM_L_X12Y146_SLICE_X16Y146_AO5;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_B1 = 1'b1;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_B2 = 1'b1;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_B3 = 1'b1;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_A1 = CLBLM_L_X12Y134_SLICE_X17Y134_AQ;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_A2 = CLBLM_R_X11Y146_SLICE_X14Y146_AQ;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_A5 = CLBLM_R_X5Y136_SLICE_X6Y136_CQ;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_A6 = CLBLM_R_X7Y134_SLICE_X8Y134_CQ;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_C1 = 1'b1;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_C2 = 1'b1;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_C3 = 1'b1;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_B1 = CLBLL_L_X4Y137_SLICE_X4Y137_CQ;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_B2 = CLBLM_R_X7Y136_SLICE_X8Y136_BQ;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_B4 = CLBLM_L_X10Y136_SLICE_X12Y136_A5Q;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_B5 = CLBLM_R_X11Y136_SLICE_X14Y136_AQ;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_B6 = CLBLM_L_X12Y135_SLICE_X17Y135_AQ;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_D1 = 1'b1;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_D2 = 1'b1;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_C1 = CLBLM_L_X8Y138_SLICE_X11Y138_AQ;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_C2 = CLBLM_R_X7Y136_SLICE_X8Y136_CQ;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_C4 = CLBLM_L_X12Y136_SLICE_X16Y136_BQ;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_C5 = 1'b1;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_C6 = CLBLM_R_X7Y144_SLICE_X9Y144_BO6;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_D3 = 1'b1;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_D4 = 1'b1;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_D5 = 1'b1;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_D6 = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_D1 = CLBLM_R_X3Y136_SLICE_X3Y136_BQ;
  assign LIOI3_SING_X0Y100_OLOGIC_X0Y100_T1 = 1'b1;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_D1 = CLBLL_L_X4Y134_SLICE_X4Y134_AQ;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_D2 = CLBLM_L_X10Y134_SLICE_X12Y134_CQ;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_D3 = CLBLM_R_X5Y142_SLICE_X6Y142_CO6;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_D4 = CLBLM_R_X7Y135_SLICE_X9Y135_CO6;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_D5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_D6 = 1'b1;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_A1 = CLBLM_L_X8Y144_SLICE_X11Y144_BO5;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_A2 = CLBLM_R_X11Y143_SLICE_X14Y143_DO6;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_A3 = CLBLM_R_X11Y144_SLICE_X14Y144_AQ;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_A4 = CLBLM_L_X8Y142_SLICE_X10Y142_D5Q;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_A5 = CLBLM_L_X10Y141_SLICE_X12Y141_C5Q;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_A6 = CLBLM_R_X7Y143_SLICE_X8Y143_BO5;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_B1 = CLBLM_L_X8Y144_SLICE_X11Y144_BO5;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_B2 = CLBLM_L_X8Y142_SLICE_X11Y142_DQ;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_B3 = CLBLM_L_X10Y142_SLICE_X12Y142_CQ;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_B4 = CLBLM_L_X8Y142_SLICE_X10Y142_D5Q;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_B5 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_B6 = CLBLM_R_X11Y144_SLICE_X14Y144_AQ;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_C1 = 1'b1;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_C2 = CLBLM_R_X7Y144_SLICE_X8Y144_BQ;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_C3 = CLBLM_R_X7Y144_SLICE_X8Y144_AQ;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_C4 = CLBLM_R_X7Y143_SLICE_X9Y143_BQ;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_C5 = 1'b1;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_C6 = 1'b1;
  assign LIOI3_X0Y153_OLOGIC_X0Y154_D1 = LIOB33_X0Y67_IOB_X0Y68_I;
  assign RIOI3_X105Y179_OLOGIC_X1Y179_T1 = 1'b1;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_D1 = 1'b1;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_D2 = 1'b1;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_D3 = 1'b1;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_D4 = 1'b1;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_D5 = 1'b1;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_D6 = 1'b1;
  assign LIOI3_X0Y153_OLOGIC_X0Y154_T1 = 1'b1;
  assign RIOI3_X105Y197_OLOGIC_X1Y198_D1 = CLBLM_R_X103Y175_SLICE_X163Y175_AO6;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_A2 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_A3 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_A4 = CLBLM_L_X10Y142_SLICE_X12Y142_CQ;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_A5 = CLBLM_R_X3Y137_SLICE_X2Y137_AQ;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_A6 = CLBLM_R_X11Y143_SLICE_X14Y143_DO6;
  assign LIOI3_X0Y153_OLOGIC_X0Y153_D1 = LIOB33_X0Y67_IOB_X0Y67_I;
  assign RIOI3_X105Y197_OLOGIC_X1Y198_T1 = 1'b1;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_B1 = CLBLM_L_X8Y140_SLICE_X10Y140_DQ;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_B2 = CLBLM_L_X8Y143_SLICE_X10Y143_BQ;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_B4 = CLBLM_L_X8Y143_SLICE_X10Y143_DO5;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_B5 = 1'b1;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_B6 = CLBLM_L_X8Y141_SLICE_X10Y141_DQ;
  assign LIOI3_X0Y153_OLOGIC_X0Y153_T1 = 1'b1;
  assign RIOI3_X105Y197_OLOGIC_X1Y197_D1 = CLBLM_R_X103Y175_SLICE_X163Y175_AO6;
  assign CLBLM_R_X37Y138_SLICE_X56Y138_B4 = 1'b1;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_C1 = CLBLL_L_X4Y133_SLICE_X5Y133_BO6;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_C2 = CLBLM_L_X8Y143_SLICE_X10Y143_CQ;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_C3 = 1'b1;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_C5 = CLBLM_R_X11Y143_SLICE_X14Y143_AQ;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_C6 = CLBLL_L_X4Y137_SLICE_X4Y137_A5Q;
  assign RIOI3_X105Y197_OLOGIC_X1Y197_T1 = 1'b1;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_D1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_D2 = CLBLM_R_X11Y136_SLICE_X14Y136_DQ;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_D3 = CLBLM_R_X11Y141_SLICE_X15Y141_AQ;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_D4 = CLBLM_R_X7Y144_SLICE_X8Y144_CQ;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_D5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_D6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_D1 = CLBLM_R_X103Y170_SLICE_X163Y170_AO6;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_C4 = CLBLM_L_X12Y140_SLICE_X17Y140_BQ;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_C5 = CLBLM_L_X12Y143_SLICE_X17Y143_CO5;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_T1 = 1'b1;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_D1 = CLBLM_R_X103Y169_SLICE_X163Y169_AO6;
  assign LIOB33_X0Y143_IOB_X0Y143_O = LIOB33_X0Y55_IOB_X0Y55_I;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_A3 = CLBLM_L_X12Y142_SLICE_X16Y142_A5Q;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_T1 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_A1 = CLBLM_L_X10Y139_SLICE_X12Y139_AQ;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_A3 = CLBLM_R_X7Y137_SLICE_X9Y137_AQ;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_A4 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_A6 = CLBLM_R_X7Y137_SLICE_X9Y137_CO6;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_B1 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_B4 = CLBLM_L_X10Y137_SLICE_X13Y137_BQ;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_B5 = CLBLM_L_X8Y138_SLICE_X11Y138_AQ;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_B6 = CLBLM_L_X10Y138_SLICE_X13Y138_DO6;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_C1 = CLBLL_L_X4Y136_SLICE_X4Y136_DQ;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_A4 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_C2 = CLBLM_R_X7Y136_SLICE_X9Y136_DO6;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_C3 = CLBLM_L_X12Y139_SLICE_X16Y139_A5Q;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_D1 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_C4 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_C5 = CLBLM_R_X7Y137_SLICE_X9Y137_DO6;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_C6 = CLBLM_L_X8Y140_SLICE_X11Y140_DO6;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_D2 = CLBLM_R_X13Y144_SLICE_X18Y144_CO6;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_D3 = CLBLM_R_X13Y141_SLICE_X18Y141_BO5;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_D1 = CLBLM_L_X10Y137_SLICE_X13Y137_AQ;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_D2 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_D3 = CLBLL_L_X4Y135_SLICE_X5Y135_BQ;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_D4 = CLBLM_R_X7Y137_SLICE_X9Y137_BQ;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_D5 = CLBLM_L_X8Y139_SLICE_X10Y139_BQ;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_D6 = CLBLM_R_X7Y133_SLICE_X8Y133_BQ;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_A5 = CLBLM_L_X12Y144_SLICE_X16Y144_AQ;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_A6 = CLBLM_L_X10Y145_SLICE_X13Y145_BO6;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_A1 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_A2 = CLBLM_L_X8Y136_SLICE_X10Y136_BQ;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_A3 = CLBLM_R_X7Y137_SLICE_X8Y137_AQ;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_A4 = CLBLM_R_X7Y133_SLICE_X8Y133_BQ;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_A6 = CLBLM_R_X7Y144_SLICE_X9Y144_BO6;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_B1 = CLBLM_R_X7Y138_SLICE_X8Y138_CQ;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_B2 = CLBLM_R_X7Y137_SLICE_X8Y137_BQ;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_B4 = CLBLM_L_X10Y141_SLICE_X13Y141_A5Q;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_B5 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_B6 = CLBLM_L_X8Y143_SLICE_X10Y143_DO5;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_C1 = CLBLM_L_X12Y136_SLICE_X16Y136_C5Q;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_A6 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_C2 = CLBLM_R_X7Y137_SLICE_X8Y137_CQ;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_B1 = CLBLM_L_X10Y145_SLICE_X13Y145_BO6;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_C3 = CLBLL_L_X4Y137_SLICE_X5Y137_AO5;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_C5 = CLBLM_R_X7Y140_SLICE_X9Y140_BQ;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_C6 = CLBLM_R_X11Y135_SLICE_X14Y135_AQ;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_B2 = CLBLM_L_X10Y142_SLICE_X13Y142_BQ;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_D = RIOB33_X105Y107_IOB_X1Y107_I;
  assign LIOB33_X0Y197_IOB_X0Y198_O = LIOB33_X0Y73_IOB_X0Y73_I;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_D1 = CLBLM_R_X3Y138_SLICE_X3Y138_AQ;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_D2 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_B4 = CLBLM_L_X8Y144_SLICE_X11Y144_CO6;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_D3 = CLBLM_R_X7Y143_SLICE_X8Y143_A5Q;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_D4 = CLBLL_L_X4Y136_SLICE_X5Y136_CQ;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_D5 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_D6 = CLBLM_R_X7Y133_SLICE_X8Y133_CQ;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_B5 = CLBLM_L_X10Y142_SLICE_X12Y142_AQ;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_B6 = CLBLM_L_X10Y133_SLICE_X12Y133_CQ;
  assign RIOB33_X105Y179_IOB_X1Y180_O = CLBLM_L_X12Y138_SLICE_X17Y138_DO6;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_D1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign RIOB33_X105Y179_IOB_X1Y179_O = CLBLM_L_X12Y144_SLICE_X17Y144_AO5;
  assign RIOI3_X105Y135_ILOGIC_X1Y136_D = RIOB33_X105Y135_IOB_X1Y136_I;
  assign RIOI3_X105Y135_ILOGIC_X1Y135_D = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_T1 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_C2 = CLBLM_L_X8Y138_SLICE_X10Y138_BQ;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_A3 = CLBLM_R_X3Y133_SLICE_X2Y133_BO6;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_C3 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_A4 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_C4 = CLBLM_R_X11Y144_SLICE_X14Y144_DO6;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_A5 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_C5 = CLBLM_L_X10Y142_SLICE_X13Y142_DO6;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_A6 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_C6 = CLBLM_L_X10Y144_SLICE_X12Y144_AO6;
  assign LIOI3_X0Y103_OLOGIC_X0Y103_T1 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_A1 = CLBLM_L_X8Y144_SLICE_X11Y144_AQ;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_B6 = CLBLM_L_X12Y143_SLICE_X17Y143_CO5;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_A5 = CLBLM_R_X7Y143_SLICE_X9Y143_BQ;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_A6 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_B1 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_A2 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_A3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_B1 = CLBLM_R_X7Y144_SLICE_X8Y144_BQ;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_B2 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_B2 = CLBLM_L_X10Y145_SLICE_X13Y145_BO6;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_B3 = CLBLM_R_X7Y143_SLICE_X9Y143_BQ;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_B4 = CLBLM_R_X7Y144_SLICE_X8Y144_AQ;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_B6 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_B3 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_B5 = CLBLM_L_X8Y142_SLICE_X11Y142_BQ;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_C1 = CLBLM_R_X7Y143_SLICE_X9Y143_BQ;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_B4 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_C2 = CLBLM_R_X7Y144_SLICE_X8Y144_AQ;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_C3 = CLBLM_L_X10Y141_SLICE_X12Y141_C5Q;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_C4 = CLBLM_R_X7Y144_SLICE_X8Y144_BQ;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_C5 = CLBLM_L_X8Y142_SLICE_X10Y142_D5Q;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_B5 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_C6 = CLBLM_L_X8Y142_SLICE_X11Y142_BQ;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_B6 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_D1 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_D2 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_D3 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_D4 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_D5 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_D6 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_D2 = CLBLM_L_X10Y142_SLICE_X13Y142_CQ;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_D3 = CLBLM_L_X10Y144_SLICE_X13Y144_DO6;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_D4 = CLBLM_L_X10Y144_SLICE_X13Y144_CO6;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_C4 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_A1 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_A2 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_A3 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_A4 = 1'b1;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_C5 = CLBLM_R_X13Y141_SLICE_X18Y141_AO6;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_B1 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_A5 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_A6 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_C1 = 1'b1;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_B1 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_B2 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_B3 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_C2 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_B5 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_B4 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_B6 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_C1 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_C2 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_C3 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_C4 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_C5 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_C6 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_C5 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_B2 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_C6 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_D1 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_D2 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_D3 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_D4 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_D5 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_D6 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_B3 = 1'b1;
  assign LIOB33_X0Y145_IOB_X0Y145_O = LIOB33_X0Y57_IOB_X0Y58_I;
  assign LIOB33_X0Y145_IOB_X0Y146_O = LIOB33_X0Y59_IOB_X0Y59_I;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_A3 = CLBLM_L_X10Y142_SLICE_X12Y142_AQ;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_A4 = CLBLM_L_X10Y143_SLICE_X12Y143_BQ;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_B4 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_D1 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_D2 = 1'b1;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_A1 = CLBLM_L_X8Y138_SLICE_X10Y138_CQ;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_A2 = 1'b1;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_A4 = CLBLM_L_X8Y138_SLICE_X11Y138_CO5;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_A6 = CLBLM_R_X11Y138_SLICE_X14Y138_DQ;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_D5 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_B5 = 1'b1;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_B1 = CLBLM_R_X7Y138_SLICE_X9Y138_DO6;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_D6 = 1'b1;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_B2 = CLBLM_R_X7Y134_SLICE_X8Y134_AQ;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_B3 = CLBLL_L_X4Y138_SLICE_X5Y138_BQ;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_B4 = CLBLM_L_X10Y134_SLICE_X13Y134_BQ;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_B5 = CLBLM_R_X11Y137_SLICE_X14Y137_AQ;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_B6 = CLBLM_L_X8Y140_SLICE_X11Y140_CO6;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_B4 = CLBLM_L_X8Y144_SLICE_X11Y144_CO6;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_C1 = CLBLM_L_X8Y138_SLICE_X10Y138_AQ;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_C2 = CLBLM_R_X7Y137_SLICE_X8Y137_CQ;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_C3 = CLBLM_R_X7Y140_SLICE_X9Y140_BQ;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_C4 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_B5 = CLBLM_L_X10Y142_SLICE_X13Y142_AQ;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_C5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_C6 = 1'b1;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_B6 = CLBLM_L_X8Y140_SLICE_X11Y140_A5Q;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_D1 = CLBLM_R_X7Y134_SLICE_X9Y134_AQ;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_D2 = 1'b1;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_D3 = CLBLM_L_X8Y140_SLICE_X10Y140_DQ;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_D4 = CLBLM_R_X5Y138_SLICE_X6Y138_CQ;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_D5 = 1'b1;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_D6 = CLBLM_R_X7Y138_SLICE_X9Y138_AQ;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_A1 = CLBLM_R_X7Y138_SLICE_X8Y138_DO6;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_A2 = CLBLM_R_X7Y138_SLICE_X9Y138_BO6;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_A3 = CLBLM_R_X7Y138_SLICE_X8Y138_AQ;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_A6 = CLBLM_L_X12Y138_SLICE_X16Y138_BQ;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_B1 = CLBLM_R_X7Y136_SLICE_X9Y136_BO5;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_B2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_B4 = CLBLM_R_X11Y139_SLICE_X15Y139_A5Q;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_B5 = 1'b1;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_B6 = CLBLM_R_X5Y138_SLICE_X6Y138_CQ;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_C2 = CLBLM_R_X5Y139_SLICE_X7Y139_BQ;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_C3 = 1'b1;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_C4 = CLBLM_R_X7Y135_SLICE_X9Y135_CO6;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_C5 = CLBLM_L_X8Y140_SLICE_X10Y140_DQ;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_C4 = CLBLM_L_X8Y133_SLICE_X10Y133_BQ;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_C6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_C5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_C6 = CLBLM_R_X11Y143_SLICE_X14Y143_BO6;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_D1 = CLBLM_L_X8Y136_SLICE_X11Y136_AQ;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_D2 = CLBLM_R_X7Y138_SLICE_X8Y138_CQ;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_D3 = CLBLM_L_X8Y138_SLICE_X10Y138_CQ;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_D4 = CLBLM_R_X5Y139_SLICE_X7Y139_BQ;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_D5 = CLBLM_R_X7Y138_SLICE_X8Y138_BQ;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_D6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign LIOI3_SING_X0Y150_OLOGIC_X0Y150_D1 = LIOB33_X0Y63_IOB_X0Y63_I;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_A1 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_A2 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_A3 = 1'b1;
  assign LIOI3_SING_X0Y150_OLOGIC_X0Y150_T1 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_A4 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_A5 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_A6 = 1'b1;
endmodule
