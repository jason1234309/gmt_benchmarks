module top(
  input LIOB33_SING_X0Y100_IOB_X0Y100_IPAD,
  input LIOB33_X0Y101_IOB_X0Y101_IPAD,
  input LIOB33_X0Y101_IOB_X0Y102_IPAD,
  input LIOB33_X0Y103_IOB_X0Y103_IPAD,
  input LIOB33_X0Y103_IOB_X0Y104_IPAD,
  input LIOB33_X0Y105_IOB_X0Y105_IPAD,
  input LIOB33_X0Y105_IOB_X0Y106_IPAD,
  input LIOB33_X0Y107_IOB_X0Y107_IPAD,
  input LIOB33_X0Y107_IOB_X0Y108_IPAD,
  input LIOB33_X0Y109_IOB_X0Y109_IPAD,
  input LIOB33_X0Y109_IOB_X0Y110_IPAD,
  input LIOB33_X0Y111_IOB_X0Y111_IPAD,
  input LIOB33_X0Y111_IOB_X0Y112_IPAD,
  input LIOB33_X0Y113_IOB_X0Y113_IPAD,
  input LIOB33_X0Y113_IOB_X0Y114_IPAD,
  input LIOB33_X0Y115_IOB_X0Y115_IPAD,
  input LIOB33_X0Y115_IOB_X0Y116_IPAD,
  input LIOB33_X0Y117_IOB_X0Y117_IPAD,
  input RIOB33_SING_X105Y100_IOB_X1Y100_IPAD,
  input RIOB33_X105Y101_IOB_X1Y101_IPAD,
  input RIOB33_X105Y101_IOB_X1Y102_IPAD,
  input RIOB33_X105Y103_IOB_X1Y103_IPAD,
  input RIOB33_X105Y103_IOB_X1Y104_IPAD,
  input RIOB33_X105Y105_IOB_X1Y105_IPAD,
  input RIOB33_X105Y105_IOB_X1Y106_IPAD,
  input RIOB33_X105Y107_IOB_X1Y107_IPAD,
  input RIOB33_X105Y107_IOB_X1Y108_IPAD,
  input RIOB33_X105Y109_IOB_X1Y109_IPAD,
  input RIOB33_X105Y109_IOB_X1Y110_IPAD,
  input RIOB33_X105Y111_IOB_X1Y111_IPAD,
  input RIOB33_X105Y111_IOB_X1Y112_IPAD,
  input RIOB33_X105Y113_IOB_X1Y113_IPAD,
  output LIOB33_SING_X0Y149_IOB_X0Y149_OPAD,
  output LIOB33_X0Y117_IOB_X0Y118_OPAD,
  output LIOB33_X0Y119_IOB_X0Y119_OPAD,
  output LIOB33_X0Y119_IOB_X0Y120_OPAD,
  output LIOB33_X0Y121_IOB_X0Y121_OPAD,
  output LIOB33_X0Y121_IOB_X0Y122_OPAD,
  output LIOB33_X0Y123_IOB_X0Y123_OPAD,
  output LIOB33_X0Y123_IOB_X0Y124_OPAD,
  output LIOB33_X0Y125_IOB_X0Y125_OPAD,
  output LIOB33_X0Y125_IOB_X0Y126_OPAD,
  output LIOB33_X0Y127_IOB_X0Y127_OPAD,
  output LIOB33_X0Y127_IOB_X0Y128_OPAD,
  output LIOB33_X0Y129_IOB_X0Y129_OPAD,
  output LIOB33_X0Y129_IOB_X0Y130_OPAD,
  output LIOB33_X0Y131_IOB_X0Y131_OPAD,
  output LIOB33_X0Y131_IOB_X0Y132_OPAD,
  output LIOB33_X0Y133_IOB_X0Y133_OPAD,
  output LIOB33_X0Y133_IOB_X0Y134_OPAD,
  output LIOB33_X0Y135_IOB_X0Y135_OPAD,
  output LIOB33_X0Y135_IOB_X0Y136_OPAD,
  output LIOB33_X0Y137_IOB_X0Y137_OPAD,
  output LIOB33_X0Y137_IOB_X0Y138_OPAD,
  output LIOB33_X0Y139_IOB_X0Y139_OPAD,
  output LIOB33_X0Y139_IOB_X0Y140_OPAD,
  output LIOB33_X0Y141_IOB_X0Y141_OPAD,
  output LIOB33_X0Y141_IOB_X0Y142_OPAD,
  output LIOB33_X0Y143_IOB_X0Y143_OPAD,
  output LIOB33_X0Y145_IOB_X0Y145_OPAD,
  output LIOB33_X0Y145_IOB_X0Y146_OPAD,
  output LIOB33_X0Y147_IOB_X0Y147_OPAD,
  output LIOB33_X0Y147_IOB_X0Y148_OPAD
  );
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_A;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_A1;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_A2;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_A3;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_A4;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_A5;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_A6;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_AO5;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_AO6;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_A_CY;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_A_XOR;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_B;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_B1;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_B2;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_B3;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_B4;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_B5;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_B6;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_BO5;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_BO6;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_B_CY;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_B_XOR;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_C;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_C1;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_C2;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_C3;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_C4;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_C5;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_C6;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_CO5;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_CO6;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_C_CY;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_C_XOR;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_D;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_D1;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_D2;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_D3;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_D4;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_D5;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_D6;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_DO5;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_DO6;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_D_CY;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X0Y102_D_XOR;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_A;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_A1;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_A2;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_A3;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_A4;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_A5;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_A6;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_AO5;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_AO6;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_A_CY;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_A_XOR;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_B;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_B1;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_B2;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_B3;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_B4;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_B5;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_B6;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_BO5;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_BO6;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_B_CY;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_B_XOR;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_C;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_C1;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_C2;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_C3;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_C4;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_C5;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_C6;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_CO5;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_CO6;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_C_CY;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_C_XOR;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_D;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_D1;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_D2;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_D3;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_D4;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_D5;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_D6;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_DO5;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_DO6;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_D_CY;
  wire [0:0] CLBLL_L_X2Y102_SLICE_X1Y102_D_XOR;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_A;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_A1;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_A2;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_A3;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_A4;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_A5;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_A6;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_AO5;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_AO6;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_A_CY;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_A_XOR;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_B;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_B1;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_B2;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_B3;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_B4;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_B5;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_B6;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_BO5;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_BO6;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_B_CY;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_B_XOR;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_C;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_C1;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_C2;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_C3;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_C4;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_C5;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_C6;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_CO5;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_CO6;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_C_CY;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_C_XOR;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_D;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_D1;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_D2;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_D3;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_D4;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_D5;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_D6;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_DO5;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_DO6;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_D_CY;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_D_XOR;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_A;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_A1;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_A2;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_A3;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_A4;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_A5;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_A6;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_AMUX;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_AO5;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_AO6;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_A_CY;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_A_XOR;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_B;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_B1;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_B2;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_B3;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_B4;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_B5;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_B6;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_BO5;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_BO6;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_B_CY;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_B_XOR;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_C;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_C1;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_C2;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_C3;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_C4;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_C5;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_C6;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_CO5;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_CO6;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_C_CY;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_C_XOR;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_D;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_D1;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_D2;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_D3;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_D4;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_D5;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_D6;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_DO5;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_DO6;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_D_CY;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_D_XOR;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_A;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_A1;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_A2;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_A3;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_A4;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_A5;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_A6;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_AMUX;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_AO5;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_AO6;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_A_CY;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_A_XOR;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_B;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_B1;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_B2;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_B3;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_B4;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_B5;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_B6;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_BMUX;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_BO5;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_BO6;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_B_CY;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_B_XOR;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_C;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_C1;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_C2;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_C3;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_C4;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_C5;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_C6;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_CO5;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_CO6;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_C_CY;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_C_XOR;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_D;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_D1;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_D2;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_D3;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_D4;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_D5;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_D6;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_DMUX;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_DO5;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_DO6;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_D_CY;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_D_XOR;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_A;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_A1;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_A2;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_A3;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_A4;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_A5;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_A6;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_AMUX;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_AO5;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_AO6;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_A_CY;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_A_XOR;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_B;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_B1;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_B2;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_B3;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_B4;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_B5;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_B6;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_BO5;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_BO6;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_B_CY;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_B_XOR;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_C;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_C1;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_C2;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_C3;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_C4;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_C5;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_C6;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_CO5;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_CO6;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_C_CY;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_C_XOR;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_D;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_D1;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_D2;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_D3;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_D4;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_D5;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_D6;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_DO5;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_DO6;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_D_CY;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_D_XOR;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_A;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_A1;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_A2;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_A3;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_A4;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_A5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_A6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_AMUX;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_AO5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_AO6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_A_CY;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_A_XOR;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_B;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_B1;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_B2;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_B3;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_B4;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_B5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_B6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_BMUX;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_BO5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_BO6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_B_CY;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_B_XOR;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_C;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_C1;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_C2;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_C3;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_C4;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_C5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_C6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_CMUX;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_CO5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_CO6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_C_CY;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_C_XOR;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_D;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_D1;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_D2;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_D3;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_D4;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_D5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_D6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_DO5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_DO6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_D_CY;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_D_XOR;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_A;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_A1;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_A2;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_A3;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_A4;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_A5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_A6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_AMUX;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_AO5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_AO6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_A_CY;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_A_XOR;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_B;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_B1;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_B2;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_B3;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_B4;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_B5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_B6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_BO5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_BO6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_B_CY;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_B_XOR;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_C;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_C1;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_C2;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_C3;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_C4;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_C5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_C6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_CO5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_CO6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_C_CY;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_C_XOR;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_D;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_D1;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_D2;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_D3;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_D4;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_D5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_D6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_DO5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_DO6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_D_CY;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_D_XOR;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_A;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_A1;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_A2;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_A3;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_A4;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_A5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_A6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_AO5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_AO6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_A_CY;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_A_XOR;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_B;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_B1;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_B2;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_B3;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_B4;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_B5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_B6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_BO5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_BO6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_B_CY;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_B_XOR;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_C;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_C1;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_C2;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_C3;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_C4;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_C5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_C6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_CO5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_CO6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_C_CY;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_C_XOR;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_D;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_D1;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_D2;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_D3;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_D4;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_D5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_D6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_DO5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_DO6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_D_CY;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_D_XOR;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_A;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_A1;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_A2;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_A3;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_A4;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_A5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_A6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_AMUX;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_AO5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_AO6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_A_CY;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_A_XOR;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_B;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_B1;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_B2;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_B3;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_B4;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_B5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_B6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_BMUX;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_BO5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_BO6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_B_CY;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_B_XOR;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_C;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_C1;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_C2;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_C3;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_C4;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_C5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_C6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_CO5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_CO6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_C_CY;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_C_XOR;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_D;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_D1;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_D2;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_D3;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_D4;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_D5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_D6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_DO5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_DO6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_D_CY;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_D_XOR;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_A;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_A1;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_A2;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_A3;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_A4;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_A5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_A6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_AO5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_AO6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_A_CY;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_A_XOR;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_B;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_B1;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_B2;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_B3;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_B4;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_B5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_B6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_BO5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_BO6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_B_CY;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_B_XOR;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_C;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_C1;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_C2;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_C3;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_C4;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_C5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_C6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_CO5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_CO6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_C_CY;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_C_XOR;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_D;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_D1;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_D2;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_D3;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_D4;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_D5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_D6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_DO5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_DO6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_D_CY;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_D_XOR;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_A;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_A1;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_A2;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_A3;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_A4;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_A5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_A6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_AO5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_AO6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_A_CY;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_A_XOR;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_B;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_B1;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_B2;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_B3;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_B4;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_B5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_B6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_BO5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_BO6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_B_CY;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_B_XOR;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_C;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_C1;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_C2;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_C3;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_C4;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_C5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_C6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_CO5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_CO6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_C_CY;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_C_XOR;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_D;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_D1;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_D2;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_D3;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_D4;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_D5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_D6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_DO5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_DO6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_D_CY;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_D_XOR;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_A;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_A1;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_A2;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_A3;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_A4;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_A5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_A6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_AMUX;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_AO5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_AO6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_A_CY;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_A_XOR;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_B;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_B1;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_B2;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_B3;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_B4;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_B5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_B6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_BO5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_BO6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_B_CY;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_B_XOR;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_C;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_C1;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_C2;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_C3;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_C4;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_C5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_C6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_CO5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_CO6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_C_CY;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_C_XOR;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_D;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_D1;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_D2;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_D3;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_D4;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_D5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_D6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_DO5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_DO6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_D_CY;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_D_XOR;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_A;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_A1;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_A2;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_A3;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_A4;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_A5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_A6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_AO5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_AO6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_A_CY;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_A_XOR;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_B;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_B1;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_B2;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_B3;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_B4;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_B5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_B6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_BO5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_BO6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_B_CY;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_B_XOR;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_C;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_C1;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_C2;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_C3;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_C4;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_C5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_C6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_CO5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_CO6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_C_CY;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_C_XOR;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_D;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_D1;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_D2;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_D3;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_D4;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_D5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_D6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_DO5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_DO6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_D_CY;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_D_XOR;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A1;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A2;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A3;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A4;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_AO5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_AO6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A_CY;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A_XOR;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B1;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B2;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B3;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B4;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_BO5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_BO6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B_CY;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B_XOR;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C1;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C2;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C3;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C4;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_CO5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_CO6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C_CY;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C_XOR;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D1;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D2;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D3;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D4;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_DO5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_DO6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D_CY;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D_XOR;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A1;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A2;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A3;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A4;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_AO5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_AO6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A_CY;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A_XOR;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B1;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B2;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B3;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B4;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_BO5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_BO6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B_CY;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B_XOR;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C1;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C2;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C3;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C4;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_CO5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_CO6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C_CY;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C_XOR;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D1;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D2;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D3;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D4;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_DO5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_DO6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D_CY;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D_XOR;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_A;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_A1;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_A2;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_A3;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_A4;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_A5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_A6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_AO5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_AO6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_A_CY;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_A_XOR;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_B;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_B1;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_B2;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_B3;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_B4;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_B5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_B6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_BO5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_BO6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_B_CY;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_B_XOR;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_C;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_C1;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_C2;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_C3;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_C4;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_C5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_C6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_CO5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_CO6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_C_CY;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_C_XOR;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_D;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_D1;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_D2;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_D3;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_D4;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_D5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_D6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_DO5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_DO6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_D_CY;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_D_XOR;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_A;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_A1;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_A2;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_A3;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_A4;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_A5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_A6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_AO5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_AO6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_A_CY;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_A_XOR;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_B;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_B1;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_B2;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_B3;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_B4;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_B5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_B6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_BO5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_BO6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_B_CY;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_B_XOR;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_C;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_C1;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_C2;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_C3;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_C4;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_C5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_C6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_CO5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_CO6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_C_CY;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_C_XOR;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_D;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_D1;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_D2;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_D3;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_D4;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_D5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_D6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_DO5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_DO6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_D_CY;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_D_XOR;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A1;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A2;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A3;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A4;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_AMUX;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_AO5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_AO6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A_CY;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A_XOR;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B1;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B2;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B3;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B4;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_BMUX;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_BO5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_BO6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B_CY;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B_XOR;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C1;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C2;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C3;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C4;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_CO5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_CO6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C_CY;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C_XOR;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D1;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D2;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D3;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D4;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_DO5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_DO6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D_CY;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D_XOR;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A1;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A2;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A3;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A4;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_AMUX;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_AO5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_AO6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A_CY;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A_XOR;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B1;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B2;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B3;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B4;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_BO5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_BO6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B_CY;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B_XOR;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C1;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C2;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C3;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C4;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_CO5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_CO6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C_CY;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C_XOR;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D1;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D2;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D3;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D4;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_DO5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_DO6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D_CY;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D_XOR;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_A;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_A1;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_A2;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_A3;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_A4;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_A5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_A6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_AMUX;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_AO5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_AO6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_A_CY;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_A_XOR;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_B;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_B1;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_B2;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_B3;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_B4;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_B5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_B6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_BMUX;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_BO5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_BO6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_B_CY;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_B_XOR;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_C;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_C1;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_C2;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_C3;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_C4;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_C5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_C6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_CO5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_CO6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_C_CY;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_C_XOR;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_D;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_D1;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_D2;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_D3;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_D4;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_D5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_D6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_DO5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_DO6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_D_CY;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_D_XOR;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_A;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_A1;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_A2;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_A3;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_A4;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_A5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_A6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_AO5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_AO6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_A_CY;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_A_XOR;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_B;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_B1;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_B2;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_B3;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_B4;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_B5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_B6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_BO5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_BO6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_B_CY;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_B_XOR;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_C;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_C1;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_C2;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_C3;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_C4;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_C5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_C6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_CO5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_CO6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_C_CY;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_C_XOR;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_D;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_D1;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_D2;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_D3;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_D4;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_D5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_D6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_DO5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_DO6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_D_CY;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_D_XOR;
  wire [0:0] CLBLL_L_X4Y100_SLICE_X4Y100_A;
  wire [0:0] CLBLL_L_X4Y100_SLICE_X4Y100_A1;
  wire [0:0] CLBLL_L_X4Y100_SLICE_X4Y100_A2;
  wire [0:0] CLBLL_L_X4Y100_SLICE_X4Y100_A3;
  wire [0:0] CLBLL_L_X4Y100_SLICE_X4Y100_A4;
  wire [0:0] CLBLL_L_X4Y100_SLICE_X4Y100_A5;
  wire [0:0] CLBLL_L_X4Y100_SLICE_X4Y100_A6;
  wire [0:0] CLBLL_L_X4Y100_SLICE_X4Y100_AMUX;
  wire [0:0] CLBLL_L_X4Y100_SLICE_X4Y100_AO5;
  wire [0:0] CLBLL_L_X4Y100_SLICE_X4Y100_AO6;
  wire [0:0] CLBLL_L_X4Y100_SLICE_X4Y100_A_CY;
  wire [0:0] CLBLL_L_X4Y100_SLICE_X4Y100_A_XOR;
  wire [0:0] CLBLL_L_X4Y100_SLICE_X4Y100_B;
  wire [0:0] CLBLL_L_X4Y100_SLICE_X4Y100_B1;
  wire [0:0] CLBLL_L_X4Y100_SLICE_X4Y100_B2;
  wire [0:0] CLBLL_L_X4Y100_SLICE_X4Y100_B3;
  wire [0:0] CLBLL_L_X4Y100_SLICE_X4Y100_B4;
  wire [0:0] CLBLL_L_X4Y100_SLICE_X4Y100_B5;
  wire [0:0] CLBLL_L_X4Y100_SLICE_X4Y100_B6;
  wire [0:0] CLBLL_L_X4Y100_SLICE_X4Y100_BO5;
  wire [0:0] CLBLL_L_X4Y100_SLICE_X4Y100_BO6;
  wire [0:0] CLBLL_L_X4Y100_SLICE_X4Y100_B_CY;
  wire [0:0] CLBLL_L_X4Y100_SLICE_X4Y100_B_XOR;
  wire [0:0] CLBLL_L_X4Y100_SLICE_X4Y100_C;
  wire [0:0] CLBLL_L_X4Y100_SLICE_X4Y100_C1;
  wire [0:0] CLBLL_L_X4Y100_SLICE_X4Y100_C2;
  wire [0:0] CLBLL_L_X4Y100_SLICE_X4Y100_C3;
  wire [0:0] CLBLL_L_X4Y100_SLICE_X4Y100_C4;
  wire [0:0] CLBLL_L_X4Y100_SLICE_X4Y100_C5;
  wire [0:0] CLBLL_L_X4Y100_SLICE_X4Y100_C6;
  wire [0:0] CLBLL_L_X4Y100_SLICE_X4Y100_CMUX;
  wire [0:0] CLBLL_L_X4Y100_SLICE_X4Y100_CO5;
  wire [0:0] CLBLL_L_X4Y100_SLICE_X4Y100_CO6;
  wire [0:0] CLBLL_L_X4Y100_SLICE_X4Y100_C_CY;
  wire [0:0] CLBLL_L_X4Y100_SLICE_X4Y100_C_XOR;
  wire [0:0] CLBLL_L_X4Y100_SLICE_X4Y100_D;
  wire [0:0] CLBLL_L_X4Y100_SLICE_X4Y100_D1;
  wire [0:0] CLBLL_L_X4Y100_SLICE_X4Y100_D2;
  wire [0:0] CLBLL_L_X4Y100_SLICE_X4Y100_D3;
  wire [0:0] CLBLL_L_X4Y100_SLICE_X4Y100_D4;
  wire [0:0] CLBLL_L_X4Y100_SLICE_X4Y100_D5;
  wire [0:0] CLBLL_L_X4Y100_SLICE_X4Y100_D6;
  wire [0:0] CLBLL_L_X4Y100_SLICE_X4Y100_DO5;
  wire [0:0] CLBLL_L_X4Y100_SLICE_X4Y100_DO6;
  wire [0:0] CLBLL_L_X4Y100_SLICE_X4Y100_D_CY;
  wire [0:0] CLBLL_L_X4Y100_SLICE_X4Y100_D_XOR;
  wire [0:0] CLBLL_L_X4Y100_SLICE_X5Y100_A;
  wire [0:0] CLBLL_L_X4Y100_SLICE_X5Y100_A1;
  wire [0:0] CLBLL_L_X4Y100_SLICE_X5Y100_A2;
  wire [0:0] CLBLL_L_X4Y100_SLICE_X5Y100_A3;
  wire [0:0] CLBLL_L_X4Y100_SLICE_X5Y100_A4;
  wire [0:0] CLBLL_L_X4Y100_SLICE_X5Y100_A5;
  wire [0:0] CLBLL_L_X4Y100_SLICE_X5Y100_A6;
  wire [0:0] CLBLL_L_X4Y100_SLICE_X5Y100_AO5;
  wire [0:0] CLBLL_L_X4Y100_SLICE_X5Y100_AO6;
  wire [0:0] CLBLL_L_X4Y100_SLICE_X5Y100_A_CY;
  wire [0:0] CLBLL_L_X4Y100_SLICE_X5Y100_A_XOR;
  wire [0:0] CLBLL_L_X4Y100_SLICE_X5Y100_B;
  wire [0:0] CLBLL_L_X4Y100_SLICE_X5Y100_B1;
  wire [0:0] CLBLL_L_X4Y100_SLICE_X5Y100_B2;
  wire [0:0] CLBLL_L_X4Y100_SLICE_X5Y100_B3;
  wire [0:0] CLBLL_L_X4Y100_SLICE_X5Y100_B4;
  wire [0:0] CLBLL_L_X4Y100_SLICE_X5Y100_B5;
  wire [0:0] CLBLL_L_X4Y100_SLICE_X5Y100_B6;
  wire [0:0] CLBLL_L_X4Y100_SLICE_X5Y100_BO5;
  wire [0:0] CLBLL_L_X4Y100_SLICE_X5Y100_BO6;
  wire [0:0] CLBLL_L_X4Y100_SLICE_X5Y100_B_CY;
  wire [0:0] CLBLL_L_X4Y100_SLICE_X5Y100_B_XOR;
  wire [0:0] CLBLL_L_X4Y100_SLICE_X5Y100_C;
  wire [0:0] CLBLL_L_X4Y100_SLICE_X5Y100_C1;
  wire [0:0] CLBLL_L_X4Y100_SLICE_X5Y100_C2;
  wire [0:0] CLBLL_L_X4Y100_SLICE_X5Y100_C3;
  wire [0:0] CLBLL_L_X4Y100_SLICE_X5Y100_C4;
  wire [0:0] CLBLL_L_X4Y100_SLICE_X5Y100_C5;
  wire [0:0] CLBLL_L_X4Y100_SLICE_X5Y100_C6;
  wire [0:0] CLBLL_L_X4Y100_SLICE_X5Y100_CO5;
  wire [0:0] CLBLL_L_X4Y100_SLICE_X5Y100_CO6;
  wire [0:0] CLBLL_L_X4Y100_SLICE_X5Y100_C_CY;
  wire [0:0] CLBLL_L_X4Y100_SLICE_X5Y100_C_XOR;
  wire [0:0] CLBLL_L_X4Y100_SLICE_X5Y100_D;
  wire [0:0] CLBLL_L_X4Y100_SLICE_X5Y100_D1;
  wire [0:0] CLBLL_L_X4Y100_SLICE_X5Y100_D2;
  wire [0:0] CLBLL_L_X4Y100_SLICE_X5Y100_D3;
  wire [0:0] CLBLL_L_X4Y100_SLICE_X5Y100_D4;
  wire [0:0] CLBLL_L_X4Y100_SLICE_X5Y100_D5;
  wire [0:0] CLBLL_L_X4Y100_SLICE_X5Y100_D6;
  wire [0:0] CLBLL_L_X4Y100_SLICE_X5Y100_DO5;
  wire [0:0] CLBLL_L_X4Y100_SLICE_X5Y100_DO6;
  wire [0:0] CLBLL_L_X4Y100_SLICE_X5Y100_D_CY;
  wire [0:0] CLBLL_L_X4Y100_SLICE_X5Y100_D_XOR;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X4Y101_A;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X4Y101_A1;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X4Y101_A2;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X4Y101_A3;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X4Y101_A4;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X4Y101_A5;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X4Y101_A6;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X4Y101_AO5;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X4Y101_AO6;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X4Y101_A_CY;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X4Y101_A_XOR;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X4Y101_B;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X4Y101_B1;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X4Y101_B2;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X4Y101_B3;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X4Y101_B4;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X4Y101_B5;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X4Y101_B6;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X4Y101_BO5;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X4Y101_BO6;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X4Y101_B_CY;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X4Y101_B_XOR;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X4Y101_C;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X4Y101_C1;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X4Y101_C2;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X4Y101_C3;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X4Y101_C4;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X4Y101_C5;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X4Y101_C6;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X4Y101_CO5;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X4Y101_CO6;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X4Y101_C_CY;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X4Y101_C_XOR;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X4Y101_D;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X4Y101_D1;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X4Y101_D2;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X4Y101_D3;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X4Y101_D4;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X4Y101_D5;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X4Y101_D6;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X4Y101_DO5;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X4Y101_DO6;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X4Y101_D_CY;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X4Y101_D_XOR;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X5Y101_A;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X5Y101_A1;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X5Y101_A2;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X5Y101_A3;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X5Y101_A4;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X5Y101_A5;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X5Y101_A6;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X5Y101_AMUX;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X5Y101_AO5;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X5Y101_AO6;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X5Y101_A_CY;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X5Y101_A_XOR;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X5Y101_B;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X5Y101_B1;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X5Y101_B2;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X5Y101_B3;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X5Y101_B4;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X5Y101_B5;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X5Y101_B6;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X5Y101_BMUX;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X5Y101_BO5;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X5Y101_BO6;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X5Y101_B_CY;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X5Y101_B_XOR;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X5Y101_C;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X5Y101_C1;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X5Y101_C2;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X5Y101_C3;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X5Y101_C4;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X5Y101_C5;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X5Y101_C6;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X5Y101_CMUX;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X5Y101_CO5;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X5Y101_CO6;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X5Y101_C_CY;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X5Y101_C_XOR;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X5Y101_D;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X5Y101_D1;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X5Y101_D2;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X5Y101_D3;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X5Y101_D4;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X5Y101_D5;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X5Y101_D6;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X5Y101_DO5;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X5Y101_DO6;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X5Y101_D_CY;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X5Y101_D_XOR;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X4Y102_A;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X4Y102_A1;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X4Y102_A2;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X4Y102_A3;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X4Y102_A4;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X4Y102_A5;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X4Y102_A6;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X4Y102_AMUX;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X4Y102_AO5;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X4Y102_AO6;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X4Y102_A_CY;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X4Y102_A_XOR;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X4Y102_B;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X4Y102_B1;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X4Y102_B2;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X4Y102_B3;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X4Y102_B4;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X4Y102_B5;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X4Y102_B6;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X4Y102_BMUX;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X4Y102_BO5;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X4Y102_BO6;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X4Y102_B_CY;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X4Y102_B_XOR;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X4Y102_C;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X4Y102_C1;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X4Y102_C2;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X4Y102_C3;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X4Y102_C4;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X4Y102_C5;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X4Y102_C6;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X4Y102_CO5;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X4Y102_CO6;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X4Y102_C_CY;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X4Y102_C_XOR;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X4Y102_D;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X4Y102_D1;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X4Y102_D2;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X4Y102_D3;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X4Y102_D4;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X4Y102_D5;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X4Y102_D6;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X4Y102_DO5;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X4Y102_DO6;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X4Y102_D_CY;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X4Y102_D_XOR;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X5Y102_A;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X5Y102_A1;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X5Y102_A2;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X5Y102_A3;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X5Y102_A4;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X5Y102_A5;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X5Y102_A6;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X5Y102_AO5;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X5Y102_AO6;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X5Y102_A_CY;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X5Y102_A_XOR;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X5Y102_B;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X5Y102_B1;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X5Y102_B2;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X5Y102_B3;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X5Y102_B4;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X5Y102_B5;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X5Y102_B6;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X5Y102_BO5;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X5Y102_BO6;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X5Y102_B_CY;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X5Y102_B_XOR;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X5Y102_C;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X5Y102_C1;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X5Y102_C2;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X5Y102_C3;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X5Y102_C4;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X5Y102_C5;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X5Y102_C6;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X5Y102_CO5;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X5Y102_CO6;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X5Y102_C_CY;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X5Y102_C_XOR;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X5Y102_D;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X5Y102_D1;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X5Y102_D2;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X5Y102_D3;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X5Y102_D4;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X5Y102_D5;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X5Y102_D6;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X5Y102_DO5;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X5Y102_DO6;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X5Y102_D_CY;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X5Y102_D_XOR;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_A;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_A1;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_A2;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_A3;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_A4;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_A5;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_A6;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_AO5;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_AO6;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_A_CY;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_A_XOR;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_B;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_B1;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_B2;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_B3;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_B4;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_B5;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_B6;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_BO5;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_BO6;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_B_CY;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_B_XOR;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_C;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_C1;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_C2;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_C3;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_C4;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_C5;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_C6;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_CO5;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_CO6;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_C_CY;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_C_XOR;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_D;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_D1;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_D2;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_D3;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_D4;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_D5;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_D6;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_DO5;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_DO6;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_D_CY;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_D_XOR;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_A;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_A1;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_A2;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_A3;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_A4;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_A5;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_A6;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_AMUX;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_AO5;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_AO6;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_A_CY;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_A_XOR;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_B;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_B1;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_B2;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_B3;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_B4;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_B5;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_B6;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_BMUX;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_BO5;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_BO6;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_B_CY;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_B_XOR;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_C;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_C1;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_C2;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_C3;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_C4;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_C5;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_C6;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_CMUX;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_CO5;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_CO6;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_C_CY;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_C_XOR;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_D;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_D1;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_D2;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_D3;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_D4;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_D5;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_D6;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_DO5;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_DO6;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_D_CY;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_D_XOR;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_A;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_A1;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_A2;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_A3;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_A4;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_A5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_A6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_AMUX;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_AO5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_AO6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_A_CY;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_A_XOR;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_B;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_B1;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_B2;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_B3;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_B4;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_B5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_B6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_BMUX;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_BO5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_BO6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_B_CY;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_B_XOR;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_C;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_C1;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_C2;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_C3;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_C4;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_C5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_C6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_CMUX;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_CO5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_CO6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_C_CY;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_C_XOR;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_D;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_D1;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_D2;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_D3;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_D4;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_D5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_D6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_DO5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_DO6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_D_CY;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_D_XOR;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_A;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_A1;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_A2;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_A3;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_A4;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_A5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_A6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_AMUX;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_AO5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_AO6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_A_CY;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_A_XOR;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_B;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_B1;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_B2;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_B3;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_B4;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_B5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_B6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_BMUX;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_BO5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_BO6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_B_CY;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_B_XOR;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_C;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_C1;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_C2;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_C3;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_C4;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_C5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_C6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_CO5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_CO6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_C_CY;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_C_XOR;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_D;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_D1;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_D2;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_D3;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_D4;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_D5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_D6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_DO5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_DO6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_D_CY;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_D_XOR;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_A;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_A1;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_A2;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_A3;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_A4;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_A5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_A6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_AMUX;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_AO5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_AO6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_A_CY;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_A_XOR;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_B;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_B1;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_B2;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_B3;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_B4;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_B5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_B6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_BO5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_BO6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_B_CY;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_B_XOR;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_C;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_C1;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_C2;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_C3;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_C4;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_C5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_C6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_CO5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_CO6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_C_CY;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_C_XOR;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_D;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_D1;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_D2;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_D3;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_D4;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_D5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_D6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_DO5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_DO6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_D_CY;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_D_XOR;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_A;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_A1;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_A2;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_A3;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_A4;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_A5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_A6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_AO5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_AO6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_A_CY;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_A_XOR;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_B;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_B1;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_B2;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_B3;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_B4;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_B5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_B6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_BMUX;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_BO5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_BO6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_B_CY;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_B_XOR;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_C;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_C1;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_C2;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_C3;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_C4;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_C5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_C6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_CMUX;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_CO5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_CO6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_C_CY;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_C_XOR;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_D;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_D1;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_D2;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_D3;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_D4;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_D5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_D6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_DO5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_DO6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_D_CY;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_D_XOR;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_A;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_A1;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_A2;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_A3;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_A4;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_A5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_A6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_AMUX;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_AO5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_AO6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_A_CY;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_A_XOR;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_B;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_B1;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_B2;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_B3;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_B4;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_B5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_B6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_BO5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_BO6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_B_CY;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_B_XOR;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_C;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_C1;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_C2;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_C3;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_C4;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_C5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_C6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_CO5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_CO6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_C_CY;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_C_XOR;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_D;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_D1;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_D2;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_D3;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_D4;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_D5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_D6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_DO5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_DO6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_D_CY;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_D_XOR;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_A;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_A1;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_A2;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_A3;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_A4;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_A5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_A6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_AO5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_AO6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_A_CY;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_A_XOR;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_B;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_B1;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_B2;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_B3;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_B4;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_B5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_B6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_BO5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_BO6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_B_CY;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_B_XOR;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_C;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_C1;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_C2;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_C3;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_C4;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_C5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_C6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_CO5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_CO6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_C_CY;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_C_XOR;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_D;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_D1;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_D2;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_D3;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_D4;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_D5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_D6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_DO5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_DO6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_D_CY;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_D_XOR;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A1;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A2;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A3;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A4;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_AMUX;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_AO5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_AO6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A_CY;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A_XOR;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B1;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B2;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B3;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B4;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_BO5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_BO6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B_CY;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B_XOR;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C1;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C2;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C3;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C4;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_CO5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_CO6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C_CY;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C_XOR;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D1;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D2;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D3;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D4;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_DO5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_DO6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D_CY;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D_XOR;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A1;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A2;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A3;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A4;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_AMUX;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_AO5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_AO6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A_CY;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A_XOR;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B1;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B2;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B3;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B4;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_BO5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_BO6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B_CY;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B_XOR;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C1;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C2;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C3;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C4;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_CO5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_CO6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C_CY;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C_XOR;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D1;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D2;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D3;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D4;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_DO5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_DO6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D_CY;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D_XOR;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A1;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A2;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A3;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A4;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_AO5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_AO6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A_CY;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A_XOR;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B1;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B2;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B3;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B4;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_BO5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_BO6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B_CY;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B_XOR;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C1;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C2;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C3;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C4;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_CO5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_CO6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C_CY;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C_XOR;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D1;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D2;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D3;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D4;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_DO5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_DO6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D_CY;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D_XOR;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A1;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A2;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A3;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A4;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_AO5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_AO6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A_CY;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A_XOR;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B1;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B2;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B3;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B4;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_BMUX;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_BO5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_BO6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B_CY;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B_XOR;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C1;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C2;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C3;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C4;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_CO5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_CO6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C_CY;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C_XOR;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D1;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D2;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D3;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D4;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_DO5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_DO6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D_CY;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_AO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_AO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_BO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_BO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_CO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_CO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_DO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_DO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_AMUX;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_AO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_AO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_BO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_BO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_CO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_CO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_DMUX;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_DO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_DO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D_XOR;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A1;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A2;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A3;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A4;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_AMUX;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_AO5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_AO6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A_CY;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A_XOR;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B1;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B2;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B3;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B4;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_BO5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_BO6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B_CY;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B_XOR;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C1;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C2;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C3;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C4;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_CO5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_CO6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C_CY;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C_XOR;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D1;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D2;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D3;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D4;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_DO5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_DO6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D_CY;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D_XOR;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A1;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A2;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A3;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A4;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_AMUX;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_AO5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_AO6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A_CY;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A_XOR;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B1;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B2;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B3;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B4;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_BO5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_BO6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B_CY;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B_XOR;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C1;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C2;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C3;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C4;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_CMUX;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_CO5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_CO6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C_CY;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C_XOR;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D1;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D2;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D3;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D4;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_DO5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_DO6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D_CY;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D_XOR;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A1;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A2;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A3;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A4;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_AO5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_AO6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A_CY;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A_XOR;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B1;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B2;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B3;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B4;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_BO5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_BO6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B_CY;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B_XOR;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C1;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C2;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C3;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C4;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_CO5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_CO6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C_CY;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C_XOR;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D1;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D2;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D3;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D4;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_DO5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_DO6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D_CY;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D_XOR;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A1;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A2;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A3;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A4;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_AO5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_AO6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A_CY;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A_XOR;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B1;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B2;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B3;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B4;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_BMUX;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_BO5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_BO6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B_CY;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B_XOR;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C1;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C2;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C3;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C4;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_CO5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_CO6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C_CY;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C_XOR;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D1;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D2;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D3;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D4;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_DO5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_DO6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D_CY;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_AMUX;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_AO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_AO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_BO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_BO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_CO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_CO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_DO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_DO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_AO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_AO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_BO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_BO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_CO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_CO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_DMUX;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_DO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_DO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_AO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_AO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_BO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_BO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_CO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_CO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_DO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_DO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_AMUX;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_AO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_AO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_BO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_BO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_CO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_CO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_DO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_DO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D_XOR;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_A;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_A1;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_A2;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_A3;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_A4;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_A5;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_A6;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_AMUX;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_AO5;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_AO6;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_A_CY;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_A_XOR;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_B;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_B1;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_B2;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_B3;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_B4;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_B5;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_B6;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_BO5;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_BO6;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_B_CY;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_B_XOR;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_C;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_C1;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_C2;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_C3;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_C4;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_C5;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_C6;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_CO5;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_CO6;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_C_CY;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_C_XOR;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_D;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_D1;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_D2;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_D3;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_D4;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_D5;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_D6;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_DO5;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_DO6;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_D_CY;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_D_XOR;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_A;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_A1;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_A2;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_A3;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_A4;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_A5;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_A6;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_AO5;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_AO6;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_A_CY;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_A_XOR;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_B;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_B1;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_B2;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_B3;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_B4;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_B5;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_B6;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_BO5;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_BO6;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_B_CY;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_B_XOR;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_C;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_C1;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_C2;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_C3;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_C4;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_C5;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_C6;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_CO5;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_CO6;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_C_CY;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_C_XOR;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_D;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_D1;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_D2;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_D3;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_D4;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_D5;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_D6;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_DO5;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_DO6;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_D_CY;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_D_XOR;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_A;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_A1;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_A2;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_A3;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_A4;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_A5;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_A6;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_AMUX;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_AO5;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_AO6;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_A_CY;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_A_XOR;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_B;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_B1;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_B2;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_B3;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_B4;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_B5;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_B6;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_BO5;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_BO6;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_B_CY;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_B_XOR;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_C;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_C1;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_C2;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_C3;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_C4;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_C5;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_C6;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_CO5;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_CO6;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_C_CY;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_C_XOR;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_D;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_D1;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_D2;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_D3;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_D4;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_D5;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_D6;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_DO5;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_DO6;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_D_CY;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_D_XOR;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_A;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_A1;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_A2;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_A3;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_A4;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_A5;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_A6;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_AO5;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_AO6;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_A_CY;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_A_XOR;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_B;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_B1;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_B2;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_B3;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_B4;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_B5;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_B6;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_BMUX;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_BO5;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_BO6;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_B_CY;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_B_XOR;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_C;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_C1;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_C2;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_C3;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_C4;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_C5;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_C6;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_CMUX;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_CO5;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_CO6;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_C_CY;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_C_XOR;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_D;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_D1;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_D2;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_D3;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_D4;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_D5;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_D6;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_DO5;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_DO6;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_D_CY;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_D_XOR;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_A;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_A1;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_A2;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_A3;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_A4;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_A5;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_A6;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_AMUX;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_AO5;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_AO6;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_A_CY;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_A_XOR;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_B;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_B1;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_B2;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_B3;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_B4;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_B5;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_B6;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_BO5;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_BO6;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_B_CY;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_B_XOR;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_C;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_C1;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_C2;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_C3;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_C4;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_C5;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_C6;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_CO5;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_CO6;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_C_CY;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_C_XOR;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_D;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_D1;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_D2;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_D3;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_D4;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_D5;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_D6;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_DO5;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_DO6;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_D_CY;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_D_XOR;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_A;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_A1;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_A2;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_A3;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_A4;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_A5;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_A6;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_AO5;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_AO6;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_A_CY;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_A_XOR;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_B;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_B1;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_B2;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_B3;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_B4;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_B5;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_B6;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_BO5;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_BO6;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_B_CY;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_B_XOR;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_C;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_C1;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_C2;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_C3;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_C4;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_C5;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_C6;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_CO5;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_CO6;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_C_CY;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_C_XOR;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_D;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_D1;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_D2;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_D3;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_D4;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_D5;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_D6;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_DO5;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_DO6;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_D_CY;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_D_XOR;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_A;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_A1;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_A2;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_A3;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_A4;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_A5;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_A6;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_AO5;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_AO6;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_A_CY;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_A_XOR;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_B;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_B1;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_B2;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_B3;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_B4;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_B5;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_B6;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_BO5;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_BO6;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_B_CY;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_B_XOR;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_C;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_C1;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_C2;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_C3;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_C4;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_C5;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_C6;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_CO5;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_CO6;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_C_CY;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_C_XOR;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_D;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_D1;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_D2;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_D3;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_D4;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_D5;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_D6;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_DO5;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_DO6;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_D_CY;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_D_XOR;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_A;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_A1;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_A2;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_A3;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_A4;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_A5;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_A6;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_AMUX;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_AO5;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_AO6;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_A_CY;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_A_XOR;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_B;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_B1;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_B2;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_B3;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_B4;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_B5;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_B6;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_BO5;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_BO6;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_B_CY;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_B_XOR;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_C;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_C1;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_C2;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_C3;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_C4;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_C5;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_C6;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_CO5;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_CO6;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_C_CY;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_C_XOR;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_D;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_D1;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_D2;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_D3;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_D4;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_D5;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_D6;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_DO5;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_DO6;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_D_CY;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_D_XOR;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_A;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_A1;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_A2;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_A3;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_A4;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_A5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_A6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_AMUX;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_AO5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_AO6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_A_CY;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_A_XOR;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_B;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_B1;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_B2;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_B3;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_B4;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_B5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_B6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_BO5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_BO6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_B_CY;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_B_XOR;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_C;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_C1;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_C2;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_C3;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_C4;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_C5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_C6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_CO5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_CO6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_C_CY;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_C_XOR;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_D;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_D1;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_D2;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_D3;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_D4;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_D5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_D6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_DO5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_DO6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_D_CY;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_D_XOR;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_A;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_A1;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_A2;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_A3;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_A4;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_A5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_A6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_AMUX;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_AO5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_AO6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_A_CY;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_A_XOR;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_B;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_B1;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_B2;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_B3;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_B4;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_B5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_B6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_BO5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_BO6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_B_CY;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_B_XOR;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_C;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_C1;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_C2;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_C3;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_C4;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_C5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_C6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_CO5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_CO6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_C_CY;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_C_XOR;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_D;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_D1;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_D2;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_D3;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_D4;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_D5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_D6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_DO5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_DO6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_D_CY;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_D_XOR;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_A;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_A1;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_A2;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_A3;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_A4;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_A5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_A6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_AMUX;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_AO5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_AO6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_A_CY;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_A_XOR;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_B;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_B1;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_B2;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_B3;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_B4;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_B5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_B6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_BO5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_BO6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_B_CY;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_B_XOR;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_C;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_C1;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_C2;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_C3;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_C4;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_C5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_C6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_CO5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_CO6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_C_CY;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_C_XOR;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_D;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_D1;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_D2;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_D3;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_D4;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_D5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_D6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_DO5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_DO6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_D_CY;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_D_XOR;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_A;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_A1;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_A2;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_A3;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_A4;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_A5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_A6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_AO5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_AO6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_A_CY;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_A_XOR;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_B;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_B1;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_B2;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_B3;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_B4;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_B5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_B6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_BMUX;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_BO5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_BO6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_B_CY;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_B_XOR;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_C;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_C1;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_C2;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_C3;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_C4;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_C5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_C6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_CO5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_CO6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_C_CY;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_C_XOR;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_D;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_D1;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_D2;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_D3;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_D4;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_D5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_D6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_DO5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_DO6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_D_CY;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_D_XOR;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_A;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_A1;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_A2;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_A3;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_A4;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_A5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_A6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_AMUX;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_AO5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_AO6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_A_CY;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_A_XOR;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_B;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_B1;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_B2;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_B3;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_B4;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_B5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_B6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_BO5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_BO6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_B_CY;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_B_XOR;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_C;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_C1;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_C2;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_C3;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_C4;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_C5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_C6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_CO5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_CO6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_C_CY;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_C_XOR;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_D;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_D1;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_D2;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_D3;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_D4;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_D5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_D6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_DO5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_DO6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_D_CY;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_D_XOR;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_A;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_A1;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_A2;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_A3;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_A4;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_A5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_A6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_AMUX;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_AO5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_AO6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_A_CY;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_A_XOR;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_B;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_B1;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_B2;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_B3;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_B4;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_B5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_B6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_BO5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_BO6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_B_CY;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_B_XOR;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_C;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_C1;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_C2;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_C3;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_C4;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_C5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_C6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_CO5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_CO6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_C_CY;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_C_XOR;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_D;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_D1;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_D2;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_D3;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_D4;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_D5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_D6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_DO5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_DO6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_D_CY;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_D_XOR;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_A;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_A1;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_A2;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_A3;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_A4;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_A5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_A6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_AMUX;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_AO5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_AO6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_A_CY;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_A_XOR;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_B;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_B1;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_B2;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_B3;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_B4;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_B5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_B6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_BO5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_BO6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_B_CY;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_B_XOR;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_C;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_C1;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_C2;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_C3;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_C4;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_C5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_C6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_CO5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_CO6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_C_CY;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_C_XOR;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_D;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_D1;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_D2;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_D3;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_D4;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_D5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_D6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_DO5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_DO6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_D_CY;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_D_XOR;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_A;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_A1;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_A2;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_A3;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_A4;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_A5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_A6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_AO5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_AO6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_A_CY;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_A_XOR;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_B;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_B1;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_B2;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_B3;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_B4;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_B5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_B6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_BO5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_BO6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_B_CY;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_B_XOR;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_C;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_C1;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_C2;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_C3;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_C4;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_C5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_C6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_CO5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_CO6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_C_CY;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_C_XOR;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_D;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_D1;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_D2;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_D3;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_D4;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_D5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_D6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_DO5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_DO6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_D_CY;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_D_XOR;
  wire [0:0] CLBLM_L_X8Y100_SLICE_X10Y100_A;
  wire [0:0] CLBLM_L_X8Y100_SLICE_X10Y100_A1;
  wire [0:0] CLBLM_L_X8Y100_SLICE_X10Y100_A2;
  wire [0:0] CLBLM_L_X8Y100_SLICE_X10Y100_A3;
  wire [0:0] CLBLM_L_X8Y100_SLICE_X10Y100_A4;
  wire [0:0] CLBLM_L_X8Y100_SLICE_X10Y100_A5;
  wire [0:0] CLBLM_L_X8Y100_SLICE_X10Y100_A6;
  wire [0:0] CLBLM_L_X8Y100_SLICE_X10Y100_AMUX;
  wire [0:0] CLBLM_L_X8Y100_SLICE_X10Y100_AO5;
  wire [0:0] CLBLM_L_X8Y100_SLICE_X10Y100_AO6;
  wire [0:0] CLBLM_L_X8Y100_SLICE_X10Y100_A_CY;
  wire [0:0] CLBLM_L_X8Y100_SLICE_X10Y100_A_XOR;
  wire [0:0] CLBLM_L_X8Y100_SLICE_X10Y100_B;
  wire [0:0] CLBLM_L_X8Y100_SLICE_X10Y100_B1;
  wire [0:0] CLBLM_L_X8Y100_SLICE_X10Y100_B2;
  wire [0:0] CLBLM_L_X8Y100_SLICE_X10Y100_B3;
  wire [0:0] CLBLM_L_X8Y100_SLICE_X10Y100_B4;
  wire [0:0] CLBLM_L_X8Y100_SLICE_X10Y100_B5;
  wire [0:0] CLBLM_L_X8Y100_SLICE_X10Y100_B6;
  wire [0:0] CLBLM_L_X8Y100_SLICE_X10Y100_BO5;
  wire [0:0] CLBLM_L_X8Y100_SLICE_X10Y100_BO6;
  wire [0:0] CLBLM_L_X8Y100_SLICE_X10Y100_B_CY;
  wire [0:0] CLBLM_L_X8Y100_SLICE_X10Y100_B_XOR;
  wire [0:0] CLBLM_L_X8Y100_SLICE_X10Y100_C;
  wire [0:0] CLBLM_L_X8Y100_SLICE_X10Y100_C1;
  wire [0:0] CLBLM_L_X8Y100_SLICE_X10Y100_C2;
  wire [0:0] CLBLM_L_X8Y100_SLICE_X10Y100_C3;
  wire [0:0] CLBLM_L_X8Y100_SLICE_X10Y100_C4;
  wire [0:0] CLBLM_L_X8Y100_SLICE_X10Y100_C5;
  wire [0:0] CLBLM_L_X8Y100_SLICE_X10Y100_C6;
  wire [0:0] CLBLM_L_X8Y100_SLICE_X10Y100_CO5;
  wire [0:0] CLBLM_L_X8Y100_SLICE_X10Y100_CO6;
  wire [0:0] CLBLM_L_X8Y100_SLICE_X10Y100_C_CY;
  wire [0:0] CLBLM_L_X8Y100_SLICE_X10Y100_C_XOR;
  wire [0:0] CLBLM_L_X8Y100_SLICE_X10Y100_D;
  wire [0:0] CLBLM_L_X8Y100_SLICE_X10Y100_D1;
  wire [0:0] CLBLM_L_X8Y100_SLICE_X10Y100_D2;
  wire [0:0] CLBLM_L_X8Y100_SLICE_X10Y100_D3;
  wire [0:0] CLBLM_L_X8Y100_SLICE_X10Y100_D4;
  wire [0:0] CLBLM_L_X8Y100_SLICE_X10Y100_D5;
  wire [0:0] CLBLM_L_X8Y100_SLICE_X10Y100_D6;
  wire [0:0] CLBLM_L_X8Y100_SLICE_X10Y100_DO5;
  wire [0:0] CLBLM_L_X8Y100_SLICE_X10Y100_DO6;
  wire [0:0] CLBLM_L_X8Y100_SLICE_X10Y100_D_CY;
  wire [0:0] CLBLM_L_X8Y100_SLICE_X10Y100_D_XOR;
  wire [0:0] CLBLM_L_X8Y100_SLICE_X11Y100_A;
  wire [0:0] CLBLM_L_X8Y100_SLICE_X11Y100_A1;
  wire [0:0] CLBLM_L_X8Y100_SLICE_X11Y100_A2;
  wire [0:0] CLBLM_L_X8Y100_SLICE_X11Y100_A3;
  wire [0:0] CLBLM_L_X8Y100_SLICE_X11Y100_A4;
  wire [0:0] CLBLM_L_X8Y100_SLICE_X11Y100_A5;
  wire [0:0] CLBLM_L_X8Y100_SLICE_X11Y100_A6;
  wire [0:0] CLBLM_L_X8Y100_SLICE_X11Y100_AO5;
  wire [0:0] CLBLM_L_X8Y100_SLICE_X11Y100_AO6;
  wire [0:0] CLBLM_L_X8Y100_SLICE_X11Y100_A_CY;
  wire [0:0] CLBLM_L_X8Y100_SLICE_X11Y100_A_XOR;
  wire [0:0] CLBLM_L_X8Y100_SLICE_X11Y100_B;
  wire [0:0] CLBLM_L_X8Y100_SLICE_X11Y100_B1;
  wire [0:0] CLBLM_L_X8Y100_SLICE_X11Y100_B2;
  wire [0:0] CLBLM_L_X8Y100_SLICE_X11Y100_B3;
  wire [0:0] CLBLM_L_X8Y100_SLICE_X11Y100_B4;
  wire [0:0] CLBLM_L_X8Y100_SLICE_X11Y100_B5;
  wire [0:0] CLBLM_L_X8Y100_SLICE_X11Y100_B6;
  wire [0:0] CLBLM_L_X8Y100_SLICE_X11Y100_BO5;
  wire [0:0] CLBLM_L_X8Y100_SLICE_X11Y100_BO6;
  wire [0:0] CLBLM_L_X8Y100_SLICE_X11Y100_B_CY;
  wire [0:0] CLBLM_L_X8Y100_SLICE_X11Y100_B_XOR;
  wire [0:0] CLBLM_L_X8Y100_SLICE_X11Y100_C;
  wire [0:0] CLBLM_L_X8Y100_SLICE_X11Y100_C1;
  wire [0:0] CLBLM_L_X8Y100_SLICE_X11Y100_C2;
  wire [0:0] CLBLM_L_X8Y100_SLICE_X11Y100_C3;
  wire [0:0] CLBLM_L_X8Y100_SLICE_X11Y100_C4;
  wire [0:0] CLBLM_L_X8Y100_SLICE_X11Y100_C5;
  wire [0:0] CLBLM_L_X8Y100_SLICE_X11Y100_C6;
  wire [0:0] CLBLM_L_X8Y100_SLICE_X11Y100_CO5;
  wire [0:0] CLBLM_L_X8Y100_SLICE_X11Y100_CO6;
  wire [0:0] CLBLM_L_X8Y100_SLICE_X11Y100_C_CY;
  wire [0:0] CLBLM_L_X8Y100_SLICE_X11Y100_C_XOR;
  wire [0:0] CLBLM_L_X8Y100_SLICE_X11Y100_D;
  wire [0:0] CLBLM_L_X8Y100_SLICE_X11Y100_D1;
  wire [0:0] CLBLM_L_X8Y100_SLICE_X11Y100_D2;
  wire [0:0] CLBLM_L_X8Y100_SLICE_X11Y100_D3;
  wire [0:0] CLBLM_L_X8Y100_SLICE_X11Y100_D4;
  wire [0:0] CLBLM_L_X8Y100_SLICE_X11Y100_D5;
  wire [0:0] CLBLM_L_X8Y100_SLICE_X11Y100_D6;
  wire [0:0] CLBLM_L_X8Y100_SLICE_X11Y100_DMUX;
  wire [0:0] CLBLM_L_X8Y100_SLICE_X11Y100_DO5;
  wire [0:0] CLBLM_L_X8Y100_SLICE_X11Y100_DO6;
  wire [0:0] CLBLM_L_X8Y100_SLICE_X11Y100_D_CY;
  wire [0:0] CLBLM_L_X8Y100_SLICE_X11Y100_D_XOR;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_A;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_A1;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_A2;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_A3;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_A4;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_A5;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_A6;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_AO5;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_AO6;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_A_CY;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_A_XOR;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_B;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_B1;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_B2;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_B3;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_B4;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_B5;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_B6;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_BO5;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_BO6;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_B_CY;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_B_XOR;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_C;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_C1;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_C2;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_C3;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_C4;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_C5;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_C6;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_CO5;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_CO6;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_C_CY;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_C_XOR;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_D;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_D1;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_D2;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_D3;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_D4;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_D5;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_D6;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_DO5;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_DO6;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_D_CY;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_D_XOR;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_A;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_A1;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_A2;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_A3;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_A4;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_A5;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_A6;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_AMUX;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_AO5;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_AO6;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_A_CY;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_A_XOR;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_B;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_B1;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_B2;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_B3;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_B4;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_B5;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_B6;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_BO5;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_BO6;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_B_CY;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_B_XOR;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_C;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_C1;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_C2;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_C3;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_C4;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_C5;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_C6;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_CO5;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_CO6;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_C_CY;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_C_XOR;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_D;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_D1;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_D2;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_D3;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_D4;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_D5;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_D6;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_DO5;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_DO6;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_D_CY;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_D_XOR;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_A;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_A1;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_A2;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_A3;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_A4;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_A5;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_A6;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_AMUX;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_AO5;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_AO6;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_A_CY;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_A_XOR;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_B;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_B1;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_B2;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_B3;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_B4;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_B5;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_B6;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_BO5;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_BO6;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_B_CY;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_B_XOR;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_C;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_C1;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_C2;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_C3;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_C4;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_C5;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_C6;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_CO5;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_CO6;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_C_CY;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_C_XOR;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_D;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_D1;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_D2;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_D3;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_D4;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_D5;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_D6;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_DO5;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_DO6;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_D_CY;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_D_XOR;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_A;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_A1;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_A2;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_A3;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_A4;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_A5;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_A6;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_AO5;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_AO6;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_A_CY;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_A_XOR;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_B;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_B1;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_B2;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_B3;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_B4;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_B5;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_B6;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_BO5;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_BO6;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_B_CY;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_B_XOR;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_C;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_C1;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_C2;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_C3;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_C4;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_C5;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_C6;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_CMUX;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_CO5;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_CO6;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_C_CY;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_C_XOR;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_D;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_D1;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_D2;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_D3;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_D4;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_D5;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_D6;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_DO5;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_DO6;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_D_CY;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_D_XOR;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_A;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_A1;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_A2;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_A3;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_A4;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_A5;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_A6;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_AMUX;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_AO5;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_AO6;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_A_CY;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_A_XOR;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_B;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_B1;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_B2;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_B3;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_B4;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_B5;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_B6;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_BO5;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_BO6;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_B_CY;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_B_XOR;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_C;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_C1;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_C2;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_C3;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_C4;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_C5;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_C6;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_CO5;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_CO6;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_C_CY;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_C_XOR;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_D;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_D1;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_D2;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_D3;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_D4;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_D5;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_D6;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_DO5;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_DO6;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_D_CY;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_D_XOR;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_A;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_A1;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_A2;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_A3;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_A4;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_A5;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_A6;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_AMUX;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_AO5;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_AO6;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_A_CY;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_A_XOR;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_B;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_B1;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_B2;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_B3;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_B4;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_B5;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_B6;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_BO5;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_BO6;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_B_CY;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_B_XOR;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_C;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_C1;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_C2;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_C3;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_C4;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_C5;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_C6;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_CO5;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_CO6;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_C_CY;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_C_XOR;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_D;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_D1;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_D2;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_D3;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_D4;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_D5;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_D6;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_DO5;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_DO6;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_D_CY;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_D_XOR;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_A;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_A1;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_A2;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_A3;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_A4;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_A5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_A6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_AMUX;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_AO5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_AO6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_A_CY;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_A_XOR;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_B;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_B1;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_B2;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_B3;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_B4;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_B5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_B6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_BO5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_BO6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_B_CY;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_B_XOR;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_C;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_C1;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_C2;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_C3;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_C4;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_C5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_C6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_CO5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_CO6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_C_CY;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_C_XOR;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_D;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_D1;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_D2;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_D3;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_D4;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_D5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_D6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_DO5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_DO6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_D_CY;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_D_XOR;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_A;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_A1;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_A2;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_A3;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_A4;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_A5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_A6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_AO5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_AO6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_A_CY;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_A_XOR;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_B;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_B1;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_B2;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_B3;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_B4;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_B5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_B6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_BO5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_BO6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_B_CY;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_B_XOR;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_C;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_C1;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_C2;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_C3;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_C4;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_C5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_C6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_CO5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_CO6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_C_CY;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_C_XOR;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_D;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_D1;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_D2;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_D3;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_D4;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_D5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_D6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_DO5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_DO6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_D_CY;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_D_XOR;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_A;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_A1;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_A2;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_A3;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_A4;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_A5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_A6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_AMUX;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_AO5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_AO6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_A_CY;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_A_XOR;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_B;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_B1;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_B2;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_B3;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_B4;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_B5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_B6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_BO5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_BO6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_B_CY;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_B_XOR;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_C;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_C1;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_C2;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_C3;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_C4;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_C5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_C6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_CO5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_CO6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_C_CY;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_C_XOR;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_D;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_D1;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_D2;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_D3;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_D4;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_D5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_D6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_DO5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_DO6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_D_CY;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_D_XOR;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_A;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_A1;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_A2;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_A3;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_A4;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_A5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_A6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_AO5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_AO6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_A_CY;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_A_XOR;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_B;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_B1;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_B2;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_B3;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_B4;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_B5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_B6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_BMUX;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_BO5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_BO6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_B_CY;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_B_XOR;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_C;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_C1;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_C2;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_C3;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_C4;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_C5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_C6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_CO5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_CO6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_C_CY;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_C_XOR;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_D;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_D1;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_D2;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_D3;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_D4;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_D5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_D6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_DMUX;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_DO5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_DO6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_D_CY;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_D_XOR;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_A;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_A1;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_A2;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_A3;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_A4;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_A5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_A6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_AMUX;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_AO5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_AO6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_A_CY;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_A_XOR;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_B;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_B1;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_B2;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_B3;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_B4;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_B5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_B6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_BO5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_BO6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_B_CY;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_B_XOR;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_C;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_C1;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_C2;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_C3;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_C4;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_C5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_C6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_CO5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_CO6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_C_CY;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_C_XOR;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_D;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_D1;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_D2;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_D3;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_D4;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_D5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_D6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_DO5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_DO6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_D_CY;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_D_XOR;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_A;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_A1;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_A2;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_A3;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_A4;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_A5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_A6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_AMUX;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_AO5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_AO6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_A_CY;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_A_XOR;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_B;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_B1;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_B2;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_B3;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_B4;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_B5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_B6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_BO5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_BO6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_B_CY;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_B_XOR;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_C;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_C1;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_C2;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_C3;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_C4;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_C5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_C6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_CO5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_CO6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_C_CY;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_C_XOR;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_D;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_D1;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_D2;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_D3;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_D4;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_D5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_D6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_DO5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_DO6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_D_CY;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_D_XOR;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_A;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_A1;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_A2;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_A3;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_A4;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_A5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_A6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_AMUX;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_AO5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_AO6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_A_CY;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_A_XOR;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_B;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_B1;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_B2;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_B3;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_B4;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_B5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_B6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_BO5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_BO6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_B_CY;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_B_XOR;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_C;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_C1;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_C2;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_C3;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_C4;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_C5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_C6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_CO5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_CO6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_C_CY;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_C_XOR;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_D;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_D1;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_D2;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_D3;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_D4;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_D5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_D6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_DO5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_DO6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_D_CY;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_D_XOR;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_A;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_A1;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_A2;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_A3;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_A4;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_A5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_A6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_AO5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_AO6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_A_CY;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_A_XOR;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_B;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_B1;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_B2;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_B3;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_B4;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_B5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_B6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_BO5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_BO6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_B_CY;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_B_XOR;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_C;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_C1;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_C2;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_C3;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_C4;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_C5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_C6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_CO5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_CO6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_C_CY;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_C_XOR;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_D;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_D1;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_D2;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_D3;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_D4;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_D5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_D6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_DO5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_DO6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_D_CY;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_D_XOR;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_A;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_A1;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_A2;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_A3;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_A4;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_A5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_A6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_AMUX;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_AO5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_AO6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_A_CY;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_A_XOR;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_B;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_B1;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_B2;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_B3;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_B4;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_B5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_B6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_BO5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_BO6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_B_CY;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_B_XOR;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_C;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_C1;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_C2;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_C3;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_C4;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_C5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_C6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_CO5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_CO6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_C_CY;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_C_XOR;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_D;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_D1;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_D2;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_D3;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_D4;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_D5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_D6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_DO5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_DO6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_D_CY;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_D_XOR;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_A;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_A1;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_A2;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_A3;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_A4;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_A5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_A6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_AO5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_AO6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_A_CY;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_A_XOR;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_B;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_B1;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_B2;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_B3;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_B4;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_B5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_B6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_BO5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_BO6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_B_CY;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_B_XOR;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_C;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_C1;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_C2;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_C3;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_C4;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_C5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_C6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_CO5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_CO6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_C_CY;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_C_XOR;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_D;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_D1;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_D2;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_D3;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_D4;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_D5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_D6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_DO5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_DO6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_D_CY;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_D_XOR;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_A;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_A1;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_A2;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_A3;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_A4;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_A5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_A6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_AMUX;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_AO5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_AO6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_A_CY;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_A_XOR;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_B;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_B1;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_B2;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_B3;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_B4;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_B5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_B6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_BO5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_BO6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_B_CY;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_B_XOR;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_C;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_C1;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_C2;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_C3;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_C4;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_C5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_C6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_CMUX;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_CO5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_CO6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_C_CY;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_C_XOR;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_D;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_D1;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_D2;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_D3;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_D4;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_D5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_D6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_DO5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_DO6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_D_CY;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_D_XOR;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_A;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_A1;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_A2;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_A3;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_A4;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_A5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_A6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_AO5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_AO6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_A_CY;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_A_XOR;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_B;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_B1;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_B2;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_B3;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_B4;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_B5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_B6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_BO5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_BO6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_B_CY;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_B_XOR;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_C;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_C1;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_C2;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_C3;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_C4;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_C5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_C6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_CO5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_CO6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_C_CY;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_C_XOR;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_D;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_D1;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_D2;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_D3;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_D4;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_D5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_D6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_DO5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_DO6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_D_CY;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_D_XOR;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A1;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A2;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A3;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A4;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_AO5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_AO6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A_CY;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A_XOR;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B1;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B2;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B3;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B4;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_BO5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_BO6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B_CY;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B_XOR;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C1;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C2;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C3;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C4;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_CO5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_CO6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C_CY;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C_XOR;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D1;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D2;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D3;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D4;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_DO5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_DO6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D_CY;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D_XOR;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A1;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A2;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A3;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A4;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_AMUX;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_AO5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_AO6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A_CY;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A_XOR;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B1;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B2;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B3;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B4;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_BO5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_BO6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B_CY;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B_XOR;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C1;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C2;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C3;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C4;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_CO5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_CO6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C_CY;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C_XOR;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D1;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D2;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D3;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D4;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_DO5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_DO6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D_CY;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D_XOR;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A1;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A2;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A3;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A4;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_AO5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_AO6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A_CY;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A_XOR;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B1;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B2;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B3;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B4;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_BO5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_BO6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B_CY;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B_XOR;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C1;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C2;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C3;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C4;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_CO5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_CO6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C_CY;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C_XOR;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D1;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D2;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D3;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D4;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_DO5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_DO6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D_CY;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D_XOR;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A1;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A2;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A3;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A4;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_AO5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_AO6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A_CY;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A_XOR;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B1;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B2;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B3;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B4;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_BO5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_BO6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B_CY;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B_XOR;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C1;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C2;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C3;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C4;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_CO5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_CO6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C_CY;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C_XOR;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D1;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D2;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D3;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D4;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_DO5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_DO6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D_CY;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D_XOR;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A1;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A2;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A3;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A4;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_AMUX;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_AO5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_AO6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A_CY;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A_XOR;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B1;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B2;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B3;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B4;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_BO5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_BO6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B_CY;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B_XOR;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C1;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C2;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C3;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C4;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_CO5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_CO6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C_CY;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C_XOR;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D1;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D2;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D3;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D4;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_DO5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_DO6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D_CY;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D_XOR;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A1;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A2;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A3;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A4;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_AO5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_AO6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A_CY;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A_XOR;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B1;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B2;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B3;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B4;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_BO5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_BO6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B_CY;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B_XOR;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C1;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C2;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C3;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C4;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_CO5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_CO6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C_CY;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C_XOR;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D1;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D2;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D3;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D4;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_DO5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_DO6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D_CY;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D_XOR;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A1;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A2;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A3;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A4;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_AO5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_AO6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A_CY;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A_XOR;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B1;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B2;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B3;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B4;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_BO5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_BO6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B_CY;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B_XOR;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C1;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C2;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C3;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C4;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_CO5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_CO6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C_CY;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C_XOR;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D1;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D2;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D3;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D4;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_DO5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_DO6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D_CY;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D_XOR;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A1;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A2;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A3;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A4;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_AMUX;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_AO5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_AO6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A_CY;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A_XOR;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B1;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B2;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B3;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B4;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_BO5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_BO6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B_CY;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B_XOR;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C1;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C2;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C3;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C4;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_CO5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_CO6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C_CY;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C_XOR;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D1;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D2;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D3;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D4;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_DO5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_DO6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D_CY;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D_XOR;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_A;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_A1;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_A2;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_A3;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_A4;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_A5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_A6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_AMUX;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_AO5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_AO6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_A_CY;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_A_XOR;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_B;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_B1;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_B2;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_B3;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_B4;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_B5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_B6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_BO5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_BO6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_B_CY;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_B_XOR;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_C;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_C1;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_C2;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_C3;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_C4;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_C5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_C6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_CO5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_CO6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_C_CY;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_C_XOR;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_D;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_D1;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_D2;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_D3;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_D4;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_D5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_D6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_DO5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_DO6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_D_CY;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_D_XOR;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_A;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_A1;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_A2;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_A3;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_A4;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_A5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_A6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_AO5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_AO6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_A_CY;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_A_XOR;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_B;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_B1;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_B2;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_B3;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_B4;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_B5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_B6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_BO5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_BO6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_B_CY;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_B_XOR;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_C;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_C1;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_C2;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_C3;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_C4;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_C5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_C6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_CO5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_CO6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_C_CY;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_C_XOR;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_D;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_D1;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_D2;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_D3;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_D4;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_D5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_D6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_DO5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_DO6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_D_CY;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_D_XOR;
  wire [0:0] CLBLM_R_X3Y100_SLICE_X2Y100_A;
  wire [0:0] CLBLM_R_X3Y100_SLICE_X2Y100_A1;
  wire [0:0] CLBLM_R_X3Y100_SLICE_X2Y100_A2;
  wire [0:0] CLBLM_R_X3Y100_SLICE_X2Y100_A3;
  wire [0:0] CLBLM_R_X3Y100_SLICE_X2Y100_A4;
  wire [0:0] CLBLM_R_X3Y100_SLICE_X2Y100_A5;
  wire [0:0] CLBLM_R_X3Y100_SLICE_X2Y100_A6;
  wire [0:0] CLBLM_R_X3Y100_SLICE_X2Y100_AO5;
  wire [0:0] CLBLM_R_X3Y100_SLICE_X2Y100_AO6;
  wire [0:0] CLBLM_R_X3Y100_SLICE_X2Y100_A_CY;
  wire [0:0] CLBLM_R_X3Y100_SLICE_X2Y100_A_XOR;
  wire [0:0] CLBLM_R_X3Y100_SLICE_X2Y100_B;
  wire [0:0] CLBLM_R_X3Y100_SLICE_X2Y100_B1;
  wire [0:0] CLBLM_R_X3Y100_SLICE_X2Y100_B2;
  wire [0:0] CLBLM_R_X3Y100_SLICE_X2Y100_B3;
  wire [0:0] CLBLM_R_X3Y100_SLICE_X2Y100_B4;
  wire [0:0] CLBLM_R_X3Y100_SLICE_X2Y100_B5;
  wire [0:0] CLBLM_R_X3Y100_SLICE_X2Y100_B6;
  wire [0:0] CLBLM_R_X3Y100_SLICE_X2Y100_BO5;
  wire [0:0] CLBLM_R_X3Y100_SLICE_X2Y100_BO6;
  wire [0:0] CLBLM_R_X3Y100_SLICE_X2Y100_B_CY;
  wire [0:0] CLBLM_R_X3Y100_SLICE_X2Y100_B_XOR;
  wire [0:0] CLBLM_R_X3Y100_SLICE_X2Y100_C;
  wire [0:0] CLBLM_R_X3Y100_SLICE_X2Y100_C1;
  wire [0:0] CLBLM_R_X3Y100_SLICE_X2Y100_C2;
  wire [0:0] CLBLM_R_X3Y100_SLICE_X2Y100_C3;
  wire [0:0] CLBLM_R_X3Y100_SLICE_X2Y100_C4;
  wire [0:0] CLBLM_R_X3Y100_SLICE_X2Y100_C5;
  wire [0:0] CLBLM_R_X3Y100_SLICE_X2Y100_C6;
  wire [0:0] CLBLM_R_X3Y100_SLICE_X2Y100_CO5;
  wire [0:0] CLBLM_R_X3Y100_SLICE_X2Y100_CO6;
  wire [0:0] CLBLM_R_X3Y100_SLICE_X2Y100_C_CY;
  wire [0:0] CLBLM_R_X3Y100_SLICE_X2Y100_C_XOR;
  wire [0:0] CLBLM_R_X3Y100_SLICE_X2Y100_D;
  wire [0:0] CLBLM_R_X3Y100_SLICE_X2Y100_D1;
  wire [0:0] CLBLM_R_X3Y100_SLICE_X2Y100_D2;
  wire [0:0] CLBLM_R_X3Y100_SLICE_X2Y100_D3;
  wire [0:0] CLBLM_R_X3Y100_SLICE_X2Y100_D4;
  wire [0:0] CLBLM_R_X3Y100_SLICE_X2Y100_D5;
  wire [0:0] CLBLM_R_X3Y100_SLICE_X2Y100_D6;
  wire [0:0] CLBLM_R_X3Y100_SLICE_X2Y100_DO5;
  wire [0:0] CLBLM_R_X3Y100_SLICE_X2Y100_DO6;
  wire [0:0] CLBLM_R_X3Y100_SLICE_X2Y100_D_CY;
  wire [0:0] CLBLM_R_X3Y100_SLICE_X2Y100_D_XOR;
  wire [0:0] CLBLM_R_X3Y100_SLICE_X3Y100_A;
  wire [0:0] CLBLM_R_X3Y100_SLICE_X3Y100_A1;
  wire [0:0] CLBLM_R_X3Y100_SLICE_X3Y100_A2;
  wire [0:0] CLBLM_R_X3Y100_SLICE_X3Y100_A3;
  wire [0:0] CLBLM_R_X3Y100_SLICE_X3Y100_A4;
  wire [0:0] CLBLM_R_X3Y100_SLICE_X3Y100_A5;
  wire [0:0] CLBLM_R_X3Y100_SLICE_X3Y100_A6;
  wire [0:0] CLBLM_R_X3Y100_SLICE_X3Y100_AMUX;
  wire [0:0] CLBLM_R_X3Y100_SLICE_X3Y100_AO5;
  wire [0:0] CLBLM_R_X3Y100_SLICE_X3Y100_AO6;
  wire [0:0] CLBLM_R_X3Y100_SLICE_X3Y100_A_CY;
  wire [0:0] CLBLM_R_X3Y100_SLICE_X3Y100_A_XOR;
  wire [0:0] CLBLM_R_X3Y100_SLICE_X3Y100_B;
  wire [0:0] CLBLM_R_X3Y100_SLICE_X3Y100_B1;
  wire [0:0] CLBLM_R_X3Y100_SLICE_X3Y100_B2;
  wire [0:0] CLBLM_R_X3Y100_SLICE_X3Y100_B3;
  wire [0:0] CLBLM_R_X3Y100_SLICE_X3Y100_B4;
  wire [0:0] CLBLM_R_X3Y100_SLICE_X3Y100_B5;
  wire [0:0] CLBLM_R_X3Y100_SLICE_X3Y100_B6;
  wire [0:0] CLBLM_R_X3Y100_SLICE_X3Y100_BO5;
  wire [0:0] CLBLM_R_X3Y100_SLICE_X3Y100_BO6;
  wire [0:0] CLBLM_R_X3Y100_SLICE_X3Y100_B_CY;
  wire [0:0] CLBLM_R_X3Y100_SLICE_X3Y100_B_XOR;
  wire [0:0] CLBLM_R_X3Y100_SLICE_X3Y100_C;
  wire [0:0] CLBLM_R_X3Y100_SLICE_X3Y100_C1;
  wire [0:0] CLBLM_R_X3Y100_SLICE_X3Y100_C2;
  wire [0:0] CLBLM_R_X3Y100_SLICE_X3Y100_C3;
  wire [0:0] CLBLM_R_X3Y100_SLICE_X3Y100_C4;
  wire [0:0] CLBLM_R_X3Y100_SLICE_X3Y100_C5;
  wire [0:0] CLBLM_R_X3Y100_SLICE_X3Y100_C6;
  wire [0:0] CLBLM_R_X3Y100_SLICE_X3Y100_CO5;
  wire [0:0] CLBLM_R_X3Y100_SLICE_X3Y100_CO6;
  wire [0:0] CLBLM_R_X3Y100_SLICE_X3Y100_C_CY;
  wire [0:0] CLBLM_R_X3Y100_SLICE_X3Y100_C_XOR;
  wire [0:0] CLBLM_R_X3Y100_SLICE_X3Y100_D;
  wire [0:0] CLBLM_R_X3Y100_SLICE_X3Y100_D1;
  wire [0:0] CLBLM_R_X3Y100_SLICE_X3Y100_D2;
  wire [0:0] CLBLM_R_X3Y100_SLICE_X3Y100_D3;
  wire [0:0] CLBLM_R_X3Y100_SLICE_X3Y100_D4;
  wire [0:0] CLBLM_R_X3Y100_SLICE_X3Y100_D5;
  wire [0:0] CLBLM_R_X3Y100_SLICE_X3Y100_D6;
  wire [0:0] CLBLM_R_X3Y100_SLICE_X3Y100_DO5;
  wire [0:0] CLBLM_R_X3Y100_SLICE_X3Y100_DO6;
  wire [0:0] CLBLM_R_X3Y100_SLICE_X3Y100_D_CY;
  wire [0:0] CLBLM_R_X3Y100_SLICE_X3Y100_D_XOR;
  wire [0:0] CLBLM_R_X3Y101_SLICE_X2Y101_A;
  wire [0:0] CLBLM_R_X3Y101_SLICE_X2Y101_A1;
  wire [0:0] CLBLM_R_X3Y101_SLICE_X2Y101_A2;
  wire [0:0] CLBLM_R_X3Y101_SLICE_X2Y101_A3;
  wire [0:0] CLBLM_R_X3Y101_SLICE_X2Y101_A4;
  wire [0:0] CLBLM_R_X3Y101_SLICE_X2Y101_A5;
  wire [0:0] CLBLM_R_X3Y101_SLICE_X2Y101_A6;
  wire [0:0] CLBLM_R_X3Y101_SLICE_X2Y101_AO5;
  wire [0:0] CLBLM_R_X3Y101_SLICE_X2Y101_AO6;
  wire [0:0] CLBLM_R_X3Y101_SLICE_X2Y101_A_CY;
  wire [0:0] CLBLM_R_X3Y101_SLICE_X2Y101_A_XOR;
  wire [0:0] CLBLM_R_X3Y101_SLICE_X2Y101_B;
  wire [0:0] CLBLM_R_X3Y101_SLICE_X2Y101_B1;
  wire [0:0] CLBLM_R_X3Y101_SLICE_X2Y101_B2;
  wire [0:0] CLBLM_R_X3Y101_SLICE_X2Y101_B3;
  wire [0:0] CLBLM_R_X3Y101_SLICE_X2Y101_B4;
  wire [0:0] CLBLM_R_X3Y101_SLICE_X2Y101_B5;
  wire [0:0] CLBLM_R_X3Y101_SLICE_X2Y101_B6;
  wire [0:0] CLBLM_R_X3Y101_SLICE_X2Y101_BO5;
  wire [0:0] CLBLM_R_X3Y101_SLICE_X2Y101_BO6;
  wire [0:0] CLBLM_R_X3Y101_SLICE_X2Y101_B_CY;
  wire [0:0] CLBLM_R_X3Y101_SLICE_X2Y101_B_XOR;
  wire [0:0] CLBLM_R_X3Y101_SLICE_X2Y101_C;
  wire [0:0] CLBLM_R_X3Y101_SLICE_X2Y101_C1;
  wire [0:0] CLBLM_R_X3Y101_SLICE_X2Y101_C2;
  wire [0:0] CLBLM_R_X3Y101_SLICE_X2Y101_C3;
  wire [0:0] CLBLM_R_X3Y101_SLICE_X2Y101_C4;
  wire [0:0] CLBLM_R_X3Y101_SLICE_X2Y101_C5;
  wire [0:0] CLBLM_R_X3Y101_SLICE_X2Y101_C6;
  wire [0:0] CLBLM_R_X3Y101_SLICE_X2Y101_CO5;
  wire [0:0] CLBLM_R_X3Y101_SLICE_X2Y101_CO6;
  wire [0:0] CLBLM_R_X3Y101_SLICE_X2Y101_C_CY;
  wire [0:0] CLBLM_R_X3Y101_SLICE_X2Y101_C_XOR;
  wire [0:0] CLBLM_R_X3Y101_SLICE_X2Y101_D;
  wire [0:0] CLBLM_R_X3Y101_SLICE_X2Y101_D1;
  wire [0:0] CLBLM_R_X3Y101_SLICE_X2Y101_D2;
  wire [0:0] CLBLM_R_X3Y101_SLICE_X2Y101_D3;
  wire [0:0] CLBLM_R_X3Y101_SLICE_X2Y101_D4;
  wire [0:0] CLBLM_R_X3Y101_SLICE_X2Y101_D5;
  wire [0:0] CLBLM_R_X3Y101_SLICE_X2Y101_D6;
  wire [0:0] CLBLM_R_X3Y101_SLICE_X2Y101_DO5;
  wire [0:0] CLBLM_R_X3Y101_SLICE_X2Y101_DO6;
  wire [0:0] CLBLM_R_X3Y101_SLICE_X2Y101_D_CY;
  wire [0:0] CLBLM_R_X3Y101_SLICE_X2Y101_D_XOR;
  wire [0:0] CLBLM_R_X3Y101_SLICE_X3Y101_A;
  wire [0:0] CLBLM_R_X3Y101_SLICE_X3Y101_A1;
  wire [0:0] CLBLM_R_X3Y101_SLICE_X3Y101_A2;
  wire [0:0] CLBLM_R_X3Y101_SLICE_X3Y101_A3;
  wire [0:0] CLBLM_R_X3Y101_SLICE_X3Y101_A4;
  wire [0:0] CLBLM_R_X3Y101_SLICE_X3Y101_A5;
  wire [0:0] CLBLM_R_X3Y101_SLICE_X3Y101_A6;
  wire [0:0] CLBLM_R_X3Y101_SLICE_X3Y101_AMUX;
  wire [0:0] CLBLM_R_X3Y101_SLICE_X3Y101_AO5;
  wire [0:0] CLBLM_R_X3Y101_SLICE_X3Y101_AO6;
  wire [0:0] CLBLM_R_X3Y101_SLICE_X3Y101_A_CY;
  wire [0:0] CLBLM_R_X3Y101_SLICE_X3Y101_A_XOR;
  wire [0:0] CLBLM_R_X3Y101_SLICE_X3Y101_B;
  wire [0:0] CLBLM_R_X3Y101_SLICE_X3Y101_B1;
  wire [0:0] CLBLM_R_X3Y101_SLICE_X3Y101_B2;
  wire [0:0] CLBLM_R_X3Y101_SLICE_X3Y101_B3;
  wire [0:0] CLBLM_R_X3Y101_SLICE_X3Y101_B4;
  wire [0:0] CLBLM_R_X3Y101_SLICE_X3Y101_B5;
  wire [0:0] CLBLM_R_X3Y101_SLICE_X3Y101_B6;
  wire [0:0] CLBLM_R_X3Y101_SLICE_X3Y101_BO5;
  wire [0:0] CLBLM_R_X3Y101_SLICE_X3Y101_BO6;
  wire [0:0] CLBLM_R_X3Y101_SLICE_X3Y101_B_CY;
  wire [0:0] CLBLM_R_X3Y101_SLICE_X3Y101_B_XOR;
  wire [0:0] CLBLM_R_X3Y101_SLICE_X3Y101_C;
  wire [0:0] CLBLM_R_X3Y101_SLICE_X3Y101_C1;
  wire [0:0] CLBLM_R_X3Y101_SLICE_X3Y101_C2;
  wire [0:0] CLBLM_R_X3Y101_SLICE_X3Y101_C3;
  wire [0:0] CLBLM_R_X3Y101_SLICE_X3Y101_C4;
  wire [0:0] CLBLM_R_X3Y101_SLICE_X3Y101_C5;
  wire [0:0] CLBLM_R_X3Y101_SLICE_X3Y101_C6;
  wire [0:0] CLBLM_R_X3Y101_SLICE_X3Y101_CO5;
  wire [0:0] CLBLM_R_X3Y101_SLICE_X3Y101_CO6;
  wire [0:0] CLBLM_R_X3Y101_SLICE_X3Y101_C_CY;
  wire [0:0] CLBLM_R_X3Y101_SLICE_X3Y101_C_XOR;
  wire [0:0] CLBLM_R_X3Y101_SLICE_X3Y101_D;
  wire [0:0] CLBLM_R_X3Y101_SLICE_X3Y101_D1;
  wire [0:0] CLBLM_R_X3Y101_SLICE_X3Y101_D2;
  wire [0:0] CLBLM_R_X3Y101_SLICE_X3Y101_D3;
  wire [0:0] CLBLM_R_X3Y101_SLICE_X3Y101_D4;
  wire [0:0] CLBLM_R_X3Y101_SLICE_X3Y101_D5;
  wire [0:0] CLBLM_R_X3Y101_SLICE_X3Y101_D6;
  wire [0:0] CLBLM_R_X3Y101_SLICE_X3Y101_DO5;
  wire [0:0] CLBLM_R_X3Y101_SLICE_X3Y101_DO6;
  wire [0:0] CLBLM_R_X3Y101_SLICE_X3Y101_D_CY;
  wire [0:0] CLBLM_R_X3Y101_SLICE_X3Y101_D_XOR;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X2Y102_A;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X2Y102_A1;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X2Y102_A2;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X2Y102_A3;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X2Y102_A4;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X2Y102_A5;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X2Y102_A6;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X2Y102_AO5;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X2Y102_AO6;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X2Y102_A_CY;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X2Y102_A_XOR;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X2Y102_B;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X2Y102_B1;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X2Y102_B2;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X2Y102_B3;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X2Y102_B4;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X2Y102_B5;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X2Y102_B6;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X2Y102_BO5;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X2Y102_BO6;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X2Y102_B_CY;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X2Y102_B_XOR;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X2Y102_C;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X2Y102_C1;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X2Y102_C2;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X2Y102_C3;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X2Y102_C4;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X2Y102_C5;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X2Y102_C6;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X2Y102_CO5;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X2Y102_CO6;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X2Y102_C_CY;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X2Y102_C_XOR;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X2Y102_D;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X2Y102_D1;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X2Y102_D2;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X2Y102_D3;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X2Y102_D4;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X2Y102_D5;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X2Y102_D6;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X2Y102_DO5;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X2Y102_DO6;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X2Y102_D_CY;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X2Y102_D_XOR;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X3Y102_A;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X3Y102_A1;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X3Y102_A2;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X3Y102_A3;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X3Y102_A4;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X3Y102_A5;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X3Y102_A6;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X3Y102_AO5;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X3Y102_AO6;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X3Y102_A_CY;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X3Y102_A_XOR;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X3Y102_B;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X3Y102_B1;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X3Y102_B2;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X3Y102_B3;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X3Y102_B4;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X3Y102_B5;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X3Y102_B6;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X3Y102_BO5;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X3Y102_BO6;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X3Y102_B_CY;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X3Y102_B_XOR;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X3Y102_C;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X3Y102_C1;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X3Y102_C2;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X3Y102_C3;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X3Y102_C4;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X3Y102_C5;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X3Y102_C6;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X3Y102_CO5;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X3Y102_CO6;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X3Y102_C_CY;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X3Y102_C_XOR;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X3Y102_D;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X3Y102_D1;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X3Y102_D2;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X3Y102_D3;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X3Y102_D4;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X3Y102_D5;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X3Y102_D6;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X3Y102_DO5;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X3Y102_DO6;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X3Y102_D_CY;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X3Y102_D_XOR;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_A;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_A1;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_A2;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_A3;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_A4;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_A5;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_A6;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_AMUX;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_AO5;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_AO6;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_A_CY;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_A_XOR;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_B;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_B1;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_B2;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_B3;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_B4;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_B5;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_B6;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_BO5;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_BO6;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_B_CY;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_B_XOR;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_C;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_C1;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_C2;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_C3;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_C4;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_C5;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_C6;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_CO5;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_CO6;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_C_CY;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_C_XOR;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_D;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_D1;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_D2;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_D3;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_D4;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_D5;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_D6;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_DO5;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_DO6;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_D_CY;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_D_XOR;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_A;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_A1;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_A2;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_A3;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_A4;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_A5;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_A6;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_AMUX;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_AO5;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_AO6;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_A_CY;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_A_XOR;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_B;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_B1;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_B2;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_B3;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_B4;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_B5;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_B6;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_BO5;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_BO6;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_B_CY;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_B_XOR;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_C;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_C1;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_C2;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_C3;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_C4;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_C5;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_C6;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_CMUX;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_CO5;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_CO6;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_C_CY;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_C_XOR;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_D;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_D1;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_D2;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_D3;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_D4;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_D5;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_D6;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_DO5;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_DO6;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_D_CY;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_D_XOR;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_A;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_A1;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_A2;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_A3;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_A4;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_A5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_A6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_AO5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_AO6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_A_CY;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_A_XOR;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_B;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_B1;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_B2;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_B3;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_B4;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_B5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_B6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_BO5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_BO6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_B_CY;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_B_XOR;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_C;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_C1;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_C2;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_C3;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_C4;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_C5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_C6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_CO5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_CO6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_C_CY;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_C_XOR;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_D;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_D1;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_D2;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_D3;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_D4;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_D5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_D6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_DO5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_DO6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_D_CY;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_D_XOR;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_A;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_A1;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_A2;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_A3;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_A4;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_A5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_A6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_AMUX;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_AO5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_AO6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_A_CY;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_A_XOR;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_B;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_B1;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_B2;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_B3;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_B4;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_B5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_B6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_BO5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_BO6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_B_CY;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_B_XOR;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_C;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_C1;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_C2;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_C3;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_C4;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_C5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_C6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_CO5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_CO6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_C_CY;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_C_XOR;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_D;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_D1;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_D2;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_D3;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_D4;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_D5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_D6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_DO5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_DO6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_D_CY;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_D_XOR;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_A;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_A1;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_A2;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_A3;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_A4;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_A5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_A6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_AMUX;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_AO5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_AO6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_A_CY;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_A_XOR;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_B;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_B1;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_B2;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_B3;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_B4;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_B5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_B6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_BO5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_BO6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_B_CY;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_B_XOR;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_C;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_C1;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_C2;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_C3;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_C4;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_C5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_C6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_CO5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_CO6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_C_CY;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_C_XOR;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_D;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_D1;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_D2;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_D3;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_D4;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_D5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_D6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_DO5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_DO6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_D_CY;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_D_XOR;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_A;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_A1;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_A2;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_A3;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_A4;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_A5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_A6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_AO5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_AO6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_A_CY;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_A_XOR;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_B;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_B1;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_B2;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_B3;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_B4;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_B5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_B6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_BO5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_BO6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_B_CY;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_B_XOR;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_C;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_C1;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_C2;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_C3;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_C4;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_C5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_C6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_CO5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_CO6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_C_CY;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_C_XOR;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_D;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_D1;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_D2;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_D3;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_D4;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_D5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_D6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_DO5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_DO6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_D_CY;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_D_XOR;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_A;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_A1;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_A2;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_A3;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_A4;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_A5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_A6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_AMUX;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_AO5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_AO6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_A_CY;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_A_XOR;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_B;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_B1;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_B2;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_B3;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_B4;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_B5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_B6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_BO5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_BO6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_B_CY;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_B_XOR;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_C;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_C1;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_C2;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_C3;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_C4;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_C5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_C6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_CO5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_CO6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_C_CY;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_C_XOR;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_D;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_D1;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_D2;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_D3;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_D4;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_D5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_D6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_DO5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_DO6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_D_CY;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_D_XOR;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_A;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_A1;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_A2;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_A3;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_A4;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_A5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_A6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_AMUX;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_AO5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_AO6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_A_CY;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_A_XOR;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_B;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_B1;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_B2;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_B3;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_B4;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_B5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_B6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_BO5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_BO6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_B_CY;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_B_XOR;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_C;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_C1;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_C2;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_C3;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_C4;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_C5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_C6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_CO5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_CO6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_C_CY;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_C_XOR;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_D;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_D1;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_D2;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_D3;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_D4;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_D5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_D6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_DO5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_DO6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_D_CY;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_D_XOR;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_A;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_A1;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_A2;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_A3;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_A4;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_A5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_A6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_AMUX;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_AO5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_AO6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_A_CY;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_A_XOR;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_B;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_B1;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_B2;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_B3;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_B4;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_B5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_B6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_BO5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_BO6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_B_CY;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_B_XOR;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_C;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_C1;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_C2;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_C3;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_C4;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_C5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_C6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_CMUX;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_CO5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_CO6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_C_CY;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_C_XOR;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_D;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_D1;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_D2;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_D3;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_D4;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_D5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_D6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_DO5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_DO6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_D_CY;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_D_XOR;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_A;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_A1;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_A2;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_A3;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_A4;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_A5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_A6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_AMUX;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_AO5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_AO6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_A_CY;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_A_XOR;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_B;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_B1;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_B2;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_B3;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_B4;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_B5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_B6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_BO5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_BO6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_B_CY;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_B_XOR;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_C;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_C1;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_C2;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_C3;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_C4;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_C5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_C6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_CO5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_CO6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_C_CY;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_C_XOR;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_D;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_D1;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_D2;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_D3;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_D4;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_D5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_D6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_DO5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_DO6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_D_CY;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_D_XOR;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_A;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_A1;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_A2;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_A3;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_A4;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_A5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_A6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_AMUX;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_AO5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_AO6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_A_CY;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_A_XOR;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_B;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_B1;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_B2;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_B3;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_B4;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_B5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_B6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_BO5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_BO6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_B_CY;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_B_XOR;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_C;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_C1;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_C2;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_C3;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_C4;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_C5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_C6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_CO5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_CO6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_C_CY;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_C_XOR;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_D;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_D1;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_D2;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_D3;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_D4;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_D5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_D6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_DO5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_DO6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_D_CY;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_D_XOR;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_A;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_A1;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_A2;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_A3;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_A4;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_A5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_A6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_AO5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_AO6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_A_CY;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_A_XOR;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_B;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_B1;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_B2;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_B3;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_B4;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_B5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_B6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_BMUX;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_BO5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_BO6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_B_CY;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_B_XOR;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_C;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_C1;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_C2;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_C3;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_C4;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_C5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_C6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_CO5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_CO6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_C_CY;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_C_XOR;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_D;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_D1;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_D2;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_D3;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_D4;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_D5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_D6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_DMUX;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_DO5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_DO6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_D_CY;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_D_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_AO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_AO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_BO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_BO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_CO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_CO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_DO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_DO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_AO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_AO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_BO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_BO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_CO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_CO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_DO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_DO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D_XOR;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A1;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A2;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A3;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A4;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_AMUX;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_AO5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_AO6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A_CY;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A_XOR;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B1;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B2;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B3;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B4;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_BMUX;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_BO5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_BO6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B_CY;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B_XOR;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C1;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C2;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C3;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C4;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_CO5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_CO6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C_CY;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C_XOR;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D1;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D2;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D3;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D4;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_DO5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_DO6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D_CY;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D_XOR;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A1;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A2;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A3;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A4;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_AO5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_AO6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A_CY;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A_XOR;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B1;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B2;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B3;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B4;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_BO5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_BO6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B_CY;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B_XOR;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C1;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C2;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C3;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C4;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_CO5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_CO6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C_CY;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C_XOR;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D1;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D2;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D3;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D4;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_DO5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_DO6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D_CY;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D_XOR;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A1;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A2;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A3;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A4;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_AO5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_AO6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A_CY;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A_XOR;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B1;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B2;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B3;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B4;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_BO5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_BO6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B_CY;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B_XOR;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C1;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C2;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C3;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C4;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_CO5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_CO6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C_CY;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C_XOR;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D1;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D2;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D3;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D4;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_DO5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_DO6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D_CY;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D_XOR;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A1;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A2;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A3;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A4;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_AMUX;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_AO5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_AO6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A_CY;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A_XOR;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B1;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B2;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B3;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B4;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_BMUX;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_BO5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_BO6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B_CY;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B_XOR;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C1;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C2;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C3;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C4;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_CMUX;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_CO5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_CO6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C_CY;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C_XOR;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D1;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D2;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D3;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D4;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_DO5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_DO6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D_CY;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_AMUX;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_AO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_AO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_BO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_BO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_CMUX;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_CO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_CO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_DO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_DO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_AMUX;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_AO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_AO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_BMUX;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_BO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_BO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_CO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_CO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_DO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_DO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D_XOR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A1;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A2;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A3;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A4;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_AMUX;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_AO5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_AO6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A_CY;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A_XOR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B1;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B2;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B3;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B4;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_BMUX;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_BO5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_BO6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B_CY;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B_XOR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C1;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C2;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C3;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C4;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_CO5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_CO6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C_CY;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C_XOR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D1;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D2;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D3;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D4;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_DO5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_DO6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D_CY;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D_XOR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A1;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A2;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A3;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A4;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_AMUX;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_AO5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_AO6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A_CY;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A_XOR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B1;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B2;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B3;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B4;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_BO5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_BO6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B_CY;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B_XOR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C1;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C2;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C3;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C4;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_CO5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_CO6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C_CY;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C_XOR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D1;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D2;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D3;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D4;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_DMUX;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_DO5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_DO6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D_CY;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D_XOR;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A1;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A2;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A3;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A4;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_AMUX;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_AO5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_AO6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A_CY;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A_XOR;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B1;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B2;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B3;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B4;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_BO5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_BO6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B_CY;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B_XOR;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C1;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C2;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C3;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C4;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_CO5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_CO6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C_CY;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C_XOR;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D1;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D2;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D3;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D4;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_DO5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_DO6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D_CY;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D_XOR;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A1;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A2;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A3;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A4;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_AO5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_AO6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A_CY;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A_XOR;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B1;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B2;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B3;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B4;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_BO5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_BO6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B_CY;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B_XOR;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C1;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C2;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C3;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C4;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_CO5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_CO6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C_CY;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C_XOR;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D1;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D2;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D3;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D4;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_DO5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_DO6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D_CY;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D_XOR;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X6Y100_A;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X6Y100_A1;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X6Y100_A2;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X6Y100_A3;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X6Y100_A4;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X6Y100_A5;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X6Y100_A6;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X6Y100_AMUX;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X6Y100_AO5;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X6Y100_AO6;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X6Y100_A_CY;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X6Y100_A_XOR;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X6Y100_B;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X6Y100_B1;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X6Y100_B2;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X6Y100_B3;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X6Y100_B4;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X6Y100_B5;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X6Y100_B6;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X6Y100_BO5;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X6Y100_BO6;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X6Y100_B_CY;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X6Y100_B_XOR;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X6Y100_C;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X6Y100_C1;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X6Y100_C2;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X6Y100_C3;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X6Y100_C4;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X6Y100_C5;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X6Y100_C6;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X6Y100_CO5;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X6Y100_CO6;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X6Y100_C_CY;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X6Y100_C_XOR;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X6Y100_D;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X6Y100_D1;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X6Y100_D2;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X6Y100_D3;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X6Y100_D4;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X6Y100_D5;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X6Y100_D6;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X6Y100_DO5;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X6Y100_DO6;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X6Y100_D_CY;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X6Y100_D_XOR;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X7Y100_A;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X7Y100_A1;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X7Y100_A2;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X7Y100_A3;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X7Y100_A4;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X7Y100_A5;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X7Y100_A6;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X7Y100_AO5;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X7Y100_AO6;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X7Y100_A_CY;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X7Y100_A_XOR;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X7Y100_B;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X7Y100_B1;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X7Y100_B2;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X7Y100_B3;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X7Y100_B4;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X7Y100_B5;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X7Y100_B6;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X7Y100_BO5;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X7Y100_BO6;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X7Y100_B_CY;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X7Y100_B_XOR;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X7Y100_C;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X7Y100_C1;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X7Y100_C2;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X7Y100_C3;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X7Y100_C4;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X7Y100_C5;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X7Y100_C6;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X7Y100_CO5;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X7Y100_CO6;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X7Y100_C_CY;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X7Y100_C_XOR;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X7Y100_D;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X7Y100_D1;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X7Y100_D2;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X7Y100_D3;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X7Y100_D4;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X7Y100_D5;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X7Y100_D6;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X7Y100_DO5;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X7Y100_DO6;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X7Y100_D_CY;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X7Y100_D_XOR;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_A;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_A1;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_A2;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_A3;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_A4;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_A5;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_A6;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_AMUX;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_AO5;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_AO6;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_A_CY;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_A_XOR;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_B;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_B1;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_B2;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_B3;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_B4;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_B5;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_B6;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_BO5;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_BO6;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_B_CY;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_B_XOR;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_C;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_C1;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_C2;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_C3;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_C4;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_C5;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_C6;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_CMUX;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_CO5;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_CO6;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_C_CY;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_C_XOR;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_D;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_D1;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_D2;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_D3;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_D4;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_D5;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_D6;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_DO5;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_DO6;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_D_CY;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_D_XOR;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_A;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_A1;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_A2;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_A3;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_A4;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_A5;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_A6;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_AMUX;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_AO5;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_AO6;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_A_CY;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_A_XOR;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_B;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_B1;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_B2;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_B3;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_B4;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_B5;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_B6;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_BO5;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_BO6;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_B_CY;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_B_XOR;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_C;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_C1;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_C2;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_C3;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_C4;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_C5;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_C6;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_CO5;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_CO6;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_C_CY;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_C_XOR;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_D;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_D1;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_D2;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_D3;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_D4;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_D5;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_D6;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_DO5;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_DO6;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_D_CY;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_D_XOR;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_A;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_A1;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_A2;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_A3;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_A4;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_A5;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_A6;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_AMUX;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_AO5;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_AO6;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_A_CY;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_A_XOR;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_B;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_B1;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_B2;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_B3;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_B4;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_B5;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_B6;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_BMUX;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_BO5;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_BO6;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_B_CY;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_B_XOR;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_C;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_C1;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_C2;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_C3;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_C4;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_C5;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_C6;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_CO5;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_CO6;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_C_CY;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_C_XOR;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_D;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_D1;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_D2;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_D3;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_D4;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_D5;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_D6;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_DMUX;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_DO5;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_DO6;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_D_CY;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_D_XOR;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_A;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_A1;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_A2;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_A3;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_A4;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_A5;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_A6;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_AO5;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_AO6;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_A_CY;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_A_XOR;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_B;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_B1;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_B2;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_B3;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_B4;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_B5;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_B6;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_BO5;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_BO6;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_B_CY;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_B_XOR;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_C;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_C1;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_C2;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_C3;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_C4;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_C5;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_C6;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_CO5;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_CO6;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_C_CY;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_C_XOR;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_D;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_D1;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_D2;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_D3;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_D4;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_D5;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_D6;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_DO5;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_DO6;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_D_CY;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_D_XOR;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_A;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_A1;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_A2;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_A3;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_A4;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_A5;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_A6;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_AMUX;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_AO5;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_AO6;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_A_CY;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_A_XOR;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_B;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_B1;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_B2;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_B3;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_B4;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_B5;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_B6;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_BO5;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_BO6;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_B_CY;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_B_XOR;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_C;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_C1;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_C2;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_C3;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_C4;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_C5;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_C6;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_CO5;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_CO6;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_C_CY;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_C_XOR;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_D;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_D1;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_D2;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_D3;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_D4;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_D5;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_D6;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_DO5;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_DO6;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_D_CY;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_D_XOR;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_A;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_A1;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_A2;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_A3;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_A4;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_A5;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_A6;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_AO5;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_AO6;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_A_CY;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_A_XOR;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_B;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_B1;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_B2;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_B3;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_B4;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_B5;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_B6;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_BO5;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_BO6;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_B_CY;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_B_XOR;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_C;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_C1;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_C2;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_C3;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_C4;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_C5;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_C6;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_CO5;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_CO6;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_C_CY;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_C_XOR;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_D;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_D1;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_D2;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_D3;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_D4;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_D5;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_D6;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_DO5;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_DO6;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_D_CY;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_D_XOR;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_A;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_A1;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_A2;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_A3;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_A4;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_A5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_A6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_AO5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_AO6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_A_CY;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_A_XOR;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_B;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_B1;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_B2;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_B3;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_B4;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_B5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_B6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_BO5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_BO6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_B_CY;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_B_XOR;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_C;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_C1;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_C2;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_C3;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_C4;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_C5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_C6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_CO5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_CO6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_C_CY;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_C_XOR;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_D;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_D1;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_D2;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_D3;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_D4;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_D5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_D6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_DO5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_DO6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_D_CY;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_D_XOR;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_A;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_A1;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_A2;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_A3;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_A4;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_A5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_A6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_AO5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_AO6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_A_CY;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_A_XOR;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_B;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_B1;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_B2;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_B3;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_B4;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_B5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_B6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_BO5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_BO6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_B_CY;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_B_XOR;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_C;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_C1;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_C2;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_C3;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_C4;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_C5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_C6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_CO5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_CO6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_C_CY;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_C_XOR;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_D;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_D1;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_D2;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_D3;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_D4;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_D5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_D6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_DO5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_DO6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_D_CY;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_D_XOR;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_A;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_A1;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_A2;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_A3;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_A4;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_A5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_A6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_AO5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_AO6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_A_CY;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_A_XOR;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_B;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_B1;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_B2;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_B3;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_B4;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_B5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_B6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_BO5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_BO6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_B_CY;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_B_XOR;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_C;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_C1;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_C2;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_C3;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_C4;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_C5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_C6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_CO5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_CO6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_C_CY;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_C_XOR;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_D;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_D1;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_D2;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_D3;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_D4;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_D5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_D6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_DO5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_DO6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_D_CY;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_D_XOR;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_A;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_A1;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_A2;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_A3;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_A4;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_A5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_A6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_AMUX;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_AO5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_AO6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_A_CY;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_A_XOR;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_B;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_B1;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_B2;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_B3;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_B4;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_B5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_B6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_BMUX;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_BO5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_BO6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_B_CY;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_B_XOR;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_C;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_C1;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_C2;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_C3;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_C4;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_C5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_C6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_CO5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_CO6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_C_CY;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_C_XOR;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_D;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_D1;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_D2;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_D3;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_D4;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_D5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_D6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_DO5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_DO6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_D_CY;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_D_XOR;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_A;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_A1;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_A2;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_A3;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_A4;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_A5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_A6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_AO5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_AO6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_A_CY;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_A_XOR;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_B;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_B1;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_B2;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_B3;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_B4;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_B5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_B6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_BO5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_BO6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_B_CY;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_B_XOR;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_C;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_C1;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_C2;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_C3;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_C4;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_C5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_C6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_CO5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_CO6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_C_CY;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_C_XOR;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_D;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_D1;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_D2;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_D3;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_D4;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_D5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_D6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_DO5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_DO6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_D_CY;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_D_XOR;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_A;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_A1;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_A2;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_A3;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_A4;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_A5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_A6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_AMUX;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_AO5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_AO6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_A_CY;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_A_XOR;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_B;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_B1;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_B2;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_B3;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_B4;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_B5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_B6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_BO5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_BO6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_B_CY;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_B_XOR;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_C;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_C1;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_C2;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_C3;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_C4;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_C5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_C6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_CO5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_CO6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_C_CY;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_C_XOR;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_D;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_D1;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_D2;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_D3;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_D4;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_D5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_D6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_DO5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_DO6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_D_CY;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_D_XOR;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_A;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_A1;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_A2;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_A3;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_A4;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_A5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_A6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_AMUX;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_AO5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_AO6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_A_CY;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_A_XOR;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_B;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_B1;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_B2;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_B3;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_B4;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_B5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_B6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_BO5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_BO6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_B_CY;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_B_XOR;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_C;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_C1;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_C2;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_C3;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_C4;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_C5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_C6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_CO5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_CO6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_C_CY;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_C_XOR;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_D;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_D1;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_D2;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_D3;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_D4;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_D5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_D6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_DO5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_DO6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_D_CY;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_D_XOR;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_A;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_A1;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_A2;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_A3;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_A4;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_A5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_A6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_AO5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_AO6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_A_CY;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_A_XOR;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_B;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_B1;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_B2;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_B3;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_B4;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_B5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_B6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_BO5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_BO6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_B_CY;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_B_XOR;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_C;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_C1;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_C2;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_C3;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_C4;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_C5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_C6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_CO5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_CO6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_C_CY;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_C_XOR;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_D;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_D1;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_D2;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_D3;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_D4;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_D5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_D6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_DO5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_DO6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_D_CY;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_D_XOR;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_A;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_A1;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_A2;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_A3;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_A4;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_A5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_A6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_AMUX;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_AO5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_AO6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_A_CY;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_A_XOR;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_B;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_B1;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_B2;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_B3;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_B4;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_B5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_B6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_BO5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_BO6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_B_CY;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_B_XOR;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_C;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_C1;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_C2;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_C3;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_C4;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_C5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_C6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_CO5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_CO6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_C_CY;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_C_XOR;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_D;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_D1;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_D2;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_D3;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_D4;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_D5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_D6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_DO5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_DO6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_D_CY;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_D_XOR;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_A;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_A1;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_A2;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_A3;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_A4;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_A5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_A6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_AMUX;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_AO5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_AO6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_A_CY;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_A_XOR;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_B;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_B1;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_B2;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_B3;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_B4;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_B5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_B6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_BO5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_BO6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_B_CY;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_B_XOR;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_C;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_C1;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_C2;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_C3;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_C4;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_C5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_C6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_CO5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_CO6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_C_CY;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_C_XOR;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_D;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_D1;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_D2;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_D3;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_D4;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_D5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_D6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_DO5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_DO6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_D_CY;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_D_XOR;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A1;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A2;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A3;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A4;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_AMUX;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_AO5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_AO6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A_CY;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A_XOR;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B1;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B2;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B3;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B4;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_BO5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_BO6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B_CY;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B_XOR;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C1;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C2;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C3;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C4;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_CO5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_CO6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C_CY;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C_XOR;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D1;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D2;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D3;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D4;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_DO5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_DO6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D_CY;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D_XOR;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A1;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A2;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A3;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A4;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_AO5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_AO6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A_CY;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A_XOR;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B1;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B2;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B3;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B4;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_BO5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_BO6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B_CY;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B_XOR;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C1;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C2;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C3;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C4;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_CO5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_CO6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C_CY;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C_XOR;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D1;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D2;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D3;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D4;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_DO5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_DO6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D_CY;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D_XOR;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A1;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A2;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A3;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A4;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_AMUX;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_AO5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_AO6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A_CY;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A_XOR;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B1;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B2;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B3;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B4;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_BO5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_BO6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B_CY;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B_XOR;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C1;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C2;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C3;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C4;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_CO5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_CO6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C_CY;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C_XOR;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D1;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D2;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D3;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D4;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_DO5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_DO6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D_CY;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D_XOR;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A1;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A2;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A3;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A4;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_AMUX;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_AO5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_AO6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A_CY;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A_XOR;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B1;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B2;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B3;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B4;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_BO5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_BO6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B_CY;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B_XOR;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C1;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C2;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C3;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C4;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_CO5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_CO6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C_CY;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C_XOR;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D1;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D2;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D3;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D4;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_DO5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_DO6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D_CY;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D_XOR;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A1;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A2;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A3;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A4;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_AO5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_AO6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A_CY;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A_XOR;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B1;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B2;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B3;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B4;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_BO5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_BO6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B_CY;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B_XOR;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C1;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C2;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C3;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C4;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_CO5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_CO6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C_CY;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C_XOR;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D1;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D2;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D3;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D4;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_DO5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_DO6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D_CY;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D_XOR;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A1;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A2;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A3;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A4;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_AMUX;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_AO5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_AO6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A_CY;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A_XOR;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B1;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B2;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B3;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B4;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_BO5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_BO6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B_CY;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B_XOR;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C1;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C2;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C3;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C4;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_CO5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_CO6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C_CY;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C_XOR;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D1;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D2;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D3;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D4;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_DO5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_DO6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D_CY;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D_XOR;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A1;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A2;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A3;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A4;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_AMUX;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_AO5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_AO6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A_CY;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A_XOR;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B1;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B2;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B3;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B4;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_BO5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_BO6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B_CY;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B_XOR;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C1;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C2;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C3;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C4;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_CO5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_CO6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C_CY;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C_XOR;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D1;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D2;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D3;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D4;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_DMUX;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_DO5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_DO6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D_CY;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D_XOR;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A1;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A2;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A3;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A4;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_AMUX;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_AO5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_AO6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A_CY;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A_XOR;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B1;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B2;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B3;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B4;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_BO5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_BO6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B_CY;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B_XOR;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C1;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C2;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C3;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C4;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_CO5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_CO6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C_CY;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C_XOR;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D1;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D2;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D3;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D4;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_DO5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_DO6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D_CY;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D_XOR;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A1;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A2;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A3;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A4;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_AO5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_AO6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A_CY;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A_XOR;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B1;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B2;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B3;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B4;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_BO5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_BO6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B_CY;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B_XOR;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C1;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C2;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C3;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C4;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_CO5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_CO6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C_CY;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C_XOR;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D1;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D2;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D3;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D4;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_DO5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_DO6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D_CY;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D_XOR;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A1;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A2;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A3;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A4;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_AMUX;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_AO5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_AO6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A_CY;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A_XOR;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B1;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B2;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B3;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B4;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_BO5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_BO6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B_CY;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B_XOR;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C1;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C2;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C3;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C4;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_CO5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_CO6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C_CY;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C_XOR;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D1;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D2;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D3;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D4;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_DO5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_DO6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D_CY;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D_XOR;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X8Y100_A;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X8Y100_A1;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X8Y100_A2;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X8Y100_A3;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X8Y100_A4;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X8Y100_A5;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X8Y100_A6;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X8Y100_AMUX;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X8Y100_AO5;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X8Y100_AO6;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X8Y100_A_CY;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X8Y100_A_XOR;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X8Y100_B;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X8Y100_B1;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X8Y100_B2;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X8Y100_B3;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X8Y100_B4;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X8Y100_B5;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X8Y100_B6;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X8Y100_BO5;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X8Y100_BO6;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X8Y100_B_CY;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X8Y100_B_XOR;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X8Y100_C;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X8Y100_C1;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X8Y100_C2;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X8Y100_C3;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X8Y100_C4;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X8Y100_C5;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X8Y100_C6;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X8Y100_CO5;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X8Y100_CO6;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X8Y100_C_CY;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X8Y100_C_XOR;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X8Y100_D;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X8Y100_D1;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X8Y100_D2;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X8Y100_D3;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X8Y100_D4;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X8Y100_D5;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X8Y100_D6;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X8Y100_DO5;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X8Y100_DO6;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X8Y100_D_CY;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X8Y100_D_XOR;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X9Y100_A;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X9Y100_A1;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X9Y100_A2;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X9Y100_A3;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X9Y100_A4;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X9Y100_A5;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X9Y100_A6;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X9Y100_AO5;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X9Y100_AO6;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X9Y100_A_CY;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X9Y100_A_XOR;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X9Y100_B;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X9Y100_B1;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X9Y100_B2;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X9Y100_B3;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X9Y100_B4;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X9Y100_B5;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X9Y100_B6;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X9Y100_BO5;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X9Y100_BO6;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X9Y100_B_CY;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X9Y100_B_XOR;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X9Y100_C;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X9Y100_C1;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X9Y100_C2;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X9Y100_C3;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X9Y100_C4;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X9Y100_C5;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X9Y100_C6;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X9Y100_CO5;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X9Y100_CO6;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X9Y100_C_CY;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X9Y100_C_XOR;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X9Y100_D;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X9Y100_D1;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X9Y100_D2;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X9Y100_D3;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X9Y100_D4;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X9Y100_D5;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X9Y100_D6;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X9Y100_DO5;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X9Y100_DO6;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X9Y100_D_CY;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X9Y100_D_XOR;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X8Y101_A;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X8Y101_A1;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X8Y101_A2;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X8Y101_A3;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X8Y101_A4;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X8Y101_A5;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X8Y101_A6;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X8Y101_AO5;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X8Y101_AO6;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X8Y101_A_CY;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X8Y101_A_XOR;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X8Y101_B;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X8Y101_B1;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X8Y101_B2;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X8Y101_B3;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X8Y101_B4;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X8Y101_B5;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X8Y101_B6;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X8Y101_BO5;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X8Y101_BO6;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X8Y101_B_CY;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X8Y101_B_XOR;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X8Y101_C;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X8Y101_C1;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X8Y101_C2;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X8Y101_C3;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X8Y101_C4;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X8Y101_C5;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X8Y101_C6;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X8Y101_CMUX;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X8Y101_CO5;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X8Y101_CO6;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X8Y101_C_CY;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X8Y101_C_XOR;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X8Y101_D;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X8Y101_D1;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X8Y101_D2;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X8Y101_D3;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X8Y101_D4;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X8Y101_D5;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X8Y101_D6;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X8Y101_DO5;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X8Y101_DO6;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X8Y101_D_CY;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X8Y101_D_XOR;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X9Y101_A;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X9Y101_A1;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X9Y101_A2;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X9Y101_A3;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X9Y101_A4;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X9Y101_A5;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X9Y101_A6;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X9Y101_AMUX;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X9Y101_AO5;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X9Y101_AO6;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X9Y101_A_CY;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X9Y101_A_XOR;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X9Y101_B;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X9Y101_B1;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X9Y101_B2;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X9Y101_B3;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X9Y101_B4;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X9Y101_B5;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X9Y101_B6;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X9Y101_BO5;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X9Y101_BO6;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X9Y101_B_CY;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X9Y101_B_XOR;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X9Y101_C;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X9Y101_C1;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X9Y101_C2;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X9Y101_C3;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X9Y101_C4;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X9Y101_C5;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X9Y101_C6;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X9Y101_CO5;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X9Y101_CO6;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X9Y101_C_CY;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X9Y101_C_XOR;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X9Y101_D;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X9Y101_D1;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X9Y101_D2;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X9Y101_D3;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X9Y101_D4;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X9Y101_D5;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X9Y101_D6;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X9Y101_DO5;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X9Y101_DO6;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X9Y101_D_CY;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X9Y101_D_XOR;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_A;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_A1;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_A2;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_A3;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_A4;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_A5;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_A6;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_AMUX;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_AO5;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_AO6;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_A_CY;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_A_XOR;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_B;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_B1;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_B2;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_B3;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_B4;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_B5;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_B6;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_BO5;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_BO6;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_B_CY;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_B_XOR;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_C;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_C1;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_C2;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_C3;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_C4;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_C5;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_C6;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_CO5;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_CO6;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_C_CY;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_C_XOR;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_D;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_D1;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_D2;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_D3;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_D4;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_D5;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_D6;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_DO5;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_DO6;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_D_CY;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_D_XOR;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_A;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_A1;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_A2;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_A3;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_A4;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_A5;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_A6;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_AMUX;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_AO5;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_AO6;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_A_CY;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_A_XOR;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_B;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_B1;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_B2;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_B3;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_B4;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_B5;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_B6;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_BO5;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_BO6;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_B_CY;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_B_XOR;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_C;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_C1;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_C2;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_C3;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_C4;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_C5;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_C6;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_CMUX;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_CO5;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_CO6;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_C_CY;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_C_XOR;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_D;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_D1;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_D2;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_D3;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_D4;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_D5;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_D6;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_DO5;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_DO6;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_D_CY;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_D_XOR;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_A;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_A1;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_A2;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_A3;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_A4;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_A5;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_A6;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_AMUX;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_AO5;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_AO6;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_A_CY;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_A_XOR;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_B;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_B1;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_B2;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_B3;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_B4;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_B5;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_B6;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_BMUX;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_BO5;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_BO6;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_B_CY;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_B_XOR;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_C;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_C1;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_C2;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_C3;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_C4;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_C5;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_C6;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_CMUX;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_CO5;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_CO6;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_C_CY;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_C_XOR;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_D;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_D1;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_D2;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_D3;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_D4;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_D5;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_D6;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_DO5;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_DO6;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_D_CY;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_D_XOR;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_A;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_A1;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_A2;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_A3;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_A4;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_A5;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_A6;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_AMUX;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_AO5;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_AO6;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_A_CY;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_A_XOR;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_B;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_B1;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_B2;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_B3;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_B4;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_B5;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_B6;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_BO5;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_BO6;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_B_CY;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_B_XOR;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_C;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_C1;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_C2;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_C3;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_C4;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_C5;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_C6;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_CO5;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_CO6;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_C_CY;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_C_XOR;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_D;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_D1;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_D2;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_D3;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_D4;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_D5;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_D6;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_DO5;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_DO6;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_D_CY;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_D_XOR;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_A;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_A1;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_A2;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_A3;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_A4;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_A5;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_A6;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_AO5;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_AO6;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_A_CY;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_A_XOR;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_B;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_B1;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_B2;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_B3;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_B4;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_B5;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_B6;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_BO5;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_BO6;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_B_CY;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_B_XOR;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_C;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_C1;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_C2;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_C3;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_C4;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_C5;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_C6;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_CO5;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_CO6;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_C_CY;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_C_XOR;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_D;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_D1;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_D2;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_D3;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_D4;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_D5;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_D6;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_DO5;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_DO6;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_D_CY;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_D_XOR;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_A;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_A1;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_A2;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_A3;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_A4;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_A5;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_A6;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_AO5;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_AO6;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_A_CY;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_A_XOR;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_B;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_B1;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_B2;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_B3;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_B4;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_B5;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_B6;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_BO5;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_BO6;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_B_CY;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_B_XOR;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_C;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_C1;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_C2;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_C3;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_C4;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_C5;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_C6;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_CO5;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_CO6;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_C_CY;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_C_XOR;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_D;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_D1;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_D2;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_D3;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_D4;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_D5;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_D6;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_DO5;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_DO6;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_D_CY;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_D_XOR;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_A;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_A1;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_A2;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_A3;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_A4;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_A5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_A6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_AO5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_AO6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_A_CY;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_A_XOR;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_B;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_B1;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_B2;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_B3;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_B4;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_B5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_B6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_BO5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_BO6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_B_CY;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_B_XOR;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_C;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_C1;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_C2;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_C3;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_C4;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_C5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_C6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_CO5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_CO6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_C_CY;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_C_XOR;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_D;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_D1;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_D2;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_D3;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_D4;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_D5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_D6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_DO5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_DO6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_D_CY;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_D_XOR;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_A;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_A1;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_A2;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_A3;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_A4;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_A5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_A6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_AMUX;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_AO5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_AO6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_A_CY;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_A_XOR;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_B;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_B1;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_B2;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_B3;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_B4;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_B5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_B6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_BO5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_BO6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_B_CY;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_B_XOR;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_C;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_C1;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_C2;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_C3;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_C4;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_C5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_C6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_CO5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_CO6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_C_CY;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_C_XOR;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_D;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_D1;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_D2;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_D3;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_D4;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_D5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_D6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_DO5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_DO6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_D_CY;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_D_XOR;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_A;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_A1;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_A2;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_A3;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_A4;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_A5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_A6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_AO5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_AO6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_A_CY;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_A_XOR;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_B;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_B1;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_B2;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_B3;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_B4;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_B5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_B6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_BO5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_BO6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_B_CY;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_B_XOR;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_C;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_C1;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_C2;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_C3;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_C4;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_C5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_C6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_CO5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_CO6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_C_CY;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_C_XOR;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_D;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_D1;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_D2;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_D3;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_D4;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_D5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_D6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_DO5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_DO6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_D_CY;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_D_XOR;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_A;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_A1;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_A2;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_A3;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_A4;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_A5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_A6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_AMUX;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_AO5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_AO6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_A_CY;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_A_XOR;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_B;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_B1;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_B2;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_B3;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_B4;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_B5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_B6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_BO5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_BO6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_B_CY;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_B_XOR;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_C;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_C1;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_C2;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_C3;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_C4;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_C5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_C6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_CO5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_CO6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_C_CY;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_C_XOR;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_D;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_D1;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_D2;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_D3;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_D4;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_D5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_D6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_DO5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_DO6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_D_CY;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_D_XOR;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_A;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_A1;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_A2;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_A3;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_A4;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_A5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_A6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_AO5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_AO6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_A_CY;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_A_XOR;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_B;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_B1;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_B2;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_B3;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_B4;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_B5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_B6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_BO5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_BO6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_B_CY;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_B_XOR;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_C;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_C1;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_C2;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_C3;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_C4;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_C5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_C6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_CO5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_CO6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_C_CY;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_C_XOR;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_D;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_D1;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_D2;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_D3;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_D4;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_D5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_D6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_DO5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_DO6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_D_CY;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_D_XOR;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_A;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_A1;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_A2;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_A3;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_A4;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_A5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_A6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_AMUX;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_AO5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_AO6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_A_CY;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_A_XOR;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_B;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_B1;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_B2;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_B3;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_B4;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_B5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_B6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_BO5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_BO6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_B_CY;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_B_XOR;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_C;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_C1;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_C2;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_C3;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_C4;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_C5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_C6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_CO5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_CO6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_C_CY;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_C_XOR;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_D;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_D1;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_D2;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_D3;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_D4;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_D5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_D6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_DO5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_DO6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_D_CY;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_D_XOR;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_A;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_A1;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_A2;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_A3;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_A4;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_A5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_A6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_AMUX;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_AO5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_AO6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_A_CY;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_A_XOR;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_B;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_B1;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_B2;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_B3;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_B4;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_B5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_B6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_BO5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_BO6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_B_CY;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_B_XOR;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_C;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_C1;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_C2;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_C3;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_C4;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_C5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_C6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_CO5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_CO6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_C_CY;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_C_XOR;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_D;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_D1;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_D2;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_D3;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_D4;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_D5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_D6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_DO5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_DO6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_D_CY;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_D_XOR;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_A;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_A1;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_A2;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_A3;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_A4;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_A5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_A6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_AO5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_AO6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_A_CY;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_A_XOR;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_B;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_B1;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_B2;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_B3;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_B4;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_B5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_B6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_BO5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_BO6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_B_CY;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_B_XOR;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_C;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_C1;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_C2;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_C3;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_C4;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_C5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_C6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_CO5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_CO6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_C_CY;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_C_XOR;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_D;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_D1;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_D2;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_D3;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_D4;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_D5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_D6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_DO5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_DO6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_D_CY;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_D_XOR;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A1;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A2;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A3;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A4;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_AO5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_AO6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A_CY;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A_XOR;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B1;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B2;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B3;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B4;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_BO5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_BO6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B_CY;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B_XOR;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C1;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C2;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C3;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C4;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_CO5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_CO6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C_CY;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C_XOR;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D1;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D2;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D3;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D4;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_DO5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_DO6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D_CY;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D_XOR;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A1;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A2;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A3;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A4;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_AO5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_AO6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A_CY;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A_XOR;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B1;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B2;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B3;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B4;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_BO5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_BO6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B_CY;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B_XOR;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C1;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C2;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C3;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C4;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_CO5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_CO6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C_CY;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C_XOR;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D1;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D2;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D3;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D4;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_DO5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_DO6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D_CY;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D_XOR;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A1;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A2;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A3;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A4;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_AO5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_AO6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A_CY;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A_XOR;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B1;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B2;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B3;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B4;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_BO5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_BO6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B_CY;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B_XOR;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C1;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C2;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C3;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C4;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_CO5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_CO6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C_CY;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C_XOR;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D1;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D2;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D3;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D4;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_DO5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_DO6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D_CY;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D_XOR;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A1;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A2;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A3;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A4;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_AMUX;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_AO5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_AO6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A_CY;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A_XOR;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B1;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B2;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B3;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B4;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_BO5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_BO6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B_CY;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B_XOR;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C1;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C2;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C3;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C4;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_CO5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_CO6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C_CY;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C_XOR;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D1;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D2;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D3;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D4;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_DO5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_DO6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D_CY;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D_XOR;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A1;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A2;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A3;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A4;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_AMUX;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_AO5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_AO6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A_CY;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A_XOR;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B1;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B2;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B3;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B4;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_BO5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_BO6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B_CY;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B_XOR;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C1;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C2;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C3;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C4;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_CO5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_CO6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C_CY;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C_XOR;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D1;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D2;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D3;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D4;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_DO5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_DO6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D_CY;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D_XOR;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A1;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A2;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A3;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A4;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_AO5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_AO6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A_CY;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A_XOR;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B1;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B2;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B3;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B4;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_BO5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_BO6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B_CY;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B_XOR;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C1;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C2;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C3;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C4;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_CO5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_CO6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C_CY;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C_XOR;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D1;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D2;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D3;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D4;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_DO5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_DO6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D_CY;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D_XOR;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A1;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A2;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A3;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A4;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_AMUX;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_AO5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_AO6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A_CY;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A_XOR;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B1;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B2;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B3;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B4;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_BO5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_BO6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B_CY;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B_XOR;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C1;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C2;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C3;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C4;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_CO5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_CO6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C_CY;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C_XOR;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D1;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D2;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D3;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D4;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_DO5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_DO6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D_CY;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D_XOR;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A1;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A2;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A3;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A4;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_AMUX;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_AO5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_AO6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A_CY;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A_XOR;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B1;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B2;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B3;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B4;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_BO5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_BO6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B_CY;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B_XOR;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C1;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C2;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C3;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C4;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_CO5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_CO6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C_CY;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C_XOR;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D1;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D2;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D3;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D4;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_DO5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_DO6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D_CY;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D_XOR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A1;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A2;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A3;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A4;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_AMUX;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_AO5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_AO6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A_CY;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A_XOR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B1;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B2;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B3;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B4;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_BMUX;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_BO5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_BO6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B_CY;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B_XOR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C1;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C2;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C3;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C4;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_CO5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_CO6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C_CY;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C_XOR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D1;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D2;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D3;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D4;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_DO5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_DO6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D_CY;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D_XOR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A1;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A2;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A3;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A4;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_AMUX;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_AO5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_AO6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A_CY;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A_XOR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B1;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B2;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B3;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B4;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_BO5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_BO6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B_CY;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B_XOR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C1;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C2;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C3;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C4;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_CO5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_CO6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C_CY;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C_XOR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D1;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D2;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D3;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D4;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_DO5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_DO6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D_CY;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D_XOR;
  wire [0:0] LIOB33_SING_X0Y100_IOB_X0Y100_I;
  wire [0:0] LIOB33_SING_X0Y149_IOB_X0Y149_O;
  wire [0:0] LIOB33_X0Y101_IOB_X0Y101_I;
  wire [0:0] LIOB33_X0Y101_IOB_X0Y102_I;
  wire [0:0] LIOB33_X0Y103_IOB_X0Y103_I;
  wire [0:0] LIOB33_X0Y103_IOB_X0Y104_I;
  wire [0:0] LIOB33_X0Y105_IOB_X0Y105_I;
  wire [0:0] LIOB33_X0Y105_IOB_X0Y106_I;
  wire [0:0] LIOB33_X0Y107_IOB_X0Y107_I;
  wire [0:0] LIOB33_X0Y107_IOB_X0Y108_I;
  wire [0:0] LIOB33_X0Y109_IOB_X0Y109_I;
  wire [0:0] LIOB33_X0Y109_IOB_X0Y110_I;
  wire [0:0] LIOB33_X0Y111_IOB_X0Y111_I;
  wire [0:0] LIOB33_X0Y111_IOB_X0Y112_I;
  wire [0:0] LIOB33_X0Y113_IOB_X0Y113_I;
  wire [0:0] LIOB33_X0Y113_IOB_X0Y114_I;
  wire [0:0] LIOB33_X0Y115_IOB_X0Y115_I;
  wire [0:0] LIOB33_X0Y115_IOB_X0Y116_I;
  wire [0:0] LIOB33_X0Y117_IOB_X0Y117_I;
  wire [0:0] LIOB33_X0Y117_IOB_X0Y118_O;
  wire [0:0] LIOB33_X0Y119_IOB_X0Y119_O;
  wire [0:0] LIOB33_X0Y119_IOB_X0Y120_O;
  wire [0:0] LIOB33_X0Y121_IOB_X0Y121_O;
  wire [0:0] LIOB33_X0Y121_IOB_X0Y122_O;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y123_O;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y124_O;
  wire [0:0] LIOB33_X0Y125_IOB_X0Y125_O;
  wire [0:0] LIOB33_X0Y125_IOB_X0Y126_O;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y127_O;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y128_O;
  wire [0:0] LIOB33_X0Y129_IOB_X0Y129_O;
  wire [0:0] LIOB33_X0Y129_IOB_X0Y130_O;
  wire [0:0] LIOB33_X0Y131_IOB_X0Y131_O;
  wire [0:0] LIOB33_X0Y131_IOB_X0Y132_O;
  wire [0:0] LIOB33_X0Y133_IOB_X0Y133_O;
  wire [0:0] LIOB33_X0Y133_IOB_X0Y134_O;
  wire [0:0] LIOB33_X0Y135_IOB_X0Y135_O;
  wire [0:0] LIOB33_X0Y135_IOB_X0Y136_O;
  wire [0:0] LIOB33_X0Y137_IOB_X0Y137_O;
  wire [0:0] LIOB33_X0Y137_IOB_X0Y138_O;
  wire [0:0] LIOB33_X0Y139_IOB_X0Y139_O;
  wire [0:0] LIOB33_X0Y139_IOB_X0Y140_O;
  wire [0:0] LIOB33_X0Y141_IOB_X0Y141_O;
  wire [0:0] LIOB33_X0Y141_IOB_X0Y142_O;
  wire [0:0] LIOB33_X0Y143_IOB_X0Y143_O;
  wire [0:0] LIOB33_X0Y145_IOB_X0Y145_O;
  wire [0:0] LIOB33_X0Y145_IOB_X0Y146_O;
  wire [0:0] LIOB33_X0Y147_IOB_X0Y147_O;
  wire [0:0] LIOB33_X0Y147_IOB_X0Y148_O;
  wire [0:0] LIOI3_SING_X0Y100_ILOGIC_X0Y100_D;
  wire [0:0] LIOI3_SING_X0Y100_ILOGIC_X0Y100_O;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_D1;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_OQ;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_T1;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y107_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y107_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y108_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y108_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y113_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y113_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y114_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y114_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_TQ;
  wire [0:0] LIOI3_X0Y101_ILOGIC_X0Y101_D;
  wire [0:0] LIOI3_X0Y101_ILOGIC_X0Y101_O;
  wire [0:0] LIOI3_X0Y101_ILOGIC_X0Y102_D;
  wire [0:0] LIOI3_X0Y101_ILOGIC_X0Y102_O;
  wire [0:0] LIOI3_X0Y103_ILOGIC_X0Y103_D;
  wire [0:0] LIOI3_X0Y103_ILOGIC_X0Y103_O;
  wire [0:0] LIOI3_X0Y103_ILOGIC_X0Y104_D;
  wire [0:0] LIOI3_X0Y103_ILOGIC_X0Y104_O;
  wire [0:0] LIOI3_X0Y105_ILOGIC_X0Y105_D;
  wire [0:0] LIOI3_X0Y105_ILOGIC_X0Y105_O;
  wire [0:0] LIOI3_X0Y105_ILOGIC_X0Y106_D;
  wire [0:0] LIOI3_X0Y105_ILOGIC_X0Y106_O;
  wire [0:0] LIOI3_X0Y109_ILOGIC_X0Y109_D;
  wire [0:0] LIOI3_X0Y109_ILOGIC_X0Y109_O;
  wire [0:0] LIOI3_X0Y109_ILOGIC_X0Y110_D;
  wire [0:0] LIOI3_X0Y109_ILOGIC_X0Y110_O;
  wire [0:0] LIOI3_X0Y111_ILOGIC_X0Y111_D;
  wire [0:0] LIOI3_X0Y111_ILOGIC_X0Y111_O;
  wire [0:0] LIOI3_X0Y111_ILOGIC_X0Y112_D;
  wire [0:0] LIOI3_X0Y111_ILOGIC_X0Y112_O;
  wire [0:0] LIOI3_X0Y115_ILOGIC_X0Y115_D;
  wire [0:0] LIOI3_X0Y115_ILOGIC_X0Y115_O;
  wire [0:0] LIOI3_X0Y115_ILOGIC_X0Y116_D;
  wire [0:0] LIOI3_X0Y115_ILOGIC_X0Y116_O;
  wire [0:0] LIOI3_X0Y117_ILOGIC_X0Y117_D;
  wire [0:0] LIOI3_X0Y117_ILOGIC_X0Y117_O;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_D1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_OQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_T1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_TQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_D1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_OQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_T1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_TQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_D1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_OQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_T1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_TQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_D1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_OQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_T1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_TQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_D1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_OQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_T1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_TQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_D1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_OQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_T1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_TQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_D1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_OQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_T1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_TQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_D1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_OQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_T1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_TQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_D1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_OQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_T1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_TQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_D1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_OQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_T1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_TQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_D1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_OQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_T1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_TQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_D1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_OQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_T1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_TQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_D1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_OQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_T1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_TQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_D1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_OQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_T1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_TQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_D1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_OQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_T1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_TQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_D1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_OQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_T1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_TQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_D1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_OQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_T1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_TQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_D1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_OQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_T1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_TQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_D1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_OQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_T1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_TQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_D1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_OQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_T1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_TQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_D1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_OQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_T1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_TQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_D1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_OQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_T1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_TQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_D1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_OQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_T1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_TQ;
  wire [0:0] RIOB33_SING_X105Y100_IOB_X1Y100_I;
  wire [0:0] RIOB33_X105Y101_IOB_X1Y101_I;
  wire [0:0] RIOB33_X105Y101_IOB_X1Y102_I;
  wire [0:0] RIOB33_X105Y103_IOB_X1Y103_I;
  wire [0:0] RIOB33_X105Y103_IOB_X1Y104_I;
  wire [0:0] RIOB33_X105Y105_IOB_X1Y105_I;
  wire [0:0] RIOB33_X105Y105_IOB_X1Y106_I;
  wire [0:0] RIOB33_X105Y107_IOB_X1Y107_I;
  wire [0:0] RIOB33_X105Y107_IOB_X1Y108_I;
  wire [0:0] RIOB33_X105Y109_IOB_X1Y109_I;
  wire [0:0] RIOB33_X105Y109_IOB_X1Y110_I;
  wire [0:0] RIOB33_X105Y111_IOB_X1Y111_I;
  wire [0:0] RIOB33_X105Y111_IOB_X1Y112_I;
  wire [0:0] RIOB33_X105Y113_IOB_X1Y113_I;
  wire [0:0] RIOI3_SING_X105Y100_ILOGIC_X1Y100_D;
  wire [0:0] RIOI3_SING_X105Y100_ILOGIC_X1Y100_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_O;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y101_D;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y101_O;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y102_D;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y102_O;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y103_D;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y103_O;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y104_D;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y104_O;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y105_D;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y105_O;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y106_D;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y106_O;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y109_D;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y109_O;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y110_D;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y110_O;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y111_D;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y111_O;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y112_D;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y112_O;


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y102_SLICE_X0Y102_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y102_SLICE_X0Y102_DO5),
.O6(CLBLL_L_X2Y102_SLICE_X0Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y102_SLICE_X0Y102_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y102_SLICE_X0Y102_CO5),
.O6(CLBLL_L_X2Y102_SLICE_X0Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y102_SLICE_X0Y102_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y102_SLICE_X0Y102_BO5),
.O6(CLBLL_L_X2Y102_SLICE_X0Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y102_SLICE_X0Y102_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y102_SLICE_X0Y102_AO5),
.O6(CLBLL_L_X2Y102_SLICE_X0Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y102_SLICE_X1Y102_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y102_SLICE_X1Y102_DO5),
.O6(CLBLL_L_X2Y102_SLICE_X1Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y102_SLICE_X1Y102_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y102_SLICE_X1Y102_CO5),
.O6(CLBLL_L_X2Y102_SLICE_X1Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h9f5fb79fdf5f975f)
  ) CLBLL_L_X2Y102_SLICE_X1Y102_BLUT (
.I0(LIOB33_X0Y109_IOB_X0Y110_I),
.I1(LIOB33_X0Y109_IOB_X0Y109_I),
.I2(RIOB33_X105Y111_IOB_X1Y111_I),
.I3(RIOB33_X105Y109_IOB_X1Y110_I),
.I4(CLBLL_L_X2Y102_SLICE_X1Y102_AO6),
.I5(LIOB33_X0Y107_IOB_X0Y108_I),
.O5(CLBLL_L_X2Y102_SLICE_X1Y102_BO5),
.O6(CLBLL_L_X2Y102_SLICE_X1Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h50f7f7ff75fff7ff)
  ) CLBLL_L_X2Y102_SLICE_X1Y102_ALUT (
.I0(RIOB33_X105Y111_IOB_X1Y111_I),
.I1(LIOB33_X0Y105_IOB_X0Y106_I),
.I2(CLBLL_L_X4Y101_SLICE_X4Y101_DO6),
.I3(LIOB33_X0Y107_IOB_X0Y107_I),
.I4(RIOB33_X105Y109_IOB_X1Y110_I),
.I5(LIOB33_X0Y107_IOB_X0Y108_I),
.O5(CLBLL_L_X2Y102_SLICE_X1Y102_AO5),
.O6(CLBLL_L_X2Y102_SLICE_X1Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y103_SLICE_X0Y103_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y103_SLICE_X0Y103_DO5),
.O6(CLBLL_L_X2Y103_SLICE_X0Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y103_SLICE_X0Y103_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y103_SLICE_X0Y103_CO5),
.O6(CLBLL_L_X2Y103_SLICE_X0Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y103_SLICE_X0Y103_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y103_SLICE_X0Y103_BO5),
.O6(CLBLL_L_X2Y103_SLICE_X0Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f0f3f0f3f0f3f0f)
  ) CLBLL_L_X2Y103_SLICE_X0Y103_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y102_SLICE_X6Y102_CO6),
.I2(CLBLL_L_X2Y103_SLICE_X1Y103_AO6),
.I3(CLBLL_L_X4Y106_SLICE_X4Y106_AO5),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y103_SLICE_X0Y103_AO5),
.O6(CLBLL_L_X2Y103_SLICE_X0Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h23bfbbff2bffffff)
  ) CLBLL_L_X2Y103_SLICE_X1Y103_DLUT (
.I0(CLBLL_L_X2Y102_SLICE_X1Y102_AO6),
.I1(RIOB33_X105Y111_IOB_X1Y111_I),
.I2(LIOB33_X0Y109_IOB_X0Y110_I),
.I3(LIOB33_X0Y109_IOB_X0Y109_I),
.I4(RIOB33_X105Y109_IOB_X1Y110_I),
.I5(LIOB33_X0Y107_IOB_X0Y108_I),
.O5(CLBLL_L_X2Y103_SLICE_X1Y103_DO5),
.O6(CLBLL_L_X2Y103_SLICE_X1Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hbc4cc434f0007888)
  ) CLBLL_L_X2Y103_SLICE_X1Y103_CLUT (
.I0(LIOB33_X0Y109_IOB_X0Y110_I),
.I1(RIOB33_X105Y111_IOB_X1Y111_I),
.I2(RIOB33_X105Y109_IOB_X1Y110_I),
.I3(LIOB33_X0Y111_IOB_X0Y112_I),
.I4(CLBLL_L_X2Y103_SLICE_X1Y103_DO6),
.I5(LIOB33_X0Y111_IOB_X0Y111_I),
.O5(CLBLL_L_X2Y103_SLICE_X1Y103_CO5),
.O6(CLBLL_L_X2Y103_SLICE_X1Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha5695a5a0fc3f0f0)
  ) CLBLL_L_X2Y103_SLICE_X1Y103_BLUT (
.I0(LIOB33_X0Y111_IOB_X0Y111_I),
.I1(CLBLL_L_X4Y106_SLICE_X4Y106_AO5),
.I2(CLBLL_L_X4Y101_SLICE_X5Y101_DO6),
.I3(CLBLM_R_X5Y102_SLICE_X6Y102_CO6),
.I4(CLBLL_L_X2Y103_SLICE_X1Y103_AO6),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLL_L_X2Y103_SLICE_X1Y103_BO5),
.O6(CLBLL_L_X2Y103_SLICE_X1Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3fc33cc3cc3cc33)
  ) CLBLL_L_X2Y103_SLICE_X1Y103_ALUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y106_SLICE_X4Y106_AO5),
.I2(RIOB33_X105Y103_IOB_X1Y104_I),
.I3(CLBLM_R_X5Y102_SLICE_X6Y102_CO6),
.I4(LIOB33_X0Y111_IOB_X0Y111_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y103_SLICE_X1Y103_AO5),
.O6(CLBLL_L_X2Y103_SLICE_X1Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00ffffffffff)
  ) CLBLL_L_X2Y104_SLICE_X0Y104_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(RIOB33_X105Y103_IOB_X1Y104_I),
.I4(1'b1),
.I5(LIOB33_X0Y115_IOB_X0Y115_I),
.O5(CLBLL_L_X2Y104_SLICE_X0Y104_DO5),
.O6(CLBLL_L_X2Y104_SLICE_X0Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff2bff002b)
  ) CLBLL_L_X2Y104_SLICE_X0Y104_CLUT (
.I0(CLBLL_L_X2Y104_SLICE_X0Y104_AO6),
.I1(CLBLL_L_X2Y105_SLICE_X1Y105_CO6),
.I2(CLBLL_L_X2Y105_SLICE_X0Y105_BO5),
.I3(CLBLL_L_X2Y104_SLICE_X0Y104_AO5),
.I4(CLBLL_L_X4Y103_SLICE_X4Y103_AO6),
.I5(CLBLL_L_X4Y104_SLICE_X4Y104_CO5),
.O5(CLBLL_L_X2Y104_SLICE_X0Y104_CO5),
.O6(CLBLL_L_X2Y104_SLICE_X0Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hbf3b3b233b232302)
  ) CLBLL_L_X2Y104_SLICE_X0Y104_BLUT (
.I0(CLBLL_L_X2Y105_SLICE_X0Y105_BO5),
.I1(CLBLL_L_X4Y103_SLICE_X4Y103_AO6),
.I2(CLBLL_L_X4Y104_SLICE_X4Y104_BO5),
.I3(CLBLL_L_X2Y104_SLICE_X0Y104_DO6),
.I4(CLBLL_L_X2Y105_SLICE_X0Y105_DO6),
.I5(CLBLL_L_X2Y105_SLICE_X1Y105_CO6),
.O5(CLBLL_L_X2Y104_SLICE_X0Y104_BO5),
.O6(CLBLL_L_X2Y104_SLICE_X0Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h69a569a571f571f5)
  ) CLBLL_L_X2Y104_SLICE_X0Y104_ALUT (
.I0(CLBLL_L_X4Y104_SLICE_X4Y104_BO5),
.I1(LIOB33_X0Y115_IOB_X0Y115_I),
.I2(CLBLL_L_X2Y105_SLICE_X0Y105_DO6),
.I3(RIOB33_X105Y103_IOB_X1Y104_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y104_SLICE_X0Y104_AO5),
.O6(CLBLL_L_X2Y104_SLICE_X0Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y104_SLICE_X1Y104_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y104_SLICE_X1Y104_DO5),
.O6(CLBLL_L_X2Y104_SLICE_X1Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5a5a5a5a5a5a5a5a)
  ) CLBLL_L_X2Y104_SLICE_X1Y104_CLUT (
.I0(CLBLL_L_X4Y104_SLICE_X4Y104_CO5),
.I1(1'b1),
.I2(CLBLL_L_X2Y104_SLICE_X0Y104_BO6),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y104_SLICE_X1Y104_CO5),
.O6(CLBLL_L_X2Y104_SLICE_X1Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h23bbbfff3bffbfff)
  ) CLBLL_L_X2Y104_SLICE_X1Y104_BLUT (
.I0(CLBLL_L_X2Y103_SLICE_X1Y103_DO6),
.I1(LIOB33_X0Y111_IOB_X0Y111_I),
.I2(LIOB33_X0Y109_IOB_X0Y110_I),
.I3(RIOB33_X105Y111_IOB_X1Y111_I),
.I4(RIOB33_X105Y109_IOB_X1Y110_I),
.I5(LIOB33_X0Y111_IOB_X0Y112_I),
.O5(CLBLL_L_X2Y104_SLICE_X1Y104_BO5),
.O6(CLBLL_L_X2Y104_SLICE_X1Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h44dddddd66999999)
  ) CLBLL_L_X2Y104_SLICE_X1Y104_ALUT (
.I0(CLBLM_R_X3Y103_SLICE_X2Y103_BO6),
.I1(CLBLL_L_X4Y104_SLICE_X4Y104_AO5),
.I2(1'b1),
.I3(LIOB33_X0Y115_IOB_X0Y115_I),
.I4(RIOB33_X105Y101_IOB_X1Y101_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y104_SLICE_X1Y104_AO5),
.O6(CLBLL_L_X2Y104_SLICE_X1Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0b0b2bbb2fbfffff)
  ) CLBLL_L_X2Y105_SLICE_X0Y105_DLUT (
.I0(CLBLL_L_X2Y103_SLICE_X0Y103_AO6),
.I1(CLBLL_L_X2Y105_SLICE_X1Y105_AO5),
.I2(RIOB33_X105Y103_IOB_X1Y104_I),
.I3(LIOB33_X0Y111_IOB_X0Y112_I),
.I4(LIOB33_X0Y113_IOB_X0Y113_I),
.I5(CLBLL_L_X4Y101_SLICE_X4Y101_BO6),
.O5(CLBLL_L_X2Y105_SLICE_X0Y105_DO5),
.O6(CLBLL_L_X2Y105_SLICE_X0Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hdb4b2bbb24b4d444)
  ) CLBLL_L_X2Y105_SLICE_X0Y105_CLUT (
.I0(CLBLL_L_X2Y103_SLICE_X0Y103_AO6),
.I1(CLBLL_L_X2Y105_SLICE_X1Y105_AO5),
.I2(RIOB33_X105Y103_IOB_X1Y104_I),
.I3(LIOB33_X0Y111_IOB_X0Y112_I),
.I4(LIOB33_X0Y113_IOB_X0Y113_I),
.I5(CLBLL_L_X4Y101_SLICE_X4Y101_BO6),
.O5(CLBLL_L_X2Y105_SLICE_X0Y105_CO5),
.O6(CLBLL_L_X2Y105_SLICE_X0Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5aaaa5550aaaafff)
  ) CLBLL_L_X2Y105_SLICE_X0Y105_BLUT (
.I0(CLBLL_L_X2Y106_SLICE_X1Y106_BO6),
.I1(1'b1),
.I2(RIOB33_X105Y103_IOB_X1Y103_I),
.I3(LIOB33_X0Y115_IOB_X0Y115_I),
.I4(CLBLL_L_X2Y105_SLICE_X0Y105_CO6),
.I5(1'b1),
.O5(CLBLL_L_X2Y105_SLICE_X0Y105_BO5),
.O6(CLBLL_L_X2Y105_SLICE_X0Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc33cc33c95a96a56)
  ) CLBLL_L_X2Y105_SLICE_X0Y105_ALUT (
.I0(CLBLL_L_X2Y105_SLICE_X0Y105_BO5),
.I1(CLBLL_L_X2Y105_SLICE_X1Y105_BO6),
.I2(CLBLM_R_X3Y106_SLICE_X3Y106_CO6),
.I3(CLBLL_L_X2Y105_SLICE_X0Y105_BO6),
.I4(CLBLL_L_X2Y104_SLICE_X0Y104_AO6),
.I5(1'b1),
.O5(CLBLL_L_X2Y105_SLICE_X0Y105_AO5),
.O6(CLBLL_L_X2Y105_SLICE_X0Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hb42db42d4bd24bd2)
  ) CLBLL_L_X2Y105_SLICE_X1Y105_DLUT (
.I0(CLBLL_L_X2Y107_SLICE_X1Y107_AO6),
.I1(CLBLL_L_X2Y104_SLICE_X1Y104_AO5),
.I2(CLBLL_L_X2Y104_SLICE_X1Y104_AO6),
.I3(CLBLM_R_X3Y105_SLICE_X2Y105_AO5),
.I4(1'b1),
.I5(CLBLM_R_X3Y106_SLICE_X3Y106_BO6),
.O5(CLBLL_L_X2Y105_SLICE_X1Y105_DO5),
.O6(CLBLL_L_X2Y105_SLICE_X1Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfd545500ff55fd54)
  ) CLBLL_L_X2Y105_SLICE_X1Y105_CLUT (
.I0(CLBLL_L_X2Y105_SLICE_X0Y105_BO6),
.I1(CLBLM_R_X3Y105_SLICE_X2Y105_CO6),
.I2(CLBLM_R_X3Y106_SLICE_X2Y106_DO6),
.I3(CLBLM_R_X3Y106_SLICE_X3Y106_CO6),
.I4(CLBLL_L_X2Y104_SLICE_X1Y104_AO6),
.I5(CLBLM_R_X3Y106_SLICE_X3Y106_BO6),
.O5(CLBLL_L_X2Y105_SLICE_X1Y105_CO5),
.O6(CLBLL_L_X2Y105_SLICE_X1Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hb3323220fbb3b332)
  ) CLBLL_L_X2Y105_SLICE_X1Y105_BLUT (
.I0(CLBLL_L_X4Y104_SLICE_X4Y104_AO5),
.I1(CLBLM_R_X3Y106_SLICE_X3Y106_BO6),
.I2(CLBLL_L_X2Y106_SLICE_X1Y106_AO6),
.I3(CLBLM_R_X3Y105_SLICE_X2Y105_AO5),
.I4(CLBLL_L_X2Y107_SLICE_X1Y107_AO6),
.I5(CLBLM_R_X3Y103_SLICE_X2Y103_BO6),
.O5(CLBLL_L_X2Y105_SLICE_X1Y105_BO5),
.O6(CLBLL_L_X2Y105_SLICE_X1Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h55ff55ffcc0033ff)
  ) CLBLL_L_X2Y105_SLICE_X1Y105_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y106_I),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(1'b1),
.I3(LIOB33_X0Y111_IOB_X0Y111_I),
.I4(CLBLL_L_X4Y101_SLICE_X5Y101_DO6),
.I5(1'b1),
.O5(CLBLL_L_X2Y105_SLICE_X1Y105_AO5),
.O6(CLBLL_L_X2Y105_SLICE_X1Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y106_SLICE_X0Y106_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y106_SLICE_X0Y106_DO5),
.O6(CLBLL_L_X2Y106_SLICE_X0Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y106_SLICE_X0Y106_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y106_SLICE_X0Y106_CO5),
.O6(CLBLL_L_X2Y106_SLICE_X0Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc33333333cccc)
  ) CLBLL_L_X2Y106_SLICE_X0Y106_BLUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y103_SLICE_X4Y103_AO6),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLL_L_X2Y106_SLICE_X0Y106_AO6),
.I5(CLBLL_L_X2Y104_SLICE_X0Y104_AO5),
.O5(CLBLL_L_X2Y106_SLICE_X0Y106_BO5),
.O6(CLBLL_L_X2Y106_SLICE_X0Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000fee8e880fffe)
  ) CLBLL_L_X2Y106_SLICE_X0Y106_ALUT (
.I0(CLBLM_R_X3Y106_SLICE_X3Y106_CO6),
.I1(CLBLL_L_X2Y106_SLICE_X1Y106_BO6),
.I2(CLBLL_L_X2Y106_SLICE_X1Y106_AO5),
.I3(CLBLL_L_X2Y105_SLICE_X1Y105_BO6),
.I4(CLBLL_L_X2Y104_SLICE_X0Y104_AO6),
.I5(CLBLL_L_X2Y105_SLICE_X0Y105_CO6),
.O5(CLBLL_L_X2Y106_SLICE_X0Y106_AO5),
.O6(CLBLL_L_X2Y106_SLICE_X0Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y106_SLICE_X1Y106_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y106_SLICE_X1Y106_DO5),
.O6(CLBLL_L_X2Y106_SLICE_X1Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y106_SLICE_X1Y106_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y106_SLICE_X1Y106_CO5),
.O6(CLBLL_L_X2Y106_SLICE_X1Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h78ffffff00787878)
  ) CLBLL_L_X2Y106_SLICE_X1Y106_BLUT (
.I0(RIOB33_X105Y103_IOB_X1Y104_I),
.I1(LIOB33_X0Y111_IOB_X0Y112_I),
.I2(CLBLL_L_X2Y103_SLICE_X1Y103_BO6),
.I3(LIOB33_X0Y113_IOB_X0Y113_I),
.I4(RIOB33_X105Y103_IOB_X1Y103_I),
.I5(CLBLM_R_X3Y103_SLICE_X2Y103_CO6),
.O5(CLBLL_L_X2Y106_SLICE_X1Y106_BO5),
.O6(CLBLL_L_X2Y106_SLICE_X1Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h55ff55ff00ffffff)
  ) CLBLL_L_X2Y106_SLICE_X1Y106_ALUT (
.I0(RIOB33_X105Y101_IOB_X1Y101_I),
.I1(1'b1),
.I2(1'b1),
.I3(LIOB33_X0Y115_IOB_X0Y115_I),
.I4(RIOB33_X105Y103_IOB_X1Y103_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y106_SLICE_X1Y106_AO5),
.O6(CLBLL_L_X2Y106_SLICE_X1Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y107_SLICE_X0Y107_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y107_SLICE_X0Y107_DO5),
.O6(CLBLL_L_X2Y107_SLICE_X0Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y107_SLICE_X0Y107_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y107_SLICE_X0Y107_CO5),
.O6(CLBLL_L_X2Y107_SLICE_X0Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hba222000b2000000)
  ) CLBLL_L_X2Y107_SLICE_X0Y107_BLUT (
.I0(RIOB33_X105Y109_IOB_X1Y110_I),
.I1(CLBLL_L_X2Y104_SLICE_X1Y104_BO6),
.I2(LIOB33_X0Y111_IOB_X0Y112_I),
.I3(RIOB33_X105Y111_IOB_X1Y111_I),
.I4(LIOB33_X0Y113_IOB_X0Y113_I),
.I5(LIOB33_X0Y115_IOB_X0Y115_I),
.O5(CLBLL_L_X2Y107_SLICE_X0Y107_BO5),
.O6(CLBLL_L_X2Y107_SLICE_X0Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'he69eaa224c340088)
  ) CLBLL_L_X2Y107_SLICE_X0Y107_ALUT (
.I0(RIOB33_X105Y109_IOB_X1Y110_I),
.I1(LIOB33_X0Y113_IOB_X0Y113_I),
.I2(LIOB33_X0Y111_IOB_X0Y112_I),
.I3(CLBLL_L_X2Y104_SLICE_X1Y104_BO6),
.I4(RIOB33_X105Y111_IOB_X1Y111_I),
.I5(LIOB33_X0Y115_IOB_X0Y115_I),
.O5(CLBLL_L_X2Y107_SLICE_X0Y107_AO5),
.O6(CLBLL_L_X2Y107_SLICE_X0Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y107_SLICE_X1Y107_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y107_SLICE_X1Y107_DO5),
.O6(CLBLL_L_X2Y107_SLICE_X1Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h55555555aaaaaaaa)
  ) CLBLL_L_X2Y107_SLICE_X1Y107_CLUT (
.I0(CLBLL_L_X2Y107_SLICE_X1Y107_AO6),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X3Y105_SLICE_X2Y105_BO6),
.O5(CLBLL_L_X2Y107_SLICE_X1Y107_CO5),
.O6(CLBLL_L_X2Y107_SLICE_X1Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h1020000000000000)
  ) CLBLL_L_X2Y107_SLICE_X1Y107_BLUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(CLBLL_L_X2Y107_SLICE_X0Y107_BO6),
.I2(RIOB33_X105Y111_IOB_X1Y111_I),
.I3(CLBLL_L_X4Y104_SLICE_X4Y104_DO6),
.I4(LIOB33_X0Y115_IOB_X0Y115_I),
.I5(CLBLL_L_X2Y108_SLICE_X1Y108_CO6),
.O5(CLBLL_L_X2Y107_SLICE_X1Y107_BO5),
.O6(CLBLL_L_X2Y107_SLICE_X1Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h4fbfdf2f040b0d02)
  ) CLBLL_L_X2Y107_SLICE_X1Y107_ALUT (
.I0(CLBLM_R_X3Y109_SLICE_X2Y109_AO6),
.I1(CLBLM_R_X3Y106_SLICE_X2Y106_BO6),
.I2(CLBLM_R_X3Y105_SLICE_X2Y105_AO6),
.I3(CLBLL_L_X2Y107_SLICE_X1Y107_BO6),
.I4(CLBLM_R_X3Y108_SLICE_X2Y108_DO6),
.I5(CLBLM_R_X3Y106_SLICE_X2Y106_CO6),
.O5(CLBLL_L_X2Y107_SLICE_X1Y107_AO5),
.O6(CLBLL_L_X2Y107_SLICE_X1Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h9696969696969696)
  ) CLBLL_L_X2Y108_SLICE_X0Y108_DLUT (
.I0(CLBLM_R_X3Y104_SLICE_X2Y104_CO6),
.I1(CLBLL_L_X2Y107_SLICE_X0Y107_AO6),
.I2(CLBLM_R_X3Y104_SLICE_X3Y104_CO6),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y108_SLICE_X0Y108_DO5),
.O6(CLBLL_L_X2Y108_SLICE_X0Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h4db2b2b2b24d4d4d)
  ) CLBLL_L_X2Y108_SLICE_X0Y108_CLUT (
.I0(CLBLM_R_X3Y104_SLICE_X2Y104_CO6),
.I1(CLBLL_L_X2Y107_SLICE_X0Y107_AO6),
.I2(CLBLM_R_X3Y104_SLICE_X3Y104_CO6),
.I3(RIOB33_X105Y111_IOB_X1Y111_I),
.I4(LIOB33_X0Y115_IOB_X0Y115_I),
.I5(CLBLL_L_X2Y107_SLICE_X0Y107_BO6),
.O5(CLBLL_L_X2Y108_SLICE_X0Y108_CO5),
.O6(CLBLL_L_X2Y108_SLICE_X0Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hba302000fbf3a200)
  ) CLBLL_L_X2Y108_SLICE_X0Y108_BLUT (
.I0(RIOB33_X105Y111_IOB_X1Y111_I),
.I1(CLBLM_R_X3Y104_SLICE_X2Y104_CO6),
.I2(CLBLL_L_X2Y107_SLICE_X0Y107_AO6),
.I3(LIOB33_X0Y115_IOB_X0Y115_I),
.I4(CLBLL_L_X2Y107_SLICE_X0Y107_BO6),
.I5(CLBLM_R_X3Y104_SLICE_X3Y104_CO6),
.O5(CLBLL_L_X2Y108_SLICE_X0Y108_BO5),
.O6(CLBLL_L_X2Y108_SLICE_X0Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0fff0fff00005f5f)
  ) CLBLL_L_X2Y108_SLICE_X0Y108_ALUT (
.I0(RIOB33_X105Y111_IOB_X1Y111_I),
.I1(1'b1),
.I2(LIOB33_X0Y115_IOB_X0Y115_I),
.I3(RIOB33_X105Y105_IOB_X1Y106_I),
.I4(CLBLL_L_X2Y107_SLICE_X0Y107_BO6),
.I5(1'b1),
.O5(CLBLL_L_X2Y108_SLICE_X0Y108_AO5),
.O6(CLBLL_L_X2Y108_SLICE_X0Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6666666699999999)
  ) CLBLL_L_X2Y108_SLICE_X1Y108_DLUT (
.I0(CLBLL_L_X2Y108_SLICE_X1Y108_AO6),
.I1(CLBLM_R_X3Y105_SLICE_X2Y105_AO6),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X3Y106_SLICE_X2Y106_CO6),
.O5(CLBLL_L_X2Y108_SLICE_X1Y108_DO5),
.O6(CLBLL_L_X2Y108_SLICE_X1Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000001000100)
  ) CLBLL_L_X2Y108_SLICE_X1Y108_CLUT (
.I0(CLBLM_R_X5Y102_SLICE_X6Y102_CO6),
.I1(CLBLL_L_X4Y106_SLICE_X4Y106_AO5),
.I2(CLBLL_L_X4Y107_SLICE_X4Y107_BO6),
.I3(CLBLM_R_X5Y110_SLICE_X6Y110_DO6),
.I4(1'b1),
.I5(CLBLM_R_X3Y110_SLICE_X2Y110_AO6),
.O5(CLBLL_L_X2Y108_SLICE_X1Y108_CO5),
.O6(CLBLL_L_X2Y108_SLICE_X1Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000002)
  ) CLBLL_L_X2Y108_SLICE_X1Y108_BLUT (
.I0(CLBLM_R_X5Y110_SLICE_X6Y110_DO6),
.I1(CLBLL_L_X4Y106_SLICE_X4Y106_AO5),
.I2(CLBLL_L_X2Y107_SLICE_X0Y107_BO6),
.I3(CLBLM_R_X3Y110_SLICE_X2Y110_AO6),
.I4(CLBLM_R_X5Y102_SLICE_X6Y102_CO6),
.I5(CLBLL_L_X4Y107_SLICE_X4Y107_BO6),
.O5(CLBLL_L_X2Y108_SLICE_X1Y108_BO5),
.O6(CLBLL_L_X2Y108_SLICE_X1Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h1100e1f0e1f0eeff)
  ) CLBLL_L_X2Y108_SLICE_X1Y108_ALUT (
.I0(CLBLL_L_X2Y108_SLICE_X0Y108_AO5),
.I1(CLBLM_R_X3Y105_SLICE_X2Y105_AO6),
.I2(CLBLM_R_X3Y106_SLICE_X2Y106_BO6),
.I3(CLBLL_L_X2Y108_SLICE_X1Y108_BO6),
.I4(CLBLM_R_X3Y109_SLICE_X2Y109_AO6),
.I5(CLBLM_R_X3Y108_SLICE_X2Y108_DO6),
.O5(CLBLL_L_X2Y108_SLICE_X1Y108_AO5),
.O6(CLBLL_L_X2Y108_SLICE_X1Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y109_SLICE_X0Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y109_SLICE_X0Y109_DO5),
.O6(CLBLL_L_X2Y109_SLICE_X0Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y109_SLICE_X0Y109_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y109_SLICE_X0Y109_CO5),
.O6(CLBLL_L_X2Y109_SLICE_X0Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y109_SLICE_X0Y109_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y109_SLICE_X0Y109_BO5),
.O6(CLBLL_L_X2Y109_SLICE_X0Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y109_SLICE_X0Y109_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y109_SLICE_X0Y109_AO5),
.O6(CLBLL_L_X2Y109_SLICE_X0Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y109_SLICE_X1Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y109_SLICE_X1Y109_DO5),
.O6(CLBLL_L_X2Y109_SLICE_X1Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y109_SLICE_X1Y109_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y109_SLICE_X1Y109_CO5),
.O6(CLBLL_L_X2Y109_SLICE_X1Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y109_SLICE_X1Y109_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y109_SLICE_X1Y109_BO5),
.O6(CLBLL_L_X2Y109_SLICE_X1Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc33cc33cc33cc33c)
  ) CLBLL_L_X2Y109_SLICE_X1Y109_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y109_SLICE_X2Y109_AO6),
.I2(CLBLM_R_X3Y108_SLICE_X2Y108_DO6),
.I3(CLBLM_R_X3Y106_SLICE_X2Y106_BO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y109_SLICE_X1Y109_AO5),
.O6(CLBLL_L_X2Y109_SLICE_X1Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y112_SLICE_X0Y112_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y112_SLICE_X0Y112_DO5),
.O6(CLBLL_L_X2Y112_SLICE_X0Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y112_SLICE_X0Y112_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y112_SLICE_X0Y112_CO5),
.O6(CLBLL_L_X2Y112_SLICE_X0Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h04f4500044345000)
  ) CLBLL_L_X2Y112_SLICE_X0Y112_BLUT (
.I0(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I1(LIOB33_X0Y103_IOB_X0Y103_I),
.I2(RIOB33_X105Y105_IOB_X1Y106_I),
.I3(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I4(RIOB33_X105Y113_IOB_X1Y113_I),
.I5(RIOB33_X105Y111_IOB_X1Y112_I),
.O5(CLBLL_L_X2Y112_SLICE_X0Y112_BO5),
.O6(CLBLL_L_X2Y112_SLICE_X0Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h03737c0c80f0b0c0)
  ) CLBLL_L_X2Y112_SLICE_X0Y112_ALUT (
.I0(RIOB33_X105Y111_IOB_X1Y112_I),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(RIOB33_X105Y113_IOB_X1Y113_I),
.I3(LIOB33_X0Y103_IOB_X0Y103_I),
.I4(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I5(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.O5(CLBLL_L_X2Y112_SLICE_X0Y112_AO5),
.O6(CLBLL_L_X2Y112_SLICE_X0Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y112_SLICE_X1Y112_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y112_SLICE_X1Y112_DO5),
.O6(CLBLL_L_X2Y112_SLICE_X1Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y112_SLICE_X1Y112_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y112_SLICE_X1Y112_CO5),
.O6(CLBLL_L_X2Y112_SLICE_X1Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y112_SLICE_X1Y112_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y112_SLICE_X1Y112_BO5),
.O6(CLBLL_L_X2Y112_SLICE_X1Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6fafffff060a66aa)
  ) CLBLL_L_X2Y112_SLICE_X1Y112_ALUT (
.I0(CLBLM_R_X3Y113_SLICE_X2Y113_CO6),
.I1(LIOB33_X0Y103_IOB_X0Y104_I),
.I2(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I3(RIOB33_X105Y105_IOB_X1Y106_I),
.I4(LIOB33_X0Y105_IOB_X0Y105_I),
.I5(CLBLL_L_X2Y113_SLICE_X1Y113_DO6),
.O5(CLBLL_L_X2Y112_SLICE_X1Y112_AO5),
.O6(CLBLL_L_X2Y112_SLICE_X1Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffdc73cc334010)
  ) CLBLL_L_X2Y113_SLICE_X0Y113_DLUT (
.I0(CLBLL_L_X2Y112_SLICE_X0Y112_AO6),
.I1(CLBLM_R_X3Y113_SLICE_X3Y113_AO5),
.I2(CLBLL_L_X2Y114_SLICE_X0Y114_BO6),
.I3(CLBLM_R_X3Y114_SLICE_X2Y114_AO6),
.I4(CLBLL_L_X2Y112_SLICE_X0Y112_BO6),
.I5(CLBLL_L_X2Y113_SLICE_X0Y113_BO6),
.O5(CLBLL_L_X2Y113_SLICE_X0Y113_DO5),
.O6(CLBLL_L_X2Y113_SLICE_X0Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0ff0f0f0e11e5a5a)
  ) CLBLL_L_X2Y113_SLICE_X0Y113_CLUT (
.I0(CLBLL_L_X2Y112_SLICE_X0Y112_AO6),
.I1(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I2(CLBLM_R_X3Y114_SLICE_X2Y114_AO6),
.I3(RIOB33_X105Y105_IOB_X1Y106_I),
.I4(LIOB33_X0Y101_IOB_X0Y101_I),
.I5(CLBLL_L_X2Y112_SLICE_X0Y112_BO6),
.O5(CLBLL_L_X2Y113_SLICE_X0Y113_CO5),
.O6(CLBLL_L_X2Y113_SLICE_X0Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555ffff99993333)
  ) CLBLL_L_X2Y113_SLICE_X0Y113_BLUT (
.I0(LIOB33_X0Y101_IOB_X0Y102_I),
.I1(CLBLL_L_X2Y113_SLICE_X0Y113_CO6),
.I2(1'b1),
.I3(1'b1),
.I4(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y113_SLICE_X0Y113_BO5),
.O6(CLBLL_L_X2Y113_SLICE_X0Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff05ff0fa5a50f0f)
  ) CLBLL_L_X2Y113_SLICE_X0Y113_ALUT (
.I0(LIOB33_X0Y101_IOB_X0Y101_I),
.I1(1'b1),
.I2(CLBLL_L_X2Y112_SLICE_X0Y112_AO6),
.I3(CLBLL_L_X2Y112_SLICE_X0Y112_BO6),
.I4(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y113_SLICE_X0Y113_AO5),
.O6(CLBLL_L_X2Y113_SLICE_X0Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h71f5f3ffd450fcf0)
  ) CLBLL_L_X2Y113_SLICE_X1Y113_DLUT (
.I0(LIOB33_X0Y103_IOB_X0Y104_I),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(CLBLL_L_X2Y113_SLICE_X0Y113_DO6),
.I3(LIOB33_X0Y101_IOB_X0Y102_I),
.I4(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I5(CLBLM_R_X3Y114_SLICE_X2Y114_BO6),
.O5(CLBLL_L_X2Y113_SLICE_X1Y113_DO5),
.O6(CLBLL_L_X2Y113_SLICE_X1Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7888877787777888)
  ) CLBLL_L_X2Y113_SLICE_X1Y113_CLUT (
.I0(LIOB33_X0Y103_IOB_X0Y104_I),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(LIOB33_X0Y105_IOB_X0Y105_I),
.I3(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I4(CLBLL_L_X2Y113_SLICE_X1Y113_DO6),
.I5(CLBLM_R_X3Y113_SLICE_X2Y113_CO6),
.O5(CLBLL_L_X2Y113_SLICE_X1Y113_CO5),
.O6(CLBLL_L_X2Y113_SLICE_X1Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h9c6339c6f00fff00)
  ) CLBLL_L_X2Y113_SLICE_X1Y113_BLUT (
.I0(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(CLBLL_L_X2Y113_SLICE_X0Y113_AO6),
.I3(CLBLM_R_X3Y114_SLICE_X2Y114_BO6),
.I4(CLBLM_R_X3Y113_SLICE_X2Y113_AO6),
.I5(LIOB33_X0Y101_IOB_X0Y102_I),
.O5(CLBLL_L_X2Y113_SLICE_X1Y113_BO5),
.O6(CLBLL_L_X2Y113_SLICE_X1Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf00f00ff3333ffff)
  ) CLBLL_L_X2Y113_SLICE_X1Y113_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I3(CLBLL_L_X2Y113_SLICE_X1Y113_BO6),
.I4(LIOB33_X0Y103_IOB_X0Y104_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y113_SLICE_X1Y113_AO5),
.O6(CLBLL_L_X2Y113_SLICE_X1Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y114_SLICE_X0Y114_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y114_SLICE_X0Y114_DO5),
.O6(CLBLL_L_X2Y114_SLICE_X0Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y114_SLICE_X0Y114_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y114_SLICE_X0Y114_CO5),
.O6(CLBLL_L_X2Y114_SLICE_X0Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555ffffaa00aa00)
  ) CLBLL_L_X2Y114_SLICE_X0Y114_BLUT (
.I0(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I1(1'b1),
.I2(1'b1),
.I3(RIOB33_X105Y111_IOB_X1Y112_I),
.I4(LIOB33_X0Y101_IOB_X0Y101_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y114_SLICE_X0Y114_BO5),
.O6(CLBLL_L_X2Y114_SLICE_X0Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hb5351f9f5f5f5f5f)
  ) CLBLL_L_X2Y114_SLICE_X0Y114_ALUT (
.I0(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(RIOB33_X105Y113_IOB_X1Y113_I),
.I3(RIOB33_X105Y111_IOB_X1Y112_I),
.I4(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y114_SLICE_X0Y114_AO5),
.O6(CLBLL_L_X2Y114_SLICE_X0Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y114_SLICE_X1Y114_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y114_SLICE_X1Y114_DO5),
.O6(CLBLL_L_X2Y114_SLICE_X1Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y114_SLICE_X1Y114_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y114_SLICE_X1Y114_CO5),
.O6(CLBLL_L_X2Y114_SLICE_X1Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y114_SLICE_X1Y114_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y114_SLICE_X1Y114_BO5),
.O6(CLBLL_L_X2Y114_SLICE_X1Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y114_SLICE_X1Y114_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y114_SLICE_X1Y114_AO5),
.O6(CLBLL_L_X2Y114_SLICE_X1Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y100_SLICE_X4Y100_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y100_SLICE_X4Y100_DO5),
.O6(CLBLL_L_X4Y100_SLICE_X4Y100_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haca06ca0906c9ca0)
  ) CLBLL_L_X4Y100_SLICE_X4Y100_CLUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(RIOB33_X105Y111_IOB_X1Y111_I),
.I2(RIOB33_X105Y109_IOB_X1Y110_I),
.I3(LIOB33_X0Y105_IOB_X0Y105_I),
.I4(LIOB33_X0Y103_IOB_X0Y104_I),
.I5(CLBLL_L_X4Y100_SLICE_X5Y100_AO6),
.O5(CLBLL_L_X4Y100_SLICE_X4Y100_CO5),
.O6(CLBLL_L_X4Y100_SLICE_X4Y100_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hce0871fff3ffffff)
  ) CLBLL_L_X4Y100_SLICE_X4Y100_BLUT (
.I0(LIOB33_X0Y103_IOB_X0Y104_I),
.I1(RIOB33_X105Y109_IOB_X1Y110_I),
.I2(CLBLL_L_X4Y100_SLICE_X5Y100_AO6),
.I3(LIOB33_X0Y105_IOB_X0Y105_I),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(RIOB33_X105Y111_IOB_X1Y111_I),
.O5(CLBLL_L_X4Y100_SLICE_X4Y100_BO5),
.O6(CLBLL_L_X4Y100_SLICE_X4Y100_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0ccccfff55ff55ff)
  ) CLBLL_L_X4Y100_SLICE_X4Y100_ALUT (
.I0(LIOB33_X0Y103_IOB_X0Y104_I),
.I1(CLBLL_L_X4Y100_SLICE_X5Y100_BO6),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(RIOB33_X105Y109_IOB_X1Y109_I),
.I4(CLBLL_L_X4Y100_SLICE_X4Y100_CO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y100_SLICE_X4Y100_AO5),
.O6(CLBLL_L_X4Y100_SLICE_X4Y100_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha7e1ff5f0f8fffff)
  ) CLBLL_L_X4Y100_SLICE_X5Y100_DLUT (
.I0(RIOB33_X105Y109_IOB_X1Y110_I),
.I1(LIOB33_X0Y101_IOB_X0Y101_I),
.I2(LIOB33_X0Y103_IOB_X0Y104_I),
.I3(CLBLM_R_X5Y103_SLICE_X6Y103_CO6),
.I4(RIOB33_X105Y111_IOB_X1Y111_I),
.I5(LIOB33_X0Y101_IOB_X0Y102_I),
.O5(CLBLL_L_X4Y100_SLICE_X5Y100_DO5),
.O6(CLBLL_L_X4Y100_SLICE_X5Y100_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h9c63c3c339c6cccc)
  ) CLBLL_L_X4Y100_SLICE_X5Y100_CLUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(CLBLL_L_X4Y100_SLICE_X4Y100_CO6),
.I2(CLBLM_R_X5Y101_SLICE_X7Y101_AO6),
.I3(LIOB33_X0Y107_IOB_X0Y107_I),
.I4(RIOB33_X105Y109_IOB_X1Y109_I),
.I5(CLBLM_R_X5Y100_SLICE_X6Y100_AO6),
.O5(CLBLL_L_X4Y100_SLICE_X5Y100_CO5),
.O6(CLBLL_L_X4Y100_SLICE_X5Y100_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7f15bf2abf2abf2a)
  ) CLBLL_L_X4Y100_SLICE_X5Y100_BLUT (
.I0(CLBLL_L_X4Y100_SLICE_X5Y100_DO6),
.I1(RIOB33_X105Y109_IOB_X1Y109_I),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(CLBLM_R_X5Y101_SLICE_X7Y101_AO6),
.I4(RIOB33_X105Y109_IOB_X1Y110_I),
.I5(LIOB33_X0Y105_IOB_X0Y105_I),
.O5(CLBLL_L_X4Y100_SLICE_X5Y100_BO5),
.O6(CLBLL_L_X4Y100_SLICE_X5Y100_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3fff7fff173f37ff)
  ) CLBLL_L_X4Y100_SLICE_X5Y100_ALUT (
.I0(LIOB33_X0Y103_IOB_X0Y104_I),
.I1(LIOB33_X0Y101_IOB_X0Y102_I),
.I2(RIOB33_X105Y111_IOB_X1Y111_I),
.I3(RIOB33_X105Y109_IOB_X1Y110_I),
.I4(LIOB33_X0Y101_IOB_X0Y101_I),
.I5(CLBLM_R_X5Y103_SLICE_X6Y103_CO6),
.O5(CLBLL_L_X4Y100_SLICE_X5Y100_AO5),
.O6(CLBLL_L_X4Y100_SLICE_X5Y100_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h37ff1377ffff3fff)
  ) CLBLL_L_X4Y101_SLICE_X4Y101_DLUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(LIOB33_X0Y105_IOB_X0Y105_I),
.I2(LIOB33_X0Y103_IOB_X0Y104_I),
.I3(RIOB33_X105Y111_IOB_X1Y111_I),
.I4(CLBLL_L_X4Y100_SLICE_X5Y100_AO6),
.I5(RIOB33_X105Y109_IOB_X1Y110_I),
.O5(CLBLL_L_X4Y101_SLICE_X4Y101_DO5),
.O6(CLBLL_L_X4Y101_SLICE_X4Y101_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h337f03077fff37ff)
  ) CLBLL_L_X4Y101_SLICE_X4Y101_CLUT (
.I0(LIOB33_X0Y111_IOB_X0Y111_I),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLL_L_X4Y101_SLICE_X5Y101_BO5),
.I3(LIOB33_X0Y111_IOB_X0Y112_I),
.I4(CLBLL_L_X4Y101_SLICE_X5Y101_CO5),
.I5(CLBLL_L_X4Y102_SLICE_X5Y102_BO6),
.O5(CLBLL_L_X4Y101_SLICE_X4Y101_CO5),
.O6(CLBLL_L_X4Y101_SLICE_X4Y101_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h9a6559a6f30cf30c)
  ) CLBLL_L_X4Y101_SLICE_X4Y101_BLUT (
.I0(LIOB33_X0Y111_IOB_X0Y112_I),
.I1(CLBLL_L_X4Y101_SLICE_X5Y101_BO5),
.I2(CLBLL_L_X4Y101_SLICE_X5Y101_CO5),
.I3(CLBLL_L_X4Y102_SLICE_X5Y102_BO6),
.I4(LIOB33_X0Y111_IOB_X0Y111_I),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLL_L_X4Y101_SLICE_X4Y101_BO5),
.O6(CLBLL_L_X4Y101_SLICE_X4Y101_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h7887877887877878)
  ) CLBLL_L_X4Y101_SLICE_X4Y101_ALUT (
.I0(RIOB33_X105Y109_IOB_X1Y109_I),
.I1(LIOB33_X0Y107_IOB_X0Y108_I),
.I2(CLBLL_L_X4Y100_SLICE_X4Y100_AO6),
.I3(LIOB33_X0Y107_IOB_X0Y107_I),
.I4(CLBLL_L_X4Y100_SLICE_X4Y100_BO6),
.I5(RIOB33_X105Y109_IOB_X1Y110_I),
.O5(CLBLL_L_X4Y101_SLICE_X4Y101_AO5),
.O6(CLBLL_L_X4Y101_SLICE_X4Y101_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hb42d4bd24bd2b42d)
  ) CLBLL_L_X4Y101_SLICE_X5Y101_DLUT (
.I0(CLBLM_R_X5Y101_SLICE_X6Y101_BO6),
.I1(CLBLM_R_X5Y102_SLICE_X6Y102_AO5),
.I2(CLBLL_L_X4Y101_SLICE_X5Y101_AO5),
.I3(CLBLL_L_X4Y101_SLICE_X5Y101_CO6),
.I4(CLBLM_R_X5Y101_SLICE_X6Y101_DO6),
.I5(CLBLL_L_X4Y101_SLICE_X5Y101_BO6),
.O5(CLBLL_L_X4Y101_SLICE_X5Y101_DO5),
.O6(CLBLL_L_X4Y101_SLICE_X5Y101_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c07f157f15)
  ) CLBLL_L_X4Y101_SLICE_X5Y101_CLUT (
.I0(CLBLM_R_X5Y101_SLICE_X6Y101_BO6),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(LIOB33_X0Y109_IOB_X0Y110_I),
.I3(CLBLM_R_X5Y102_SLICE_X6Y102_AO5),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y101_SLICE_X5Y101_CO5),
.O6(CLBLL_L_X4Y101_SLICE_X5Y101_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ffffff66999999)
  ) CLBLL_L_X4Y101_SLICE_X5Y101_BLUT (
.I0(CLBLM_R_X5Y101_SLICE_X6Y101_DO6),
.I1(CLBLL_L_X4Y101_SLICE_X5Y101_AO5),
.I2(1'b1),
.I3(LIOB33_X0Y109_IOB_X0Y110_I),
.I4(RIOB33_X105Y107_IOB_X1Y107_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y101_SLICE_X5Y101_BO5),
.O6(CLBLL_L_X4Y101_SLICE_X5Y101_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333ffff78877887)
  ) CLBLL_L_X4Y101_SLICE_X5Y101_ALUT (
.I0(LIOB33_X0Y109_IOB_X0Y109_I),
.I1(RIOB33_X105Y107_IOB_X1Y108_I),
.I2(CLBLL_L_X4Y101_SLICE_X4Y101_AO6),
.I3(CLBLM_R_X5Y100_SLICE_X6Y100_BO6),
.I4(LIOB33_X0Y101_IOB_X0Y101_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y101_SLICE_X5Y101_AO5),
.O6(CLBLL_L_X4Y101_SLICE_X5Y101_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h9a6559a6a5a5aaaa)
  ) CLBLL_L_X4Y102_SLICE_X4Y102_DLUT (
.I0(CLBLM_R_X3Y102_SLICE_X3Y102_BO6),
.I1(LIOB33_X0Y111_IOB_X0Y111_I),
.I2(CLBLL_L_X4Y102_SLICE_X5Y102_DO6),
.I3(LIOB33_X0Y111_IOB_X0Y112_I),
.I4(CLBLM_R_X3Y102_SLICE_X3Y102_CO6),
.I5(RIOB33_X105Y107_IOB_X1Y108_I),
.O5(CLBLL_L_X4Y102_SLICE_X4Y102_DO5),
.O6(CLBLL_L_X4Y102_SLICE_X4Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996969669696996)
  ) CLBLL_L_X4Y102_SLICE_X4Y102_CLUT (
.I0(CLBLL_L_X4Y102_SLICE_X4Y102_AO6),
.I1(CLBLM_R_X5Y102_SLICE_X6Y102_CO6),
.I2(CLBLL_L_X4Y106_SLICE_X4Y106_AO5),
.I3(CLBLL_L_X4Y102_SLICE_X4Y102_AO5),
.I4(CLBLM_R_X5Y103_SLICE_X6Y103_DO6),
.I5(CLBLL_L_X4Y102_SLICE_X4Y102_BO6),
.O5(CLBLL_L_X4Y102_SLICE_X4Y102_CO5),
.O6(CLBLL_L_X4Y102_SLICE_X4Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3cc3f00f96695aa5)
  ) CLBLL_L_X4Y102_SLICE_X4Y102_BLUT (
.I0(CLBLM_R_X5Y103_SLICE_X6Y103_DO6),
.I1(RIOB33_X105Y103_IOB_X1Y104_I),
.I2(CLBLM_R_X5Y102_SLICE_X6Y102_DO6),
.I3(CLBLM_R_X7Y102_SLICE_X9Y102_AO5),
.I4(LIOB33_X0Y109_IOB_X0Y110_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y102_SLICE_X4Y102_BO5),
.O6(CLBLL_L_X4Y102_SLICE_X4Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5f5f5f5f3f3f3f3f)
  ) CLBLL_L_X4Y102_SLICE_X4Y102_ALUT (
.I0(RIOB33_X105Y103_IOB_X1Y104_I),
.I1(RIOB33_X105Y103_IOB_X1Y103_I),
.I2(LIOB33_X0Y111_IOB_X0Y111_I),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y102_SLICE_X4Y102_AO5),
.O6(CLBLL_L_X4Y102_SLICE_X4Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h17ff03773fff1777)
  ) CLBLL_L_X4Y102_SLICE_X5Y102_DLUT (
.I0(CLBLL_L_X4Y101_SLICE_X4Y101_AO6),
.I1(CLBLM_R_X3Y101_SLICE_X3Y101_CO6),
.I2(LIOB33_X0Y109_IOB_X0Y110_I),
.I3(RIOB33_X105Y107_IOB_X1Y108_I),
.I4(CLBLM_R_X5Y100_SLICE_X6Y100_BO6),
.I5(LIOB33_X0Y109_IOB_X0Y109_I),
.O5(CLBLL_L_X4Y102_SLICE_X5Y102_DO5),
.O6(CLBLL_L_X4Y102_SLICE_X5Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8778e11eff0055aa)
  ) CLBLL_L_X4Y102_SLICE_X5Y102_CLUT (
.I0(CLBLL_L_X4Y101_SLICE_X4Y101_AO6),
.I1(LIOB33_X0Y109_IOB_X0Y109_I),
.I2(LIOB33_X0Y109_IOB_X0Y110_I),
.I3(CLBLM_R_X3Y101_SLICE_X3Y101_CO6),
.I4(CLBLM_R_X5Y100_SLICE_X6Y100_BO6),
.I5(RIOB33_X105Y107_IOB_X1Y108_I),
.O5(CLBLL_L_X4Y102_SLICE_X5Y102_CO5),
.O6(CLBLL_L_X4Y102_SLICE_X5Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hb4cc2dff4b33d200)
  ) CLBLL_L_X4Y102_SLICE_X5Y102_BLUT (
.I0(LIOB33_X0Y109_IOB_X0Y110_I),
.I1(CLBLM_R_X5Y101_SLICE_X6Y101_DO6),
.I2(LIOB33_X0Y111_IOB_X0Y111_I),
.I3(RIOB33_X105Y107_IOB_X1Y107_I),
.I4(CLBLL_L_X4Y101_SLICE_X5Y101_AO5),
.I5(CLBLL_L_X4Y102_SLICE_X5Y102_CO6),
.O5(CLBLL_L_X4Y102_SLICE_X5Y102_BO5),
.O6(CLBLL_L_X4Y102_SLICE_X5Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h04cc0dff4fffdfff)
  ) CLBLL_L_X4Y102_SLICE_X5Y102_ALUT (
.I0(LIOB33_X0Y109_IOB_X0Y110_I),
.I1(CLBLM_R_X5Y101_SLICE_X6Y101_DO6),
.I2(LIOB33_X0Y111_IOB_X0Y111_I),
.I3(RIOB33_X105Y107_IOB_X1Y107_I),
.I4(CLBLL_L_X4Y101_SLICE_X5Y101_AO5),
.I5(CLBLL_L_X4Y102_SLICE_X5Y102_CO6),
.O5(CLBLL_L_X4Y102_SLICE_X5Y102_AO5),
.O6(CLBLL_L_X4Y102_SLICE_X5Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f037f137f1fffff)
  ) CLBLL_L_X4Y103_SLICE_X4Y103_DLUT (
.I0(LIOB33_X0Y113_IOB_X0Y113_I),
.I1(CLBLL_L_X4Y103_SLICE_X5Y103_AO5),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLL_L_X4Y101_SLICE_X4Y101_CO6),
.I4(LIOB33_X0Y115_IOB_X0Y115_I),
.I5(CLBLL_L_X4Y103_SLICE_X4Y103_BO6),
.O5(CLBLL_L_X4Y103_SLICE_X4Y103_DO5),
.O6(CLBLL_L_X4Y103_SLICE_X4Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h233b2bff23bfafff)
  ) CLBLL_L_X4Y103_SLICE_X4Y103_CLUT (
.I0(CLBLL_L_X4Y102_SLICE_X5Y102_AO6),
.I1(RIOB33_X105Y107_IOB_X1Y107_I),
.I2(CLBLL_L_X4Y103_SLICE_X5Y103_BO5),
.I3(CLBLL_L_X4Y102_SLICE_X4Y102_DO6),
.I4(LIOB33_X0Y113_IOB_X0Y113_I),
.I5(LIOB33_X0Y111_IOB_X0Y112_I),
.O5(CLBLL_L_X4Y103_SLICE_X4Y103_CO5),
.O6(CLBLL_L_X4Y103_SLICE_X4Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h9f5fa39360a05c6c)
  ) CLBLL_L_X4Y103_SLICE_X4Y103_BLUT (
.I0(LIOB33_X0Y113_IOB_X0Y113_I),
.I1(CLBLL_L_X4Y103_SLICE_X5Y103_BO5),
.I2(RIOB33_X105Y107_IOB_X1Y107_I),
.I3(LIOB33_X0Y111_IOB_X0Y112_I),
.I4(CLBLL_L_X4Y102_SLICE_X5Y102_AO6),
.I5(CLBLL_L_X4Y102_SLICE_X4Y102_DO6),
.O5(CLBLL_L_X4Y103_SLICE_X4Y103_BO5),
.O6(CLBLL_L_X4Y103_SLICE_X4Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hb74877888b748778)
  ) CLBLL_L_X4Y103_SLICE_X4Y103_ALUT (
.I0(LIOB33_X0Y115_IOB_X0Y115_I),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLL_L_X4Y103_SLICE_X5Y103_AO5),
.I3(CLBLL_L_X4Y103_SLICE_X4Y103_BO6),
.I4(LIOB33_X0Y113_IOB_X0Y113_I),
.I5(CLBLL_L_X4Y101_SLICE_X4Y101_CO6),
.O5(CLBLL_L_X4Y103_SLICE_X4Y103_AO5),
.O6(CLBLL_L_X4Y103_SLICE_X4Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7bf31230ffff5af0)
  ) CLBLL_L_X4Y103_SLICE_X5Y103_DLUT (
.I0(LIOB33_X0Y111_IOB_X0Y111_I),
.I1(RIOB33_X105Y101_IOB_X1Y102_I),
.I2(CLBLL_L_X4Y102_SLICE_X4Y102_BO5),
.I3(RIOB33_X105Y103_IOB_X1Y103_I),
.I4(CLBLM_R_X5Y103_SLICE_X6Y103_AO6),
.I5(LIOB33_X0Y111_IOB_X0Y112_I),
.O5(CLBLL_L_X4Y103_SLICE_X5Y103_DO5),
.O6(CLBLL_L_X4Y103_SLICE_X5Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h69c3963ca50f5af0)
  ) CLBLL_L_X4Y103_SLICE_X5Y103_CLUT (
.I0(LIOB33_X0Y111_IOB_X0Y111_I),
.I1(RIOB33_X105Y101_IOB_X1Y102_I),
.I2(CLBLL_L_X4Y102_SLICE_X4Y102_BO5),
.I3(RIOB33_X105Y103_IOB_X1Y103_I),
.I4(CLBLM_R_X5Y103_SLICE_X6Y103_AO6),
.I5(LIOB33_X0Y111_IOB_X0Y112_I),
.O5(CLBLL_L_X4Y103_SLICE_X5Y103_CO5),
.O6(CLBLL_L_X4Y103_SLICE_X5Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h33ff33ff5aa5a5a5)
  ) CLBLL_L_X4Y103_SLICE_X5Y103_BLUT (
.I0(CLBLL_L_X4Y102_SLICE_X5Y102_DO6),
.I1(LIOB33_X0Y101_IOB_X0Y102_I),
.I2(CLBLM_R_X3Y102_SLICE_X3Y102_CO6),
.I3(RIOB33_X105Y107_IOB_X1Y108_I),
.I4(LIOB33_X0Y111_IOB_X0Y111_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y103_SLICE_X5Y103_BO5),
.O6(CLBLL_L_X4Y103_SLICE_X5Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ffffff69a569a5)
  ) CLBLL_L_X4Y103_SLICE_X5Y103_ALUT (
.I0(CLBLL_L_X4Y103_SLICE_X5Y103_BO5),
.I1(RIOB33_X105Y107_IOB_X1Y107_I),
.I2(CLBLL_L_X4Y102_SLICE_X5Y102_AO6),
.I3(LIOB33_X0Y111_IOB_X0Y112_I),
.I4(LIOB33_X0Y103_IOB_X0Y103_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y103_SLICE_X5Y103_AO5),
.O6(CLBLL_L_X4Y103_SLICE_X5Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5a96a56996a5695a)
  ) CLBLL_L_X4Y104_SLICE_X4Y104_DLUT (
.I0(CLBLL_L_X4Y103_SLICE_X5Y103_CO6),
.I1(CLBLL_L_X4Y104_SLICE_X5Y104_CO6),
.I2(CLBLL_L_X4Y104_SLICE_X5Y104_BO6),
.I3(CLBLL_L_X4Y105_SLICE_X4Y105_AO5),
.I4(CLBLM_R_X3Y103_SLICE_X3Y103_AO6),
.I5(CLBLL_L_X4Y104_SLICE_X4Y104_BO6),
.O5(CLBLL_L_X4Y104_SLICE_X4Y104_DO5),
.O6(CLBLL_L_X4Y104_SLICE_X4Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8778000087787887)
  ) CLBLL_L_X4Y104_SLICE_X4Y104_CLUT (
.I0(RIOB33_X105Y107_IOB_X1Y107_I),
.I1(LIOB33_X0Y115_IOB_X0Y115_I),
.I2(CLBLL_L_X4Y103_SLICE_X4Y103_CO6),
.I3(CLBLM_R_X3Y103_SLICE_X3Y103_AO5),
.I4(CLBLL_L_X4Y103_SLICE_X4Y103_DO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y104_SLICE_X4Y104_CO5),
.O6(CLBLL_L_X4Y104_SLICE_X4Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555ffff3cc3c3c3)
  ) CLBLL_L_X4Y104_SLICE_X4Y104_BLUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(CLBLL_L_X4Y103_SLICE_X5Y103_AO5),
.I2(CLBLL_L_X4Y101_SLICE_X4Y101_CO6),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(LIOB33_X0Y113_IOB_X0Y113_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y104_SLICE_X4Y104_BO5),
.O6(CLBLL_L_X4Y104_SLICE_X4Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h66cc993344ccddff)
  ) CLBLL_L_X4Y104_SLICE_X4Y104_ALUT (
.I0(LIOB33_X0Y113_IOB_X0Y113_I),
.I1(CLBLL_L_X4Y104_SLICE_X5Y104_BO6),
.I2(1'b1),
.I3(RIOB33_X105Y101_IOB_X1Y101_I),
.I4(CLBLL_L_X4Y103_SLICE_X5Y103_CO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y104_SLICE_X4Y104_AO5),
.O6(CLBLL_L_X4Y104_SLICE_X4Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y104_SLICE_X5Y104_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y104_SLICE_X5Y104_DO5),
.O6(CLBLL_L_X4Y104_SLICE_X5Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h718e8e718e71718e)
  ) CLBLL_L_X4Y104_SLICE_X5Y104_CLUT (
.I0(CLBLL_L_X4Y104_SLICE_X5Y104_AO6),
.I1(CLBLM_R_X5Y105_SLICE_X6Y105_AO6),
.I2(CLBLM_R_X7Y104_SLICE_X8Y104_AO6),
.I3(CLBLL_L_X4Y104_SLICE_X5Y104_AO5),
.I4(CLBLL_L_X4Y104_SLICE_X5Y104_BO5),
.I5(CLBLM_R_X5Y105_SLICE_X7Y105_CO6),
.O5(CLBLL_L_X4Y104_SLICE_X5Y104_CO5),
.O6(CLBLL_L_X4Y104_SLICE_X5Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h77ff007777777777)
  ) CLBLL_L_X4Y104_SLICE_X5Y104_BLUT (
.I0(RIOB33_X105Y101_IOB_X1Y101_I),
.I1(LIOB33_X0Y111_IOB_X0Y112_I),
.I2(1'b1),
.I3(CLBLM_R_X5Y104_SLICE_X6Y104_AO6),
.I4(CLBLM_R_X5Y104_SLICE_X6Y104_BO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y104_SLICE_X5Y104_BO5),
.O6(CLBLL_L_X4Y104_SLICE_X5Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h55ff55ff0fff0fff)
  ) CLBLL_L_X4Y104_SLICE_X5Y104_ALUT (
.I0(RIOB33_X105Y101_IOB_X1Y101_I),
.I1(1'b1),
.I2(RIOB33_X105Y101_IOB_X1Y102_I),
.I3(LIOB33_X0Y111_IOB_X0Y111_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y104_SLICE_X5Y104_AO5),
.O6(CLBLL_L_X4Y104_SLICE_X5Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hbc43708f3bc4f708)
  ) CLBLL_L_X4Y105_SLICE_X4Y105_DLUT (
.I0(LIOB33_X0Y111_IOB_X0Y112_I),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(CLBLL_L_X4Y105_SLICE_X5Y105_BO6),
.I3(CLBLL_L_X4Y104_SLICE_X5Y104_CO6),
.I4(LIOB33_X0Y113_IOB_X0Y113_I),
.I5(CLBLM_R_X5Y105_SLICE_X6Y105_CO6),
.O5(CLBLL_L_X4Y105_SLICE_X4Y105_DO5),
.O6(CLBLL_L_X4Y105_SLICE_X4Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6f06ff66cf0cffcc)
  ) CLBLL_L_X4Y105_SLICE_X4Y105_CLUT (
.I0(LIOB33_X0Y111_IOB_X0Y112_I),
.I1(CLBLL_L_X4Y105_SLICE_X5Y105_CO6),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(CLBLL_L_X4Y105_SLICE_X4Y105_AO5),
.I4(LIOB33_X0Y113_IOB_X0Y113_I),
.I5(RIOB33_X105Y101_IOB_X1Y101_I),
.O5(CLBLL_L_X4Y105_SLICE_X4Y105_CO5),
.O6(CLBLL_L_X4Y105_SLICE_X4Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hb44bc3c32dd2f0f0)
  ) CLBLL_L_X4Y105_SLICE_X4Y105_BLUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(CLBLL_L_X4Y105_SLICE_X5Y105_BO6),
.I2(CLBLL_L_X4Y105_SLICE_X5Y105_CO6),
.I3(RIOB33_X105Y101_IOB_X1Y101_I),
.I4(LIOB33_X0Y111_IOB_X0Y112_I),
.I5(CLBLM_R_X5Y105_SLICE_X6Y105_CO6),
.O5(CLBLL_L_X4Y105_SLICE_X4Y105_BO5),
.O6(CLBLL_L_X4Y105_SLICE_X4Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555ffff44ddccff)
  ) CLBLL_L_X4Y105_SLICE_X4Y105_ALUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(CLBLL_L_X4Y105_SLICE_X5Y105_BO6),
.I2(1'b1),
.I3(CLBLM_R_X5Y105_SLICE_X6Y105_CO6),
.I4(LIOB33_X0Y111_IOB_X0Y112_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y105_SLICE_X4Y105_AO5),
.O6(CLBLL_L_X4Y105_SLICE_X4Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y105_SLICE_X5Y105_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y105_SLICE_X5Y105_DO5),
.O6(CLBLL_L_X4Y105_SLICE_X5Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hd4bb2b442bbbd444)
  ) CLBLL_L_X4Y105_SLICE_X5Y105_CLUT (
.I0(CLBLM_R_X5Y105_SLICE_X6Y105_AO6),
.I1(CLBLM_R_X7Y104_SLICE_X8Y104_AO6),
.I2(RIOB33_X105Y101_IOB_X1Y101_I),
.I3(LIOB33_X0Y111_IOB_X0Y111_I),
.I4(CLBLM_R_X5Y105_SLICE_X7Y105_CO6),
.I5(RIOB33_X105Y101_IOB_X1Y102_I),
.O5(CLBLL_L_X4Y105_SLICE_X5Y105_CO5),
.O6(CLBLL_L_X4Y105_SLICE_X5Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7f13ff5fdf4c5f00)
  ) CLBLL_L_X4Y105_SLICE_X5Y105_BLUT (
.I0(LIOB33_X0Y111_IOB_X0Y111_I),
.I1(RIOB33_X105Y101_IOB_X1Y101_I),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(CLBLM_R_X5Y106_SLICE_X6Y106_BO6),
.I4(LIOB33_X0Y109_IOB_X0Y110_I),
.I5(CLBLM_R_X5Y106_SLICE_X6Y106_CO6),
.O5(CLBLL_L_X4Y105_SLICE_X5Y105_BO5),
.O6(CLBLL_L_X4Y105_SLICE_X5Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6c939393936c6c6c)
  ) CLBLL_L_X4Y105_SLICE_X5Y105_ALUT (
.I0(LIOB33_X0Y111_IOB_X0Y111_I),
.I1(CLBLM_R_X5Y106_SLICE_X6Y106_BO6),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(RIOB33_X105Y101_IOB_X1Y101_I),
.I4(LIOB33_X0Y109_IOB_X0Y110_I),
.I5(CLBLM_R_X5Y106_SLICE_X6Y106_CO6),
.O5(CLBLL_L_X4Y105_SLICE_X5Y105_AO5),
.O6(CLBLL_L_X4Y105_SLICE_X5Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y106_SLICE_X4Y106_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y106_SLICE_X4Y106_DO5),
.O6(CLBLL_L_X4Y106_SLICE_X4Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fbfbfbf152a2a2a)
  ) CLBLL_L_X4Y106_SLICE_X4Y106_CLUT (
.I0(CLBLM_R_X5Y106_SLICE_X7Y106_BO6),
.I1(LIOB33_X0Y115_IOB_X0Y116_I),
.I2(LIOB33_X0Y111_IOB_X0Y111_I),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(LIOB33_X0Y109_IOB_X0Y110_I),
.I5(CLBLM_R_X7Y106_SLICE_X8Y106_CO6),
.O5(CLBLL_L_X4Y106_SLICE_X4Y106_CO5),
.O6(CLBLL_L_X4Y106_SLICE_X4Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6c939393936c6c6c)
  ) CLBLL_L_X4Y106_SLICE_X4Y106_BLUT (
.I0(LIOB33_X0Y111_IOB_X0Y111_I),
.I1(CLBLM_R_X5Y106_SLICE_X7Y106_BO6),
.I2(LIOB33_X0Y115_IOB_X0Y116_I),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(LIOB33_X0Y109_IOB_X0Y110_I),
.I5(CLBLM_R_X7Y106_SLICE_X8Y106_CO6),
.O5(CLBLL_L_X4Y106_SLICE_X4Y106_BO5),
.O6(CLBLL_L_X4Y106_SLICE_X4Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0fffff7f137f13)
  ) CLBLL_L_X4Y106_SLICE_X4Y106_ALUT (
.I0(RIOB33_X105Y103_IOB_X1Y104_I),
.I1(CLBLM_R_X5Y102_SLICE_X6Y102_DO6),
.I2(LIOB33_X0Y109_IOB_X0Y110_I),
.I3(CLBLM_R_X7Y102_SLICE_X9Y102_AO5),
.I4(LIOB33_X0Y103_IOB_X0Y103_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y106_SLICE_X4Y106_AO5),
.O6(CLBLL_L_X4Y106_SLICE_X4Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y106_SLICE_X5Y106_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y106_SLICE_X5Y106_DO5),
.O6(CLBLL_L_X4Y106_SLICE_X5Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y106_SLICE_X5Y106_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y106_SLICE_X5Y106_CO5),
.O6(CLBLL_L_X4Y106_SLICE_X5Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y106_SLICE_X5Y106_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y106_SLICE_X5Y106_BO5),
.O6(CLBLL_L_X4Y106_SLICE_X5Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y106_SLICE_X5Y106_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y106_SLICE_X5Y106_AO5),
.O6(CLBLL_L_X4Y106_SLICE_X5Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y107_SLICE_X4Y107_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y107_SLICE_X4Y107_DO5),
.O6(CLBLL_L_X4Y107_SLICE_X4Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h373f7fff11153f7f)
  ) CLBLL_L_X4Y107_SLICE_X4Y107_CLUT (
.I0(CLBLL_L_X4Y106_SLICE_X4Y106_BO6),
.I1(LIOB33_X0Y113_IOB_X0Y114_I),
.I2(LIOB33_X0Y113_IOB_X0Y113_I),
.I3(LIOB33_X0Y111_IOB_X0Y112_I),
.I4(CLBLM_R_X5Y108_SLICE_X6Y108_DO6),
.I5(CLBLL_L_X4Y108_SLICE_X5Y108_BO6),
.O5(CLBLL_L_X4Y107_SLICE_X4Y107_CO5),
.O6(CLBLL_L_X4Y107_SLICE_X4Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h69963cc3c33c6996)
  ) CLBLL_L_X4Y107_SLICE_X4Y107_BLUT (
.I0(CLBLL_L_X2Y105_SLICE_X1Y105_AO6),
.I1(CLBLL_L_X4Y107_SLICE_X5Y107_BO6),
.I2(CLBLM_R_X3Y106_SLICE_X3Y106_AO6),
.I3(CLBLL_L_X4Y107_SLICE_X5Y107_AO6),
.I4(CLBLL_L_X4Y108_SLICE_X4Y108_AO6),
.I5(CLBLL_L_X4Y109_SLICE_X4Y109_CO6),
.O5(CLBLL_L_X4Y107_SLICE_X4Y107_BO5),
.O6(CLBLL_L_X4Y107_SLICE_X4Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h995599553f3f3f3f)
  ) CLBLL_L_X4Y107_SLICE_X4Y107_ALUT (
.I0(CLBLL_L_X4Y110_SLICE_X4Y110_BO6),
.I1(LIOB33_X0Y109_IOB_X0Y110_I),
.I2(LIOB33_X0Y113_IOB_X0Y114_I),
.I3(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y107_SLICE_X4Y107_AO5),
.O6(CLBLL_L_X4Y107_SLICE_X4Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h39c69c63c639639c)
  ) CLBLL_L_X4Y107_SLICE_X5Y107_DLUT (
.I0(CLBLM_R_X5Y107_SLICE_X6Y107_BO6),
.I1(CLBLM_R_X5Y107_SLICE_X7Y107_DO6),
.I2(CLBLL_L_X4Y107_SLICE_X5Y107_AO6),
.I3(CLBLL_L_X4Y107_SLICE_X5Y107_AO5),
.I4(CLBLL_L_X4Y108_SLICE_X4Y108_BO6),
.I5(CLBLL_L_X4Y103_SLICE_X5Y103_AO6),
.O5(CLBLL_L_X4Y107_SLICE_X5Y107_DO5),
.O6(CLBLL_L_X4Y107_SLICE_X5Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h2dd2b44bd22d4bb4)
  ) CLBLL_L_X4Y107_SLICE_X5Y107_CLUT (
.I0(CLBLM_R_X5Y107_SLICE_X6Y107_BO6),
.I1(CLBLL_L_X4Y107_SLICE_X5Y107_AO6),
.I2(CLBLM_R_X7Y106_SLICE_X8Y106_BO6),
.I3(CLBLL_L_X4Y107_SLICE_X5Y107_AO5),
.I4(CLBLL_L_X4Y108_SLICE_X4Y108_BO6),
.I5(CLBLM_R_X5Y107_SLICE_X7Y107_BO6),
.O5(CLBLL_L_X4Y107_SLICE_X5Y107_CO5),
.O6(CLBLL_L_X4Y107_SLICE_X5Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h2dd2b44bd22d4bb4)
  ) CLBLL_L_X4Y107_SLICE_X5Y107_BLUT (
.I0(CLBLM_R_X7Y108_SLICE_X8Y108_DO6),
.I1(CLBLL_L_X4Y109_SLICE_X5Y109_BO6),
.I2(CLBLM_R_X7Y107_SLICE_X8Y107_AO6),
.I3(CLBLL_L_X4Y107_SLICE_X4Y107_AO5),
.I4(CLBLL_L_X4Y106_SLICE_X4Y106_AO6),
.I5(CLBLM_R_X7Y108_SLICE_X8Y108_CO6),
.O5(CLBLL_L_X4Y107_SLICE_X5Y107_BO5),
.O6(CLBLL_L_X4Y107_SLICE_X5Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h33ff33ff00ffffff)
  ) CLBLL_L_X4Y107_SLICE_X5Y107_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y103_IOB_X0Y103_I),
.I2(1'b1),
.I3(LIOB33_X0Y111_IOB_X0Y111_I),
.I4(LIOB33_X0Y113_IOB_X0Y114_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y107_SLICE_X5Y107_AO5),
.O6(CLBLL_L_X4Y107_SLICE_X5Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h9c6339c6f50af50a)
  ) CLBLL_L_X4Y108_SLICE_X4Y108_DLUT (
.I0(CLBLL_L_X4Y106_SLICE_X4Y106_BO6),
.I1(LIOB33_X0Y115_IOB_X0Y116_I),
.I2(CLBLL_L_X4Y108_SLICE_X5Y108_BO6),
.I3(CLBLM_R_X5Y107_SLICE_X6Y107_CO6),
.I4(LIOB33_X0Y113_IOB_X0Y114_I),
.I5(LIOB33_X0Y111_IOB_X0Y112_I),
.O5(CLBLL_L_X4Y108_SLICE_X4Y108_DO5),
.O6(CLBLL_L_X4Y108_SLICE_X4Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fbfbfbf152a2a2a)
  ) CLBLL_L_X4Y108_SLICE_X4Y108_CLUT (
.I0(CLBLM_R_X5Y107_SLICE_X7Y107_AO6),
.I1(LIOB33_X0Y103_IOB_X0Y103_I),
.I2(LIOB33_X0Y111_IOB_X0Y111_I),
.I3(LIOB33_X0Y109_IOB_X0Y110_I),
.I4(LIOB33_X0Y113_IOB_X0Y114_I),
.I5(CLBLL_L_X4Y108_SLICE_X4Y108_BO6),
.O5(CLBLL_L_X4Y108_SLICE_X4Y108_CO5),
.O6(CLBLL_L_X4Y108_SLICE_X4Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h105175f7f7f7f7f7)
  ) CLBLL_L_X4Y108_SLICE_X4Y108_BLUT (
.I0(CLBLM_R_X7Y108_SLICE_X8Y108_DO6),
.I1(CLBLM_R_X5Y108_SLICE_X7Y108_BO6),
.I2(CLBLM_R_X5Y109_SLICE_X6Y109_DO6),
.I3(LIOB33_X0Y109_IOB_X0Y109_I),
.I4(LIOB33_X0Y109_IOB_X0Y110_I),
.I5(LIOB33_X0Y103_IOB_X0Y103_I),
.O5(CLBLL_L_X4Y108_SLICE_X4Y108_BO5),
.O6(CLBLL_L_X4Y108_SLICE_X4Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h9a5965a6a6a6a6a6)
  ) CLBLL_L_X4Y108_SLICE_X4Y108_ALUT (
.I0(CLBLM_R_X7Y108_SLICE_X8Y108_DO6),
.I1(CLBLM_R_X5Y108_SLICE_X7Y108_BO6),
.I2(CLBLM_R_X5Y109_SLICE_X6Y109_DO6),
.I3(LIOB33_X0Y109_IOB_X0Y109_I),
.I4(LIOB33_X0Y109_IOB_X0Y110_I),
.I5(LIOB33_X0Y103_IOB_X0Y103_I),
.O5(CLBLL_L_X4Y108_SLICE_X4Y108_AO5),
.O6(CLBLL_L_X4Y108_SLICE_X4Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h9cc663c639c6c6c6)
  ) CLBLL_L_X4Y108_SLICE_X5Y108_DLUT (
.I0(CLBLL_L_X4Y108_SLICE_X5Y108_AO6),
.I1(CLBLL_L_X4Y107_SLICE_X5Y107_DO6),
.I2(CLBLL_L_X4Y109_SLICE_X5Y109_CO6),
.I3(RIOB33_X105Y105_IOB_X1Y106_I),
.I4(LIOB33_X0Y113_IOB_X0Y113_I),
.I5(LIOB33_X0Y111_IOB_X0Y112_I),
.O5(CLBLL_L_X4Y108_SLICE_X5Y108_DO5),
.O6(CLBLL_L_X4Y108_SLICE_X5Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h69c39933963c66cc)
  ) CLBLL_L_X4Y108_SLICE_X5Y108_CLUT (
.I0(LIOB33_X0Y109_IOB_X0Y110_I),
.I1(CLBLM_R_X5Y107_SLICE_X7Y107_BO6),
.I2(LIOB33_X0Y111_IOB_X0Y111_I),
.I3(LIOB33_X0Y115_IOB_X0Y116_I),
.I4(LIOB33_X0Y113_IOB_X0Y114_I),
.I5(CLBLM_R_X7Y106_SLICE_X8Y106_DO6),
.O5(CLBLL_L_X4Y108_SLICE_X5Y108_CO5),
.O6(CLBLL_L_X4Y108_SLICE_X5Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6fffcfff06660ccc)
  ) CLBLL_L_X4Y108_SLICE_X5Y108_BLUT (
.I0(LIOB33_X0Y115_IOB_X0Y116_I),
.I1(CLBLM_R_X7Y106_SLICE_X8Y106_DO6),
.I2(LIOB33_X0Y111_IOB_X0Y111_I),
.I3(LIOB33_X0Y113_IOB_X0Y114_I),
.I4(LIOB33_X0Y109_IOB_X0Y110_I),
.I5(CLBLM_R_X5Y107_SLICE_X7Y107_BO6),
.O5(CLBLL_L_X4Y108_SLICE_X5Y108_BO5),
.O6(CLBLL_L_X4Y108_SLICE_X5Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h69969696c33c3c3c)
  ) CLBLL_L_X4Y108_SLICE_X5Y108_ALUT (
.I0(LIOB33_X0Y111_IOB_X0Y111_I),
.I1(CLBLL_L_X4Y108_SLICE_X4Y108_BO6),
.I2(CLBLM_R_X5Y107_SLICE_X7Y107_AO6),
.I3(LIOB33_X0Y113_IOB_X0Y114_I),
.I4(LIOB33_X0Y109_IOB_X0Y110_I),
.I5(LIOB33_X0Y103_IOB_X0Y103_I),
.O5(CLBLL_L_X4Y108_SLICE_X5Y108_AO5),
.O6(CLBLL_L_X4Y108_SLICE_X5Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hb4dd2ddd4b22d222)
  ) CLBLL_L_X4Y109_SLICE_X4Y109_DLUT (
.I0(CLBLL_L_X4Y108_SLICE_X5Y108_AO6),
.I1(CLBLL_L_X4Y109_SLICE_X5Y109_CO6),
.I2(LIOB33_X0Y103_IOB_X0Y103_I),
.I3(LIOB33_X0Y111_IOB_X0Y112_I),
.I4(RIOB33_X105Y105_IOB_X1Y106_I),
.I5(CLBLL_L_X4Y107_SLICE_X5Y107_CO6),
.O5(CLBLL_L_X4Y109_SLICE_X4Y109_DO5),
.O6(CLBLL_L_X4Y109_SLICE_X4Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h1171f3f37177ffff)
  ) CLBLL_L_X4Y109_SLICE_X4Y109_CLUT (
.I0(LIOB33_X0Y109_IOB_X0Y110_I),
.I1(CLBLL_L_X4Y109_SLICE_X5Y109_AO6),
.I2(CLBLL_L_X4Y110_SLICE_X4Y110_DO6),
.I3(LIOB33_X0Y109_IOB_X0Y109_I),
.I4(RIOB33_X105Y105_IOB_X1Y106_I),
.I5(CLBLM_R_X5Y109_SLICE_X6Y109_CO6),
.O5(CLBLL_L_X4Y109_SLICE_X4Y109_CO5),
.O6(CLBLL_L_X4Y109_SLICE_X4Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h69c39933963c66cc)
  ) CLBLL_L_X4Y109_SLICE_X4Y109_BLUT (
.I0(LIOB33_X0Y111_IOB_X0Y111_I),
.I1(CLBLM_R_X5Y108_SLICE_X6Y108_BO6),
.I2(LIOB33_X0Y109_IOB_X0Y110_I),
.I3(RIOB33_X105Y105_IOB_X1Y106_I),
.I4(LIOB33_X0Y103_IOB_X0Y103_I),
.I5(CLBLL_L_X4Y109_SLICE_X4Y109_CO6),
.O5(CLBLL_L_X4Y109_SLICE_X4Y109_BO5),
.O6(CLBLL_L_X4Y109_SLICE_X4Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hd24b2db4a5f0a5f0)
  ) CLBLL_L_X4Y109_SLICE_X4Y109_ALUT (
.I0(CLBLL_L_X4Y110_SLICE_X4Y110_DO6),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(CLBLM_R_X5Y109_SLICE_X6Y109_BO6),
.I3(CLBLM_R_X5Y109_SLICE_X6Y109_CO6),
.I4(LIOB33_X0Y103_IOB_X0Y103_I),
.I5(LIOB33_X0Y109_IOB_X0Y109_I),
.O5(CLBLL_L_X4Y109_SLICE_X4Y109_AO5),
.O6(CLBLL_L_X4Y109_SLICE_X4Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f057f157f1fffff)
  ) CLBLL_L_X4Y109_SLICE_X5Y109_DLUT (
.I0(CLBLL_L_X4Y108_SLICE_X5Y108_AO6),
.I1(LIOB33_X0Y111_IOB_X0Y112_I),
.I2(RIOB33_X105Y105_IOB_X1Y106_I),
.I3(CLBLL_L_X4Y109_SLICE_X5Y109_CO6),
.I4(LIOB33_X0Y113_IOB_X0Y113_I),
.I5(CLBLL_L_X4Y107_SLICE_X5Y107_DO6),
.O5(CLBLL_L_X4Y109_SLICE_X5Y109_DO5),
.O6(CLBLL_L_X4Y109_SLICE_X5Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h4dddcfff8eee0ccc)
  ) CLBLL_L_X4Y109_SLICE_X5Y109_CLUT (
.I0(LIOB33_X0Y109_IOB_X0Y110_I),
.I1(CLBLL_L_X4Y109_SLICE_X4Y109_CO6),
.I2(LIOB33_X0Y111_IOB_X0Y111_I),
.I3(RIOB33_X105Y105_IOB_X1Y106_I),
.I4(LIOB33_X0Y103_IOB_X0Y103_I),
.I5(CLBLM_R_X5Y108_SLICE_X6Y108_BO6),
.O5(CLBLL_L_X4Y109_SLICE_X5Y109_CO5),
.O6(CLBLL_L_X4Y109_SLICE_X5Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbf2b020b020fbf2)
  ) CLBLL_L_X4Y109_SLICE_X5Y109_BLUT (
.I0(CLBLM_R_X5Y110_SLICE_X6Y110_CO6),
.I1(CLBLM_R_X5Y110_SLICE_X7Y110_BO6),
.I2(CLBLM_R_X5Y108_SLICE_X6Y108_AO6),
.I3(CLBLM_R_X5Y109_SLICE_X6Y109_AO6),
.I4(CLBLM_R_X7Y108_SLICE_X8Y108_AO6),
.I5(CLBLM_R_X5Y111_SLICE_X7Y111_DO6),
.O5(CLBLL_L_X4Y109_SLICE_X5Y109_BO5),
.O6(CLBLL_L_X4Y109_SLICE_X5Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h4bd2b42db42d4bd2)
  ) CLBLL_L_X4Y109_SLICE_X5Y109_ALUT (
.I0(CLBLM_R_X5Y110_SLICE_X6Y110_CO6),
.I1(CLBLM_R_X5Y110_SLICE_X7Y110_BO6),
.I2(CLBLM_R_X7Y108_SLICE_X8Y108_AO6),
.I3(CLBLM_R_X5Y109_SLICE_X6Y109_AO6),
.I4(CLBLM_R_X5Y108_SLICE_X6Y108_AO6),
.I5(CLBLM_R_X5Y111_SLICE_X7Y111_DO6),
.O5(CLBLL_L_X4Y109_SLICE_X5Y109_AO5),
.O6(CLBLL_L_X4Y109_SLICE_X5Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7f13df4cdf4cdf4c)
  ) CLBLL_L_X4Y110_SLICE_X4Y110_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y106_I),
.I1(CLBLM_R_X5Y110_SLICE_X6Y110_AO6),
.I2(LIOB33_X0Y107_IOB_X0Y108_I),
.I3(CLBLL_L_X4Y111_SLICE_X4Y111_CO6),
.I4(LIOB33_X0Y103_IOB_X0Y103_I),
.I5(LIOB33_X0Y107_IOB_X0Y107_I),
.O5(CLBLL_L_X4Y110_SLICE_X4Y110_DO5),
.O6(CLBLL_L_X4Y110_SLICE_X4Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h577f5fff151f173f)
  ) CLBLL_L_X4Y110_SLICE_X4Y110_CLUT (
.I0(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I1(CLBLL_L_X4Y110_SLICE_X5Y110_AO6),
.I2(CLBLL_L_X4Y110_SLICE_X5Y110_DO6),
.I3(LIOB33_X0Y109_IOB_X0Y110_I),
.I4(LIOB33_X0Y109_IOB_X0Y109_I),
.I5(CLBLM_R_X3Y110_SLICE_X3Y110_AO6),
.O5(CLBLL_L_X4Y110_SLICE_X4Y110_CO5),
.O6(CLBLL_L_X4Y110_SLICE_X4Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h96cc66cc993c963c)
  ) CLBLL_L_X4Y110_SLICE_X4Y110_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y106_I),
.I1(CLBLL_L_X4Y110_SLICE_X5Y110_BO6),
.I2(CLBLL_L_X4Y110_SLICE_X5Y110_AO6),
.I3(LIOB33_X0Y109_IOB_X0Y109_I),
.I4(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I5(CLBLM_R_X3Y110_SLICE_X3Y110_AO6),
.O5(CLBLL_L_X4Y110_SLICE_X4Y110_BO5),
.O6(CLBLL_L_X4Y110_SLICE_X4Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h777777773cc3f00f)
  ) CLBLL_L_X4Y110_SLICE_X4Y110_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y106_I),
.I1(LIOB33_X0Y109_IOB_X0Y109_I),
.I2(CLBLL_L_X4Y110_SLICE_X5Y110_AO6),
.I3(CLBLM_R_X3Y110_SLICE_X3Y110_AO6),
.I4(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y110_SLICE_X4Y110_AO5),
.O6(CLBLL_L_X4Y110_SLICE_X4Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h399cc663c663399c)
  ) CLBLL_L_X4Y110_SLICE_X5Y110_DLUT (
.I0(CLBLL_L_X4Y110_SLICE_X5Y110_CO6),
.I1(CLBLM_R_X5Y111_SLICE_X7Y111_CO6),
.I2(CLBLM_R_X5Y109_SLICE_X6Y109_AO5),
.I3(CLBLL_L_X4Y111_SLICE_X4Y111_CO6),
.I4(CLBLM_R_X5Y109_SLICE_X6Y109_AO6),
.I5(CLBLL_L_X4Y110_SLICE_X4Y110_AO6),
.O5(CLBLL_L_X4Y110_SLICE_X5Y110_DO5),
.O6(CLBLL_L_X4Y110_SLICE_X5Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966999666699)
  ) CLBLL_L_X4Y110_SLICE_X5Y110_CLUT (
.I0(CLBLM_R_X5Y112_SLICE_X6Y112_DO6),
.I1(CLBLM_R_X3Y111_SLICE_X3Y111_AO5),
.I2(LIOB33_X0Y113_IOB_X0Y114_I),
.I3(CLBLM_R_X7Y111_SLICE_X8Y111_BO6),
.I4(CLBLL_L_X4Y111_SLICE_X5Y111_DO6),
.I5(LIOB33_X0Y105_IOB_X0Y106_I),
.O5(CLBLL_L_X4Y110_SLICE_X5Y110_CO5),
.O6(CLBLL_L_X4Y110_SLICE_X5Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h69965aa5a55a6996)
  ) CLBLL_L_X4Y110_SLICE_X5Y110_BLUT (
.I0(CLBLM_R_X5Y110_SLICE_X6Y110_CO6),
.I1(CLBLM_R_X5Y109_SLICE_X6Y109_AO5),
.I2(CLBLM_R_X5Y109_SLICE_X6Y109_AO6),
.I3(CLBLM_R_X5Y110_SLICE_X7Y110_BO6),
.I4(CLBLL_L_X4Y110_SLICE_X5Y110_CO6),
.I5(CLBLL_L_X4Y111_SLICE_X4Y111_CO6),
.O5(CLBLL_L_X4Y110_SLICE_X5Y110_BO5),
.O6(CLBLL_L_X4Y110_SLICE_X5Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6c939393936c6c6c)
  ) CLBLL_L_X4Y110_SLICE_X5Y110_ALUT (
.I0(LIOB33_X0Y107_IOB_X0Y108_I),
.I1(CLBLM_R_X5Y110_SLICE_X6Y110_AO6),
.I2(RIOB33_X105Y105_IOB_X1Y106_I),
.I3(LIOB33_X0Y103_IOB_X0Y103_I),
.I4(LIOB33_X0Y107_IOB_X0Y107_I),
.I5(CLBLL_L_X4Y111_SLICE_X4Y111_CO6),
.O5(CLBLL_L_X4Y110_SLICE_X5Y110_AO5),
.O6(CLBLL_L_X4Y110_SLICE_X5Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff8e8eff8e00008e)
  ) CLBLL_L_X4Y111_SLICE_X4Y111_DLUT (
.I0(CLBLM_R_X3Y112_SLICE_X3Y112_DO6),
.I1(CLBLM_R_X3Y111_SLICE_X3Y111_BO6),
.I2(CLBLL_L_X4Y112_SLICE_X5Y112_BO6),
.I3(CLBLL_L_X4Y112_SLICE_X5Y112_AO6),
.I4(CLBLM_R_X3Y111_SLICE_X3Y111_BO5),
.I5(CLBLM_R_X3Y111_SLICE_X3Y111_CO5),
.O5(CLBLL_L_X4Y111_SLICE_X4Y111_DO5),
.O6(CLBLL_L_X4Y111_SLICE_X4Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7dff143cf5ff50f0)
  ) CLBLL_L_X4Y111_SLICE_X4Y111_CLUT (
.I0(LIOB33_X0Y107_IOB_X0Y107_I),
.I1(LIOB33_X0Y103_IOB_X0Y103_I),
.I2(CLBLL_L_X4Y111_SLICE_X5Y111_BO6),
.I3(RIOB33_X105Y105_IOB_X1Y106_I),
.I4(CLBLL_L_X4Y111_SLICE_X4Y111_DO6),
.I5(LIOB33_X0Y105_IOB_X0Y106_I),
.O5(CLBLL_L_X4Y111_SLICE_X4Y111_CO5),
.O6(CLBLL_L_X4Y111_SLICE_X4Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h69969696c33c3c3c)
  ) CLBLL_L_X4Y111_SLICE_X4Y111_BLUT (
.I0(LIOB33_X0Y103_IOB_X0Y104_I),
.I1(CLBLL_L_X4Y112_SLICE_X5Y112_DO6),
.I2(CLBLL_L_X4Y111_SLICE_X5Y111_AO6),
.I3(LIOB33_X0Y103_IOB_X0Y103_I),
.I4(LIOB33_X0Y105_IOB_X0Y105_I),
.I5(LIOB33_X0Y113_IOB_X0Y114_I),
.O5(CLBLL_L_X4Y111_SLICE_X4Y111_BO5),
.O6(CLBLL_L_X4Y111_SLICE_X4Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc96c399c693c99cc)
  ) CLBLL_L_X4Y111_SLICE_X4Y111_ALUT (
.I0(CLBLL_L_X4Y112_SLICE_X4Y112_DO6),
.I1(CLBLL_L_X4Y111_SLICE_X5Y111_BO6),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(CLBLL_L_X4Y111_SLICE_X4Y111_BO6),
.I4(LIOB33_X0Y103_IOB_X0Y103_I),
.I5(RIOB33_X105Y105_IOB_X1Y106_I),
.O5(CLBLL_L_X4Y111_SLICE_X4Y111_AO5),
.O6(CLBLL_L_X4Y111_SLICE_X4Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'heafe80a880a8eafe)
  ) CLBLL_L_X4Y111_SLICE_X5Y111_DLUT (
.I0(CLBLM_R_X3Y111_SLICE_X3Y111_CO6),
.I1(CLBLL_L_X4Y112_SLICE_X5Y112_DO6),
.I2(CLBLM_R_X3Y111_SLICE_X3Y111_BO5),
.I3(CLBLL_L_X4Y111_SLICE_X5Y111_CO6),
.I4(CLBLM_R_X5Y112_SLICE_X7Y112_AO6),
.I5(CLBLM_R_X5Y112_SLICE_X6Y112_BO6),
.O5(CLBLL_L_X4Y111_SLICE_X5Y111_DO5),
.O6(CLBLL_L_X4Y111_SLICE_X5Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6c939393936c6c6c)
  ) CLBLL_L_X4Y111_SLICE_X5Y111_CLUT (
.I0(LIOB33_X0Y115_IOB_X0Y116_I),
.I1(CLBLM_R_X5Y111_SLICE_X6Y111_BO6),
.I2(LIOB33_X0Y101_IOB_X0Y102_I),
.I3(LIOB33_X0Y113_IOB_X0Y114_I),
.I4(LIOB33_X0Y103_IOB_X0Y104_I),
.I5(CLBLM_R_X5Y110_SLICE_X6Y110_BO6),
.O5(CLBLL_L_X4Y111_SLICE_X5Y111_CO5),
.O6(CLBLL_L_X4Y111_SLICE_X5Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h96c3cc333c96cccc)
  ) CLBLL_L_X4Y111_SLICE_X5Y111_BLUT (
.I0(LIOB33_X0Y103_IOB_X0Y103_I),
.I1(CLBLM_R_X5Y112_SLICE_X6Y112_BO6),
.I2(LIOB33_X0Y113_IOB_X0Y114_I),
.I3(CLBLL_L_X4Y112_SLICE_X5Y112_DO6),
.I4(LIOB33_X0Y105_IOB_X0Y105_I),
.I5(CLBLL_L_X4Y111_SLICE_X5Y111_CO6),
.O5(CLBLL_L_X4Y111_SLICE_X5Y111_BO5),
.O6(CLBLL_L_X4Y111_SLICE_X5Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc9396c9c69993ccc)
  ) CLBLL_L_X4Y111_SLICE_X5Y111_ALUT (
.I0(CLBLL_L_X4Y113_SLICE_X5Y113_AO5),
.I1(CLBLM_R_X5Y110_SLICE_X6Y110_BO6),
.I2(LIOB33_X0Y101_IOB_X0Y102_I),
.I3(LIOB33_X0Y115_IOB_X0Y116_I),
.I4(CLBLM_R_X5Y112_SLICE_X6Y112_AO6),
.I5(LIOB33_X0Y113_IOB_X0Y114_I),
.O5(CLBLL_L_X4Y111_SLICE_X5Y111_AO5),
.O6(CLBLL_L_X4Y111_SLICE_X5Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6c00ff6cff6cff6c)
  ) CLBLL_L_X4Y112_SLICE_X4Y112_DLUT (
.I0(LIOB33_X0Y103_IOB_X0Y104_I),
.I1(CLBLL_L_X4Y112_SLICE_X5Y112_CO6),
.I2(LIOB33_X0Y103_IOB_X0Y103_I),
.I3(CLBLM_R_X3Y112_SLICE_X3Y112_DO6),
.I4(LIOB33_X0Y105_IOB_X0Y105_I),
.I5(RIOB33_X105Y105_IOB_X1Y106_I),
.O5(CLBLL_L_X4Y112_SLICE_X4Y112_DO5),
.O6(CLBLL_L_X4Y112_SLICE_X4Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6c93936c936c936c)
  ) CLBLL_L_X4Y112_SLICE_X4Y112_CLUT (
.I0(LIOB33_X0Y103_IOB_X0Y104_I),
.I1(CLBLL_L_X4Y112_SLICE_X5Y112_CO6),
.I2(LIOB33_X0Y103_IOB_X0Y103_I),
.I3(CLBLM_R_X3Y112_SLICE_X3Y112_DO6),
.I4(LIOB33_X0Y105_IOB_X0Y105_I),
.I5(RIOB33_X105Y105_IOB_X1Y106_I),
.O5(CLBLL_L_X4Y112_SLICE_X4Y112_CO5),
.O6(CLBLL_L_X4Y112_SLICE_X4Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hd25a78f0b4961e3c)
  ) CLBLL_L_X4Y112_SLICE_X4Y112_BLUT (
.I0(LIOB33_X0Y105_IOB_X0Y105_I),
.I1(CLBLL_L_X4Y112_SLICE_X5Y112_BO6),
.I2(CLBLL_L_X4Y112_SLICE_X5Y112_AO6),
.I3(RIOB33_X105Y105_IOB_X1Y106_I),
.I4(LIOB33_X0Y103_IOB_X0Y103_I),
.I5(CLBLM_R_X3Y112_SLICE_X3Y112_DO6),
.O5(CLBLL_L_X4Y112_SLICE_X4Y112_BO5),
.O6(CLBLL_L_X4Y112_SLICE_X4Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0fff0fff55ff55ff)
  ) CLBLL_L_X4Y112_SLICE_X4Y112_ALUT (
.I0(LIOB33_X0Y113_IOB_X0Y114_I),
.I1(1'b1),
.I2(LIOB33_X0Y103_IOB_X0Y103_I),
.I3(LIOB33_X0Y103_IOB_X0Y104_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y112_SLICE_X4Y112_AO5),
.O6(CLBLL_L_X4Y112_SLICE_X4Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7ddd1444ffff3ccc)
  ) CLBLL_L_X4Y112_SLICE_X5Y112_DLUT (
.I0(LIOB33_X0Y103_IOB_X0Y103_I),
.I1(CLBLM_R_X5Y111_SLICE_X6Y111_CO6),
.I2(LIOB33_X0Y113_IOB_X0Y114_I),
.I3(LIOB33_X0Y101_IOB_X0Y102_I),
.I4(CLBLM_R_X3Y113_SLICE_X3Y113_CO6),
.I5(LIOB33_X0Y103_IOB_X0Y104_I),
.O5(CLBLL_L_X4Y112_SLICE_X5Y112_DO5),
.O6(CLBLL_L_X4Y112_SLICE_X5Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h9c6339c6c6c6c6c6)
  ) CLBLL_L_X4Y112_SLICE_X5Y112_CLUT (
.I0(CLBLL_L_X4Y113_SLICE_X5Y113_AO6),
.I1(CLBLM_R_X5Y111_SLICE_X6Y111_CO6),
.I2(CLBLM_R_X3Y113_SLICE_X2Y113_BO5),
.I3(LIOB33_X0Y113_IOB_X0Y114_I),
.I4(LIOB33_X0Y103_IOB_X0Y103_I),
.I5(LIOB33_X0Y101_IOB_X0Y102_I),
.O5(CLBLL_L_X4Y112_SLICE_X5Y112_CO5),
.O6(CLBLL_L_X4Y112_SLICE_X5Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6c939393936c6c6c)
  ) CLBLL_L_X4Y112_SLICE_X5Y112_BLUT (
.I0(LIOB33_X0Y101_IOB_X0Y102_I),
.I1(CLBLM_R_X5Y111_SLICE_X6Y111_CO6),
.I2(LIOB33_X0Y113_IOB_X0Y114_I),
.I3(LIOB33_X0Y103_IOB_X0Y104_I),
.I4(LIOB33_X0Y103_IOB_X0Y103_I),
.I5(CLBLM_R_X3Y113_SLICE_X3Y113_CO6),
.O5(CLBLL_L_X4Y112_SLICE_X5Y112_BO5),
.O6(CLBLL_L_X4Y112_SLICE_X5Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6966969999696696)
  ) CLBLL_L_X4Y112_SLICE_X5Y112_ALUT (
.I0(CLBLL_L_X4Y112_SLICE_X4Y112_AO5),
.I1(CLBLM_R_X5Y113_SLICE_X6Y113_BO6),
.I2(CLBLL_L_X4Y112_SLICE_X4Y112_AO6),
.I3(CLBLM_R_X5Y111_SLICE_X6Y111_AO6),
.I4(CLBLM_R_X5Y111_SLICE_X6Y111_BO6),
.I5(CLBLM_R_X3Y113_SLICE_X3Y113_CO6),
.O5(CLBLL_L_X4Y112_SLICE_X5Y112_AO5),
.O6(CLBLL_L_X4Y112_SLICE_X5Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y113_SLICE_X4Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y113_SLICE_X4Y113_DO5),
.O6(CLBLL_L_X4Y113_SLICE_X4Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y113_SLICE_X4Y113_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y113_SLICE_X4Y113_CO5),
.O6(CLBLL_L_X4Y113_SLICE_X4Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y113_SLICE_X4Y113_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y113_SLICE_X4Y113_BO5),
.O6(CLBLL_L_X4Y113_SLICE_X4Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3545303040404040)
  ) CLBLL_L_X4Y113_SLICE_X4Y113_ALUT (
.I0(LIOB33_X0Y103_IOB_X0Y103_I),
.I1(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I2(LIOB33_X0Y113_IOB_X0Y114_I),
.I3(RIOB33_X105Y111_IOB_X1Y112_I),
.I4(LIOB33_X0Y115_IOB_X0Y116_I),
.I5(RIOB33_X105Y113_IOB_X1Y113_I),
.O5(CLBLL_L_X4Y113_SLICE_X4Y113_AO5),
.O6(CLBLL_L_X4Y113_SLICE_X4Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y113_SLICE_X5Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y113_SLICE_X5Y113_DO5),
.O6(CLBLL_L_X4Y113_SLICE_X5Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y113_SLICE_X5Y113_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y113_SLICE_X5Y113_CO5),
.O6(CLBLL_L_X4Y113_SLICE_X5Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y113_SLICE_X5Y113_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y113_SLICE_X5Y113_BO5),
.O6(CLBLL_L_X4Y113_SLICE_X5Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa555555f0f5f5f5)
  ) CLBLL_L_X4Y113_SLICE_X5Y113_ALUT (
.I0(CLBLM_R_X3Y111_SLICE_X2Y111_AO6),
.I1(1'b1),
.I2(CLBLM_R_X3Y111_SLICE_X3Y111_DO6),
.I3(LIOB33_X0Y101_IOB_X0Y101_I),
.I4(LIOB33_X0Y113_IOB_X0Y114_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y113_SLICE_X5Y113_AO5),
.O6(CLBLL_L_X4Y113_SLICE_X5Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6969666996969996)
  ) CLBLM_L_X8Y100_SLICE_X10Y100_DLUT (
.I0(CLBLL_L_X4Y103_SLICE_X5Y103_BO6),
.I1(CLBLM_L_X8Y100_SLICE_X11Y100_CO6),
.I2(CLBLM_L_X8Y100_SLICE_X11Y100_DO6),
.I3(CLBLL_L_X4Y101_SLICE_X5Y101_AO6),
.I4(CLBLM_L_X8Y102_SLICE_X10Y102_DO6),
.I5(CLBLM_R_X3Y100_SLICE_X3Y100_AO6),
.O5(CLBLM_L_X8Y100_SLICE_X10Y100_DO5),
.O6(CLBLM_L_X8Y100_SLICE_X10Y100_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'he8e8eee8b2b2bbb2)
  ) CLBLM_L_X8Y100_SLICE_X10Y100_CLUT (
.I0(CLBLL_L_X4Y103_SLICE_X5Y103_BO6),
.I1(CLBLM_L_X8Y100_SLICE_X11Y100_CO6),
.I2(CLBLM_L_X8Y100_SLICE_X11Y100_DO6),
.I3(CLBLL_L_X4Y101_SLICE_X5Y101_AO6),
.I4(CLBLM_L_X8Y102_SLICE_X10Y102_DO6),
.I5(CLBLM_R_X3Y100_SLICE_X3Y100_AO6),
.O5(CLBLM_L_X8Y100_SLICE_X10Y100_CO5),
.O6(CLBLM_L_X8Y100_SLICE_X10Y100_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha569695ac3c3f0f0)
  ) CLBLM_L_X8Y100_SLICE_X10Y100_BLUT (
.I0(RIOB33_X105Y107_IOB_X1Y108_I),
.I1(CLBLM_L_X8Y102_SLICE_X10Y102_AO5),
.I2(CLBLM_L_X8Y100_SLICE_X11Y100_AO6),
.I3(RIOB33_X105Y107_IOB_X1Y107_I),
.I4(CLBLM_L_X8Y100_SLICE_X10Y100_AO6),
.I5(LIOB33_X0Y101_IOB_X0Y102_I),
.O5(CLBLM_L_X8Y100_SLICE_X10Y100_BO5),
.O6(CLBLM_L_X8Y100_SLICE_X10Y100_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa5500ffccddccff)
  ) CLBLM_L_X8Y100_SLICE_X10Y100_ALUT (
.I0(RIOB33_X105Y107_IOB_X1Y108_I),
.I1(CLBLM_L_X8Y100_SLICE_X11Y100_DO6),
.I2(1'b1),
.I3(CLBLM_L_X8Y102_SLICE_X10Y102_DO6),
.I4(LIOB33_X0Y101_IOB_X0Y101_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y100_SLICE_X10Y100_AO5),
.O6(CLBLM_L_X8Y100_SLICE_X10Y100_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00006e448088a288)
  ) CLBLM_L_X8Y100_SLICE_X11Y100_DLUT (
.I0(RIOB33_X105Y113_IOB_X1Y113_I),
.I1(RIOB33_X105Y109_IOB_X1Y109_I),
.I2(RIOB33_X105Y111_IOB_X1Y112_I),
.I3(RIOB33_X105Y109_IOB_X1Y110_I),
.I4(RIOB33_X105Y107_IOB_X1Y108_I),
.I5(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.O5(CLBLM_L_X8Y100_SLICE_X11Y100_DO5),
.O6(CLBLM_L_X8Y100_SLICE_X11Y100_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hec99e6335fdd5577)
  ) CLBLM_L_X8Y100_SLICE_X11Y100_CLUT (
.I0(RIOB33_X105Y113_IOB_X1Y113_I),
.I1(RIOB33_X105Y109_IOB_X1Y109_I),
.I2(RIOB33_X105Y111_IOB_X1Y112_I),
.I3(RIOB33_X105Y109_IOB_X1Y110_I),
.I4(RIOB33_X105Y111_IOB_X1Y111_I),
.I5(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.O5(CLBLM_L_X8Y100_SLICE_X11Y100_CO5),
.O6(CLBLM_L_X8Y100_SLICE_X11Y100_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha05f030fb00f333f)
  ) CLBLM_L_X8Y100_SLICE_X11Y100_BLUT (
.I0(RIOB33_X105Y111_IOB_X1Y112_I),
.I1(RIOB33_X105Y109_IOB_X1Y109_I),
.I2(RIOB33_X105Y113_IOB_X1Y113_I),
.I3(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I4(RIOB33_X105Y109_IOB_X1Y110_I),
.I5(RIOB33_X105Y111_IOB_X1Y111_I),
.O5(CLBLM_L_X8Y100_SLICE_X11Y100_BO5),
.O6(CLBLM_L_X8Y100_SLICE_X11Y100_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0fe3ff13f01c00ec)
  ) CLBLM_L_X8Y100_SLICE_X11Y100_ALUT (
.I0(RIOB33_X105Y107_IOB_X1Y108_I),
.I1(CLBLM_L_X8Y102_SLICE_X10Y102_DO6),
.I2(LIOB33_X0Y101_IOB_X0Y101_I),
.I3(CLBLM_L_X8Y100_SLICE_X11Y100_DO6),
.I4(RIOB33_X105Y109_IOB_X1Y109_I),
.I5(CLBLM_L_X8Y100_SLICE_X11Y100_CO6),
.O5(CLBLM_L_X8Y100_SLICE_X11Y100_AO5),
.O6(CLBLM_L_X8Y100_SLICE_X11Y100_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996969699666666)
  ) CLBLM_L_X8Y101_SLICE_X10Y101_DLUT (
.I0(CLBLM_L_X8Y100_SLICE_X11Y100_AO6),
.I1(CLBLM_L_X10Y102_SLICE_X12Y102_DO6),
.I2(RIOB33_X105Y107_IOB_X1Y107_I),
.I3(LIOB33_X0Y101_IOB_X0Y102_I),
.I4(RIOB33_X105Y107_IOB_X1Y108_I),
.I5(LIOB33_X0Y103_IOB_X0Y104_I),
.O5(CLBLM_L_X8Y101_SLICE_X10Y101_DO5),
.O6(CLBLM_L_X8Y101_SLICE_X10Y101_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h48dedede88eeeeee)
  ) CLBLM_L_X8Y101_SLICE_X10Y101_CLUT (
.I0(CLBLM_L_X8Y100_SLICE_X11Y100_AO6),
.I1(CLBLM_L_X10Y102_SLICE_X12Y102_DO6),
.I2(RIOB33_X105Y107_IOB_X1Y108_I),
.I3(LIOB33_X0Y103_IOB_X0Y104_I),
.I4(RIOB33_X105Y107_IOB_X1Y107_I),
.I5(LIOB33_X0Y101_IOB_X0Y102_I),
.O5(CLBLM_L_X8Y101_SLICE_X10Y101_CO5),
.O6(CLBLM_L_X8Y101_SLICE_X10Y101_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'he74d18b265cf9a30)
  ) CLBLM_L_X8Y101_SLICE_X10Y101_BLUT (
.I0(RIOB33_X105Y107_IOB_X1Y108_I),
.I1(CLBLM_L_X8Y100_SLICE_X10Y100_AO5),
.I2(CLBLM_L_X8Y101_SLICE_X11Y101_AO6),
.I3(LIOB33_X0Y103_IOB_X0Y104_I),
.I4(CLBLM_L_X8Y101_SLICE_X11Y101_CO6),
.I5(LIOB33_X0Y101_IOB_X0Y102_I),
.O5(CLBLM_L_X8Y101_SLICE_X10Y101_BO5),
.O6(CLBLM_L_X8Y101_SLICE_X10Y101_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h008c0000738cc0c0)
  ) CLBLM_L_X8Y101_SLICE_X10Y101_ALUT (
.I0(RIOB33_X105Y111_IOB_X1Y112_I),
.I1(RIOB33_X105Y113_IOB_X1Y113_I),
.I2(RIOB33_X105Y109_IOB_X1Y109_I),
.I3(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I4(RIOB33_X105Y107_IOB_X1Y108_I),
.I5(RIOB33_X105Y107_IOB_X1Y107_I),
.O5(CLBLM_L_X8Y101_SLICE_X10Y101_AO5),
.O6(CLBLM_L_X8Y101_SLICE_X10Y101_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h9966f708cccc0000)
  ) CLBLM_L_X8Y101_SLICE_X11Y101_DLUT (
.I0(RIOB33_X105Y113_IOB_X1Y113_I),
.I1(RIOB33_X105Y111_IOB_X1Y111_I),
.I2(RIOB33_X105Y111_IOB_X1Y112_I),
.I3(LIOB33_X0Y101_IOB_X0Y101_I),
.I4(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I5(RIOB33_X105Y109_IOB_X1Y110_I),
.O5(CLBLM_L_X8Y101_SLICE_X11Y101_DO5),
.O6(CLBLM_L_X8Y101_SLICE_X11Y101_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h33c9cc36ff5500aa)
  ) CLBLM_L_X8Y101_SLICE_X11Y101_CLUT (
.I0(CLBLM_L_X8Y100_SLICE_X11Y100_CO6),
.I1(LIOB33_X0Y101_IOB_X0Y102_I),
.I2(LIOB33_X0Y101_IOB_X0Y101_I),
.I3(CLBLM_L_X8Y100_SLICE_X11Y100_BO6),
.I4(CLBLM_L_X8Y101_SLICE_X11Y101_DO6),
.I5(RIOB33_X105Y109_IOB_X1Y109_I),
.O5(CLBLM_L_X8Y101_SLICE_X11Y101_CO5),
.O6(CLBLM_L_X8Y101_SLICE_X11Y101_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h50f551fff5f5f7ff)
  ) CLBLM_L_X8Y101_SLICE_X11Y101_BLUT (
.I0(CLBLM_L_X8Y101_SLICE_X11Y101_DO6),
.I1(LIOB33_X0Y101_IOB_X0Y101_I),
.I2(CLBLM_L_X8Y100_SLICE_X11Y100_BO6),
.I3(RIOB33_X105Y109_IOB_X1Y109_I),
.I4(CLBLM_L_X8Y100_SLICE_X11Y100_CO6),
.I5(LIOB33_X0Y101_IOB_X0Y102_I),
.O5(CLBLM_L_X8Y101_SLICE_X11Y101_BO5),
.O6(CLBLM_L_X8Y101_SLICE_X11Y101_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf00f00ff95959595)
  ) CLBLM_L_X8Y101_SLICE_X11Y101_ALUT (
.I0(CLBLM_L_X10Y104_SLICE_X13Y104_AO6),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(LIOB33_X0Y101_IOB_X0Y101_I),
.I3(CLBLM_L_X8Y100_SLICE_X11Y100_CO6),
.I4(RIOB33_X105Y109_IOB_X1Y109_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y101_SLICE_X11Y101_AO5),
.O6(CLBLM_L_X8Y101_SLICE_X11Y101_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h075a8d00705afa00)
  ) CLBLM_L_X8Y102_SLICE_X10Y102_DLUT (
.I0(RIOB33_X105Y109_IOB_X1Y109_I),
.I1(RIOB33_X105Y111_IOB_X1Y112_I),
.I2(RIOB33_X105Y107_IOB_X1Y108_I),
.I3(RIOB33_X105Y113_IOB_X1Y113_I),
.I4(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I5(RIOB33_X105Y109_IOB_X1Y110_I),
.O5(CLBLM_L_X8Y102_SLICE_X10Y102_DO5),
.O6(CLBLM_L_X8Y102_SLICE_X10Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h639cc6399c6339c6)
  ) CLBLM_L_X8Y102_SLICE_X10Y102_CLUT (
.I0(CLBLM_L_X10Y102_SLICE_X12Y102_AO5),
.I1(CLBLM_L_X8Y101_SLICE_X11Y101_CO6),
.I2(CLBLM_L_X8Y100_SLICE_X10Y100_DO6),
.I3(CLBLM_L_X8Y103_SLICE_X11Y103_AO5),
.I4(CLBLM_L_X10Y102_SLICE_X12Y102_DO6),
.I5(CLBLM_L_X8Y100_SLICE_X10Y100_CO6),
.O5(CLBLM_L_X8Y102_SLICE_X10Y102_CO5),
.O6(CLBLM_L_X8Y102_SLICE_X10Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h60f6f6f6c0fcfcfc)
  ) CLBLM_L_X8Y102_SLICE_X10Y102_BLUT (
.I0(LIOB33_X0Y103_IOB_X0Y104_I),
.I1(CLBLM_L_X8Y100_SLICE_X10Y100_BO6),
.I2(CLBLM_L_X8Y102_SLICE_X11Y102_CO6),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(LIOB33_X0Y105_IOB_X0Y105_I),
.I5(RIOB33_X105Y107_IOB_X1Y107_I),
.O5(CLBLM_L_X8Y102_SLICE_X10Y102_BO5),
.O6(CLBLM_L_X8Y102_SLICE_X10Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc30fc30fffff030f)
  ) CLBLM_L_X8Y102_SLICE_X10Y102_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y101_IOB_X0Y101_I),
.I2(CLBLM_L_X10Y102_SLICE_X13Y102_AO6),
.I3(RIOB33_X105Y107_IOB_X1Y107_I),
.I4(CLBLM_L_X8Y101_SLICE_X10Y101_AO6),
.I5(1'b1),
.O5(CLBLM_L_X8Y102_SLICE_X10Y102_AO5),
.O6(CLBLM_L_X8Y102_SLICE_X10Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6969a5a5783cb4f0)
  ) CLBLM_L_X8Y102_SLICE_X11Y102_DLUT (
.I0(CLBLM_L_X8Y101_SLICE_X10Y101_AO6),
.I1(LIOB33_X0Y101_IOB_X0Y101_I),
.I2(CLBLM_L_X8Y102_SLICE_X10Y102_DO6),
.I3(RIOB33_X105Y107_IOB_X1Y107_I),
.I4(RIOB33_X105Y107_IOB_X1Y108_I),
.I5(CLBLM_L_X10Y102_SLICE_X13Y102_AO6),
.O5(CLBLM_L_X8Y102_SLICE_X11Y102_DO5),
.O6(CLBLM_L_X8Y102_SLICE_X11Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h4cdfdf4cdfdf4c4c)
  ) CLBLM_L_X8Y102_SLICE_X11Y102_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X10Y103_SLICE_X13Y103_CO6),
.I2(LIOB33_X0Y103_IOB_X0Y104_I),
.I3(RIOB33_X105Y107_IOB_X1Y107_I),
.I4(CLBLM_L_X8Y102_SLICE_X11Y102_DO6),
.I5(LIOB33_X0Y101_IOB_X0Y102_I),
.O5(CLBLM_L_X8Y102_SLICE_X11Y102_CO5),
.O6(CLBLM_L_X8Y102_SLICE_X11Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h95a9aa5a6a56aa5a)
  ) CLBLM_L_X8Y102_SLICE_X11Y102_BLUT (
.I0(CLBLM_L_X8Y102_SLICE_X11Y102_DO6),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_L_X8Y102_SLICE_X10Y102_AO6),
.I3(CLBLM_L_X8Y103_SLICE_X11Y103_BO6),
.I4(LIOB33_X0Y101_IOB_X0Y102_I),
.I5(RIOB33_X105Y107_IOB_X1Y107_I),
.O5(CLBLM_L_X8Y102_SLICE_X11Y102_BO5),
.O6(CLBLM_L_X8Y102_SLICE_X11Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6999966696669666)
  ) CLBLM_L_X8Y102_SLICE_X11Y102_ALUT (
.I0(CLBLM_L_X8Y102_SLICE_X11Y102_DO6),
.I1(CLBLM_L_X10Y103_SLICE_X13Y103_CO6),
.I2(RIOB33_X105Y107_IOB_X1Y107_I),
.I3(LIOB33_X0Y101_IOB_X0Y102_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(LIOB33_X0Y103_IOB_X0Y104_I),
.O5(CLBLM_L_X8Y102_SLICE_X11Y102_AO5),
.O6(CLBLM_L_X8Y102_SLICE_X11Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hee8e8e88bb2b2b22)
  ) CLBLM_L_X8Y103_SLICE_X10Y103_DLUT (
.I0(CLBLM_L_X8Y103_SLICE_X10Y103_AO6),
.I1(CLBLM_L_X8Y102_SLICE_X10Y102_CO6),
.I2(CLBLM_L_X8Y101_SLICE_X10Y101_DO6),
.I3(CLBLM_L_X8Y103_SLICE_X10Y103_AO5),
.I4(CLBLM_L_X8Y102_SLICE_X11Y102_CO6),
.I5(CLBLM_R_X7Y100_SLICE_X8Y100_AO5),
.O5(CLBLM_L_X8Y103_SLICE_X10Y103_DO5),
.O6(CLBLM_L_X8Y103_SLICE_X10Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hc639639caf50af50)
  ) CLBLM_L_X8Y103_SLICE_X10Y103_CLUT (
.I0(CLBLM_L_X8Y102_SLICE_X11Y102_CO6),
.I1(RIOB33_X105Y107_IOB_X1Y107_I),
.I2(CLBLM_L_X8Y101_SLICE_X10Y101_DO6),
.I3(CLBLM_L_X8Y102_SLICE_X10Y102_CO6),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(LIOB33_X0Y105_IOB_X0Y105_I),
.O5(CLBLM_L_X8Y103_SLICE_X10Y103_CO5),
.O6(CLBLM_L_X8Y103_SLICE_X10Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h39c6c6399c63639c)
  ) CLBLM_L_X8Y103_SLICE_X10Y103_BLUT (
.I0(CLBLM_L_X8Y101_SLICE_X10Y101_DO6),
.I1(CLBLM_R_X7Y100_SLICE_X8Y100_AO5),
.I2(CLBLM_L_X8Y102_SLICE_X11Y102_CO6),
.I3(CLBLM_L_X8Y102_SLICE_X10Y102_CO6),
.I4(CLBLM_L_X8Y103_SLICE_X10Y103_AO6),
.I5(CLBLM_L_X8Y103_SLICE_X10Y103_AO5),
.O5(CLBLM_L_X8Y103_SLICE_X10Y103_BO5),
.O6(CLBLM_L_X8Y103_SLICE_X10Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f3f3f3f33ff33ff)
  ) CLBLM_L_X8Y103_SLICE_X10Y103_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(LIOB33_X0Y105_IOB_X0Y105_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y103_SLICE_X10Y103_AO5),
.O6(CLBLM_L_X8Y103_SLICE_X10Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hdf0fdf0f5f5f5f5f)
  ) CLBLM_L_X8Y103_SLICE_X11Y103_DLUT (
.I0(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I1(RIOB33_X105Y111_IOB_X1Y112_I),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(RIOB33_X105Y107_IOB_X1Y107_I),
.I4(1'b1),
.I5(RIOB33_X105Y113_IOB_X1Y113_I),
.O5(CLBLM_L_X8Y103_SLICE_X11Y103_DO5),
.O6(CLBLM_L_X8Y103_SLICE_X11Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h69a59955965a66aa)
  ) CLBLM_L_X8Y103_SLICE_X11Y103_CLUT (
.I0(CLBLM_L_X8Y102_SLICE_X11Y102_CO6),
.I1(LIOB33_X0Y105_IOB_X0Y105_I),
.I2(RIOB33_X105Y107_IOB_X1Y107_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(LIOB33_X0Y103_IOB_X0Y104_I),
.I5(CLBLM_L_X8Y100_SLICE_X10Y100_BO6),
.O5(CLBLM_L_X8Y103_SLICE_X11Y103_CO5),
.O6(CLBLM_L_X8Y103_SLICE_X11Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h2bbbafff8eee0aaa)
  ) CLBLM_L_X8Y103_SLICE_X11Y103_BLUT (
.I0(CLBLM_L_X8Y103_SLICE_X11Y103_DO6),
.I1(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I2(LIOB33_X0Y101_IOB_X0Y101_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(RIOB33_X105Y107_IOB_X1Y107_I),
.I5(CLBLM_L_X8Y103_SLICE_X11Y103_AO6),
.O5(CLBLM_L_X8Y103_SLICE_X11Y103_BO5),
.O6(CLBLM_L_X8Y103_SLICE_X11Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcf00f0005f5f5f5f)
  ) CLBLM_L_X8Y103_SLICE_X11Y103_ALUT (
.I0(LIOB33_X0Y103_IOB_X0Y104_I),
.I1(RIOB33_X105Y111_IOB_X1Y112_I),
.I2(RIOB33_X105Y107_IOB_X1Y108_I),
.I3(RIOB33_X105Y113_IOB_X1Y113_I),
.I4(RIOB33_X105Y107_IOB_X1Y107_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y103_SLICE_X11Y103_AO5),
.O6(CLBLM_L_X8Y103_SLICE_X11Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y104_SLICE_X10Y104_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y104_SLICE_X10Y104_DO5),
.O6(CLBLM_L_X8Y104_SLICE_X10Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y104_SLICE_X10Y104_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y104_SLICE_X10Y104_CO5),
.O6(CLBLM_L_X8Y104_SLICE_X10Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc96939996c3c9ccc)
  ) CLBLM_L_X8Y104_SLICE_X10Y104_BLUT (
.I0(CLBLM_L_X10Y104_SLICE_X12Y104_DO6),
.I1(CLBLM_L_X8Y103_SLICE_X10Y103_CO6),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(RIOB33_X105Y103_IOB_X1Y104_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_L_X8Y103_SLICE_X11Y103_CO6),
.O5(CLBLM_L_X8Y104_SLICE_X10Y104_BO5),
.O6(CLBLM_L_X8Y104_SLICE_X10Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0fffff5f5f5f5f)
  ) CLBLM_L_X8Y104_SLICE_X10Y104_ALUT (
.I0(LIOB33_X0Y107_IOB_X0Y108_I),
.I1(1'b1),
.I2(RIOB33_X105Y103_IOB_X1Y104_I),
.I3(1'b1),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y104_SLICE_X10Y104_AO5),
.O6(CLBLM_L_X8Y104_SLICE_X10Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y104_SLICE_X11Y104_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y104_SLICE_X11Y104_DO5),
.O6(CLBLM_L_X8Y104_SLICE_X11Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y104_SLICE_X11Y104_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y104_SLICE_X11Y104_CO5),
.O6(CLBLM_L_X8Y104_SLICE_X11Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h02bb3bbb23ffbfff)
  ) CLBLM_L_X8Y104_SLICE_X11Y104_BLUT (
.I0(CLBLM_L_X10Y105_SLICE_X13Y105_BO6),
.I1(CLBLM_L_X10Y103_SLICE_X12Y103_CO6),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(RIOB33_X105Y103_IOB_X1Y103_I),
.I4(LIOB33_X0Y107_IOB_X0Y107_I),
.I5(CLBLM_L_X10Y104_SLICE_X12Y104_CO6),
.O5(CLBLM_L_X8Y104_SLICE_X11Y104_BO5),
.O6(CLBLM_L_X8Y104_SLICE_X11Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8f707f80e51a15ea)
  ) CLBLM_L_X8Y104_SLICE_X11Y104_ALUT (
.I0(CLBLM_L_X10Y104_SLICE_X12Y104_CO6),
.I1(RIOB33_X105Y103_IOB_X1Y103_I),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(CLBLM_L_X10Y103_SLICE_X12Y103_DO6),
.I4(RIOB33_X105Y103_IOB_X1Y104_I),
.I5(CLBLM_L_X10Y105_SLICE_X13Y105_BO6),
.O5(CLBLM_L_X8Y104_SLICE_X11Y104_AO5),
.O6(CLBLM_L_X8Y104_SLICE_X11Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6999c33396663ccc)
  ) CLBLM_L_X8Y105_SLICE_X10Y105_DLUT (
.I0(RIOB33_X105Y103_IOB_X1Y103_I),
.I1(CLBLM_L_X10Y105_SLICE_X12Y105_CO6),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(RIOB33_X105Y101_IOB_X1Y102_I),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(CLBLM_L_X10Y107_SLICE_X13Y107_CO6),
.O5(CLBLM_L_X8Y105_SLICE_X10Y105_DO5),
.O6(CLBLM_L_X8Y105_SLICE_X10Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6699966996699966)
  ) CLBLM_L_X8Y105_SLICE_X10Y105_CLUT (
.I0(CLBLM_L_X10Y105_SLICE_X12Y105_BO6),
.I1(CLBLM_L_X10Y103_SLICE_X12Y103_CO6),
.I2(CLBLM_L_X10Y105_SLICE_X12Y105_AO6),
.I3(CLBLM_L_X8Y105_SLICE_X10Y105_AO5),
.I4(CLBLM_L_X10Y107_SLICE_X13Y107_CO6),
.I5(CLBLM_R_X7Y105_SLICE_X9Y105_AO6),
.O5(CLBLM_L_X8Y105_SLICE_X10Y105_CO5),
.O6(CLBLM_L_X8Y105_SLICE_X10Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6699966996699966)
  ) CLBLM_L_X8Y105_SLICE_X10Y105_BLUT (
.I0(CLBLM_R_X7Y105_SLICE_X9Y105_AO5),
.I1(CLBLM_L_X8Y103_SLICE_X10Y103_BO6),
.I2(CLBLM_L_X10Y103_SLICE_X12Y103_CO6),
.I3(CLBLM_L_X10Y103_SLICE_X12Y103_BO6),
.I4(CLBLM_L_X10Y105_SLICE_X12Y105_BO6),
.I5(CLBLM_L_X8Y105_SLICE_X10Y105_AO5),
.O5(CLBLM_L_X8Y105_SLICE_X10Y105_BO5),
.O6(CLBLM_L_X8Y105_SLICE_X10Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h55ff55ff33ff33ff)
  ) CLBLM_L_X8Y105_SLICE_X10Y105_ALUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(LIOB33_X0Y107_IOB_X0Y107_I),
.I2(1'b1),
.I3(RIOB33_X105Y103_IOB_X1Y103_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y105_SLICE_X10Y105_AO5),
.O6(CLBLM_L_X8Y105_SLICE_X10Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7b12bb22ff5affaa)
  ) CLBLM_L_X8Y105_SLICE_X11Y105_DLUT (
.I0(CLBLM_L_X8Y104_SLICE_X11Y104_AO6),
.I1(LIOB33_X0Y107_IOB_X0Y108_I),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(CLBLM_L_X8Y105_SLICE_X11Y105_CO6),
.I4(RIOB33_X105Y103_IOB_X1Y103_I),
.I5(RIOB33_X105Y101_IOB_X1Y102_I),
.O5(CLBLM_L_X8Y105_SLICE_X11Y105_DO5),
.O6(CLBLM_L_X8Y105_SLICE_X11Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fbfff3f152a3f00)
  ) CLBLM_L_X8Y105_SLICE_X11Y105_CLUT (
.I0(RIOB33_X105Y103_IOB_X1Y103_I),
.I1(RIOB33_X105Y101_IOB_X1Y102_I),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(CLBLM_L_X10Y105_SLICE_X12Y105_CO6),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(CLBLM_L_X10Y107_SLICE_X13Y107_CO6),
.O5(CLBLM_L_X8Y105_SLICE_X11Y105_CO5),
.O6(CLBLM_L_X8Y105_SLICE_X11Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hb24d4db2cf30cf30)
  ) CLBLM_L_X8Y105_SLICE_X11Y105_BLUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(CLBLM_L_X10Y105_SLICE_X13Y105_BO6),
.I2(CLBLM_L_X10Y104_SLICE_X12Y104_CO6),
.I3(CLBLM_L_X10Y103_SLICE_X12Y103_CO6),
.I4(LIOB33_X0Y107_IOB_X0Y107_I),
.I5(RIOB33_X105Y103_IOB_X1Y103_I),
.O5(CLBLM_L_X8Y105_SLICE_X11Y105_BO5),
.O6(CLBLM_L_X8Y105_SLICE_X11Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6ac0953f953f6ac0)
  ) CLBLM_L_X8Y105_SLICE_X11Y105_ALUT (
.I0(RIOB33_X105Y103_IOB_X1Y103_I),
.I1(RIOB33_X105Y101_IOB_X1Y102_I),
.I2(LIOB33_X0Y107_IOB_X0Y108_I),
.I3(LIOB33_X0Y107_IOB_X0Y107_I),
.I4(CLBLM_L_X8Y104_SLICE_X11Y104_AO6),
.I5(CLBLM_L_X8Y105_SLICE_X11Y105_CO6),
.O5(CLBLM_L_X8Y105_SLICE_X11Y105_AO5),
.O6(CLBLM_L_X8Y105_SLICE_X11Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf9909900ff99f990)
  ) CLBLM_L_X8Y106_SLICE_X10Y106_DLUT (
.I0(CLBLM_L_X8Y105_SLICE_X10Y105_CO6),
.I1(CLBLM_L_X8Y106_SLICE_X11Y106_AO5),
.I2(CLBLM_L_X8Y107_SLICE_X10Y107_DO6),
.I3(CLBLM_L_X8Y106_SLICE_X10Y106_AO5),
.I4(CLBLM_R_X7Y106_SLICE_X9Y106_AO5),
.I5(CLBLM_L_X8Y105_SLICE_X10Y105_DO6),
.O5(CLBLM_L_X8Y106_SLICE_X10Y106_DO5),
.O6(CLBLM_L_X8Y106_SLICE_X10Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha96a65a66966a5aa)
  ) CLBLM_L_X8Y106_SLICE_X10Y106_CLUT (
.I0(CLBLM_L_X8Y105_SLICE_X10Y105_CO6),
.I1(LIOB33_X0Y107_IOB_X0Y108_I),
.I2(CLBLM_L_X8Y107_SLICE_X10Y107_DO6),
.I3(CLBLM_L_X8Y105_SLICE_X10Y105_DO6),
.I4(RIOB33_X105Y101_IOB_X1Y102_I),
.I5(RIOB33_X105Y101_IOB_X1Y101_I),
.O5(CLBLM_L_X8Y106_SLICE_X10Y106_CO5),
.O6(CLBLM_L_X8Y106_SLICE_X10Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h781e87e187e1781e)
  ) CLBLM_L_X8Y106_SLICE_X10Y106_BLUT (
.I0(CLBLM_R_X7Y106_SLICE_X9Y106_AO5),
.I1(CLBLM_L_X8Y107_SLICE_X10Y107_DO6),
.I2(CLBLM_L_X8Y106_SLICE_X11Y106_AO5),
.I3(CLBLM_L_X8Y105_SLICE_X10Y105_DO6),
.I4(CLBLM_L_X8Y105_SLICE_X10Y105_CO6),
.I5(CLBLM_L_X8Y106_SLICE_X10Y106_AO5),
.O5(CLBLM_L_X8Y106_SLICE_X10Y106_BO5),
.O6(CLBLM_L_X8Y106_SLICE_X10Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h7777777733ff33ff)
  ) CLBLM_L_X8Y106_SLICE_X10Y106_ALUT (
.I0(RIOB33_X105Y101_IOB_X1Y102_I),
.I1(LIOB33_X0Y109_IOB_X0Y109_I),
.I2(1'b1),
.I3(RIOB33_X105Y101_IOB_X1Y101_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y106_SLICE_X10Y106_AO5),
.O6(CLBLM_L_X8Y106_SLICE_X10Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff9f99099f990900)
  ) CLBLM_L_X8Y106_SLICE_X11Y106_DLUT (
.I0(CLBLM_L_X8Y106_SLICE_X11Y106_AO6),
.I1(CLBLM_L_X8Y105_SLICE_X10Y105_BO6),
.I2(CLBLM_L_X8Y105_SLICE_X11Y105_BO6),
.I3(CLBLM_L_X8Y105_SLICE_X11Y105_CO6),
.I4(CLBLM_L_X8Y106_SLICE_X10Y106_AO6),
.I5(CLBLM_L_X8Y106_SLICE_X11Y106_AO5),
.O5(CLBLM_L_X8Y106_SLICE_X11Y106_DO5),
.O6(CLBLM_L_X8Y106_SLICE_X11Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hc69966c66c33cc6c)
  ) CLBLM_L_X8Y106_SLICE_X11Y106_CLUT (
.I0(LIOB33_X0Y107_IOB_X0Y108_I),
.I1(CLBLM_L_X8Y105_SLICE_X10Y105_BO6),
.I2(RIOB33_X105Y101_IOB_X1Y102_I),
.I3(CLBLM_L_X8Y105_SLICE_X11Y105_CO6),
.I4(CLBLM_L_X8Y105_SLICE_X11Y105_BO6),
.I5(RIOB33_X105Y103_IOB_X1Y103_I),
.O5(CLBLM_L_X8Y106_SLICE_X11Y106_CO5),
.O6(CLBLM_L_X8Y106_SLICE_X11Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h2dd2d22db44b4bb4)
  ) CLBLM_L_X8Y106_SLICE_X11Y106_BLUT (
.I0(CLBLM_L_X8Y105_SLICE_X11Y105_BO6),
.I1(CLBLM_L_X8Y106_SLICE_X11Y106_AO5),
.I2(CLBLM_L_X8Y106_SLICE_X10Y106_AO6),
.I3(CLBLM_L_X8Y105_SLICE_X10Y105_BO6),
.I4(CLBLM_L_X8Y106_SLICE_X11Y106_AO6),
.I5(CLBLM_L_X8Y105_SLICE_X11Y105_CO6),
.O5(CLBLM_L_X8Y106_SLICE_X11Y106_BO5),
.O6(CLBLM_L_X8Y106_SLICE_X11Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h777777775555ffff)
  ) CLBLM_L_X8Y106_SLICE_X11Y106_ALUT (
.I0(LIOB33_X0Y107_IOB_X0Y108_I),
.I1(RIOB33_X105Y103_IOB_X1Y103_I),
.I2(1'b1),
.I3(1'b1),
.I4(RIOB33_X105Y101_IOB_X1Y102_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y106_SLICE_X11Y106_AO5),
.O6(CLBLM_L_X8Y106_SLICE_X11Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fff8fff07770888)
  ) CLBLM_L_X8Y107_SLICE_X10Y107_DLUT (
.I0(RIOB33_X105Y101_IOB_X1Y102_I),
.I1(LIOB33_X0Y105_IOB_X0Y106_I),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(RIOB33_X105Y101_IOB_X1Y101_I),
.I4(CLBLM_L_X10Y107_SLICE_X13Y107_DO6),
.I5(CLBLM_L_X10Y108_SLICE_X12Y108_CO6),
.O5(CLBLM_L_X8Y107_SLICE_X10Y107_DO5),
.O6(CLBLM_L_X8Y107_SLICE_X10Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6c93936c93936c6c)
  ) CLBLM_L_X8Y107_SLICE_X10Y107_CLUT (
.I0(RIOB33_X105Y101_IOB_X1Y102_I),
.I1(CLBLM_L_X10Y106_SLICE_X12Y106_DO6),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(LIOB33_X0Y107_IOB_X0Y108_I),
.I4(CLBLM_L_X8Y107_SLICE_X10Y107_DO6),
.I5(RIOB33_X105Y101_IOB_X1Y101_I),
.O5(CLBLM_L_X8Y107_SLICE_X10Y107_CO5),
.O6(CLBLM_L_X8Y107_SLICE_X10Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h28be88eebebeeeee)
  ) CLBLM_L_X8Y107_SLICE_X10Y107_BLUT (
.I0(CLBLM_L_X8Y107_SLICE_X10Y107_DO6),
.I1(CLBLM_L_X10Y106_SLICE_X12Y106_DO6),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(RIOB33_X105Y101_IOB_X1Y101_I),
.I4(RIOB33_X105Y101_IOB_X1Y102_I),
.I5(LIOB33_X0Y107_IOB_X0Y108_I),
.O5(CLBLM_L_X8Y107_SLICE_X10Y107_BO5),
.O6(CLBLM_L_X8Y107_SLICE_X10Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6696996996996966)
  ) CLBLM_L_X8Y107_SLICE_X10Y107_ALUT (
.I0(CLBLM_R_X7Y105_SLICE_X9Y105_AO6),
.I1(CLBLM_L_X10Y107_SLICE_X13Y107_CO6),
.I2(CLBLM_L_X10Y107_SLICE_X13Y107_AO6),
.I3(CLBLM_L_X10Y108_SLICE_X12Y108_CO6),
.I4(CLBLM_L_X10Y105_SLICE_X12Y105_AO6),
.I5(CLBLM_L_X8Y108_SLICE_X10Y108_AO5),
.O5(CLBLM_L_X8Y107_SLICE_X10Y107_AO5),
.O6(CLBLM_L_X8Y107_SLICE_X10Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6a00ff6aff6aff6a)
  ) CLBLM_L_X8Y107_SLICE_X11Y107_DLUT (
.I0(CLBLM_L_X8Y108_SLICE_X11Y108_AO6),
.I1(RIOB33_X105Y101_IOB_X1Y101_I),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(CLBLM_L_X8Y107_SLICE_X11Y107_CO6),
.I4(LIOB33_X0Y107_IOB_X0Y108_I),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLM_L_X8Y107_SLICE_X11Y107_DO5),
.O6(CLBLM_L_X8Y107_SLICE_X11Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7d14f550ff3cfff0)
  ) CLBLM_L_X8Y107_SLICE_X11Y107_CLUT (
.I0(LIOB33_X0Y107_IOB_X0Y107_I),
.I1(RIOB33_X105Y101_IOB_X1Y101_I),
.I2(CLBLM_L_X10Y108_SLICE_X12Y108_DO6),
.I3(CLBLM_R_X7Y110_SLICE_X9Y110_CO6),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLM_L_X8Y107_SLICE_X11Y107_CO5),
.O6(CLBLM_L_X8Y107_SLICE_X11Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h69c3a50f963c5af0)
  ) CLBLM_L_X8Y107_SLICE_X11Y107_BLUT (
.I0(LIOB33_X0Y107_IOB_X0Y108_I),
.I1(RIOB33_X105Y101_IOB_X1Y101_I),
.I2(CLBLM_L_X8Y108_SLICE_X11Y108_AO6),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(LIOB33_X0Y107_IOB_X0Y107_I),
.I5(CLBLM_L_X8Y107_SLICE_X11Y107_CO6),
.O5(CLBLM_L_X8Y107_SLICE_X11Y107_BO5),
.O6(CLBLM_L_X8Y107_SLICE_X11Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h69c3a50f963c5af0)
  ) CLBLM_L_X8Y107_SLICE_X11Y107_ALUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(CLBLM_L_X10Y108_SLICE_X12Y108_DO6),
.I3(RIOB33_X105Y101_IOB_X1Y101_I),
.I4(LIOB33_X0Y107_IOB_X0Y107_I),
.I5(CLBLM_R_X7Y110_SLICE_X9Y110_CO6),
.O5(CLBLM_L_X8Y107_SLICE_X11Y107_AO5),
.O6(CLBLM_L_X8Y107_SLICE_X11Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y108_SLICE_X10Y108_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y108_SLICE_X10Y108_DO5),
.O6(CLBLM_L_X8Y108_SLICE_X10Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h69a59955965a66aa)
  ) CLBLM_L_X8Y108_SLICE_X10Y108_CLUT (
.I0(CLBLM_L_X10Y107_SLICE_X13Y107_DO6),
.I1(RIOB33_X105Y101_IOB_X1Y102_I),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(LIOB33_X0Y105_IOB_X0Y106_I),
.I4(RIOB33_X105Y101_IOB_X1Y101_I),
.I5(CLBLM_L_X10Y108_SLICE_X12Y108_CO6),
.O5(CLBLM_L_X8Y108_SLICE_X10Y108_CO5),
.O6(CLBLM_L_X8Y108_SLICE_X10Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h693cc36996c33c96)
  ) CLBLM_L_X8Y108_SLICE_X10Y108_BLUT (
.I0(CLBLM_R_X7Y110_SLICE_X9Y110_CO6),
.I1(CLBLM_L_X10Y107_SLICE_X13Y107_AO6),
.I2(CLBLM_L_X10Y108_SLICE_X12Y108_CO6),
.I3(CLBLM_L_X10Y108_SLICE_X12Y108_BO6),
.I4(CLBLM_L_X8Y108_SLICE_X10Y108_AO6),
.I5(CLBLM_L_X8Y108_SLICE_X10Y108_AO5),
.O5(CLBLM_L_X8Y108_SLICE_X10Y108_BO5),
.O6(CLBLM_L_X8Y108_SLICE_X10Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h55ff55ff5f5f5f5f)
  ) CLBLM_L_X8Y108_SLICE_X10Y108_ALUT (
.I0(LIOB33_X0Y107_IOB_X0Y107_I),
.I1(1'b1),
.I2(RIOB33_X105Y101_IOB_X1Y101_I),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y108_SLICE_X10Y108_AO5),
.O6(CLBLM_L_X8Y108_SLICE_X10Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6999a55596665aaa)
  ) CLBLM_L_X8Y108_SLICE_X11Y108_DLUT (
.I0(CLBLM_L_X8Y109_SLICE_X11Y109_AO6),
.I1(LIOB33_X0Y103_IOB_X0Y104_I),
.I2(LIOB33_X0Y105_IOB_X0Y105_I),
.I3(RIOB33_X105Y101_IOB_X1Y101_I),
.I4(RIOB33_X105Y101_IOB_X1Y102_I),
.I5(CLBLM_L_X8Y110_SLICE_X10Y110_BO6),
.O5(CLBLM_L_X8Y108_SLICE_X11Y108_DO5),
.O6(CLBLM_L_X8Y108_SLICE_X11Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fdfdfdf134c4c4c)
  ) CLBLM_L_X8Y108_SLICE_X11Y108_CLUT (
.I0(RIOB33_X105Y101_IOB_X1Y101_I),
.I1(CLBLM_L_X8Y109_SLICE_X11Y109_AO6),
.I2(LIOB33_X0Y105_IOB_X0Y105_I),
.I3(LIOB33_X0Y103_IOB_X0Y104_I),
.I4(RIOB33_X105Y101_IOB_X1Y102_I),
.I5(CLBLM_L_X8Y110_SLICE_X10Y110_BO6),
.O5(CLBLM_L_X8Y108_SLICE_X11Y108_CO5),
.O6(CLBLM_L_X8Y108_SLICE_X11Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hb73f48c0d1952e6a)
  ) CLBLM_L_X8Y108_SLICE_X11Y108_BLUT (
.I0(CLBLM_L_X8Y108_SLICE_X11Y108_DO6),
.I1(LIOB33_X0Y105_IOB_X0Y106_I),
.I2(RIOB33_X105Y101_IOB_X1Y101_I),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(CLBLM_L_X10Y108_SLICE_X12Y108_DO6),
.I5(CLBLM_L_X8Y111_SLICE_X10Y111_BO6),
.O5(CLBLM_L_X8Y108_SLICE_X11Y108_BO5),
.O6(CLBLM_L_X8Y108_SLICE_X11Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hb43c78f0d2961e5a)
  ) CLBLM_L_X8Y108_SLICE_X11Y108_ALUT (
.I0(CLBLM_L_X10Y106_SLICE_X12Y106_CO6),
.I1(LIOB33_X0Y105_IOB_X0Y106_I),
.I2(CLBLM_L_X10Y107_SLICE_X13Y107_DO6),
.I3(RIOB33_X105Y101_IOB_X1Y101_I),
.I4(RIOB33_X105Y101_IOB_X1Y102_I),
.I5(CLBLM_L_X8Y108_SLICE_X11Y108_CO6),
.O5(CLBLM_L_X8Y108_SLICE_X11Y108_AO5),
.O6(CLBLM_L_X8Y108_SLICE_X11Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y109_SLICE_X10Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y109_SLICE_X10Y109_DO5),
.O6(CLBLM_L_X8Y109_SLICE_X10Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h07050a0088aa0a00)
  ) CLBLM_L_X8Y109_SLICE_X10Y109_CLUT (
.I0(RIOB33_X105Y113_IOB_X1Y113_I),
.I1(RIOB33_X105Y111_IOB_X1Y112_I),
.I2(RIOB33_X105Y101_IOB_X1Y102_I),
.I3(RIOB33_X105Y103_IOB_X1Y104_I),
.I4(RIOB33_X105Y103_IOB_X1Y103_I),
.I5(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.O5(CLBLM_L_X8Y109_SLICE_X10Y109_CO5),
.O6(CLBLM_L_X8Y109_SLICE_X10Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h03737c0c80f0b0c0)
  ) CLBLM_L_X8Y109_SLICE_X10Y109_BLUT (
.I0(RIOB33_X105Y111_IOB_X1Y112_I),
.I1(RIOB33_X105Y103_IOB_X1Y103_I),
.I2(RIOB33_X105Y113_IOB_X1Y113_I),
.I3(RIOB33_X105Y103_IOB_X1Y104_I),
.I4(RIOB33_X105Y101_IOB_X1Y102_I),
.I5(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.O5(CLBLM_L_X8Y109_SLICE_X10Y109_BO5),
.O6(CLBLM_L_X8Y109_SLICE_X10Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff005fa05fa05f)
  ) CLBLM_L_X8Y109_SLICE_X10Y109_ALUT (
.I0(LIOB33_X0Y101_IOB_X0Y101_I),
.I1(1'b1),
.I2(RIOB33_X105Y101_IOB_X1Y102_I),
.I3(CLBLM_L_X8Y109_SLICE_X10Y109_BO6),
.I4(CLBLM_L_X8Y109_SLICE_X10Y109_CO6),
.I5(1'b1),
.O5(CLBLM_L_X8Y109_SLICE_X10Y109_AO5),
.O6(CLBLM_L_X8Y109_SLICE_X10Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y109_SLICE_X11Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y109_SLICE_X11Y109_DO5),
.O6(CLBLM_L_X8Y109_SLICE_X11Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y109_SLICE_X11Y109_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y109_SLICE_X11Y109_CO5),
.O6(CLBLM_L_X8Y109_SLICE_X11Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y109_SLICE_X11Y109_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y109_SLICE_X11Y109_BO5),
.O6(CLBLM_L_X8Y109_SLICE_X11Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h99696966a5aaa5aa)
  ) CLBLM_L_X8Y109_SLICE_X11Y109_ALUT (
.I0(CLBLM_L_X10Y109_SLICE_X12Y109_CO6),
.I1(RIOB33_X105Y103_IOB_X1Y103_I),
.I2(CLBLM_L_X8Y109_SLICE_X10Y109_AO6),
.I3(CLBLM_L_X10Y109_SLICE_X12Y109_AO6),
.I4(RIOB33_X105Y101_IOB_X1Y102_I),
.I5(LIOB33_X0Y101_IOB_X0Y102_I),
.O5(CLBLM_L_X8Y109_SLICE_X11Y109_AO5),
.O6(CLBLM_L_X8Y109_SLICE_X11Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y110_SLICE_X10Y110_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y110_SLICE_X10Y110_DO5),
.O6(CLBLM_L_X8Y110_SLICE_X10Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3cc3f00f3c96f0f0)
  ) CLBLM_L_X8Y110_SLICE_X10Y110_CLUT (
.I0(RIOB33_X105Y101_IOB_X1Y102_I),
.I1(RIOB33_X105Y103_IOB_X1Y103_I),
.I2(CLBLM_L_X10Y109_SLICE_X12Y109_DO6),
.I3(CLBLM_L_X8Y109_SLICE_X10Y109_CO6),
.I4(LIOB33_X0Y101_IOB_X0Y101_I),
.I5(CLBLM_L_X8Y109_SLICE_X10Y109_BO6),
.O5(CLBLM_L_X8Y110_SLICE_X10Y110_CO5),
.O6(CLBLM_L_X8Y110_SLICE_X10Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h4dcfddffd4fc44cc)
  ) CLBLM_L_X8Y110_SLICE_X10Y110_BLUT (
.I0(RIOB33_X105Y101_IOB_X1Y101_I),
.I1(CLBLM_L_X8Y112_SLICE_X11Y112_CO6),
.I2(RIOB33_X105Y101_IOB_X1Y102_I),
.I3(LIOB33_X0Y103_IOB_X0Y104_I),
.I4(LIOB33_X0Y101_IOB_X0Y102_I),
.I5(CLBLM_L_X8Y110_SLICE_X10Y110_CO6),
.O5(CLBLM_L_X8Y110_SLICE_X10Y110_BO5),
.O6(CLBLM_L_X8Y110_SLICE_X10Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h69c39933963c66cc)
  ) CLBLM_L_X8Y110_SLICE_X10Y110_ALUT (
.I0(RIOB33_X105Y101_IOB_X1Y101_I),
.I1(CLBLM_L_X8Y112_SLICE_X11Y112_CO6),
.I2(RIOB33_X105Y101_IOB_X1Y102_I),
.I3(LIOB33_X0Y103_IOB_X0Y104_I),
.I4(LIOB33_X0Y101_IOB_X0Y102_I),
.I5(CLBLM_L_X8Y110_SLICE_X10Y110_CO6),
.O5(CLBLM_L_X8Y110_SLICE_X10Y110_AO5),
.O6(CLBLM_L_X8Y110_SLICE_X10Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'he8e88e8efae8af8e)
  ) CLBLM_L_X8Y110_SLICE_X11Y110_DLUT (
.I0(CLBLM_L_X8Y110_SLICE_X11Y110_AO6),
.I1(CLBLM_L_X8Y109_SLICE_X10Y109_CO6),
.I2(CLBLM_L_X10Y109_SLICE_X12Y109_DO6),
.I3(CLBLM_L_X8Y110_SLICE_X11Y110_AO5),
.I4(CLBLM_L_X10Y108_SLICE_X13Y108_AO6),
.I5(CLBLM_L_X8Y109_SLICE_X10Y109_BO6),
.O5(CLBLM_L_X8Y110_SLICE_X11Y110_DO5),
.O6(CLBLM_L_X8Y110_SLICE_X11Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6999966666699996)
  ) CLBLM_L_X8Y110_SLICE_X11Y110_CLUT (
.I0(CLBLM_L_X10Y108_SLICE_X13Y108_BO6),
.I1(CLBLM_L_X10Y107_SLICE_X12Y107_AO6),
.I2(CLBLM_R_X7Y112_SLICE_X9Y112_AO5),
.I3(CLBLM_L_X8Y112_SLICE_X11Y112_CO6),
.I4(CLBLM_L_X8Y110_SLICE_X11Y110_DO6),
.I5(CLBLM_L_X8Y110_SLICE_X11Y110_BO6),
.O5(CLBLM_L_X8Y110_SLICE_X11Y110_CO5),
.O6(CLBLM_L_X8Y110_SLICE_X11Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5a96a5695aa5a55a)
  ) CLBLM_L_X8Y110_SLICE_X11Y110_BLUT (
.I0(CLBLM_L_X10Y109_SLICE_X12Y109_DO6),
.I1(CLBLM_L_X8Y109_SLICE_X10Y109_BO6),
.I2(CLBLM_L_X10Y108_SLICE_X13Y108_AO6),
.I3(CLBLM_L_X8Y109_SLICE_X10Y109_CO6),
.I4(CLBLM_L_X8Y110_SLICE_X11Y110_AO6),
.I5(CLBLM_L_X8Y110_SLICE_X11Y110_AO5),
.O5(CLBLM_L_X8Y110_SLICE_X11Y110_BO5),
.O6(CLBLM_L_X8Y110_SLICE_X11Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0fffff5555ffff)
  ) CLBLM_L_X8Y110_SLICE_X11Y110_ALUT (
.I0(LIOB33_X0Y101_IOB_X0Y101_I),
.I1(1'b1),
.I2(LIOB33_X0Y101_IOB_X0Y102_I),
.I3(1'b1),
.I4(RIOB33_X105Y101_IOB_X1Y102_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y110_SLICE_X11Y110_AO5),
.O6(CLBLM_L_X8Y110_SLICE_X11Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y111_SLICE_X10Y111_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y111_SLICE_X10Y111_DO5),
.O6(CLBLM_L_X8Y111_SLICE_X10Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h446c00006c6c446c)
  ) CLBLM_L_X8Y111_SLICE_X10Y111_CLUT (
.I0(LIOB33_X0Y101_IOB_X0Y102_I),
.I1(CLBLM_L_X8Y110_SLICE_X10Y110_CO6),
.I2(RIOB33_X105Y101_IOB_X1Y102_I),
.I3(RIOB33_X105Y101_IOB_X1Y101_I),
.I4(CLBLM_L_X8Y112_SLICE_X10Y112_AO5),
.I5(CLBLM_L_X8Y109_SLICE_X10Y109_AO5),
.O5(CLBLM_L_X8Y111_SLICE_X10Y111_CO5),
.O6(CLBLM_L_X8Y111_SLICE_X10Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h2abf80eabfbfeaea)
  ) CLBLM_L_X8Y111_SLICE_X10Y111_BLUT (
.I0(CLBLM_L_X8Y112_SLICE_X10Y112_DO6),
.I1(LIOB33_X0Y103_IOB_X0Y104_I),
.I2(RIOB33_X105Y101_IOB_X1Y101_I),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(CLBLM_L_X8Y111_SLICE_X10Y111_AO6),
.I5(LIOB33_X0Y105_IOB_X0Y105_I),
.O5(CLBLM_L_X8Y111_SLICE_X10Y111_BO5),
.O6(CLBLM_L_X8Y111_SLICE_X10Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc96939996c3c9ccc)
  ) CLBLM_L_X8Y111_SLICE_X10Y111_ALUT (
.I0(CLBLM_L_X8Y112_SLICE_X10Y112_AO5),
.I1(CLBLM_L_X8Y110_SLICE_X10Y110_CO6),
.I2(LIOB33_X0Y101_IOB_X0Y102_I),
.I3(RIOB33_X105Y101_IOB_X1Y101_I),
.I4(RIOB33_X105Y101_IOB_X1Y102_I),
.I5(CLBLM_L_X8Y109_SLICE_X10Y109_AO5),
.O5(CLBLM_L_X8Y111_SLICE_X10Y111_AO5),
.O6(CLBLM_L_X8Y111_SLICE_X10Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y111_SLICE_X11Y111_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y111_SLICE_X11Y111_DO5),
.O6(CLBLM_L_X8Y111_SLICE_X11Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y111_SLICE_X11Y111_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y111_SLICE_X11Y111_CO5),
.O6(CLBLM_L_X8Y111_SLICE_X11Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y111_SLICE_X11Y111_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y111_SLICE_X11Y111_BO5),
.O6(CLBLM_L_X8Y111_SLICE_X11Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y111_SLICE_X11Y111_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y111_SLICE_X11Y111_AO5),
.O6(CLBLM_L_X8Y111_SLICE_X11Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fff07778fff0888)
  ) CLBLM_L_X8Y112_SLICE_X10Y112_DLUT (
.I0(LIOB33_X0Y101_IOB_X0Y102_I),
.I1(RIOB33_X105Y101_IOB_X1Y101_I),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(LIOB33_X0Y103_IOB_X0Y104_I),
.I4(CLBLM_R_X7Y113_SLICE_X9Y113_DO6),
.I5(CLBLM_L_X8Y112_SLICE_X10Y112_BO6),
.O5(CLBLM_L_X8Y112_SLICE_X10Y112_DO5),
.O6(CLBLM_L_X8Y112_SLICE_X10Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h63c69c399c3963c6)
  ) CLBLM_L_X8Y112_SLICE_X10Y112_CLUT (
.I0(CLBLM_R_X7Y113_SLICE_X9Y113_DO6),
.I1(CLBLM_L_X8Y112_SLICE_X11Y112_CO6),
.I2(CLBLM_L_X8Y112_SLICE_X11Y112_DO6),
.I3(CLBLM_R_X7Y113_SLICE_X9Y113_AO5),
.I4(CLBLM_R_X7Y112_SLICE_X9Y112_AO5),
.I5(CLBLM_L_X8Y110_SLICE_X11Y110_BO6),
.O5(CLBLM_L_X8Y112_SLICE_X10Y112_CO5),
.O6(CLBLM_L_X8Y112_SLICE_X10Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h67cd983265cf9a30)
  ) CLBLM_L_X8Y112_SLICE_X10Y112_BLUT (
.I0(LIOB33_X0Y101_IOB_X0Y101_I),
.I1(CLBLM_L_X8Y112_SLICE_X11Y112_BO6),
.I2(CLBLM_L_X8Y112_SLICE_X11Y112_AO6),
.I3(RIOB33_X105Y101_IOB_X1Y102_I),
.I4(CLBLM_L_X8Y109_SLICE_X10Y109_BO6),
.I5(RIOB33_X105Y101_IOB_X1Y101_I),
.O5(CLBLM_L_X8Y112_SLICE_X10Y112_BO5),
.O6(CLBLM_L_X8Y112_SLICE_X10Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha50fa50fcdcfcdcf)
  ) CLBLM_L_X8Y112_SLICE_X10Y112_ALUT (
.I0(LIOB33_X0Y101_IOB_X0Y101_I),
.I1(CLBLM_L_X8Y112_SLICE_X11Y112_BO6),
.I2(CLBLM_L_X8Y112_SLICE_X11Y112_AO6),
.I3(RIOB33_X105Y101_IOB_X1Y101_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y112_SLICE_X10Y112_AO5),
.O6(CLBLM_L_X8Y112_SLICE_X10Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3c3cc3c3c3693c96)
  ) CLBLM_L_X8Y112_SLICE_X11Y112_DLUT (
.I0(CLBLM_L_X8Y113_SLICE_X11Y113_AO6),
.I1(CLBLM_L_X8Y110_SLICE_X11Y110_AO5),
.I2(CLBLM_L_X8Y113_SLICE_X11Y113_AO5),
.I3(CLBLM_L_X8Y112_SLICE_X11Y112_AO6),
.I4(CLBLM_L_X8Y109_SLICE_X10Y109_BO6),
.I5(CLBLM_L_X8Y112_SLICE_X11Y112_BO6),
.O5(CLBLM_L_X8Y112_SLICE_X11Y112_DO5),
.O6(CLBLM_L_X8Y112_SLICE_X11Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcf3fcf3c030e8b2)
  ) CLBLM_L_X8Y112_SLICE_X11Y112_CLUT (
.I0(CLBLM_L_X8Y113_SLICE_X11Y113_AO6),
.I1(CLBLM_L_X8Y109_SLICE_X10Y109_BO6),
.I2(CLBLM_L_X8Y113_SLICE_X11Y113_AO5),
.I3(CLBLM_L_X8Y110_SLICE_X11Y110_AO5),
.I4(CLBLM_L_X8Y112_SLICE_X11Y112_AO6),
.I5(CLBLM_L_X8Y112_SLICE_X11Y112_BO6),
.O5(CLBLM_L_X8Y112_SLICE_X11Y112_CO5),
.O6(CLBLM_L_X8Y112_SLICE_X11Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h002cc0e000ac4060)
  ) CLBLM_L_X8Y112_SLICE_X11Y112_BLUT (
.I0(RIOB33_X105Y103_IOB_X1Y103_I),
.I1(RIOB33_X105Y101_IOB_X1Y102_I),
.I2(RIOB33_X105Y113_IOB_X1Y113_I),
.I3(RIOB33_X105Y101_IOB_X1Y101_I),
.I4(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I5(RIOB33_X105Y111_IOB_X1Y112_I),
.O5(CLBLM_L_X8Y112_SLICE_X11Y112_BO5),
.O6(CLBLM_L_X8Y112_SLICE_X11Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h132cd0e053ac5060)
  ) CLBLM_L_X8Y112_SLICE_X11Y112_ALUT (
.I0(RIOB33_X105Y103_IOB_X1Y103_I),
.I1(RIOB33_X105Y101_IOB_X1Y102_I),
.I2(RIOB33_X105Y113_IOB_X1Y113_I),
.I3(RIOB33_X105Y101_IOB_X1Y101_I),
.I4(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I5(RIOB33_X105Y111_IOB_X1Y112_I),
.O5(CLBLM_L_X8Y112_SLICE_X11Y112_AO5),
.O6(CLBLM_L_X8Y112_SLICE_X11Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y113_SLICE_X10Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y113_SLICE_X10Y113_DO5),
.O6(CLBLM_L_X8Y113_SLICE_X10Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y113_SLICE_X10Y113_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y113_SLICE_X10Y113_CO5),
.O6(CLBLM_L_X8Y113_SLICE_X10Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y113_SLICE_X10Y113_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y113_SLICE_X10Y113_BO5),
.O6(CLBLM_L_X8Y113_SLICE_X10Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y113_SLICE_X10Y113_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y113_SLICE_X10Y113_AO5),
.O6(CLBLM_L_X8Y113_SLICE_X10Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y113_SLICE_X11Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y113_SLICE_X11Y113_DO5),
.O6(CLBLM_L_X8Y113_SLICE_X11Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y113_SLICE_X11Y113_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y113_SLICE_X11Y113_CO5),
.O6(CLBLM_L_X8Y113_SLICE_X11Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y113_SLICE_X11Y113_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y113_SLICE_X11Y113_BO5),
.O6(CLBLM_L_X8Y113_SLICE_X11Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h55ff55ff0fff0fff)
  ) CLBLM_L_X8Y113_SLICE_X11Y113_ALUT (
.I0(LIOB33_X0Y101_IOB_X0Y101_I),
.I1(1'b1),
.I2(LIOB33_X0Y101_IOB_X0Y102_I),
.I3(RIOB33_X105Y101_IOB_X1Y101_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y113_SLICE_X11Y113_AO5),
.O6(CLBLM_L_X8Y113_SLICE_X11Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbfaa2a0a2a0fbfa)
  ) CLBLM_L_X10Y102_SLICE_X12Y102_DLUT (
.I0(CLBLM_L_X10Y102_SLICE_X12Y102_AO6),
.I1(CLBLM_L_X10Y102_SLICE_X13Y102_AO6),
.I2(CLBLM_L_X8Y101_SLICE_X10Y101_AO6),
.I3(CLBLM_R_X5Y102_SLICE_X6Y102_BO6),
.I4(CLBLM_L_X8Y102_SLICE_X10Y102_DO6),
.I5(CLBLL_L_X4Y101_SLICE_X5Y101_AO6),
.O5(CLBLM_L_X10Y102_SLICE_X12Y102_DO5),
.O6(CLBLM_L_X10Y102_SLICE_X12Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h788787781ee1e11e)
  ) CLBLM_L_X10Y102_SLICE_X12Y102_CLUT (
.I0(CLBLM_L_X10Y103_SLICE_X13Y103_CO6),
.I1(CLBLM_L_X10Y103_SLICE_X12Y103_AO5),
.I2(CLBLM_L_X8Y100_SLICE_X10Y100_DO6),
.I3(CLBLM_L_X10Y102_SLICE_X12Y102_AO5),
.I4(CLBLM_L_X10Y102_SLICE_X12Y102_DO6),
.I5(CLBLM_L_X10Y102_SLICE_X12Y102_BO6),
.O5(CLBLM_L_X10Y102_SLICE_X12Y102_CO5),
.O6(CLBLM_L_X10Y102_SLICE_X12Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h65669a999a996566)
  ) CLBLM_L_X10Y102_SLICE_X12Y102_BLUT (
.I0(CLBLM_L_X8Y102_SLICE_X10Y102_DO6),
.I1(CLBLM_L_X8Y101_SLICE_X10Y101_AO6),
.I2(CLBLM_L_X10Y102_SLICE_X13Y102_AO6),
.I3(CLBLM_R_X5Y102_SLICE_X6Y102_BO6),
.I4(CLBLM_L_X10Y102_SLICE_X12Y102_AO6),
.I5(CLBLL_L_X4Y101_SLICE_X5Y101_AO6),
.O5(CLBLM_L_X10Y102_SLICE_X12Y102_BO5),
.O6(CLBLM_L_X10Y102_SLICE_X12Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0fff0fff55ff55ff)
  ) CLBLM_L_X10Y102_SLICE_X12Y102_ALUT (
.I0(LIOB33_X0Y103_IOB_X0Y104_I),
.I1(1'b1),
.I2(LIOB33_X0Y101_IOB_X0Y102_I),
.I3(RIOB33_X105Y107_IOB_X1Y107_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y102_SLICE_X12Y102_AO5),
.O6(CLBLM_L_X10Y102_SLICE_X12Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y102_SLICE_X13Y102_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y102_SLICE_X13Y102_DO5),
.O6(CLBLM_L_X10Y102_SLICE_X13Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y102_SLICE_X13Y102_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y102_SLICE_X13Y102_CO5),
.O6(CLBLM_L_X10Y102_SLICE_X13Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y102_SLICE_X13Y102_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y102_SLICE_X13Y102_BO5),
.O6(CLBLM_L_X10Y102_SLICE_X13Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h55223c882d223c88)
  ) CLBLM_L_X10Y102_SLICE_X13Y102_ALUT (
.I0(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I1(RIOB33_X105Y107_IOB_X1Y107_I),
.I2(RIOB33_X105Y109_IOB_X1Y109_I),
.I3(RIOB33_X105Y113_IOB_X1Y113_I),
.I4(RIOB33_X105Y107_IOB_X1Y108_I),
.I5(RIOB33_X105Y111_IOB_X1Y112_I),
.O5(CLBLM_L_X10Y102_SLICE_X13Y102_AO5),
.O6(CLBLM_L_X10Y102_SLICE_X13Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h9f60c53a3fc0956a)
  ) CLBLM_L_X10Y103_SLICE_X12Y103_DLUT (
.I0(CLBLM_L_X8Y102_SLICE_X11Y102_AO6),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(LIOB33_X0Y105_IOB_X0Y105_I),
.I3(CLBLM_L_X10Y102_SLICE_X12Y102_CO6),
.I4(CLBLM_L_X10Y104_SLICE_X13Y104_CO6),
.I5(RIOB33_X105Y103_IOB_X1Y104_I),
.O5(CLBLM_L_X10Y103_SLICE_X12Y103_DO5),
.O6(CLBLM_L_X10Y103_SLICE_X12Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3c9696c3c369693c)
  ) CLBLM_L_X10Y103_SLICE_X12Y103_CLUT (
.I0(CLBLM_L_X8Y102_SLICE_X11Y102_AO6),
.I1(CLBLM_L_X10Y102_SLICE_X12Y102_CO6),
.I2(CLBLM_L_X8Y103_SLICE_X10Y103_AO5),
.I3(CLBLM_L_X10Y104_SLICE_X12Y104_AO5),
.I4(CLBLM_L_X10Y104_SLICE_X13Y104_CO6),
.I5(CLBLM_L_X8Y104_SLICE_X10Y104_AO6),
.O5(CLBLM_L_X10Y103_SLICE_X12Y103_CO5),
.O6(CLBLM_L_X10Y103_SLICE_X12Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'heb82ffc3c300eb82)
  ) CLBLM_L_X10Y103_SLICE_X12Y103_BLUT (
.I0(CLBLM_L_X10Y104_SLICE_X13Y104_CO6),
.I1(CLBLM_L_X8Y103_SLICE_X10Y103_AO5),
.I2(CLBLM_L_X10Y102_SLICE_X12Y102_CO6),
.I3(CLBLM_L_X8Y104_SLICE_X10Y104_AO6),
.I4(CLBLM_L_X8Y102_SLICE_X11Y102_AO6),
.I5(CLBLM_L_X10Y104_SLICE_X12Y104_AO5),
.O5(CLBLM_L_X10Y103_SLICE_X12Y103_BO5),
.O6(CLBLM_L_X10Y103_SLICE_X12Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h55ff55ff77777777)
  ) CLBLM_L_X10Y103_SLICE_X12Y103_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(LIOB33_X0Y103_IOB_X0Y104_I),
.I2(1'b1),
.I3(LIOB33_X0Y101_IOB_X0Y102_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y103_SLICE_X12Y103_AO5),
.O6(CLBLM_L_X10Y103_SLICE_X12Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3ccc3cccc3669666)
  ) CLBLM_L_X10Y103_SLICE_X13Y103_DLUT (
.I0(CLBLM_L_X10Y104_SLICE_X13Y104_AO6),
.I1(CLBLM_L_X10Y102_SLICE_X13Y102_AO6),
.I2(RIOB33_X105Y107_IOB_X1Y107_I),
.I3(LIOB33_X0Y101_IOB_X0Y101_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_L_X10Y103_SLICE_X13Y103_BO6),
.O5(CLBLM_L_X10Y103_SLICE_X13Y103_DO5),
.O6(CLBLM_L_X10Y103_SLICE_X13Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff999999f90090)
  ) CLBLM_L_X10Y103_SLICE_X13Y103_CLUT (
.I0(CLBLM_R_X5Y102_SLICE_X6Y102_BO6),
.I1(CLBLM_L_X10Y102_SLICE_X13Y102_AO6),
.I2(CLBLM_R_X5Y102_SLICE_X6Y102_AO6),
.I3(CLBLM_L_X10Y104_SLICE_X13Y104_AO6),
.I4(CLBLM_L_X10Y103_SLICE_X12Y103_AO6),
.I5(CLBLM_L_X10Y103_SLICE_X13Y103_BO6),
.O5(CLBLM_L_X10Y103_SLICE_X13Y103_CO5),
.O6(CLBLM_L_X10Y103_SLICE_X13Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h1d0c4040510c4040)
  ) CLBLM_L_X10Y103_SLICE_X13Y103_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(RIOB33_X105Y107_IOB_X1Y107_I),
.I2(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I3(RIOB33_X105Y107_IOB_X1Y108_I),
.I4(RIOB33_X105Y113_IOB_X1Y113_I),
.I5(RIOB33_X105Y111_IOB_X1Y112_I),
.O5(CLBLM_L_X10Y103_SLICE_X13Y103_BO5),
.O6(CLBLM_L_X10Y103_SLICE_X13Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h639c66999c639966)
  ) CLBLM_L_X10Y103_SLICE_X13Y103_ALUT (
.I0(CLBLM_L_X10Y103_SLICE_X13Y103_BO6),
.I1(CLBLM_L_X10Y102_SLICE_X13Y102_AO6),
.I2(CLBLM_L_X10Y104_SLICE_X13Y104_AO6),
.I3(CLBLM_R_X5Y102_SLICE_X6Y102_BO6),
.I4(CLBLM_R_X5Y102_SLICE_X6Y102_AO6),
.I5(CLBLM_L_X10Y103_SLICE_X12Y103_AO6),
.O5(CLBLM_L_X10Y103_SLICE_X13Y103_AO5),
.O6(CLBLM_L_X10Y103_SLICE_X13Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h4dcfddffd4fc44cc)
  ) CLBLM_L_X10Y104_SLICE_X12Y104_DLUT (
.I0(RIOB33_X105Y103_IOB_X1Y104_I),
.I1(CLBLM_L_X10Y104_SLICE_X13Y104_CO6),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(LIOB33_X0Y105_IOB_X0Y105_I),
.I4(LIOB33_X0Y103_IOB_X0Y104_I),
.I5(CLBLM_L_X8Y102_SLICE_X11Y102_BO6),
.O5(CLBLM_L_X10Y104_SLICE_X12Y104_DO5),
.O6(CLBLM_L_X10Y104_SLICE_X12Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h69c39933963c66cc)
  ) CLBLM_L_X10Y104_SLICE_X12Y104_CLUT (
.I0(RIOB33_X105Y103_IOB_X1Y104_I),
.I1(CLBLM_L_X10Y104_SLICE_X13Y104_CO6),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(LIOB33_X0Y105_IOB_X0Y105_I),
.I4(LIOB33_X0Y103_IOB_X0Y104_I),
.I5(CLBLM_L_X8Y102_SLICE_X11Y102_BO6),
.O5(CLBLM_L_X10Y104_SLICE_X12Y104_CO5),
.O6(CLBLM_L_X10Y104_SLICE_X12Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3c9696c3c369693c)
  ) CLBLM_L_X10Y104_SLICE_X12Y104_BLUT (
.I0(CLBLM_L_X10Y103_SLICE_X13Y103_AO6),
.I1(CLBLM_L_X10Y102_SLICE_X12Y102_BO6),
.I2(CLBLM_L_X10Y103_SLICE_X13Y103_CO6),
.I3(CLBLM_R_X11Y106_SLICE_X14Y106_CO6),
.I4(CLBLM_L_X10Y104_SLICE_X12Y104_AO6),
.I5(CLBLM_L_X10Y103_SLICE_X12Y103_AO5),
.O5(CLBLM_L_X10Y104_SLICE_X12Y104_BO5),
.O6(CLBLM_L_X10Y104_SLICE_X12Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5f5f5f5f0f0fffff)
  ) CLBLM_L_X10Y104_SLICE_X12Y104_ALUT (
.I0(LIOB33_X0Y103_IOB_X0Y104_I),
.I1(1'b1),
.I2(RIOB33_X105Y103_IOB_X1Y104_I),
.I3(1'b1),
.I4(LIOB33_X0Y105_IOB_X0Y105_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y104_SLICE_X12Y104_AO5),
.O6(CLBLM_L_X10Y104_SLICE_X12Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y104_SLICE_X13Y104_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y104_SLICE_X13Y104_DO5),
.O6(CLBLM_L_X10Y104_SLICE_X13Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7d14ff3cdd44ffcc)
  ) CLBLM_L_X10Y104_SLICE_X13Y104_CLUT (
.I0(RIOB33_X105Y103_IOB_X1Y104_I),
.I1(CLBLM_L_X10Y103_SLICE_X13Y103_DO6),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X11Y106_SLICE_X14Y106_CO6),
.I4(LIOB33_X0Y103_IOB_X0Y104_I),
.I5(LIOB33_X0Y101_IOB_X0Y102_I),
.O5(CLBLM_L_X10Y104_SLICE_X13Y104_CO5),
.O6(CLBLM_L_X10Y104_SLICE_X13Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6c939393936c6c6c)
  ) CLBLM_L_X10Y104_SLICE_X13Y104_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X10Y103_SLICE_X13Y103_DO6),
.I2(LIOB33_X0Y101_IOB_X0Y102_I),
.I3(LIOB33_X0Y103_IOB_X0Y104_I),
.I4(RIOB33_X105Y103_IOB_X1Y104_I),
.I5(CLBLM_R_X11Y106_SLICE_X14Y106_CO6),
.O5(CLBLM_L_X10Y104_SLICE_X13Y104_BO5),
.O6(CLBLM_L_X10Y104_SLICE_X13Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h155ac05025aaf0a0)
  ) CLBLM_L_X10Y104_SLICE_X13Y104_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(RIOB33_X105Y111_IOB_X1Y112_I),
.I2(RIOB33_X105Y113_IOB_X1Y113_I),
.I3(RIOB33_X105Y107_IOB_X1Y107_I),
.I4(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I5(RIOB33_X105Y107_IOB_X1Y108_I),
.O5(CLBLM_L_X10Y104_SLICE_X13Y104_AO5),
.O6(CLBLM_L_X10Y104_SLICE_X13Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y105_SLICE_X12Y105_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y105_SLICE_X12Y105_DO5),
.O6(CLBLM_L_X10Y105_SLICE_X12Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h936cccccc9366666)
  ) CLBLM_L_X10Y105_SLICE_X12Y105_CLUT (
.I0(CLBLM_L_X10Y104_SLICE_X13Y104_BO6),
.I1(CLBLM_L_X10Y104_SLICE_X12Y104_BO6),
.I2(RIOB33_X105Y103_IOB_X1Y103_I),
.I3(RIOB33_X105Y103_IOB_X1Y104_I),
.I4(LIOB33_X0Y105_IOB_X0Y105_I),
.I5(CLBLM_L_X10Y106_SLICE_X13Y106_BO6),
.O5(CLBLM_L_X10Y105_SLICE_X12Y105_CO5),
.O6(CLBLM_L_X10Y105_SLICE_X12Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'heb82ebeb8282eb82)
  ) CLBLM_L_X10Y105_SLICE_X12Y105_BLUT (
.I0(CLBLM_L_X8Y105_SLICE_X10Y105_AO6),
.I1(CLBLM_L_X10Y104_SLICE_X12Y104_BO6),
.I2(CLBLM_L_X10Y104_SLICE_X12Y104_AO5),
.I3(CLBLM_L_X10Y106_SLICE_X13Y106_BO6),
.I4(CLBLM_L_X10Y104_SLICE_X13Y104_BO6),
.I5(CLBLM_L_X10Y106_SLICE_X12Y106_AO5),
.O5(CLBLM_L_X10Y105_SLICE_X12Y105_BO5),
.O6(CLBLM_L_X10Y105_SLICE_X12Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h69965aa5a55a6996)
  ) CLBLM_L_X10Y105_SLICE_X12Y105_ALUT (
.I0(CLBLM_L_X8Y105_SLICE_X10Y105_AO6),
.I1(CLBLM_L_X10Y106_SLICE_X13Y106_BO6),
.I2(CLBLM_L_X10Y104_SLICE_X12Y104_AO5),
.I3(CLBLM_L_X10Y104_SLICE_X12Y104_BO6),
.I4(CLBLM_L_X10Y104_SLICE_X13Y104_BO6),
.I5(CLBLM_L_X10Y106_SLICE_X12Y106_AO5),
.O5(CLBLM_L_X10Y105_SLICE_X12Y105_AO5),
.O6(CLBLM_L_X10Y105_SLICE_X12Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hda255da2708ff708)
  ) CLBLM_L_X10Y105_SLICE_X13Y105_DLUT (
.I0(LIOB33_X0Y101_IOB_X0Y102_I),
.I1(RIOB33_X105Y103_IOB_X1Y104_I),
.I2(CLBLM_L_X10Y106_SLICE_X13Y106_AO5),
.I3(CLBLM_L_X10Y103_SLICE_X13Y103_DO6),
.I4(CLBLM_L_X8Y101_SLICE_X11Y101_AO5),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X10Y105_SLICE_X13Y105_DO5),
.O6(CLBLM_L_X10Y105_SLICE_X13Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6ca0935f935f6ca0)
  ) CLBLM_L_X10Y105_SLICE_X13Y105_CLUT (
.I0(RIOB33_X105Y103_IOB_X1Y104_I),
.I1(LIOB33_X0Y105_IOB_X0Y105_I),
.I2(LIOB33_X0Y103_IOB_X0Y104_I),
.I3(RIOB33_X105Y103_IOB_X1Y103_I),
.I4(CLBLM_L_X10Y105_SLICE_X13Y105_DO6),
.I5(CLBLM_L_X10Y106_SLICE_X13Y106_BO6),
.O5(CLBLM_L_X10Y105_SLICE_X13Y105_CO5),
.O6(CLBLM_L_X10Y105_SLICE_X13Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7b12ff5abb22ffaa)
  ) CLBLM_L_X10Y105_SLICE_X13Y105_BLUT (
.I0(CLBLM_L_X10Y105_SLICE_X13Y105_DO6),
.I1(LIOB33_X0Y105_IOB_X0Y105_I),
.I2(LIOB33_X0Y103_IOB_X0Y104_I),
.I3(CLBLM_L_X10Y106_SLICE_X13Y106_BO6),
.I4(RIOB33_X105Y103_IOB_X1Y103_I),
.I5(RIOB33_X105Y103_IOB_X1Y104_I),
.O5(CLBLM_L_X10Y105_SLICE_X13Y105_BO5),
.O6(CLBLM_L_X10Y105_SLICE_X13Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h4500000065aaf000)
  ) CLBLM_L_X10Y105_SLICE_X13Y105_ALUT (
.I0(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I1(RIOB33_X105Y111_IOB_X1Y112_I),
.I2(RIOB33_X105Y107_IOB_X1Y107_I),
.I3(RIOB33_X105Y113_IOB_X1Y113_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(RIOB33_X105Y103_IOB_X1Y104_I),
.O5(CLBLM_L_X10Y105_SLICE_X13Y105_AO5),
.O6(CLBLM_L_X10Y105_SLICE_X13Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h9a65a6a659a6a6a6)
  ) CLBLM_L_X10Y106_SLICE_X12Y106_DLUT (
.I0(CLBLM_L_X10Y105_SLICE_X12Y105_CO6),
.I1(CLBLM_L_X10Y105_SLICE_X13Y105_CO6),
.I2(CLBLM_L_X10Y106_SLICE_X13Y106_DO6),
.I3(RIOB33_X105Y103_IOB_X1Y103_I),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(RIOB33_X105Y101_IOB_X1Y102_I),
.O5(CLBLM_L_X10Y106_SLICE_X12Y106_DO5),
.O6(CLBLM_L_X10Y106_SLICE_X12Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h69969696c33c3c3c)
  ) CLBLM_L_X10Y106_SLICE_X12Y106_CLUT (
.I0(LIOB33_X0Y105_IOB_X0Y105_I),
.I1(CLBLM_L_X10Y106_SLICE_X13Y106_CO6),
.I2(CLBLM_L_X10Y107_SLICE_X12Y107_DO6),
.I3(RIOB33_X105Y103_IOB_X1Y103_I),
.I4(LIOB33_X0Y103_IOB_X0Y104_I),
.I5(RIOB33_X105Y101_IOB_X1Y102_I),
.O5(CLBLM_L_X10Y106_SLICE_X12Y106_CO5),
.O6(CLBLM_L_X10Y106_SLICE_X12Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5a9696a5a569695a)
  ) CLBLM_L_X10Y106_SLICE_X12Y106_BLUT (
.I0(CLBLM_L_X10Y103_SLICE_X13Y103_AO6),
.I1(CLBLM_R_X11Y106_SLICE_X14Y106_BO6),
.I2(CLBLM_L_X10Y104_SLICE_X12Y104_AO6),
.I3(CLBLM_L_X10Y108_SLICE_X13Y108_DO6),
.I4(CLBLM_L_X10Y106_SLICE_X12Y106_AO6),
.I5(CLBLM_R_X11Y106_SLICE_X14Y106_CO6),
.O5(CLBLM_L_X10Y106_SLICE_X12Y106_BO5),
.O6(CLBLM_L_X10Y106_SLICE_X12Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h33ff33ff3333ffff)
  ) CLBLM_L_X10Y106_SLICE_X12Y106_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y103_IOB_X1Y103_I),
.I2(1'b1),
.I3(LIOB33_X0Y103_IOB_X0Y104_I),
.I4(LIOB33_X0Y105_IOB_X0Y105_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y106_SLICE_X12Y106_AO5),
.O6(CLBLM_L_X10Y106_SLICE_X12Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fd51540ffff3fc0)
  ) CLBLM_L_X10Y106_SLICE_X13Y106_DLUT (
.I0(RIOB33_X105Y101_IOB_X1Y102_I),
.I1(RIOB33_X105Y103_IOB_X1Y103_I),
.I2(LIOB33_X0Y103_IOB_X0Y104_I),
.I3(CLBLM_L_X10Y106_SLICE_X13Y106_CO6),
.I4(CLBLM_L_X10Y107_SLICE_X12Y107_DO6),
.I5(LIOB33_X0Y105_IOB_X0Y105_I),
.O5(CLBLM_L_X10Y106_SLICE_X13Y106_DO5),
.O6(CLBLM_L_X10Y106_SLICE_X13Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8e71f50a718ef50a)
  ) CLBLM_L_X10Y106_SLICE_X13Y106_CLUT (
.I0(CLBLM_L_X10Y106_SLICE_X13Y106_AO6),
.I1(RIOB33_X105Y103_IOB_X1Y103_I),
.I2(CLBLM_L_X10Y109_SLICE_X12Y109_AO5),
.I3(CLBLM_R_X11Y106_SLICE_X14Y106_DO6),
.I4(LIOB33_X0Y101_IOB_X0Y102_I),
.I5(RIOB33_X105Y103_IOB_X1Y104_I),
.O5(CLBLM_L_X10Y106_SLICE_X13Y106_CO5),
.O6(CLBLM_L_X10Y106_SLICE_X13Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7f15ff3fbf2a3f00)
  ) CLBLM_L_X10Y106_SLICE_X13Y106_BLUT (
.I0(LIOB33_X0Y101_IOB_X0Y102_I),
.I1(LIOB33_X0Y103_IOB_X0Y104_I),
.I2(RIOB33_X105Y103_IOB_X1Y103_I),
.I3(CLBLM_L_X10Y108_SLICE_X13Y108_DO6),
.I4(RIOB33_X105Y103_IOB_X1Y104_I),
.I5(CLBLM_R_X11Y106_SLICE_X14Y106_DO6),
.O5(CLBLM_L_X10Y106_SLICE_X13Y106_BO5),
.O6(CLBLM_L_X10Y106_SLICE_X13Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h99995555ff11ff55)
  ) CLBLM_L_X10Y106_SLICE_X13Y106_ALUT (
.I0(CLBLM_L_X10Y109_SLICE_X12Y109_BO6),
.I1(RIOB33_X105Y103_IOB_X1Y104_I),
.I2(1'b1),
.I3(CLBLM_L_X10Y105_SLICE_X13Y105_AO6),
.I4(LIOB33_X0Y101_IOB_X0Y101_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y106_SLICE_X13Y106_AO5),
.O6(CLBLM_L_X10Y106_SLICE_X13Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h70f7f770f770f770)
  ) CLBLM_L_X10Y107_SLICE_X12Y107_DLUT (
.I0(RIOB33_X105Y101_IOB_X1Y102_I),
.I1(LIOB33_X0Y103_IOB_X0Y104_I),
.I2(CLBLM_L_X8Y110_SLICE_X11Y110_DO6),
.I3(CLBLM_L_X10Y109_SLICE_X12Y109_CO6),
.I4(LIOB33_X0Y101_IOB_X0Y102_I),
.I5(RIOB33_X105Y103_IOB_X1Y103_I),
.O5(CLBLM_L_X10Y107_SLICE_X12Y107_DO5),
.O6(CLBLM_L_X10Y107_SLICE_X12Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7887877887788778)
  ) CLBLM_L_X10Y107_SLICE_X12Y107_CLUT (
.I0(RIOB33_X105Y101_IOB_X1Y102_I),
.I1(LIOB33_X0Y103_IOB_X0Y104_I),
.I2(CLBLM_L_X8Y110_SLICE_X11Y110_DO6),
.I3(CLBLM_L_X10Y109_SLICE_X12Y109_CO6),
.I4(LIOB33_X0Y101_IOB_X0Y102_I),
.I5(RIOB33_X105Y103_IOB_X1Y103_I),
.O5(CLBLM_L_X10Y107_SLICE_X12Y107_CO5),
.O6(CLBLM_L_X10Y107_SLICE_X12Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h693cc36996c33c96)
  ) CLBLM_L_X10Y107_SLICE_X12Y107_BLUT (
.I0(CLBLM_L_X8Y110_SLICE_X11Y110_DO6),
.I1(CLBLM_R_X11Y106_SLICE_X14Y106_BO6),
.I2(CLBLM_L_X10Y106_SLICE_X12Y106_AO6),
.I3(CLBLM_L_X10Y108_SLICE_X13Y108_BO6),
.I4(CLBLM_L_X10Y107_SLICE_X12Y107_AO6),
.I5(CLBLM_L_X10Y108_SLICE_X13Y108_DO6),
.O5(CLBLM_L_X10Y107_SLICE_X12Y107_BO5),
.O6(CLBLM_L_X10Y107_SLICE_X12Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f3f3f3f5f5f5f5f)
  ) CLBLM_L_X10Y107_SLICE_X12Y107_ALUT (
.I0(LIOB33_X0Y105_IOB_X0Y105_I),
.I1(LIOB33_X0Y103_IOB_X0Y104_I),
.I2(RIOB33_X105Y101_IOB_X1Y102_I),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y107_SLICE_X12Y107_AO5),
.O6(CLBLM_L_X10Y107_SLICE_X12Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hbc70438f3bf7c408)
  ) CLBLM_L_X10Y107_SLICE_X13Y107_DLUT (
.I0(RIOB33_X105Y101_IOB_X1Y102_I),
.I1(LIOB33_X0Y105_IOB_X0Y105_I),
.I2(CLBLM_L_X10Y107_SLICE_X12Y107_DO6),
.I3(RIOB33_X105Y103_IOB_X1Y103_I),
.I4(CLBLM_L_X10Y106_SLICE_X12Y106_BO6),
.I5(CLBLM_L_X10Y107_SLICE_X13Y107_BO6),
.O5(CLBLM_L_X10Y107_SLICE_X13Y107_DO5),
.O6(CLBLM_L_X10Y107_SLICE_X13Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hec80b320fec8fb32)
  ) CLBLM_L_X10Y107_SLICE_X13Y107_CLUT (
.I0(CLBLM_L_X10Y107_SLICE_X12Y107_AO5),
.I1(CLBLM_L_X10Y106_SLICE_X12Y106_AO5),
.I2(CLBLM_L_X10Y107_SLICE_X12Y107_DO6),
.I3(CLBLM_L_X10Y108_SLICE_X12Y108_AO5),
.I4(CLBLM_L_X10Y106_SLICE_X12Y106_BO6),
.I5(CLBLM_L_X10Y107_SLICE_X13Y107_BO6),
.O5(CLBLM_L_X10Y107_SLICE_X13Y107_CO5),
.O6(CLBLM_L_X10Y107_SLICE_X13Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996c33c96963c3c)
  ) CLBLM_L_X10Y107_SLICE_X13Y107_BLUT (
.I0(LIOB33_X0Y103_IOB_X0Y104_I),
.I1(CLBLM_L_X10Y108_SLICE_X13Y108_DO6),
.I2(CLBLM_R_X11Y106_SLICE_X14Y106_DO6),
.I3(LIOB33_X0Y101_IOB_X0Y102_I),
.I4(RIOB33_X105Y103_IOB_X1Y103_I),
.I5(RIOB33_X105Y103_IOB_X1Y104_I),
.O5(CLBLM_L_X10Y107_SLICE_X13Y107_BO5),
.O6(CLBLM_L_X10Y107_SLICE_X13Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3c9696c3c369693c)
  ) CLBLM_L_X10Y107_SLICE_X13Y107_ALUT (
.I0(CLBLM_L_X10Y107_SLICE_X13Y107_BO6),
.I1(CLBLM_L_X10Y108_SLICE_X12Y108_AO5),
.I2(CLBLM_L_X10Y106_SLICE_X12Y106_BO6),
.I3(CLBLM_L_X10Y107_SLICE_X12Y107_AO5),
.I4(CLBLM_L_X10Y107_SLICE_X12Y107_DO6),
.I5(CLBLM_L_X10Y106_SLICE_X12Y106_AO5),
.O5(CLBLM_L_X10Y107_SLICE_X13Y107_AO5),
.O6(CLBLM_L_X10Y107_SLICE_X13Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hb73f48c0c0b73f48)
  ) CLBLM_L_X10Y108_SLICE_X12Y108_DLUT (
.I0(RIOB33_X105Y101_IOB_X1Y101_I),
.I1(LIOB33_X0Y105_IOB_X0Y105_I),
.I2(RIOB33_X105Y101_IOB_X1Y102_I),
.I3(CLBLM_L_X10Y107_SLICE_X12Y107_CO6),
.I4(CLBLM_L_X10Y107_SLICE_X12Y107_BO6),
.I5(CLBLM_L_X8Y110_SLICE_X10Y110_BO6),
.O5(CLBLM_L_X10Y108_SLICE_X12Y108_DO5),
.O6(CLBLM_L_X10Y108_SLICE_X12Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf9f990f990f99090)
  ) CLBLM_L_X10Y108_SLICE_X12Y108_CLUT (
.I0(CLBLM_L_X10Y107_SLICE_X12Y107_AO5),
.I1(CLBLM_L_X10Y107_SLICE_X12Y107_BO6),
.I2(CLBLM_L_X10Y108_SLICE_X12Y108_AO6),
.I3(CLBLM_L_X10Y107_SLICE_X12Y107_CO6),
.I4(CLBLM_R_X7Y110_SLICE_X9Y110_AO5),
.I5(CLBLM_L_X8Y110_SLICE_X10Y110_BO6),
.O5(CLBLM_L_X10Y108_SLICE_X12Y108_CO5),
.O6(CLBLM_L_X10Y108_SLICE_X12Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h69c3963c3c69c396)
  ) CLBLM_L_X10Y108_SLICE_X12Y108_BLUT (
.I0(CLBLM_R_X7Y110_SLICE_X9Y110_AO5),
.I1(CLBLM_L_X10Y107_SLICE_X12Y107_BO6),
.I2(CLBLM_L_X10Y107_SLICE_X12Y107_AO5),
.I3(CLBLM_L_X8Y110_SLICE_X10Y110_BO6),
.I4(CLBLM_L_X10Y108_SLICE_X12Y108_AO6),
.I5(CLBLM_L_X10Y107_SLICE_X12Y107_CO6),
.O5(CLBLM_L_X10Y108_SLICE_X12Y108_BO5),
.O6(CLBLM_L_X10Y108_SLICE_X12Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f3f3f3f0f0fffff)
  ) CLBLM_L_X10Y108_SLICE_X12Y108_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y101_IOB_X1Y101_I),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(1'b1),
.I4(RIOB33_X105Y101_IOB_X1Y102_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y108_SLICE_X12Y108_AO5),
.O6(CLBLM_L_X10Y108_SLICE_X12Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffccce08ff333b02)
  ) CLBLM_L_X10Y108_SLICE_X13Y108_DLUT (
.I0(CLBLM_L_X10Y108_SLICE_X13Y108_AO6),
.I1(CLBLM_R_X11Y106_SLICE_X14Y106_AO6),
.I2(CLBLM_L_X10Y109_SLICE_X12Y109_DO6),
.I3(CLBLM_L_X10Y108_SLICE_X13Y108_AO5),
.I4(CLBLM_L_X10Y108_SLICE_X13Y108_CO6),
.I5(CLBLM_L_X10Y109_SLICE_X12Y109_BO6),
.O5(CLBLM_L_X10Y108_SLICE_X13Y108_DO5),
.O6(CLBLM_L_X10Y108_SLICE_X13Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h1131aa0a20202020)
  ) CLBLM_L_X10Y108_SLICE_X13Y108_CLUT (
.I0(RIOB33_X105Y113_IOB_X1Y113_I),
.I1(RIOB33_X105Y103_IOB_X1Y103_I),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(RIOB33_X105Y111_IOB_X1Y112_I),
.I4(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I5(RIOB33_X105Y103_IOB_X1Y104_I),
.O5(CLBLM_L_X10Y108_SLICE_X13Y108_CO5),
.O6(CLBLM_L_X10Y108_SLICE_X13Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h695a696996a59696)
  ) CLBLM_L_X10Y108_SLICE_X13Y108_BLUT (
.I0(CLBLM_L_X10Y109_SLICE_X12Y109_BO6),
.I1(CLBLM_L_X10Y108_SLICE_X13Y108_CO6),
.I2(CLBLM_R_X11Y106_SLICE_X14Y106_AO6),
.I3(CLBLM_L_X10Y109_SLICE_X12Y109_DO6),
.I4(CLBLM_L_X10Y108_SLICE_X13Y108_AO6),
.I5(CLBLM_L_X10Y108_SLICE_X13Y108_AO5),
.O5(CLBLM_L_X10Y108_SLICE_X13Y108_BO5),
.O6(CLBLM_L_X10Y108_SLICE_X13Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ffffff0fff0fff)
  ) CLBLM_L_X10Y108_SLICE_X13Y108_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(LIOB33_X0Y101_IOB_X0Y102_I),
.I3(RIOB33_X105Y103_IOB_X1Y103_I),
.I4(LIOB33_X0Y101_IOB_X0Y101_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y108_SLICE_X13Y108_AO5),
.O6(CLBLM_L_X10Y108_SLICE_X13Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h13a019aa6622cc88)
  ) CLBLM_L_X10Y109_SLICE_X12Y109_DLUT (
.I0(RIOB33_X105Y113_IOB_X1Y113_I),
.I1(RIOB33_X105Y103_IOB_X1Y103_I),
.I2(RIOB33_X105Y111_IOB_X1Y112_I),
.I3(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(RIOB33_X105Y103_IOB_X1Y104_I),
.O5(CLBLM_L_X10Y109_SLICE_X12Y109_DO5),
.O6(CLBLM_L_X10Y109_SLICE_X12Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5aaa4fbfa555b040)
  ) CLBLM_L_X10Y109_SLICE_X12Y109_CLUT (
.I0(CLBLM_L_X10Y108_SLICE_X13Y108_CO6),
.I1(RIOB33_X105Y103_IOB_X1Y103_I),
.I2(LIOB33_X0Y101_IOB_X0Y101_I),
.I3(RIOB33_X105Y103_IOB_X1Y104_I),
.I4(CLBLM_L_X10Y109_SLICE_X12Y109_DO6),
.I5(CLBLM_L_X10Y109_SLICE_X12Y109_BO6),
.O5(CLBLM_L_X10Y109_SLICE_X12Y109_CO5),
.O6(CLBLM_L_X10Y109_SLICE_X12Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h13b355004ce6aa00)
  ) CLBLM_L_X10Y109_SLICE_X12Y109_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(RIOB33_X105Y107_IOB_X1Y107_I),
.I2(RIOB33_X105Y111_IOB_X1Y112_I),
.I3(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I4(RIOB33_X105Y113_IOB_X1Y113_I),
.I5(RIOB33_X105Y103_IOB_X1Y104_I),
.O5(CLBLM_L_X10Y109_SLICE_X12Y109_BO5),
.O6(CLBLM_L_X10Y109_SLICE_X12Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha5a55555cdcddddd)
  ) CLBLM_L_X10Y109_SLICE_X12Y109_ALUT (
.I0(CLBLM_L_X10Y109_SLICE_X12Y109_DO6),
.I1(CLBLM_L_X10Y108_SLICE_X13Y108_CO6),
.I2(LIOB33_X0Y101_IOB_X0Y101_I),
.I3(1'b1),
.I4(RIOB33_X105Y103_IOB_X1Y103_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y109_SLICE_X12Y109_AO5),
.O6(CLBLM_L_X10Y109_SLICE_X12Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y109_SLICE_X13Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y109_SLICE_X13Y109_DO5),
.O6(CLBLM_L_X10Y109_SLICE_X13Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y109_SLICE_X13Y109_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y109_SLICE_X13Y109_CO5),
.O6(CLBLM_L_X10Y109_SLICE_X13Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y109_SLICE_X13Y109_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y109_SLICE_X13Y109_BO5),
.O6(CLBLM_L_X10Y109_SLICE_X13Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y109_SLICE_X13Y109_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y109_SLICE_X13Y109_AO5),
.O6(CLBLM_L_X10Y109_SLICE_X13Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y100_SLICE_X2Y100_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y100_SLICE_X2Y100_DO5),
.O6(CLBLM_R_X3Y100_SLICE_X2Y100_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y100_SLICE_X2Y100_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y100_SLICE_X2Y100_CO5),
.O6(CLBLM_R_X3Y100_SLICE_X2Y100_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y100_SLICE_X2Y100_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y100_SLICE_X2Y100_BO5),
.O6(CLBLM_R_X3Y100_SLICE_X2Y100_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y100_SLICE_X2Y100_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y100_SLICE_X2Y100_AO5),
.O6(CLBLM_R_X3Y100_SLICE_X2Y100_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y100_SLICE_X3Y100_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y100_SLICE_X3Y100_DO5),
.O6(CLBLM_R_X3Y100_SLICE_X3Y100_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y100_SLICE_X3Y100_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y100_SLICE_X3Y100_CO5),
.O6(CLBLM_R_X3Y100_SLICE_X3Y100_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7f13b320ff5fffa0)
  ) CLBLM_R_X3Y100_SLICE_X3Y100_BLUT (
.I0(LIOB33_X0Y107_IOB_X0Y107_I),
.I1(RIOB33_X105Y109_IOB_X1Y109_I),
.I2(RIOB33_X105Y109_IOB_X1Y110_I),
.I3(CLBLL_L_X4Y100_SLICE_X4Y100_AO6),
.I4(CLBLL_L_X4Y100_SLICE_X4Y100_BO6),
.I5(LIOB33_X0Y107_IOB_X0Y108_I),
.O5(CLBLM_R_X3Y100_SLICE_X3Y100_BO5),
.O6(CLBLM_R_X3Y100_SLICE_X3Y100_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f3f3f3f7711ff55)
  ) CLBLM_R_X3Y100_SLICE_X3Y100_ALUT (
.I0(CLBLM_R_X3Y101_SLICE_X3Y101_DO6),
.I1(RIOB33_X105Y109_IOB_X1Y109_I),
.I2(LIOB33_X0Y101_IOB_X0Y101_I),
.I3(CLBLM_R_X3Y100_SLICE_X3Y100_BO6),
.I4(LIOB33_X0Y109_IOB_X0Y109_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y100_SLICE_X3Y100_AO5),
.O6(CLBLM_R_X3Y100_SLICE_X3Y100_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y101_SLICE_X2Y101_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y101_SLICE_X2Y101_DO5),
.O6(CLBLM_R_X3Y101_SLICE_X2Y101_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y101_SLICE_X2Y101_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y101_SLICE_X2Y101_CO5),
.O6(CLBLM_R_X3Y101_SLICE_X2Y101_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y101_SLICE_X2Y101_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y101_SLICE_X2Y101_BO5),
.O6(CLBLM_R_X3Y101_SLICE_X2Y101_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y101_SLICE_X2Y101_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y101_SLICE_X2Y101_AO5),
.O6(CLBLM_R_X3Y101_SLICE_X2Y101_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hd887882878d88828)
  ) CLBLM_R_X3Y101_SLICE_X3Y101_DLUT (
.I0(RIOB33_X105Y109_IOB_X1Y110_I),
.I1(LIOB33_X0Y107_IOB_X0Y108_I),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(CLBLL_L_X4Y101_SLICE_X4Y101_DO6),
.I4(RIOB33_X105Y111_IOB_X1Y111_I),
.I5(LIOB33_X0Y105_IOB_X0Y106_I),
.O5(CLBLM_R_X3Y101_SLICE_X3Y101_DO5),
.O6(CLBLM_R_X3Y101_SLICE_X3Y101_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hda4f25b02abfd540)
  ) CLBLM_R_X3Y101_SLICE_X3Y101_CLUT (
.I0(CLBLL_L_X4Y100_SLICE_X4Y100_AO6),
.I1(LIOB33_X0Y107_IOB_X0Y108_I),
.I2(RIOB33_X105Y109_IOB_X1Y109_I),
.I3(CLBLM_R_X3Y101_SLICE_X3Y101_AO5),
.I4(CLBLM_R_X3Y101_SLICE_X3Y101_DO6),
.I5(LIOB33_X0Y109_IOB_X0Y109_I),
.O5(CLBLM_R_X3Y101_SLICE_X3Y101_CO5),
.O6(CLBLM_R_X3Y101_SLICE_X3Y101_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcbeb6f3f7f3f3f3f)
  ) CLBLM_R_X3Y101_SLICE_X3Y101_BLUT (
.I0(CLBLL_L_X4Y101_SLICE_X4Y101_DO6),
.I1(LIOB33_X0Y107_IOB_X0Y108_I),
.I2(RIOB33_X105Y111_IOB_X1Y111_I),
.I3(LIOB33_X0Y105_IOB_X0Y106_I),
.I4(RIOB33_X105Y109_IOB_X1Y110_I),
.I5(LIOB33_X0Y107_IOB_X0Y107_I),
.O5(CLBLM_R_X3Y101_SLICE_X3Y101_BO5),
.O6(CLBLM_R_X3Y101_SLICE_X3Y101_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa5500ffc3c30f0f)
  ) CLBLM_R_X3Y101_SLICE_X3Y101_ALUT (
.I0(LIOB33_X0Y109_IOB_X0Y109_I),
.I1(LIOB33_X0Y107_IOB_X0Y107_I),
.I2(CLBLL_L_X4Y100_SLICE_X4Y100_BO6),
.I3(CLBLM_R_X3Y101_SLICE_X3Y101_BO6),
.I4(RIOB33_X105Y109_IOB_X1Y110_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y101_SLICE_X3Y101_AO5),
.O6(CLBLM_R_X3Y101_SLICE_X3Y101_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y102_SLICE_X2Y102_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y102_SLICE_X2Y102_DO5),
.O6(CLBLM_R_X3Y102_SLICE_X2Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h69969696c33c3c3c)
  ) CLBLM_R_X3Y102_SLICE_X2Y102_CLUT (
.I0(LIOB33_X0Y111_IOB_X0Y111_I),
.I1(CLBLM_R_X3Y102_SLICE_X3Y102_AO6),
.I2(CLBLL_L_X2Y102_SLICE_X1Y102_BO6),
.I3(LIOB33_X0Y111_IOB_X0Y112_I),
.I4(RIOB33_X105Y109_IOB_X1Y109_I),
.I5(RIOB33_X105Y109_IOB_X1Y110_I),
.O5(CLBLM_R_X3Y102_SLICE_X2Y102_CO5),
.O6(CLBLM_R_X3Y102_SLICE_X2Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h9cccf000c63c5a00)
  ) CLBLM_R_X3Y102_SLICE_X2Y102_BLUT (
.I0(LIOB33_X0Y107_IOB_X0Y108_I),
.I1(LIOB33_X0Y109_IOB_X0Y110_I),
.I2(LIOB33_X0Y109_IOB_X0Y109_I),
.I3(RIOB33_X105Y111_IOB_X1Y111_I),
.I4(RIOB33_X105Y109_IOB_X1Y110_I),
.I5(CLBLL_L_X2Y102_SLICE_X1Y102_AO6),
.O5(CLBLM_R_X3Y102_SLICE_X2Y102_BO5),
.O6(CLBLM_R_X3Y102_SLICE_X2Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h71f5b2faf3ff30f0)
  ) CLBLM_R_X3Y102_SLICE_X2Y102_ALUT (
.I0(LIOB33_X0Y111_IOB_X0Y111_I),
.I1(RIOB33_X105Y109_IOB_X1Y109_I),
.I2(CLBLM_R_X3Y102_SLICE_X3Y102_AO6),
.I3(LIOB33_X0Y111_IOB_X0Y112_I),
.I4(CLBLL_L_X2Y102_SLICE_X1Y102_BO6),
.I5(RIOB33_X105Y109_IOB_X1Y110_I),
.O5(CLBLM_R_X3Y102_SLICE_X2Y102_AO5),
.O6(CLBLM_R_X3Y102_SLICE_X2Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h303370f773f7ffff)
  ) CLBLM_R_X3Y102_SLICE_X3Y102_DLUT (
.I0(LIOB33_X0Y111_IOB_X0Y111_I),
.I1(RIOB33_X105Y107_IOB_X1Y108_I),
.I2(CLBLL_L_X4Y102_SLICE_X5Y102_DO6),
.I3(CLBLM_R_X3Y102_SLICE_X3Y102_CO6),
.I4(LIOB33_X0Y111_IOB_X0Y112_I),
.I5(CLBLM_R_X3Y102_SLICE_X3Y102_BO6),
.O5(CLBLM_R_X3Y102_SLICE_X3Y102_DO5),
.O6(CLBLM_R_X3Y102_SLICE_X3Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6c93a05f936c5fa0)
  ) CLBLM_R_X3Y102_SLICE_X3Y102_CLUT (
.I0(RIOB33_X105Y109_IOB_X1Y109_I),
.I1(RIOB33_X105Y109_IOB_X1Y110_I),
.I2(LIOB33_X0Y109_IOB_X0Y110_I),
.I3(CLBLM_R_X3Y100_SLICE_X3Y100_AO5),
.I4(LIOB33_X0Y109_IOB_X0Y109_I),
.I5(CLBLM_R_X3Y101_SLICE_X3Y101_BO6),
.O5(CLBLM_R_X3Y102_SLICE_X3Y102_CO5),
.O6(CLBLM_R_X3Y102_SLICE_X3Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h93cc6cccc93c363c)
  ) CLBLM_R_X3Y102_SLICE_X3Y102_BLUT (
.I0(LIOB33_X0Y109_IOB_X0Y110_I),
.I1(CLBLM_R_X3Y102_SLICE_X2Y102_BO6),
.I2(CLBLM_R_X3Y101_SLICE_X3Y101_AO6),
.I3(RIOB33_X105Y109_IOB_X1Y109_I),
.I4(LIOB33_X0Y111_IOB_X0Y111_I),
.I5(CLBLM_R_X3Y100_SLICE_X3Y100_AO5),
.O5(CLBLM_R_X3Y102_SLICE_X3Y102_BO5),
.O6(CLBLM_R_X3Y102_SLICE_X3Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h13ff7fff013f373f)
  ) CLBLM_R_X3Y102_SLICE_X3Y102_ALUT (
.I0(LIOB33_X0Y109_IOB_X0Y110_I),
.I1(CLBLM_R_X3Y102_SLICE_X2Y102_BO6),
.I2(CLBLM_R_X3Y101_SLICE_X3Y101_AO6),
.I3(RIOB33_X105Y109_IOB_X1Y109_I),
.I4(LIOB33_X0Y111_IOB_X0Y111_I),
.I5(CLBLM_R_X3Y100_SLICE_X3Y100_AO5),
.O5(CLBLM_R_X3Y102_SLICE_X3Y102_AO5),
.O6(CLBLM_R_X3Y102_SLICE_X3Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y103_SLICE_X2Y103_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y103_SLICE_X2Y103_DO5),
.O6(CLBLM_R_X3Y103_SLICE_X2Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h377713177fff575f)
  ) CLBLM_R_X3Y103_SLICE_X2Y103_CLUT (
.I0(CLBLL_L_X2Y103_SLICE_X1Y103_AO5),
.I1(RIOB33_X105Y103_IOB_X1Y103_I),
.I2(CLBLL_L_X4Y102_SLICE_X4Y102_BO6),
.I3(LIOB33_X0Y111_IOB_X0Y111_I),
.I4(CLBLM_R_X5Y103_SLICE_X6Y103_DO6),
.I5(LIOB33_X0Y111_IOB_X0Y112_I),
.O5(CLBLM_R_X3Y103_SLICE_X2Y103_CO5),
.O6(CLBLM_R_X3Y103_SLICE_X2Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6a95c03f956a3fc0)
  ) CLBLM_R_X3Y103_SLICE_X2Y103_BLUT (
.I0(LIOB33_X0Y113_IOB_X0Y113_I),
.I1(RIOB33_X105Y103_IOB_X1Y103_I),
.I2(LIOB33_X0Y111_IOB_X0Y112_I),
.I3(CLBLL_L_X4Y102_SLICE_X4Y102_CO6),
.I4(RIOB33_X105Y101_IOB_X1Y102_I),
.I5(CLBLL_L_X4Y103_SLICE_X5Y103_DO6),
.O5(CLBLM_R_X3Y103_SLICE_X2Y103_BO5),
.O6(CLBLM_R_X3Y103_SLICE_X2Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5aa5f00f50f5f0ff)
  ) CLBLM_R_X3Y103_SLICE_X2Y103_ALUT (
.I0(LIOB33_X0Y113_IOB_X0Y113_I),
.I1(1'b1),
.I2(CLBLM_R_X3Y102_SLICE_X2Y102_AO6),
.I3(CLBLL_L_X2Y103_SLICE_X1Y103_CO6),
.I4(RIOB33_X105Y109_IOB_X1Y109_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y103_SLICE_X2Y103_AO5),
.O6(CLBLM_R_X3Y103_SLICE_X2Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h007171fff3f3ffff)
  ) CLBLM_R_X3Y103_SLICE_X3Y103_DLUT (
.I0(LIOB33_X0Y113_IOB_X0Y113_I),
.I1(CLBLM_R_X3Y102_SLICE_X2Y102_CO6),
.I2(CLBLM_R_X3Y102_SLICE_X3Y102_DO6),
.I3(LIOB33_X0Y115_IOB_X0Y115_I),
.I4(CLBLM_R_X3Y103_SLICE_X2Y103_AO6),
.I5(RIOB33_X105Y107_IOB_X1Y108_I),
.O5(CLBLM_R_X3Y103_SLICE_X3Y103_DO5),
.O6(CLBLM_R_X3Y103_SLICE_X3Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hb24d4db2dddd2222)
  ) CLBLM_R_X3Y103_SLICE_X3Y103_CLUT (
.I0(CLBLM_R_X3Y102_SLICE_X2Y102_CO6),
.I1(CLBLM_R_X3Y102_SLICE_X3Y102_DO6),
.I2(LIOB33_X0Y113_IOB_X0Y113_I),
.I3(LIOB33_X0Y115_IOB_X0Y115_I),
.I4(CLBLM_R_X3Y103_SLICE_X2Y103_AO6),
.I5(RIOB33_X105Y107_IOB_X1Y108_I),
.O5(CLBLM_R_X3Y103_SLICE_X3Y103_CO5),
.O6(CLBLM_R_X3Y103_SLICE_X3Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h2888beeebeeebeee)
  ) CLBLM_R_X3Y103_SLICE_X3Y103_BLUT (
.I0(CLBLL_L_X4Y103_SLICE_X5Y103_DO6),
.I1(CLBLL_L_X4Y102_SLICE_X4Y102_CO6),
.I2(LIOB33_X0Y111_IOB_X0Y112_I),
.I3(RIOB33_X105Y103_IOB_X1Y103_I),
.I4(RIOB33_X105Y101_IOB_X1Y102_I),
.I5(LIOB33_X0Y113_IOB_X0Y113_I),
.O5(CLBLM_R_X3Y103_SLICE_X3Y103_BO5),
.O6(CLBLM_R_X3Y103_SLICE_X3Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0fffff6a956a95)
  ) CLBLM_R_X3Y103_SLICE_X3Y103_ALUT (
.I0(CLBLM_R_X3Y102_SLICE_X3Y102_DO6),
.I1(RIOB33_X105Y107_IOB_X1Y108_I),
.I2(LIOB33_X0Y113_IOB_X0Y113_I),
.I3(CLBLM_R_X3Y102_SLICE_X2Y102_CO6),
.I4(RIOB33_X105Y101_IOB_X1Y101_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y103_SLICE_X3Y103_AO5),
.O6(CLBLM_R_X3Y103_SLICE_X3Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y104_SLICE_X2Y104_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y104_SLICE_X2Y104_DO5),
.O6(CLBLM_R_X3Y104_SLICE_X2Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h4dcfddff8e0ceecc)
  ) CLBLM_R_X3Y104_SLICE_X2Y104_CLUT (
.I0(LIOB33_X0Y113_IOB_X0Y113_I),
.I1(CLBLM_R_X3Y103_SLICE_X2Y103_AO5),
.I2(LIOB33_X0Y115_IOB_X0Y115_I),
.I3(RIOB33_X105Y109_IOB_X1Y110_I),
.I4(RIOB33_X105Y109_IOB_X1Y109_I),
.I5(CLBLM_R_X3Y104_SLICE_X2Y104_BO6),
.O5(CLBLM_R_X3Y104_SLICE_X2Y104_CO5),
.O6(CLBLM_R_X3Y104_SLICE_X2Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hba205ddfddffffff)
  ) CLBLM_R_X3Y104_SLICE_X2Y104_BLUT (
.I0(LIOB33_X0Y111_IOB_X0Y111_I),
.I1(CLBLL_L_X2Y103_SLICE_X1Y103_DO6),
.I2(LIOB33_X0Y109_IOB_X0Y110_I),
.I3(RIOB33_X105Y109_IOB_X1Y110_I),
.I4(LIOB33_X0Y111_IOB_X0Y112_I),
.I5(RIOB33_X105Y111_IOB_X1Y111_I),
.O5(CLBLM_R_X3Y104_SLICE_X2Y104_BO5),
.O6(CLBLM_R_X3Y104_SLICE_X2Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6c93a05f936c5fa0)
  ) CLBLM_R_X3Y104_SLICE_X2Y104_ALUT (
.I0(RIOB33_X105Y109_IOB_X1Y110_I),
.I1(RIOB33_X105Y109_IOB_X1Y109_I),
.I2(LIOB33_X0Y113_IOB_X0Y113_I),
.I3(CLBLM_R_X3Y104_SLICE_X2Y104_BO6),
.I4(LIOB33_X0Y115_IOB_X0Y115_I),
.I5(CLBLM_R_X3Y103_SLICE_X2Y103_AO5),
.O5(CLBLM_R_X3Y104_SLICE_X2Y104_AO5),
.O6(CLBLM_R_X3Y104_SLICE_X2Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haa5555aaaa55aa55)
  ) CLBLM_R_X3Y104_SLICE_X3Y104_DLUT (
.I0(CLBLM_R_X3Y103_SLICE_X3Y103_CO6),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X3Y104_SLICE_X3Y104_AO5),
.I4(CLBLL_L_X4Y104_SLICE_X4Y104_CO6),
.I5(CLBLL_L_X2Y104_SLICE_X0Y104_CO6),
.O5(CLBLM_R_X3Y104_SLICE_X3Y104_DO5),
.O6(CLBLM_R_X3Y104_SLICE_X3Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hc440fddccc44ffdd)
  ) CLBLM_R_X3Y104_SLICE_X3Y104_CLUT (
.I0(CLBLM_R_X3Y103_SLICE_X3Y103_CO6),
.I1(CLBLM_R_X3Y103_SLICE_X3Y103_DO6),
.I2(CLBLL_L_X4Y104_SLICE_X4Y104_CO6),
.I3(CLBLM_R_X3Y104_SLICE_X3Y104_AO5),
.I4(CLBLM_R_X3Y104_SLICE_X2Y104_AO6),
.I5(CLBLL_L_X2Y104_SLICE_X0Y104_CO6),
.O5(CLBLM_R_X3Y104_SLICE_X3Y104_CO5),
.O6(CLBLM_R_X3Y104_SLICE_X3Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h96c3c3c33c3c96c3)
  ) CLBLM_R_X3Y104_SLICE_X3Y104_BLUT (
.I0(CLBLL_L_X4Y104_SLICE_X4Y104_CO6),
.I1(CLBLM_R_X3Y103_SLICE_X3Y103_DO6),
.I2(CLBLM_R_X3Y104_SLICE_X2Y104_AO6),
.I3(CLBLL_L_X2Y104_SLICE_X0Y104_CO6),
.I4(CLBLM_R_X3Y103_SLICE_X3Y103_CO6),
.I5(CLBLM_R_X3Y104_SLICE_X3Y104_AO5),
.O5(CLBLM_R_X3Y104_SLICE_X3Y104_BO5),
.O6(CLBLM_R_X3Y104_SLICE_X3Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5f5f5f5f44ccddff)
  ) CLBLM_R_X3Y104_SLICE_X3Y104_ALUT (
.I0(LIOB33_X0Y115_IOB_X0Y115_I),
.I1(CLBLL_L_X4Y103_SLICE_X4Y103_CO6),
.I2(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I3(RIOB33_X105Y107_IOB_X1Y107_I),
.I4(CLBLM_R_X3Y103_SLICE_X3Y103_AO5),
.I5(1'b1),
.O5(CLBLM_R_X3Y104_SLICE_X3Y104_AO5),
.O6(CLBLM_R_X3Y104_SLICE_X3Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y105_SLICE_X2Y105_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y105_SLICE_X2Y105_DO5),
.O6(CLBLM_R_X3Y105_SLICE_X2Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3110c440c4403110)
  ) CLBLM_R_X3Y105_SLICE_X2Y105_CLUT (
.I0(CLBLL_L_X4Y104_SLICE_X4Y104_AO6),
.I1(CLBLM_R_X3Y103_SLICE_X2Y103_BO6),
.I2(CLBLL_L_X4Y105_SLICE_X4Y105_CO6),
.I3(CLBLM_R_X3Y106_SLICE_X2Y106_AO6),
.I4(CLBLL_L_X4Y104_SLICE_X4Y104_AO5),
.I5(CLBLL_L_X2Y106_SLICE_X1Y106_AO6),
.O5(CLBLM_R_X3Y105_SLICE_X2Y105_CO5),
.O6(CLBLM_R_X3Y105_SLICE_X2Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h69c33c69963cc396)
  ) CLBLM_R_X3Y105_SLICE_X2Y105_BLUT (
.I0(CLBLL_L_X4Y105_SLICE_X4Y105_CO6),
.I1(CLBLM_R_X3Y103_SLICE_X2Y103_BO6),
.I2(CLBLL_L_X4Y104_SLICE_X4Y104_AO5),
.I3(CLBLM_R_X3Y106_SLICE_X2Y106_AO6),
.I4(CLBLL_L_X4Y104_SLICE_X4Y104_AO6),
.I5(CLBLL_L_X2Y106_SLICE_X1Y106_AO6),
.O5(CLBLM_R_X3Y105_SLICE_X2Y105_BO5),
.O6(CLBLM_R_X3Y105_SLICE_X2Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h66aa995522aabbff)
  ) CLBLM_R_X3Y105_SLICE_X2Y105_ALUT (
.I0(CLBLL_L_X4Y105_SLICE_X4Y105_CO6),
.I1(LIOB33_X0Y115_IOB_X0Y115_I),
.I2(1'b1),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(CLBLL_L_X4Y104_SLICE_X4Y104_AO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y105_SLICE_X2Y105_AO5),
.O6(CLBLM_R_X3Y105_SLICE_X2Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y105_SLICE_X3Y105_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y105_SLICE_X3Y105_DO5),
.O6(CLBLM_R_X3Y105_SLICE_X3Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hb487788778b47878)
  ) CLBLM_R_X3Y105_SLICE_X3Y105_CLUT (
.I0(LIOB33_X0Y113_IOB_X0Y113_I),
.I1(LIOB33_X0Y115_IOB_X0Y116_I),
.I2(CLBLM_R_X5Y105_SLICE_X6Y105_DO6),
.I3(CLBLL_L_X4Y106_SLICE_X4Y106_CO6),
.I4(LIOB33_X0Y111_IOB_X0Y112_I),
.I5(CLBLL_L_X4Y105_SLICE_X5Y105_AO6),
.O5(CLBLM_R_X3Y105_SLICE_X3Y105_CO5),
.O6(CLBLM_R_X3Y105_SLICE_X3Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h022f0bbfbbffbbff)
  ) CLBLM_R_X3Y105_SLICE_X3Y105_BLUT (
.I0(CLBLL_L_X4Y106_SLICE_X4Y106_CO6),
.I1(CLBLL_L_X4Y105_SLICE_X5Y105_AO6),
.I2(LIOB33_X0Y113_IOB_X0Y113_I),
.I3(CLBLM_R_X5Y105_SLICE_X6Y105_DO6),
.I4(LIOB33_X0Y111_IOB_X0Y112_I),
.I5(LIOB33_X0Y115_IOB_X0Y116_I),
.O5(CLBLM_R_X3Y105_SLICE_X3Y105_BO5),
.O6(CLBLM_R_X3Y105_SLICE_X3Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h963cccccc39633cc)
  ) CLBLM_R_X3Y105_SLICE_X3Y105_ALUT (
.I0(LIOB33_X0Y115_IOB_X0Y116_I),
.I1(CLBLM_R_X5Y105_SLICE_X6Y105_BO6),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(CLBLL_L_X4Y105_SLICE_X5Y105_AO6),
.I4(LIOB33_X0Y111_IOB_X0Y112_I),
.I5(CLBLL_L_X4Y106_SLICE_X4Y106_CO6),
.O5(CLBLM_R_X3Y105_SLICE_X3Y105_AO5),
.O6(CLBLM_R_X3Y105_SLICE_X3Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000007510df45)
  ) CLBLM_R_X3Y106_SLICE_X2Y106_DLUT (
.I0(CLBLM_R_X3Y105_SLICE_X2Y105_AO6),
.I1(CLBLM_R_X3Y107_SLICE_X3Y107_BO6),
.I2(CLBLM_R_X3Y107_SLICE_X2Y107_DO6),
.I3(CLBLM_R_X3Y106_SLICE_X2Y106_CO6),
.I4(CLBLL_L_X2Y107_SLICE_X1Y107_BO6),
.I5(CLBLM_R_X3Y105_SLICE_X2Y105_BO6),
.O5(CLBLM_R_X3Y106_SLICE_X2Y106_DO5),
.O6(CLBLM_R_X3Y106_SLICE_X2Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h2b8e8e8ebbeeeeee)
  ) CLBLM_R_X3Y106_SLICE_X2Y106_CLUT (
.I0(CLBLM_R_X3Y105_SLICE_X3Y105_BO6),
.I1(CLBLL_L_X4Y105_SLICE_X4Y105_BO6),
.I2(LIOB33_X0Y115_IOB_X0Y115_I),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(LIOB33_X0Y113_IOB_X0Y113_I),
.I5(LIOB33_X0Y115_IOB_X0Y116_I),
.O5(CLBLM_R_X3Y106_SLICE_X2Y106_CO5),
.O6(CLBLM_R_X3Y106_SLICE_X2Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6c93936c93936c6c)
  ) CLBLM_R_X3Y106_SLICE_X2Y106_BLUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(CLBLL_L_X4Y105_SLICE_X4Y105_BO6),
.I2(LIOB33_X0Y113_IOB_X0Y113_I),
.I3(LIOB33_X0Y115_IOB_X0Y116_I),
.I4(CLBLM_R_X3Y105_SLICE_X3Y105_BO6),
.I5(LIOB33_X0Y115_IOB_X0Y115_I),
.O5(CLBLM_R_X3Y106_SLICE_X2Y106_BO5),
.O6(CLBLM_R_X3Y106_SLICE_X2Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f3f3f3f33ff33ff)
  ) CLBLM_R_X3Y106_SLICE_X2Y106_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y115_IOB_X0Y115_I),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(LIOB33_X0Y115_IOB_X0Y116_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y106_SLICE_X2Y106_AO5),
.O6(CLBLM_R_X3Y106_SLICE_X2Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y106_SLICE_X3Y106_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y106_SLICE_X3Y106_DO5),
.O6(CLBLM_R_X3Y106_SLICE_X3Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fd51540ffff3fc0)
  ) CLBLM_R_X3Y106_SLICE_X3Y106_CLUT (
.I0(RIOB33_X105Y101_IOB_X1Y102_I),
.I1(RIOB33_X105Y103_IOB_X1Y103_I),
.I2(LIOB33_X0Y113_IOB_X0Y113_I),
.I3(CLBLM_R_X3Y106_SLICE_X3Y106_AO5),
.I4(CLBLM_R_X3Y103_SLICE_X3Y103_BO6),
.I5(LIOB33_X0Y115_IOB_X0Y115_I),
.O5(CLBLM_R_X3Y106_SLICE_X3Y106_CO5),
.O6(CLBLM_R_X3Y106_SLICE_X3Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h69c3a50f963c5af0)
  ) CLBLM_R_X3Y106_SLICE_X3Y106_BLUT (
.I0(LIOB33_X0Y115_IOB_X0Y115_I),
.I1(RIOB33_X105Y103_IOB_X1Y103_I),
.I2(CLBLM_R_X3Y103_SLICE_X3Y103_BO6),
.I3(RIOB33_X105Y101_IOB_X1Y102_I),
.I4(LIOB33_X0Y113_IOB_X0Y113_I),
.I5(CLBLM_R_X3Y106_SLICE_X3Y106_AO5),
.O5(CLBLM_R_X3Y106_SLICE_X3Y106_BO5),
.O6(CLBLM_R_X3Y106_SLICE_X3Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5f5f5f5f3cc3cc33)
  ) CLBLM_R_X3Y106_SLICE_X3Y106_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y106_I),
.I1(CLBLL_L_X2Y103_SLICE_X1Y103_BO6),
.I2(LIOB33_X0Y111_IOB_X0Y112_I),
.I3(CLBLM_R_X3Y103_SLICE_X2Y103_CO6),
.I4(RIOB33_X105Y103_IOB_X1Y104_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y106_SLICE_X3Y106_AO5),
.O6(CLBLM_R_X3Y106_SLICE_X3Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdffccfddcffccdc)
  ) CLBLM_R_X3Y107_SLICE_X2Y107_DLUT (
.I0(CLBLM_R_X3Y108_SLICE_X2Y108_BO6),
.I1(CLBLM_R_X3Y107_SLICE_X3Y107_CO6),
.I2(CLBLM_R_X3Y108_SLICE_X3Y108_BO6),
.I3(CLBLM_R_X3Y107_SLICE_X2Y107_CO6),
.I4(CLBLM_R_X3Y108_SLICE_X2Y108_CO6),
.I5(CLBLM_R_X3Y107_SLICE_X2Y107_BO6),
.O5(CLBLM_R_X3Y107_SLICE_X2Y107_DO5),
.O6(CLBLM_R_X3Y107_SLICE_X2Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h4ddd8eeecfff0ccc)
  ) CLBLM_R_X3Y107_SLICE_X2Y107_CLUT (
.I0(LIOB33_X0Y113_IOB_X0Y113_I),
.I1(CLBLM_R_X3Y108_SLICE_X3Y108_CO6),
.I2(LIOB33_X0Y103_IOB_X0Y103_I),
.I3(LIOB33_X0Y115_IOB_X0Y115_I),
.I4(CLBLL_L_X4Y108_SLICE_X4Y108_DO6),
.I5(LIOB33_X0Y113_IOB_X0Y114_I),
.O5(CLBLM_R_X3Y107_SLICE_X2Y107_CO5),
.O6(CLBLM_R_X3Y107_SLICE_X2Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6a959595956a6a6a)
  ) CLBLM_R_X3Y107_SLICE_X2Y107_BLUT (
.I0(CLBLL_L_X4Y108_SLICE_X4Y108_DO6),
.I1(LIOB33_X0Y113_IOB_X0Y114_I),
.I2(LIOB33_X0Y113_IOB_X0Y113_I),
.I3(LIOB33_X0Y115_IOB_X0Y115_I),
.I4(LIOB33_X0Y103_IOB_X0Y103_I),
.I5(CLBLM_R_X3Y108_SLICE_X3Y108_CO6),
.O5(CLBLM_R_X3Y107_SLICE_X2Y107_BO5),
.O6(CLBLM_R_X3Y107_SLICE_X2Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h4bd2b42d66996699)
  ) CLBLM_R_X3Y107_SLICE_X2Y107_ALUT (
.I0(CLBLM_R_X3Y108_SLICE_X3Y108_BO6),
.I1(CLBLM_R_X3Y108_SLICE_X2Y108_BO6),
.I2(CLBLM_R_X3Y108_SLICE_X2Y108_CO6),
.I3(CLBLM_R_X3Y107_SLICE_X2Y107_BO6),
.I4(CLBLM_R_X3Y107_SLICE_X2Y107_CO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y107_SLICE_X2Y107_AO5),
.O6(CLBLM_R_X3Y107_SLICE_X2Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y107_SLICE_X3Y107_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y107_SLICE_X3Y107_DO5),
.O6(CLBLM_R_X3Y107_SLICE_X3Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6999966666699996)
  ) CLBLM_R_X3Y107_SLICE_X3Y107_CLUT (
.I0(CLBLM_R_X3Y105_SLICE_X3Y105_BO6),
.I1(CLBLL_L_X4Y105_SLICE_X4Y105_DO6),
.I2(CLBLL_L_X4Y107_SLICE_X4Y107_CO6),
.I3(CLBLM_R_X3Y107_SLICE_X3Y107_AO5),
.I4(CLBLM_R_X3Y106_SLICE_X2Y106_AO5),
.I5(CLBLM_R_X3Y105_SLICE_X3Y105_CO6),
.O5(CLBLM_R_X3Y107_SLICE_X3Y107_CO5),
.O6(CLBLM_R_X3Y107_SLICE_X3Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6066909900600090)
  ) CLBLM_R_X3Y107_SLICE_X3Y107_BLUT (
.I0(CLBLM_R_X3Y106_SLICE_X2Y106_AO5),
.I1(CLBLL_L_X4Y105_SLICE_X4Y105_DO6),
.I2(CLBLL_L_X4Y107_SLICE_X4Y107_CO6),
.I3(CLBLM_R_X3Y105_SLICE_X3Y105_CO6),
.I4(CLBLM_R_X3Y105_SLICE_X3Y105_BO6),
.I5(CLBLM_R_X3Y107_SLICE_X3Y107_AO5),
.O5(CLBLM_R_X3Y107_SLICE_X3Y107_BO5),
.O6(CLBLM_R_X3Y107_SLICE_X3Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5f5f5f5f55ff55ff)
  ) CLBLM_R_X3Y107_SLICE_X3Y107_ALUT (
.I0(LIOB33_X0Y115_IOB_X0Y115_I),
.I1(1'b1),
.I2(LIOB33_X0Y103_IOB_X0Y103_I),
.I3(LIOB33_X0Y113_IOB_X0Y114_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y107_SLICE_X3Y107_AO5),
.O6(CLBLM_R_X3Y107_SLICE_X3Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h4dff04df04df004d)
  ) CLBLM_R_X3Y108_SLICE_X2Y108_DLUT (
.I0(CLBLM_R_X3Y108_SLICE_X2Y108_AO6),
.I1(CLBLM_R_X3Y108_SLICE_X3Y108_CO6),
.I2(CLBLM_R_X3Y108_SLICE_X3Y108_BO6),
.I3(CLBLM_R_X3Y108_SLICE_X2Y108_CO6),
.I4(CLBLM_R_X3Y107_SLICE_X3Y107_AO6),
.I5(CLBLM_R_X3Y108_SLICE_X2Y108_BO6),
.O5(CLBLM_R_X3Y108_SLICE_X2Y108_DO5),
.O6(CLBLM_R_X3Y108_SLICE_X2Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6a95956ac03f3fc0)
  ) CLBLM_R_X3Y108_SLICE_X2Y108_CLUT (
.I0(LIOB33_X0Y113_IOB_X0Y113_I),
.I1(LIOB33_X0Y113_IOB_X0Y114_I),
.I2(LIOB33_X0Y115_IOB_X0Y115_I),
.I3(CLBLL_L_X4Y107_SLICE_X4Y107_CO6),
.I4(CLBLM_R_X3Y105_SLICE_X3Y105_AO6),
.I5(LIOB33_X0Y115_IOB_X0Y116_I),
.O5(CLBLM_R_X3Y108_SLICE_X2Y108_CO5),
.O6(CLBLM_R_X3Y108_SLICE_X2Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h2bbb8eee8eee8eee)
  ) CLBLM_R_X3Y108_SLICE_X2Y108_BLUT (
.I0(CLBLL_L_X4Y109_SLICE_X5Y109_DO6),
.I1(CLBLM_R_X3Y108_SLICE_X3Y108_DO6),
.I2(RIOB33_X105Y105_IOB_X1Y106_I),
.I3(LIOB33_X0Y115_IOB_X0Y115_I),
.I4(LIOB33_X0Y113_IOB_X0Y113_I),
.I5(LIOB33_X0Y103_IOB_X0Y103_I),
.O5(CLBLM_R_X3Y108_SLICE_X2Y108_BO5),
.O6(CLBLM_R_X3Y108_SLICE_X2Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha5a555553333ffff)
  ) CLBLM_R_X3Y108_SLICE_X2Y108_ALUT (
.I0(CLBLL_L_X4Y108_SLICE_X4Y108_DO6),
.I1(LIOB33_X0Y101_IOB_X0Y101_I),
.I2(LIOB33_X0Y113_IOB_X0Y113_I),
.I3(1'b1),
.I4(LIOB33_X0Y113_IOB_X0Y114_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y108_SLICE_X2Y108_AO5),
.O6(CLBLM_R_X3Y108_SLICE_X2Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h9f605fa0a05f9f60)
  ) CLBLM_R_X3Y108_SLICE_X3Y108_DLUT (
.I0(LIOB33_X0Y113_IOB_X0Y114_I),
.I1(LIOB33_X0Y103_IOB_X0Y103_I),
.I2(LIOB33_X0Y111_IOB_X0Y112_I),
.I3(CLBLM_R_X5Y108_SLICE_X6Y108_CO6),
.I4(CLBLL_L_X4Y108_SLICE_X5Y108_CO6),
.I5(CLBLL_L_X4Y108_SLICE_X4Y108_CO6),
.O5(CLBLM_R_X3Y108_SLICE_X3Y108_DO5),
.O6(CLBLM_R_X3Y108_SLICE_X3Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h04cc45ff5dffdfff)
  ) CLBLM_R_X3Y108_SLICE_X3Y108_CLUT (
.I0(LIOB33_X0Y113_IOB_X0Y113_I),
.I1(CLBLL_L_X4Y108_SLICE_X4Y108_CO6),
.I2(LIOB33_X0Y111_IOB_X0Y112_I),
.I3(LIOB33_X0Y103_IOB_X0Y103_I),
.I4(CLBLL_L_X4Y108_SLICE_X5Y108_CO6),
.I5(CLBLM_R_X5Y108_SLICE_X7Y108_DO6),
.O5(CLBLM_R_X3Y108_SLICE_X3Y108_CO5),
.O6(CLBLM_R_X3Y108_SLICE_X3Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h936c6c93c93636c9)
  ) CLBLM_R_X3Y108_SLICE_X3Y108_BLUT (
.I0(CLBLM_R_X3Y110_SLICE_X2Y110_DO6),
.I1(CLBLL_L_X2Y108_SLICE_X0Y108_AO6),
.I2(CLBLM_R_X3Y104_SLICE_X3Y104_AO6),
.I3(CLBLL_L_X4Y109_SLICE_X5Y109_DO6),
.I4(CLBLM_R_X3Y108_SLICE_X3Y108_AO6),
.I5(CLBLL_L_X4Y108_SLICE_X5Y108_DO6),
.O5(CLBLM_R_X3Y108_SLICE_X3Y108_BO5),
.O6(CLBLM_R_X3Y108_SLICE_X3Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hb42d4bd2dddd2222)
  ) CLBLM_R_X3Y108_SLICE_X3Y108_ALUT (
.I0(CLBLL_L_X4Y108_SLICE_X5Y108_CO6),
.I1(CLBLL_L_X4Y108_SLICE_X4Y108_CO6),
.I2(LIOB33_X0Y113_IOB_X0Y113_I),
.I3(LIOB33_X0Y111_IOB_X0Y112_I),
.I4(CLBLM_R_X5Y108_SLICE_X7Y108_DO6),
.I5(LIOB33_X0Y103_IOB_X0Y103_I),
.O5(CLBLM_R_X3Y108_SLICE_X3Y108_AO5),
.O6(CLBLM_R_X3Y108_SLICE_X3Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y109_SLICE_X2Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y109_SLICE_X2Y109_DO5),
.O6(CLBLM_R_X3Y109_SLICE_X2Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y109_SLICE_X2Y109_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y109_SLICE_X2Y109_CO5),
.O6(CLBLM_R_X3Y109_SLICE_X2Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y109_SLICE_X2Y109_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y109_SLICE_X2Y109_BO5),
.O6(CLBLM_R_X3Y109_SLICE_X2Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fffd5ff153f40c0)
  ) CLBLM_R_X3Y109_SLICE_X2Y109_ALUT (
.I0(LIOB33_X0Y113_IOB_X0Y114_I),
.I1(LIOB33_X0Y115_IOB_X0Y116_I),
.I2(LIOB33_X0Y113_IOB_X0Y113_I),
.I3(LIOB33_X0Y115_IOB_X0Y115_I),
.I4(CLBLM_R_X3Y105_SLICE_X3Y105_AO6),
.I5(CLBLL_L_X4Y107_SLICE_X4Y107_CO6),
.O5(CLBLM_R_X3Y109_SLICE_X2Y109_AO5),
.O6(CLBLM_R_X3Y109_SLICE_X2Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y109_SLICE_X3Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y109_SLICE_X3Y109_DO5),
.O6(CLBLM_R_X3Y109_SLICE_X3Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y109_SLICE_X3Y109_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y109_SLICE_X3Y109_CO5),
.O6(CLBLM_R_X3Y109_SLICE_X3Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y109_SLICE_X3Y109_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y109_SLICE_X3Y109_BO5),
.O6(CLBLM_R_X3Y109_SLICE_X3Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y109_SLICE_X3Y109_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y109_SLICE_X3Y109_AO5),
.O6(CLBLM_R_X3Y109_SLICE_X3Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0445ccff5ddfffff)
  ) CLBLM_R_X3Y110_SLICE_X2Y110_DLUT (
.I0(LIOB33_X0Y113_IOB_X0Y113_I),
.I1(CLBLM_R_X3Y110_SLICE_X3Y110_CO6),
.I2(LIOB33_X0Y111_IOB_X0Y112_I),
.I3(CLBLL_L_X4Y109_SLICE_X4Y109_BO6),
.I4(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I5(CLBLL_L_X4Y107_SLICE_X4Y107_BO6),
.O5(CLBLM_R_X3Y110_SLICE_X2Y110_DO5),
.O6(CLBLM_R_X3Y110_SLICE_X2Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h69c3963ca50f5af0)
  ) CLBLM_R_X3Y110_SLICE_X2Y110_CLUT (
.I0(LIOB33_X0Y113_IOB_X0Y113_I),
.I1(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I2(CLBLL_L_X4Y109_SLICE_X4Y109_DO6),
.I3(RIOB33_X105Y105_IOB_X1Y106_I),
.I4(CLBLM_R_X3Y110_SLICE_X2Y110_DO6),
.I5(LIOB33_X0Y115_IOB_X0Y115_I),
.O5(CLBLM_R_X3Y110_SLICE_X2Y110_CO5),
.O6(CLBLM_R_X3Y110_SLICE_X2Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'he6192ad5738cbf40)
  ) CLBLM_R_X3Y110_SLICE_X2Y110_BLUT (
.I0(CLBLM_R_X3Y110_SLICE_X3Y110_CO6),
.I1(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I2(LIOB33_X0Y111_IOB_X0Y112_I),
.I3(CLBLL_L_X4Y107_SLICE_X4Y107_BO6),
.I4(LIOB33_X0Y113_IOB_X0Y113_I),
.I5(CLBLL_L_X4Y109_SLICE_X4Y109_BO6),
.O5(CLBLM_R_X3Y110_SLICE_X2Y110_BO5),
.O6(CLBLM_R_X3Y110_SLICE_X2Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h2bbb2bbb69996999)
  ) CLBLM_R_X3Y110_SLICE_X2Y110_ALUT (
.I0(CLBLM_R_X3Y110_SLICE_X3Y110_CO6),
.I1(CLBLL_L_X4Y109_SLICE_X4Y109_BO6),
.I2(LIOB33_X0Y111_IOB_X0Y112_I),
.I3(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y110_SLICE_X2Y110_AO5),
.O6(CLBLM_R_X3Y110_SLICE_X2Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000965a965a965a)
  ) CLBLM_R_X3Y110_SLICE_X3Y110_DLUT (
.I0(CLBLL_L_X4Y111_SLICE_X4Y111_AO6),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(CLBLM_R_X3Y111_SLICE_X2Y111_CO6),
.I3(LIOB33_X0Y107_IOB_X0Y107_I),
.I4(LIOB33_X0Y107_IOB_X0Y108_I),
.I5(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.O5(CLBLM_R_X3Y110_SLICE_X3Y110_DO5),
.O6(CLBLM_R_X3Y110_SLICE_X3Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fdf134cdfdf4c4c)
  ) CLBLM_R_X3Y110_SLICE_X3Y110_CLUT (
.I0(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I1(CLBLL_L_X4Y109_SLICE_X4Y109_AO6),
.I2(LIOB33_X0Y111_IOB_X0Y111_I),
.I3(RIOB33_X105Y105_IOB_X1Y106_I),
.I4(CLBLL_L_X4Y110_SLICE_X4Y110_CO6),
.I5(LIOB33_X0Y109_IOB_X0Y110_I),
.O5(CLBLM_R_X3Y110_SLICE_X3Y110_CO5),
.O6(CLBLM_R_X3Y110_SLICE_X3Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996c33ca55a0ff0)
  ) CLBLM_R_X3Y110_SLICE_X3Y110_BLUT (
.I0(LIOB33_X0Y111_IOB_X0Y111_I),
.I1(LIOB33_X0Y109_IOB_X0Y110_I),
.I2(CLBLL_L_X4Y109_SLICE_X4Y109_AO6),
.I3(CLBLL_L_X4Y110_SLICE_X4Y110_CO6),
.I4(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I5(RIOB33_X105Y105_IOB_X1Y106_I),
.O5(CLBLM_R_X3Y110_SLICE_X3Y110_BO5),
.O6(CLBLM_R_X3Y110_SLICE_X3Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h7f15bf2aff3f3f00)
  ) CLBLM_R_X3Y110_SLICE_X3Y110_ALUT (
.I0(LIOB33_X0Y107_IOB_X0Y107_I),
.I1(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I2(LIOB33_X0Y107_IOB_X0Y108_I),
.I3(CLBLM_R_X3Y111_SLICE_X2Y111_CO6),
.I4(CLBLL_L_X4Y111_SLICE_X4Y111_AO6),
.I5(RIOB33_X105Y105_IOB_X1Y106_I),
.O5(CLBLM_R_X3Y110_SLICE_X3Y110_AO5),
.O6(CLBLM_R_X3Y110_SLICE_X3Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y111_SLICE_X2Y111_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y111_SLICE_X2Y111_DO5),
.O6(CLBLM_R_X3Y111_SLICE_X2Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h71d4f3fcf550fff0)
  ) CLBLM_R_X3Y111_SLICE_X2Y111_CLUT (
.I0(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(CLBLM_R_X3Y112_SLICE_X2Y112_DO6),
.I3(CLBLL_L_X4Y112_SLICE_X4Y112_BO6),
.I4(LIOB33_X0Y107_IOB_X0Y107_I),
.I5(LIOB33_X0Y105_IOB_X0Y106_I),
.O5(CLBLM_R_X3Y111_SLICE_X2Y111_CO5),
.O6(CLBLM_R_X3Y111_SLICE_X2Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h69c39933963c66cc)
  ) CLBLM_R_X3Y111_SLICE_X2Y111_BLUT (
.I0(LIOB33_X0Y107_IOB_X0Y107_I),
.I1(CLBLL_L_X4Y111_SLICE_X4Y111_AO6),
.I2(LIOB33_X0Y107_IOB_X0Y108_I),
.I3(RIOB33_X105Y105_IOB_X1Y106_I),
.I4(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I5(CLBLM_R_X3Y111_SLICE_X2Y111_CO6),
.O5(CLBLM_R_X3Y111_SLICE_X2Y111_BO5),
.O6(CLBLM_R_X3Y111_SLICE_X2Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h353a45ba48484848)
  ) CLBLM_R_X3Y111_SLICE_X2Y111_ALUT (
.I0(LIOB33_X0Y113_IOB_X0Y114_I),
.I1(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I2(LIOB33_X0Y115_IOB_X0Y116_I),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(RIOB33_X105Y111_IOB_X1Y112_I),
.I5(RIOB33_X105Y113_IOB_X1Y113_I),
.O5(CLBLM_R_X3Y111_SLICE_X2Y111_AO5),
.O6(CLBLM_R_X3Y111_SLICE_X2Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h07000a0a8daa0000)
  ) CLBLM_R_X3Y111_SLICE_X3Y111_DLUT (
.I0(LIOB33_X0Y115_IOB_X0Y116_I),
.I1(RIOB33_X105Y111_IOB_X1Y112_I),
.I2(LIOB33_X0Y113_IOB_X0Y114_I),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(RIOB33_X105Y113_IOB_X1Y113_I),
.I5(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.O5(CLBLM_R_X3Y111_SLICE_X3Y111_DO5),
.O6(CLBLM_R_X3Y111_SLICE_X3Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h33ff33ff00ffffff)
  ) CLBLM_R_X3Y111_SLICE_X3Y111_CLUT (
.I0(1'b1),
.I1(LIOB33_X0Y103_IOB_X0Y103_I),
.I2(1'b1),
.I3(LIOB33_X0Y105_IOB_X0Y106_I),
.I4(RIOB33_X105Y105_IOB_X1Y106_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y111_SLICE_X3Y111_CO5),
.O6(CLBLM_R_X3Y111_SLICE_X3Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h55ff55ff33ff33ff)
  ) CLBLM_R_X3Y111_SLICE_X3Y111_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y106_I),
.I1(LIOB33_X0Y103_IOB_X0Y103_I),
.I2(1'b1),
.I3(LIOB33_X0Y105_IOB_X0Y105_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y111_SLICE_X3Y111_BO5),
.O6(CLBLM_R_X3Y111_SLICE_X3Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha05fa05f77777777)
  ) CLBLM_R_X3Y111_SLICE_X3Y111_ALUT (
.I0(LIOB33_X0Y107_IOB_X0Y107_I),
.I1(LIOB33_X0Y103_IOB_X0Y103_I),
.I2(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I3(CLBLM_R_X3Y112_SLICE_X3Y112_CO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y111_SLICE_X3Y111_AO5),
.O6(CLBLM_R_X3Y111_SLICE_X3Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdd0f440df0d4f04)
  ) CLBLM_R_X3Y112_SLICE_X2Y112_DLUT (
.I0(CLBLM_R_X3Y112_SLICE_X2Y112_CO6),
.I1(CLBLM_R_X5Y101_SLICE_X7Y101_AO5),
.I2(CLBLM_R_X3Y112_SLICE_X3Y112_BO6),
.I3(CLBLM_R_X3Y112_SLICE_X2Y112_AO5),
.I4(CLBLL_L_X2Y113_SLICE_X1Y113_DO6),
.I5(CLBLM_R_X3Y111_SLICE_X3Y111_BO6),
.O5(CLBLM_R_X3Y112_SLICE_X2Y112_DO5),
.O6(CLBLM_R_X3Y112_SLICE_X2Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h69a5c30f965a3cf0)
  ) CLBLM_R_X3Y112_SLICE_X2Y112_CLUT (
.I0(LIOB33_X0Y103_IOB_X0Y103_I),
.I1(LIOB33_X0Y103_IOB_X0Y104_I),
.I2(CLBLM_R_X3Y113_SLICE_X2Y113_DO6),
.I3(RIOB33_X105Y105_IOB_X1Y106_I),
.I4(LIOB33_X0Y101_IOB_X0Y102_I),
.I5(CLBLM_R_X3Y113_SLICE_X3Y113_BO6),
.O5(CLBLM_R_X3Y112_SLICE_X2Y112_CO5),
.O6(CLBLM_R_X3Y112_SLICE_X2Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc6399999639ccccc)
  ) CLBLM_R_X3Y112_SLICE_X2Y112_BLUT (
.I0(CLBLL_L_X2Y113_SLICE_X1Y113_DO6),
.I1(CLBLM_R_X3Y112_SLICE_X3Y112_BO6),
.I2(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I3(RIOB33_X105Y105_IOB_X1Y106_I),
.I4(LIOB33_X0Y105_IOB_X0Y105_I),
.I5(CLBLM_R_X3Y112_SLICE_X2Y112_CO6),
.O5(CLBLM_R_X3Y112_SLICE_X2Y112_BO5),
.O6(CLBLM_R_X3Y112_SLICE_X2Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc3300ff3333ffff)
  ) CLBLM_R_X3Y112_SLICE_X2Y112_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y105_IOB_X0Y106_I),
.I2(1'b1),
.I3(CLBLM_R_X3Y112_SLICE_X2Y112_BO6),
.I4(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y112_SLICE_X2Y112_AO5),
.O6(CLBLM_R_X3Y112_SLICE_X2Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fffb3ff135f20a0)
  ) CLBLM_R_X3Y112_SLICE_X3Y112_DLUT (
.I0(LIOB33_X0Y101_IOB_X0Y102_I),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(LIOB33_X0Y103_IOB_X0Y103_I),
.I3(LIOB33_X0Y103_IOB_X0Y104_I),
.I4(CLBLM_R_X3Y113_SLICE_X2Y113_DO6),
.I5(CLBLM_R_X3Y113_SLICE_X3Y113_BO6),
.O5(CLBLM_R_X3Y112_SLICE_X3Y112_DO5),
.O6(CLBLM_R_X3Y112_SLICE_X3Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h956aaaaaa9566666)
  ) CLBLM_R_X3Y112_SLICE_X3Y112_CLUT (
.I0(CLBLL_L_X4Y112_SLICE_X4Y112_BO6),
.I1(CLBLL_L_X4Y112_SLICE_X4Y112_CO6),
.I2(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I3(RIOB33_X105Y105_IOB_X1Y106_I),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(CLBLL_L_X2Y112_SLICE_X1Y112_AO6),
.O5(CLBLM_R_X3Y112_SLICE_X3Y112_CO5),
.O6(CLBLM_R_X3Y112_SLICE_X3Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h2db4d24bd24b2db4)
  ) CLBLM_R_X3Y112_SLICE_X3Y112_BLUT (
.I0(CLBLM_R_X3Y113_SLICE_X3Y113_DO6),
.I1(CLBLM_R_X3Y113_SLICE_X3Y113_BO6),
.I2(CLBLL_L_X4Y112_SLICE_X4Y112_AO6),
.I3(CLBLL_L_X2Y113_SLICE_X1Y113_AO5),
.I4(CLBLM_R_X5Y111_SLICE_X6Y111_AO6),
.I5(CLBLM_R_X3Y113_SLICE_X3Y113_CO6),
.O5(CLBLM_R_X3Y112_SLICE_X3Y112_BO5),
.O6(CLBLM_R_X3Y112_SLICE_X3Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0fff0fff33ff33ff)
  ) CLBLM_R_X3Y112_SLICE_X3Y112_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(LIOB33_X0Y103_IOB_X0Y103_I),
.I3(LIOB33_X0Y101_IOB_X0Y102_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y112_SLICE_X3Y112_AO5),
.O6(CLBLM_R_X3Y112_SLICE_X3Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3cc33c96cc33cccc)
  ) CLBLM_R_X3Y113_SLICE_X2Y113_DLUT (
.I0(LIOB33_X0Y103_IOB_X0Y103_I),
.I1(CLBLM_R_X3Y111_SLICE_X2Y111_AO6),
.I2(LIOB33_X0Y113_IOB_X0Y114_I),
.I3(CLBLL_L_X4Y113_SLICE_X4Y113_AO6),
.I4(CLBLM_R_X3Y114_SLICE_X2Y114_CO6),
.I5(LIOB33_X0Y101_IOB_X0Y101_I),
.O5(CLBLM_R_X3Y113_SLICE_X2Y113_DO5),
.O6(CLBLM_R_X3Y113_SLICE_X2Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h9fa0605f5f9fa060)
  ) CLBLM_R_X3Y113_SLICE_X2Y113_CLUT (
.I0(LIOB33_X0Y103_IOB_X0Y103_I),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(LIOB33_X0Y101_IOB_X0Y102_I),
.I3(CLBLM_R_X3Y113_SLICE_X2Y113_AO5),
.I4(CLBLM_R_X3Y113_SLICE_X2Y113_DO6),
.I5(CLBLM_R_X3Y113_SLICE_X2Y113_BO6),
.O5(CLBLM_R_X3Y113_SLICE_X2Y113_CO5),
.O6(CLBLM_R_X3Y113_SLICE_X2Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha555a555cdddcddd)
  ) CLBLM_R_X3Y113_SLICE_X2Y113_BLUT (
.I0(CLBLM_R_X3Y114_SLICE_X2Y114_CO6),
.I1(CLBLL_L_X4Y113_SLICE_X4Y113_AO6),
.I2(LIOB33_X0Y103_IOB_X0Y103_I),
.I3(LIOB33_X0Y101_IOB_X0Y101_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y113_SLICE_X2Y113_BO5),
.O6(CLBLM_R_X3Y113_SLICE_X2Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc30fc30fabafabaf)
  ) CLBLM_R_X3Y113_SLICE_X2Y113_ALUT (
.I0(CLBLM_R_X3Y114_SLICE_X2Y114_DO6),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(CLBLM_R_X3Y114_SLICE_X2Y114_AO6),
.I3(LIOB33_X0Y101_IOB_X0Y101_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y113_SLICE_X2Y113_AO5),
.O6(CLBLM_R_X3Y113_SLICE_X2Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3cc3c33c1ee1e11e)
  ) CLBLM_R_X3Y113_SLICE_X3Y113_DLUT (
.I0(CLBLM_R_X3Y113_SLICE_X3Y113_AO6),
.I1(CLBLL_L_X4Y113_SLICE_X4Y113_AO6),
.I2(CLBLM_R_X3Y112_SLICE_X3Y112_AO6),
.I3(CLBLM_R_X3Y108_SLICE_X2Y108_AO5),
.I4(CLBLM_R_X3Y111_SLICE_X2Y111_AO6),
.I5(CLBLM_R_X3Y114_SLICE_X2Y114_CO6),
.O5(CLBLM_R_X3Y113_SLICE_X3Y113_DO5),
.O6(CLBLM_R_X3Y113_SLICE_X3Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcc0c0fcfee0e0fe)
  ) CLBLM_R_X3Y113_SLICE_X3Y113_CLUT (
.I0(CLBLM_R_X3Y113_SLICE_X3Y113_AO6),
.I1(CLBLL_L_X4Y113_SLICE_X4Y113_AO6),
.I2(CLBLM_R_X3Y112_SLICE_X3Y112_AO6),
.I3(CLBLM_R_X3Y108_SLICE_X2Y108_AO5),
.I4(CLBLM_R_X3Y111_SLICE_X2Y111_AO6),
.I5(CLBLM_R_X3Y114_SLICE_X2Y114_CO6),
.O5(CLBLM_R_X3Y113_SLICE_X3Y113_CO5),
.O6(CLBLM_R_X3Y113_SLICE_X3Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaeaeffae0000ae)
  ) CLBLM_R_X3Y113_SLICE_X3Y113_BLUT (
.I0(CLBLM_R_X3Y114_SLICE_X2Y114_DO6),
.I1(CLBLM_R_X3Y113_SLICE_X3Y113_AO5),
.I2(CLBLM_R_X3Y114_SLICE_X2Y114_AO6),
.I3(CLBLM_R_X3Y114_SLICE_X2Y114_CO6),
.I4(CLBLM_R_X3Y113_SLICE_X3Y113_AO6),
.I5(CLBLM_R_X3Y112_SLICE_X3Y112_AO5),
.O5(CLBLM_R_X3Y113_SLICE_X3Y113_BO5),
.O6(CLBLM_R_X3Y113_SLICE_X3Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f3f3f3f3333ffff)
  ) CLBLM_R_X3Y113_SLICE_X3Y113_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y101_IOB_X0Y101_I),
.I2(LIOB33_X0Y103_IOB_X0Y103_I),
.I3(1'b1),
.I4(RIOB33_X105Y105_IOB_X1Y106_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y113_SLICE_X3Y113_AO5),
.O6(CLBLM_R_X3Y113_SLICE_X3Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3455330044004400)
  ) CLBLM_R_X3Y114_SLICE_X2Y114_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y106_I),
.I1(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I2(RIOB33_X105Y111_IOB_X1Y112_I),
.I3(LIOB33_X0Y103_IOB_X0Y103_I),
.I4(LIOB33_X0Y113_IOB_X0Y114_I),
.I5(RIOB33_X105Y113_IOB_X1Y113_I),
.O5(CLBLM_R_X3Y114_SLICE_X2Y114_DO5),
.O6(CLBLM_R_X3Y114_SLICE_X2Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h353955aa00cccc00)
  ) CLBLM_R_X3Y114_SLICE_X2Y114_CLUT (
.I0(LIOB33_X0Y115_IOB_X0Y116_I),
.I1(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I2(RIOB33_X105Y111_IOB_X1Y112_I),
.I3(LIOB33_X0Y103_IOB_X0Y103_I),
.I4(LIOB33_X0Y113_IOB_X0Y114_I),
.I5(RIOB33_X105Y113_IOB_X1Y113_I),
.O5(CLBLM_R_X3Y114_SLICE_X2Y114_CO5),
.O6(CLBLM_R_X3Y114_SLICE_X2Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6a6a7b3f959584c0)
  ) CLBLM_R_X3Y114_SLICE_X2Y114_BLUT (
.I0(CLBLM_R_X3Y114_SLICE_X2Y114_DO6),
.I1(LIOB33_X0Y101_IOB_X0Y101_I),
.I2(LIOB33_X0Y103_IOB_X0Y103_I),
.I3(RIOB33_X105Y105_IOB_X1Y106_I),
.I4(CLBLM_R_X3Y114_SLICE_X2Y114_AO6),
.I5(CLBLM_R_X3Y114_SLICE_X2Y114_CO6),
.O5(CLBLM_R_X3Y114_SLICE_X2Y114_BO5),
.O6(CLBLM_R_X3Y114_SLICE_X2Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h1d552ea63030c0c0)
  ) CLBLM_R_X3Y114_SLICE_X2Y114_ALUT (
.I0(LIOB33_X0Y113_IOB_X0Y114_I),
.I1(LIOB33_X0Y103_IOB_X0Y103_I),
.I2(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I3(RIOB33_X105Y111_IOB_X1Y112_I),
.I4(RIOB33_X105Y105_IOB_X1Y106_I),
.I5(RIOB33_X105Y113_IOB_X1Y113_I),
.O5(CLBLM_R_X3Y114_SLICE_X2Y114_AO5),
.O6(CLBLM_R_X3Y114_SLICE_X2Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y114_SLICE_X3Y114_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y114_SLICE_X3Y114_DO5),
.O6(CLBLM_R_X3Y114_SLICE_X3Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y114_SLICE_X3Y114_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y114_SLICE_X3Y114_CO5),
.O6(CLBLM_R_X3Y114_SLICE_X3Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y114_SLICE_X3Y114_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y114_SLICE_X3Y114_BO5),
.O6(CLBLM_R_X3Y114_SLICE_X3Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y114_SLICE_X3Y114_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y114_SLICE_X3Y114_AO5),
.O6(CLBLM_R_X3Y114_SLICE_X3Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hb50faf0f5fffffff)
  ) CLBLM_R_X5Y100_SLICE_X6Y100_DLUT (
.I0(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I1(RIOB33_X105Y111_IOB_X1Y112_I),
.I2(LIOB33_X0Y101_IOB_X0Y101_I),
.I3(RIOB33_X105Y109_IOB_X1Y110_I),
.I4(RIOB33_X105Y113_IOB_X1Y113_I),
.I5(RIOB33_X105Y111_IOB_X1Y111_I),
.O5(CLBLM_R_X5Y100_SLICE_X6Y100_DO5),
.O6(CLBLM_R_X5Y100_SLICE_X6Y100_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996a55a996655aa)
  ) CLBLM_R_X5Y100_SLICE_X6Y100_CLUT (
.I0(CLBLM_R_X5Y101_SLICE_X7Y101_AO6),
.I1(RIOB33_X105Y109_IOB_X1Y110_I),
.I2(RIOB33_X105Y109_IOB_X1Y109_I),
.I3(CLBLL_L_X4Y100_SLICE_X5Y100_DO6),
.I4(LIOB33_X0Y105_IOB_X0Y105_I),
.I5(LIOB33_X0Y105_IOB_X0Y106_I),
.O5(CLBLM_R_X5Y100_SLICE_X6Y100_CO5),
.O6(CLBLM_R_X5Y100_SLICE_X6Y100_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h57137f137f577f7f)
  ) CLBLM_R_X5Y100_SLICE_X6Y100_BLUT (
.I0(RIOB33_X105Y107_IOB_X1Y108_I),
.I1(CLBLL_L_X4Y100_SLICE_X5Y100_CO6),
.I2(LIOB33_X0Y107_IOB_X0Y108_I),
.I3(CLBLM_R_X5Y102_SLICE_X7Y102_AO6),
.I4(LIOB33_X0Y107_IOB_X0Y107_I),
.I5(CLBLM_R_X5Y100_SLICE_X6Y100_CO6),
.O5(CLBLM_R_X5Y100_SLICE_X6Y100_BO5),
.O6(CLBLM_R_X5Y100_SLICE_X6Y100_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0000fff95959595)
  ) CLBLM_R_X5Y100_SLICE_X6Y100_ALUT (
.I0(CLBLM_R_X5Y100_SLICE_X6Y100_DO6),
.I1(LIOB33_X0Y101_IOB_X0Y102_I),
.I2(RIOB33_X105Y109_IOB_X1Y110_I),
.I3(LIOB33_X0Y105_IOB_X0Y105_I),
.I4(CLBLL_L_X4Y100_SLICE_X5Y100_DO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y100_SLICE_X6Y100_AO5),
.O6(CLBLM_R_X5Y100_SLICE_X6Y100_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y100_SLICE_X7Y100_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y100_SLICE_X7Y100_DO5),
.O6(CLBLM_R_X5Y100_SLICE_X7Y100_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y100_SLICE_X7Y100_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y100_SLICE_X7Y100_CO5),
.O6(CLBLM_R_X5Y100_SLICE_X7Y100_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y100_SLICE_X7Y100_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y100_SLICE_X7Y100_BO5),
.O6(CLBLM_R_X5Y100_SLICE_X7Y100_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y100_SLICE_X7Y100_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y100_SLICE_X7Y100_AO5),
.O6(CLBLM_R_X5Y100_SLICE_X7Y100_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h317375f77177f5ff)
  ) CLBLM_R_X5Y101_SLICE_X6Y101_DLUT (
.I0(CLBLM_R_X5Y101_SLICE_X6Y101_CO6),
.I1(RIOB33_X105Y107_IOB_X1Y107_I),
.I2(CLBLM_R_X7Y102_SLICE_X8Y102_BO6),
.I3(CLBLM_R_X5Y101_SLICE_X6Y101_AO5),
.I4(LIOB33_X0Y109_IOB_X0Y109_I),
.I5(LIOB33_X0Y107_IOB_X0Y108_I),
.O5(CLBLM_R_X5Y101_SLICE_X6Y101_DO5),
.O6(CLBLM_R_X5Y101_SLICE_X6Y101_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hd42bbbbb2bd44444)
  ) CLBLM_R_X5Y101_SLICE_X6Y101_CLUT (
.I0(CLBLM_R_X5Y102_SLICE_X7Y102_AO6),
.I1(CLBLM_R_X5Y100_SLICE_X6Y100_CO6),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(LIOB33_X0Y107_IOB_X0Y108_I),
.I4(RIOB33_X105Y107_IOB_X1Y108_I),
.I5(CLBLL_L_X4Y100_SLICE_X5Y100_CO6),
.O5(CLBLM_R_X5Y101_SLICE_X6Y101_CO5),
.O6(CLBLM_R_X5Y101_SLICE_X6Y101_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hca6a35956f3f90c0)
  ) CLBLM_R_X5Y101_SLICE_X6Y101_BLUT (
.I0(CLBLM_R_X7Y102_SLICE_X8Y102_BO6),
.I1(LIOB33_X0Y109_IOB_X0Y109_I),
.I2(RIOB33_X105Y107_IOB_X1Y107_I),
.I3(LIOB33_X0Y107_IOB_X0Y108_I),
.I4(CLBLM_R_X5Y101_SLICE_X6Y101_CO6),
.I5(CLBLM_R_X5Y101_SLICE_X6Y101_AO5),
.O5(CLBLM_R_X5Y101_SLICE_X6Y101_BO5),
.O6(CLBLM_R_X5Y101_SLICE_X6Y101_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h965a69a53cf0c30f)
  ) CLBLM_R_X5Y101_SLICE_X6Y101_ALUT (
.I0(CLBLM_R_X7Y102_SLICE_X8Y102_BO6),
.I1(RIOB33_X105Y107_IOB_X1Y108_I),
.I2(CLBLM_R_X5Y100_SLICE_X6Y100_CO6),
.I3(LIOB33_X0Y107_IOB_X0Y107_I),
.I4(CLBLM_R_X5Y102_SLICE_X7Y102_AO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y101_SLICE_X6Y101_AO5),
.O6(CLBLM_R_X5Y101_SLICE_X6Y101_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h48c0defcdefcdefc)
  ) CLBLM_R_X5Y101_SLICE_X7Y101_DLUT (
.I0(RIOB33_X105Y109_IOB_X1Y110_I),
.I1(CLBLM_L_X8Y101_SLICE_X11Y101_BO6),
.I2(CLBLM_R_X5Y100_SLICE_X6Y100_DO6),
.I3(LIOB33_X0Y101_IOB_X0Y102_I),
.I4(LIOB33_X0Y103_IOB_X0Y104_I),
.I5(RIOB33_X105Y109_IOB_X1Y109_I),
.O5(CLBLM_R_X5Y101_SLICE_X7Y101_DO5),
.O6(CLBLM_R_X5Y101_SLICE_X7Y101_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'he482a06c6cc6a0a0)
  ) CLBLM_R_X5Y101_SLICE_X7Y101_CLUT (
.I0(RIOB33_X105Y109_IOB_X1Y110_I),
.I1(RIOB33_X105Y111_IOB_X1Y111_I),
.I2(LIOB33_X0Y103_IOB_X0Y104_I),
.I3(CLBLM_R_X5Y103_SLICE_X6Y103_CO6),
.I4(LIOB33_X0Y101_IOB_X0Y102_I),
.I5(LIOB33_X0Y101_IOB_X0Y101_I),
.O5(CLBLM_R_X5Y101_SLICE_X7Y101_CO5),
.O6(CLBLM_R_X5Y101_SLICE_X7Y101_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h963cccccc39633cc)
  ) CLBLM_R_X5Y101_SLICE_X7Y101_BLUT (
.I0(LIOB33_X0Y103_IOB_X0Y104_I),
.I1(CLBLM_R_X5Y101_SLICE_X7Y101_CO6),
.I2(LIOB33_X0Y105_IOB_X0Y105_I),
.I3(CLBLM_R_X5Y100_SLICE_X6Y100_AO5),
.I4(RIOB33_X105Y109_IOB_X1Y109_I),
.I5(CLBLM_L_X8Y101_SLICE_X11Y101_BO6),
.O5(CLBLM_R_X5Y101_SLICE_X7Y101_BO5),
.O6(CLBLM_R_X5Y101_SLICE_X7Y101_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h2bbb2bbb0f0fffff)
  ) CLBLM_R_X5Y101_SLICE_X7Y101_ALUT (
.I0(CLBLM_R_X5Y101_SLICE_X7Y101_DO6),
.I1(CLBLM_R_X5Y101_SLICE_X7Y101_CO6),
.I2(LIOB33_X0Y105_IOB_X0Y105_I),
.I3(RIOB33_X105Y109_IOB_X1Y109_I),
.I4(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y101_SLICE_X7Y101_AO5),
.O6(CLBLM_R_X5Y101_SLICE_X7Y101_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996996696966666)
  ) CLBLM_R_X5Y102_SLICE_X6Y102_DLUT (
.I0(CLBLM_R_X5Y101_SLICE_X6Y101_AO6),
.I1(CLBLM_R_X7Y103_SLICE_X8Y103_AO6),
.I2(RIOB33_X105Y107_IOB_X1Y107_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(LIOB33_X0Y107_IOB_X0Y108_I),
.I5(LIOB33_X0Y109_IOB_X0Y109_I),
.O5(CLBLM_R_X5Y102_SLICE_X6Y102_DO5),
.O6(CLBLM_R_X5Y102_SLICE_X6Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha9656aa669a566aa)
  ) CLBLM_R_X5Y102_SLICE_X6Y102_CLUT (
.I0(CLBLM_R_X5Y101_SLICE_X6Y101_BO6),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X7Y103_SLICE_X8Y103_AO6),
.I3(LIOB33_X0Y109_IOB_X0Y110_I),
.I4(CLBLM_R_X5Y102_SLICE_X6Y102_BO5),
.I5(LIOB33_X0Y109_IOB_X0Y109_I),
.O5(CLBLM_R_X5Y102_SLICE_X6Y102_CO5),
.O6(CLBLM_R_X5Y102_SLICE_X6Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h33ff33ff87878787)
  ) CLBLM_R_X5Y102_SLICE_X6Y102_BLUT (
.I0(LIOB33_X0Y107_IOB_X0Y108_I),
.I1(RIOB33_X105Y107_IOB_X1Y107_I),
.I2(CLBLM_R_X5Y101_SLICE_X6Y101_AO6),
.I3(LIOB33_X0Y101_IOB_X0Y101_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y102_SLICE_X6Y102_BO5),
.O6(CLBLM_R_X5Y102_SLICE_X6Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333ffff71f571f5)
  ) CLBLM_R_X5Y102_SLICE_X6Y102_ALUT (
.I0(CLBLM_R_X5Y102_SLICE_X6Y102_BO5),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X7Y103_SLICE_X8Y103_AO6),
.I3(LIOB33_X0Y109_IOB_X0Y109_I),
.I4(LIOB33_X0Y101_IOB_X0Y101_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y102_SLICE_X6Y102_AO5),
.O6(CLBLM_R_X5Y102_SLICE_X6Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y102_SLICE_X7Y102_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y102_SLICE_X7Y102_DO5),
.O6(CLBLM_R_X5Y102_SLICE_X7Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y102_SLICE_X7Y102_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y102_SLICE_X7Y102_CO5),
.O6(CLBLM_R_X5Y102_SLICE_X7Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6c93936c93936c6c)
  ) CLBLM_R_X5Y102_SLICE_X7Y102_BLUT (
.I0(LIOB33_X0Y103_IOB_X0Y104_I),
.I1(CLBLM_R_X5Y100_SLICE_X6Y100_DO6),
.I2(RIOB33_X105Y109_IOB_X1Y109_I),
.I3(LIOB33_X0Y101_IOB_X0Y102_I),
.I4(CLBLM_L_X8Y101_SLICE_X11Y101_BO6),
.I5(RIOB33_X105Y109_IOB_X1Y110_I),
.O5(CLBLM_R_X5Y102_SLICE_X7Y102_BO5),
.O6(CLBLM_R_X5Y102_SLICE_X7Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0c0f4cdf4fdfffff)
  ) CLBLM_R_X5Y102_SLICE_X7Y102_ALUT (
.I0(LIOB33_X0Y105_IOB_X0Y105_I),
.I1(CLBLM_R_X7Y101_SLICE_X9Y101_CO6),
.I2(RIOB33_X105Y107_IOB_X1Y108_I),
.I3(CLBLM_R_X5Y102_SLICE_X7Y102_BO6),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(CLBLM_R_X5Y101_SLICE_X7Y101_BO6),
.O5(CLBLM_R_X5Y102_SLICE_X7Y102_AO5),
.O6(CLBLM_R_X5Y102_SLICE_X7Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h1703ff5f3f17ff5f)
  ) CLBLM_R_X5Y103_SLICE_X6Y103_DLUT (
.I0(CLBLM_R_X7Y102_SLICE_X9Y102_DO6),
.I1(LIOB33_X0Y109_IOB_X0Y110_I),
.I2(CLBLM_R_X7Y103_SLICE_X9Y103_CO6),
.I3(CLBLM_R_X7Y104_SLICE_X8Y104_DO6),
.I4(RIOB33_X105Y103_IOB_X1Y103_I),
.I5(LIOB33_X0Y109_IOB_X0Y109_I),
.O5(CLBLM_R_X5Y103_SLICE_X6Y103_DO5),
.O6(CLBLM_R_X5Y103_SLICE_X6Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h337777fff7ffffff)
  ) CLBLM_R_X5Y103_SLICE_X6Y103_CLUT (
.I0(LIOB33_X0Y101_IOB_X0Y101_I),
.I1(RIOB33_X105Y109_IOB_X1Y110_I),
.I2(RIOB33_X105Y111_IOB_X1Y112_I),
.I3(RIOB33_X105Y113_IOB_X1Y113_I),
.I4(RIOB33_X105Y111_IOB_X1Y111_I),
.I5(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.O5(CLBLM_R_X5Y103_SLICE_X6Y103_CO5),
.O6(CLBLM_R_X5Y103_SLICE_X6Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h96a55a96aa55aaaa)
  ) CLBLM_R_X5Y103_SLICE_X6Y103_BLUT (
.I0(CLBLM_R_X7Y103_SLICE_X8Y103_DO6),
.I1(RIOB33_X105Y103_IOB_X1Y103_I),
.I2(RIOB33_X105Y103_IOB_X1Y104_I),
.I3(CLBLM_R_X7Y104_SLICE_X8Y104_DO6),
.I4(CLBLM_R_X7Y102_SLICE_X9Y102_DO6),
.I5(LIOB33_X0Y109_IOB_X0Y109_I),
.O5(CLBLM_R_X5Y103_SLICE_X6Y103_BO5),
.O6(CLBLM_R_X5Y103_SLICE_X6Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fdfff5f134c5f00)
  ) CLBLM_R_X5Y103_SLICE_X6Y103_ALUT (
.I0(LIOB33_X0Y111_IOB_X0Y111_I),
.I1(RIOB33_X105Y103_IOB_X1Y103_I),
.I2(RIOB33_X105Y101_IOB_X1Y102_I),
.I3(CLBLM_R_X5Y103_SLICE_X6Y103_BO6),
.I4(LIOB33_X0Y109_IOB_X0Y110_I),
.I5(CLBLM_R_X7Y104_SLICE_X8Y104_CO6),
.O5(CLBLM_R_X5Y103_SLICE_X6Y103_AO5),
.O6(CLBLM_R_X5Y103_SLICE_X6Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y103_SLICE_X7Y103_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y103_SLICE_X7Y103_DO5),
.O6(CLBLM_R_X5Y103_SLICE_X7Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y103_SLICE_X7Y103_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y103_SLICE_X7Y103_CO5),
.O6(CLBLM_R_X5Y103_SLICE_X7Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y103_SLICE_X7Y103_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y103_SLICE_X7Y103_BO5),
.O6(CLBLM_R_X5Y103_SLICE_X7Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y103_SLICE_X7Y103_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y103_SLICE_X7Y103_AO5),
.O6(CLBLM_R_X5Y103_SLICE_X7Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y104_SLICE_X6Y104_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y104_SLICE_X6Y104_DO5),
.O6(CLBLM_R_X5Y104_SLICE_X6Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y104_SLICE_X6Y104_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y104_SLICE_X6Y104_CO5),
.O6(CLBLM_R_X5Y104_SLICE_X6Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fff153fd5ff40c0)
  ) CLBLM_R_X5Y104_SLICE_X6Y104_BLUT (
.I0(LIOB33_X0Y111_IOB_X0Y111_I),
.I1(RIOB33_X105Y101_IOB_X1Y102_I),
.I2(LIOB33_X0Y109_IOB_X0Y110_I),
.I3(RIOB33_X105Y101_IOB_X1Y101_I),
.I4(CLBLM_R_X5Y105_SLICE_X6Y105_AO6),
.I5(CLBLM_R_X7Y105_SLICE_X8Y105_BO6),
.O5(CLBLM_R_X5Y104_SLICE_X6Y104_BO5),
.O6(CLBLM_R_X5Y104_SLICE_X6Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h69c3963c993366cc)
  ) CLBLM_R_X5Y104_SLICE_X6Y104_ALUT (
.I0(LIOB33_X0Y111_IOB_X0Y111_I),
.I1(CLBLM_R_X7Y104_SLICE_X8Y104_CO6),
.I2(LIOB33_X0Y109_IOB_X0Y110_I),
.I3(RIOB33_X105Y101_IOB_X1Y102_I),
.I4(CLBLM_R_X5Y103_SLICE_X6Y103_BO6),
.I5(RIOB33_X105Y103_IOB_X1Y103_I),
.O5(CLBLM_R_X5Y104_SLICE_X6Y104_AO5),
.O6(CLBLM_R_X5Y104_SLICE_X6Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y104_SLICE_X7Y104_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y104_SLICE_X7Y104_DO5),
.O6(CLBLM_R_X5Y104_SLICE_X7Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y104_SLICE_X7Y104_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y104_SLICE_X7Y104_CO5),
.O6(CLBLM_R_X5Y104_SLICE_X7Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y104_SLICE_X7Y104_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y104_SLICE_X7Y104_BO5),
.O6(CLBLM_R_X5Y104_SLICE_X7Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y104_SLICE_X7Y104_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y104_SLICE_X7Y104_AO5),
.O6(CLBLM_R_X5Y104_SLICE_X7Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h695aa56996a55a96)
  ) CLBLM_R_X5Y105_SLICE_X6Y105_DLUT (
.I0(CLBLL_L_X4Y104_SLICE_X5Y104_AO6),
.I1(CLBLM_R_X5Y106_SLICE_X6Y106_BO6),
.I2(CLBLM_R_X5Y105_SLICE_X7Y105_DO6),
.I3(CLBLM_R_X5Y106_SLICE_X6Y106_AO6),
.I4(CLBLM_R_X5Y107_SLICE_X6Y107_AO6),
.I5(CLBLL_L_X4Y105_SLICE_X4Y105_AO6),
.O5(CLBLM_R_X5Y105_SLICE_X6Y105_DO5),
.O6(CLBLM_R_X5Y105_SLICE_X6Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h69969966a55a55aa)
  ) CLBLM_R_X5Y105_SLICE_X6Y105_CLUT (
.I0(CLBLM_R_X5Y105_SLICE_X6Y105_AO6),
.I1(RIOB33_X105Y101_IOB_X1Y102_I),
.I2(RIOB33_X105Y101_IOB_X1Y101_I),
.I3(CLBLM_R_X7Y105_SLICE_X8Y105_BO6),
.I4(LIOB33_X0Y111_IOB_X0Y111_I),
.I5(LIOB33_X0Y109_IOB_X0Y110_I),
.O5(CLBLM_R_X5Y105_SLICE_X6Y105_CO5),
.O6(CLBLM_R_X5Y105_SLICE_X6Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h693c96c3c3693c96)
  ) CLBLM_R_X5Y105_SLICE_X6Y105_BLUT (
.I0(CLBLM_R_X5Y107_SLICE_X6Y107_AO6),
.I1(CLBLM_R_X7Y104_SLICE_X8Y104_AO6),
.I2(CLBLL_L_X4Y104_SLICE_X5Y104_AO6),
.I3(CLBLM_R_X5Y106_SLICE_X6Y106_AO6),
.I4(CLBLM_R_X5Y105_SLICE_X6Y105_AO6),
.I5(CLBLM_R_X5Y106_SLICE_X6Y106_BO6),
.O5(CLBLM_R_X5Y105_SLICE_X6Y105_BO5),
.O6(CLBLM_R_X5Y105_SLICE_X6Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h515171f375f7ffff)
  ) CLBLM_R_X5Y105_SLICE_X6Y105_ALUT (
.I0(RIOB33_X105Y101_IOB_X1Y101_I),
.I1(CLBLM_L_X8Y105_SLICE_X11Y105_AO6),
.I2(CLBLM_L_X8Y107_SLICE_X10Y107_BO6),
.I3(LIOB33_X0Y109_IOB_X0Y109_I),
.I4(LIOB33_X0Y109_IOB_X0Y110_I),
.I5(CLBLM_L_X8Y106_SLICE_X11Y106_BO6),
.O5(CLBLM_R_X5Y105_SLICE_X6Y105_AO5),
.O6(CLBLM_R_X5Y105_SLICE_X6Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6c93936c36c9c936)
  ) CLBLM_R_X5Y105_SLICE_X7Y105_DLUT (
.I0(CLBLM_R_X5Y105_SLICE_X7Y105_AO6),
.I1(CLBLM_R_X7Y105_SLICE_X8Y105_AO6),
.I2(CLBLM_L_X8Y106_SLICE_X10Y106_DO6),
.I3(CLBLM_R_X5Y105_SLICE_X7Y105_AO5),
.I4(CLBLM_L_X8Y106_SLICE_X11Y106_DO6),
.I5(CLBLM_L_X8Y106_SLICE_X11Y106_BO6),
.O5(CLBLM_R_X5Y105_SLICE_X7Y105_DO5),
.O6(CLBLM_R_X5Y105_SLICE_X7Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h399cc663c663399c)
  ) CLBLM_R_X5Y105_SLICE_X7Y105_CLUT (
.I0(CLBLM_R_X7Y105_SLICE_X8Y105_AO6),
.I1(CLBLM_R_X7Y105_SLICE_X8Y105_CO6),
.I2(CLBLM_L_X8Y106_SLICE_X11Y106_DO6),
.I3(CLBLM_R_X5Y105_SLICE_X7Y105_AO5),
.I4(CLBLM_R_X7Y103_SLICE_X9Y103_CO6),
.I5(CLBLM_R_X5Y105_SLICE_X7Y105_BO5),
.O5(CLBLM_R_X5Y105_SLICE_X7Y105_CO5),
.O6(CLBLM_R_X5Y105_SLICE_X7Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ffffff0f0fffff)
  ) CLBLM_R_X5Y105_SLICE_X7Y105_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(LIOB33_X0Y109_IOB_X0Y110_I),
.I3(LIOB33_X0Y109_IOB_X0Y109_I),
.I4(RIOB33_X105Y103_IOB_X1Y103_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y105_SLICE_X7Y105_BO5),
.O6(CLBLM_R_X5Y105_SLICE_X7Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555ffff0f0fffff)
  ) CLBLM_R_X5Y105_SLICE_X7Y105_ALUT (
.I0(RIOB33_X105Y101_IOB_X1Y101_I),
.I1(1'b1),
.I2(RIOB33_X105Y101_IOB_X1Y102_I),
.I3(1'b1),
.I4(LIOB33_X0Y109_IOB_X0Y110_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y105_SLICE_X7Y105_AO5),
.O6(CLBLM_R_X5Y105_SLICE_X7Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y106_SLICE_X6Y106_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y106_SLICE_X6Y106_DO5),
.O6(CLBLM_R_X5Y106_SLICE_X6Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8778f0f0e11e5a5a)
  ) CLBLM_R_X5Y106_SLICE_X6Y106_CLUT (
.I0(CLBLM_L_X8Y105_SLICE_X11Y105_AO6),
.I1(RIOB33_X105Y101_IOB_X1Y101_I),
.I2(CLBLM_L_X8Y106_SLICE_X11Y106_CO6),
.I3(RIOB33_X105Y101_IOB_X1Y102_I),
.I4(LIOB33_X0Y109_IOB_X0Y109_I),
.I5(CLBLM_L_X8Y107_SLICE_X10Y107_BO6),
.O5(CLBLM_R_X5Y106_SLICE_X6Y106_CO5),
.O6(CLBLM_R_X5Y106_SLICE_X6Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0a2f2aff0fbfbfff)
  ) CLBLM_R_X5Y106_SLICE_X6Y106_BLUT (
.I0(CLBLM_L_X8Y107_SLICE_X11Y107_DO6),
.I1(LIOB33_X0Y109_IOB_X0Y109_I),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(CLBLM_L_X8Y106_SLICE_X10Y106_BO6),
.I4(LIOB33_X0Y109_IOB_X0Y110_I),
.I5(CLBLM_L_X8Y107_SLICE_X10Y107_CO6),
.O5(CLBLM_R_X5Y106_SLICE_X6Y106_BO5),
.O6(CLBLM_R_X5Y106_SLICE_X6Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hd25a78f0b4961e3c)
  ) CLBLM_R_X5Y106_SLICE_X6Y106_ALUT (
.I0(RIOB33_X105Y101_IOB_X1Y101_I),
.I1(CLBLM_L_X8Y105_SLICE_X11Y105_AO6),
.I2(CLBLM_L_X8Y106_SLICE_X11Y106_BO6),
.I3(LIOB33_X0Y109_IOB_X0Y109_I),
.I4(LIOB33_X0Y109_IOB_X0Y110_I),
.I5(CLBLM_L_X8Y107_SLICE_X10Y107_BO6),
.O5(CLBLM_R_X5Y106_SLICE_X6Y106_AO5),
.O6(CLBLM_R_X5Y106_SLICE_X6Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y106_SLICE_X7Y106_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y106_SLICE_X7Y106_DO5),
.O6(CLBLM_R_X5Y106_SLICE_X7Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h4db2b24db24d4db2)
  ) CLBLM_R_X5Y106_SLICE_X7Y106_CLUT (
.I0(CLBLM_R_X5Y106_SLICE_X7Y106_AO6),
.I1(CLBLM_L_X8Y106_SLICE_X10Y106_BO6),
.I2(CLBLM_R_X7Y107_SLICE_X9Y107_DO6),
.I3(CLBLM_L_X8Y106_SLICE_X10Y106_DO6),
.I4(CLBLM_R_X5Y105_SLICE_X7Y105_AO6),
.I5(CLBLM_L_X8Y106_SLICE_X11Y106_BO6),
.O5(CLBLM_R_X5Y106_SLICE_X7Y106_CO5),
.O6(CLBLM_R_X5Y106_SLICE_X7Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h9c936c936c9c6c6c)
  ) CLBLM_R_X5Y106_SLICE_X7Y106_BLUT (
.I0(RIOB33_X105Y101_IOB_X1Y101_I),
.I1(CLBLM_L_X8Y106_SLICE_X10Y106_CO6),
.I2(LIOB33_X0Y109_IOB_X0Y109_I),
.I3(CLBLM_L_X8Y107_SLICE_X11Y107_DO6),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(CLBLM_L_X8Y107_SLICE_X10Y107_CO6),
.O5(CLBLM_R_X5Y106_SLICE_X7Y106_BO5),
.O6(CLBLM_R_X5Y106_SLICE_X7Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h55ff55ff77777777)
  ) CLBLM_R_X5Y106_SLICE_X7Y106_ALUT (
.I0(LIOB33_X0Y109_IOB_X0Y110_I),
.I1(LIOB33_X0Y115_IOB_X0Y116_I),
.I2(1'b1),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y106_SLICE_X7Y106_AO5),
.O6(CLBLM_R_X5Y106_SLICE_X7Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hc6936c936cc66c6c)
  ) CLBLM_R_X5Y107_SLICE_X6Y107_DLUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(CLBLM_L_X8Y106_SLICE_X10Y106_BO6),
.I2(LIOB33_X0Y109_IOB_X0Y110_I),
.I3(CLBLM_L_X8Y107_SLICE_X11Y107_DO6),
.I4(LIOB33_X0Y109_IOB_X0Y109_I),
.I5(CLBLM_L_X8Y107_SLICE_X10Y107_CO6),
.O5(CLBLM_R_X5Y107_SLICE_X6Y107_DO5),
.O6(CLBLM_R_X5Y107_SLICE_X6Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h69a55a69965aa596)
  ) CLBLM_R_X5Y107_SLICE_X6Y107_CLUT (
.I0(CLBLM_R_X5Y107_SLICE_X6Y107_AO6),
.I1(CLBLM_R_X7Y106_SLICE_X8Y106_CO6),
.I2(CLBLM_R_X5Y106_SLICE_X6Y106_AO6),
.I3(CLBLM_R_X5Y107_SLICE_X6Y107_AO5),
.I4(CLBLM_R_X5Y107_SLICE_X6Y107_DO6),
.I5(CLBLM_R_X5Y106_SLICE_X6Y106_BO6),
.O5(CLBLM_R_X5Y107_SLICE_X6Y107_CO5),
.O6(CLBLM_R_X5Y107_SLICE_X6Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hd25a78f0a5d20f78)
  ) CLBLM_R_X5Y107_SLICE_X6Y107_BLUT (
.I0(LIOB33_X0Y113_IOB_X0Y114_I),
.I1(LIOB33_X0Y109_IOB_X0Y109_I),
.I2(CLBLM_R_X7Y107_SLICE_X8Y107_AO6),
.I3(CLBLM_R_X7Y107_SLICE_X8Y107_BO6),
.I4(LIOB33_X0Y109_IOB_X0Y110_I),
.I5(CLBLM_R_X5Y108_SLICE_X7Y108_CO6),
.O5(CLBLM_R_X5Y107_SLICE_X6Y107_BO5),
.O6(CLBLM_R_X5Y107_SLICE_X6Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333ffff33ff33ff)
  ) CLBLM_R_X5Y107_SLICE_X6Y107_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y111_IOB_X0Y111_I),
.I2(1'b1),
.I3(LIOB33_X0Y115_IOB_X0Y116_I),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y107_SLICE_X6Y107_AO5),
.O6(CLBLM_R_X5Y107_SLICE_X6Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h39c6c6399c63639c)
  ) CLBLM_R_X5Y107_SLICE_X7Y107_DLUT (
.I0(CLBLM_R_X7Y107_SLICE_X8Y107_AO6),
.I1(CLBLM_R_X7Y107_SLICE_X8Y107_DO6),
.I2(CLBLL_L_X4Y107_SLICE_X4Y107_AO5),
.I3(CLBLM_R_X5Y106_SLICE_X7Y106_AO5),
.I4(CLBLM_R_X7Y107_SLICE_X9Y107_BO6),
.I5(CLBLM_R_X7Y108_SLICE_X8Y108_CO6),
.O5(CLBLM_R_X5Y107_SLICE_X7Y107_DO5),
.O6(CLBLM_R_X5Y107_SLICE_X7Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h69a55a69965aa596)
  ) CLBLM_R_X5Y107_SLICE_X7Y107_CLUT (
.I0(CLBLM_R_X5Y106_SLICE_X7Y106_AO6),
.I1(CLBLM_R_X5Y106_SLICE_X7Y106_AO5),
.I2(CLBLM_R_X7Y107_SLICE_X9Y107_DO6),
.I3(CLBLM_R_X7Y107_SLICE_X8Y107_DO6),
.I4(CLBLM_R_X7Y107_SLICE_X9Y107_BO6),
.I5(CLBLM_L_X8Y106_SLICE_X10Y106_BO6),
.O5(CLBLM_R_X5Y107_SLICE_X7Y107_CO5),
.O6(CLBLM_R_X5Y107_SLICE_X7Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h575f7fff11135f7f)
  ) CLBLM_R_X5Y107_SLICE_X7Y107_BLUT (
.I0(LIOB33_X0Y113_IOB_X0Y114_I),
.I1(CLBLM_R_X7Y107_SLICE_X8Y107_BO6),
.I2(LIOB33_X0Y109_IOB_X0Y110_I),
.I3(LIOB33_X0Y109_IOB_X0Y109_I),
.I4(CLBLM_R_X7Y107_SLICE_X8Y107_AO6),
.I5(CLBLM_R_X5Y108_SLICE_X7Y108_CO6),
.O5(CLBLM_R_X5Y107_SLICE_X7Y107_BO5),
.O6(CLBLM_R_X5Y107_SLICE_X7Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h87ff7800e1331ecc)
  ) CLBLM_R_X5Y107_SLICE_X7Y107_ALUT (
.I0(LIOB33_X0Y113_IOB_X0Y114_I),
.I1(CLBLM_R_X7Y107_SLICE_X8Y107_BO6),
.I2(LIOB33_X0Y115_IOB_X0Y116_I),
.I3(LIOB33_X0Y109_IOB_X0Y109_I),
.I4(CLBLM_R_X7Y107_SLICE_X8Y107_CO6),
.I5(CLBLM_R_X5Y108_SLICE_X7Y108_CO6),
.O5(CLBLM_R_X5Y107_SLICE_X7Y107_AO5),
.O6(CLBLM_R_X5Y107_SLICE_X7Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6999666996669996)
  ) CLBLM_R_X5Y108_SLICE_X6Y108_DLUT (
.I0(CLBLM_R_X5Y107_SLICE_X6Y107_AO6),
.I1(CLBLM_R_X5Y108_SLICE_X7Y108_AO5),
.I2(CLBLM_R_X7Y106_SLICE_X8Y106_CO6),
.I3(CLBLM_R_X5Y107_SLICE_X6Y107_AO5),
.I4(CLBLM_R_X5Y107_SLICE_X6Y107_DO6),
.I5(CLBLM_R_X5Y106_SLICE_X7Y106_CO6),
.O5(CLBLM_R_X5Y108_SLICE_X6Y108_DO5),
.O6(CLBLM_R_X5Y108_SLICE_X6Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3c96c36996c3693c)
  ) CLBLM_R_X5Y108_SLICE_X6Y108_CLUT (
.I0(CLBLM_R_X7Y106_SLICE_X8Y106_BO6),
.I1(CLBLM_R_X5Y107_SLICE_X6Y107_AO5),
.I2(CLBLM_R_X7Y106_SLICE_X8Y106_CO6),
.I3(CLBLL_L_X4Y107_SLICE_X5Y107_AO5),
.I4(CLBLM_R_X5Y107_SLICE_X6Y107_DO6),
.I5(CLBLM_R_X5Y107_SLICE_X7Y107_BO6),
.O5(CLBLM_R_X5Y108_SLICE_X6Y108_CO5),
.O6(CLBLM_R_X5Y108_SLICE_X6Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h9af359f3650ca60c)
  ) CLBLM_R_X5Y108_SLICE_X6Y108_BLUT (
.I0(LIOB33_X0Y113_IOB_X0Y114_I),
.I1(CLBLM_R_X5Y108_SLICE_X7Y108_BO6),
.I2(CLBLM_R_X5Y109_SLICE_X6Y109_DO6),
.I3(LIOB33_X0Y109_IOB_X0Y109_I),
.I4(LIOB33_X0Y103_IOB_X0Y103_I),
.I5(CLBLM_R_X7Y108_SLICE_X8Y108_BO6),
.O5(CLBLM_R_X5Y108_SLICE_X6Y108_BO5),
.O6(CLBLM_R_X5Y108_SLICE_X6Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h33ff33ff55ff55ff)
  ) CLBLM_R_X5Y108_SLICE_X6Y108_ALUT (
.I0(LIOB33_X0Y113_IOB_X0Y114_I),
.I1(LIOB33_X0Y103_IOB_X0Y103_I),
.I2(1'b1),
.I3(LIOB33_X0Y109_IOB_X0Y109_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y108_SLICE_X6Y108_AO5),
.O6(CLBLM_R_X5Y108_SLICE_X6Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6a9556a9956aa956)
  ) CLBLM_R_X5Y108_SLICE_X7Y108_DLUT (
.I0(CLBLM_R_X5Y108_SLICE_X7Y108_AO6),
.I1(CLBLL_L_X4Y107_SLICE_X5Y107_AO5),
.I2(CLBLM_R_X5Y107_SLICE_X7Y107_BO6),
.I3(CLBLM_R_X5Y107_SLICE_X6Y107_AO5),
.I4(CLBLM_R_X7Y106_SLICE_X8Y106_BO6),
.I5(CLBLM_R_X5Y107_SLICE_X7Y107_CO6),
.O5(CLBLM_R_X5Y108_SLICE_X7Y108_DO5),
.O6(CLBLM_R_X5Y108_SLICE_X7Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7f13ff5fdf4c5f00)
  ) CLBLM_R_X5Y108_SLICE_X7Y108_CLUT (
.I0(LIOB33_X0Y107_IOB_X0Y108_I),
.I1(LIOB33_X0Y107_IOB_X0Y107_I),
.I2(LIOB33_X0Y113_IOB_X0Y114_I),
.I3(CLBLM_R_X5Y110_SLICE_X7Y110_CO6),
.I4(LIOB33_X0Y115_IOB_X0Y116_I),
.I5(CLBLM_R_X7Y111_SLICE_X9Y111_AO6),
.O5(CLBLM_R_X5Y108_SLICE_X7Y108_CO5),
.O6(CLBLM_R_X5Y108_SLICE_X7Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h69969696a55a5a5a)
  ) CLBLM_R_X5Y108_SLICE_X7Y108_BLUT (
.I0(CLBLM_R_X5Y110_SLICE_X7Y110_CO6),
.I1(LIOB33_X0Y107_IOB_X0Y107_I),
.I2(CLBLM_R_X7Y111_SLICE_X9Y111_AO6),
.I3(LIOB33_X0Y113_IOB_X0Y114_I),
.I4(LIOB33_X0Y107_IOB_X0Y108_I),
.I5(LIOB33_X0Y115_IOB_X0Y116_I),
.O5(CLBLM_R_X5Y108_SLICE_X7Y108_BO5),
.O6(CLBLM_R_X5Y108_SLICE_X7Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0fff0fff3f3f3f3f)
  ) CLBLM_R_X5Y108_SLICE_X7Y108_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y115_IOB_X0Y116_I),
.I2(LIOB33_X0Y111_IOB_X0Y112_I),
.I3(LIOB33_X0Y113_IOB_X0Y114_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y108_SLICE_X7Y108_AO5),
.O6(CLBLM_R_X5Y108_SLICE_X7Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7f13b320ff5fffa0)
  ) CLBLM_R_X5Y109_SLICE_X6Y109_DLUT (
.I0(LIOB33_X0Y107_IOB_X0Y107_I),
.I1(LIOB33_X0Y107_IOB_X0Y108_I),
.I2(LIOB33_X0Y113_IOB_X0Y114_I),
.I3(CLBLM_R_X5Y110_SLICE_X6Y110_CO6),
.I4(CLBLM_R_X5Y110_SLICE_X7Y110_DO6),
.I5(LIOB33_X0Y103_IOB_X0Y103_I),
.O5(CLBLM_R_X5Y109_SLICE_X6Y109_DO5),
.O6(CLBLM_R_X5Y109_SLICE_X6Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6c93936ca05f5fa0)
  ) CLBLM_R_X5Y109_SLICE_X6Y109_CLUT (
.I0(LIOB33_X0Y107_IOB_X0Y107_I),
.I1(LIOB33_X0Y107_IOB_X0Y108_I),
.I2(LIOB33_X0Y113_IOB_X0Y114_I),
.I3(CLBLM_R_X5Y110_SLICE_X6Y110_CO6),
.I4(CLBLM_R_X5Y110_SLICE_X7Y110_DO6),
.I5(LIOB33_X0Y103_IOB_X0Y103_I),
.O5(CLBLM_R_X5Y109_SLICE_X6Y109_CO5),
.O6(CLBLM_R_X5Y109_SLICE_X6Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6969966996699696)
  ) CLBLM_R_X5Y109_SLICE_X6Y109_BLUT (
.I0(CLBLM_R_X5Y110_SLICE_X7Y110_CO6),
.I1(CLBLM_R_X7Y108_SLICE_X8Y108_AO6),
.I2(CLBLM_R_X7Y109_SLICE_X8Y109_AO6),
.I3(CLBLM_R_X5Y110_SLICE_X7Y110_BO6),
.I4(CLBLM_R_X5Y109_SLICE_X6Y109_AO6),
.I5(CLBLM_R_X5Y110_SLICE_X6Y110_CO6),
.O5(CLBLM_R_X5Y109_SLICE_X6Y109_BO5),
.O6(CLBLM_R_X5Y109_SLICE_X6Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f3f3f3f0fff0fff)
  ) CLBLM_R_X5Y109_SLICE_X6Y109_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y103_IOB_X0Y103_I),
.I2(LIOB33_X0Y107_IOB_X0Y108_I),
.I3(RIOB33_X105Y105_IOB_X1Y106_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y109_SLICE_X6Y109_AO5),
.O6(CLBLM_R_X5Y109_SLICE_X6Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y109_SLICE_X7Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y109_SLICE_X7Y109_DO5),
.O6(CLBLM_R_X5Y109_SLICE_X7Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y109_SLICE_X7Y109_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y109_SLICE_X7Y109_CO5),
.O6(CLBLM_R_X5Y109_SLICE_X7Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y109_SLICE_X7Y109_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y109_SLICE_X7Y109_BO5),
.O6(CLBLM_R_X5Y109_SLICE_X7Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000040000000c00)
  ) CLBLM_R_X5Y109_SLICE_X7Y109_ALUT (
.I0(LIOB33_X0Y109_IOB_X0Y110_I),
.I1(RIOB33_X105Y107_IOB_X1Y107_I),
.I2(CLBLM_R_X5Y110_SLICE_X7Y110_AO6),
.I3(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I4(CLBLM_L_X8Y103_SLICE_X11Y103_AO6),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X5Y109_SLICE_X7Y109_AO5),
.O6(CLBLM_R_X5Y109_SLICE_X7Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000002000000)
  ) CLBLM_R_X5Y110_SLICE_X6Y110_DLUT (
.I0(CLBLM_R_X5Y109_SLICE_X7Y109_AO6),
.I1(CLBLL_L_X4Y101_SLICE_X4Y101_AO6),
.I2(CLBLM_R_X5Y113_SLICE_X6Y113_DO6),
.I3(CLBLM_L_X8Y111_SLICE_X10Y111_CO6),
.I4(CLBLM_R_X3Y110_SLICE_X3Y110_DO6),
.I5(CLBLM_R_X5Y112_SLICE_X6Y112_DO6),
.O5(CLBLM_R_X5Y110_SLICE_X6Y110_DO5),
.O6(CLBLM_R_X5Y110_SLICE_X6Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h4d8eddee8e4deedd)
  ) CLBLM_R_X5Y110_SLICE_X6Y110_CLUT (
.I0(CLBLM_R_X7Y111_SLICE_X8Y111_BO6),
.I1(CLBLL_L_X4Y111_SLICE_X5Y111_DO6),
.I2(LIOB33_X0Y103_IOB_X0Y103_I),
.I3(CLBLM_R_X5Y110_SLICE_X6Y110_AO5),
.I4(LIOB33_X0Y107_IOB_X0Y107_I),
.I5(CLBLM_R_X5Y112_SLICE_X6Y112_DO6),
.O5(CLBLM_R_X5Y110_SLICE_X6Y110_CO5),
.O6(CLBLM_R_X5Y110_SLICE_X6Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc36999cc693c99cc)
  ) CLBLM_R_X5Y110_SLICE_X6Y110_BLUT (
.I0(CLBLM_R_X5Y113_SLICE_X6Y113_DO6),
.I1(CLBLM_R_X5Y111_SLICE_X7Y111_BO6),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(CLBLM_R_X5Y110_SLICE_X7Y110_AO5),
.I4(LIOB33_X0Y101_IOB_X0Y101_I),
.I5(LIOB33_X0Y115_IOB_X0Y116_I),
.O5(CLBLM_R_X5Y110_SLICE_X6Y110_BO5),
.O6(CLBLM_R_X5Y110_SLICE_X6Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8778788777777777)
  ) CLBLM_R_X5Y110_SLICE_X6Y110_ALUT (
.I0(LIOB33_X0Y113_IOB_X0Y114_I),
.I1(LIOB33_X0Y105_IOB_X0Y106_I),
.I2(CLBLM_R_X7Y111_SLICE_X8Y111_BO6),
.I3(CLBLM_R_X5Y112_SLICE_X6Y112_DO6),
.I4(CLBLL_L_X4Y111_SLICE_X5Y111_DO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y110_SLICE_X6Y110_AO5),
.O6(CLBLM_R_X5Y110_SLICE_X6Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h96cc3cccc3669666)
  ) CLBLM_R_X5Y110_SLICE_X7Y110_DLUT (
.I0(CLBLM_R_X7Y111_SLICE_X8Y111_BO6),
.I1(CLBLM_R_X7Y112_SLICE_X8Y112_CO6),
.I2(LIOB33_X0Y115_IOB_X0Y116_I),
.I3(LIOB33_X0Y105_IOB_X0Y106_I),
.I4(LIOB33_X0Y113_IOB_X0Y114_I),
.I5(CLBLM_R_X5Y112_SLICE_X6Y112_DO6),
.O5(CLBLM_R_X5Y110_SLICE_X7Y110_DO5),
.O6(CLBLM_R_X5Y110_SLICE_X7Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0d4d0ddd4fffdfff)
  ) CLBLM_R_X5Y110_SLICE_X7Y110_CLUT (
.I0(CLBLM_R_X7Y111_SLICE_X8Y111_BO6),
.I1(CLBLM_R_X5Y112_SLICE_X6Y112_DO6),
.I2(LIOB33_X0Y113_IOB_X0Y114_I),
.I3(LIOB33_X0Y107_IOB_X0Y107_I),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(CLBLM_R_X7Y111_SLICE_X8Y111_CO6),
.O5(CLBLM_R_X5Y110_SLICE_X7Y110_CO5),
.O6(CLBLM_R_X5Y110_SLICE_X7Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'he74d18b265cf9a30)
  ) CLBLM_R_X5Y110_SLICE_X7Y110_BLUT (
.I0(LIOB33_X0Y113_IOB_X0Y114_I),
.I1(CLBLM_R_X5Y112_SLICE_X6Y112_DO6),
.I2(CLBLM_R_X7Y111_SLICE_X8Y111_BO6),
.I3(LIOB33_X0Y107_IOB_X0Y107_I),
.I4(CLBLM_R_X7Y111_SLICE_X8Y111_CO6),
.I5(LIOB33_X0Y105_IOB_X0Y106_I),
.O5(CLBLM_R_X5Y110_SLICE_X7Y110_BO5),
.O6(CLBLM_R_X5Y110_SLICE_X7Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555ffff99395f5f)
  ) CLBLM_R_X5Y110_SLICE_X7Y110_ALUT (
.I0(RIOB33_X105Y113_IOB_X1Y113_I),
.I1(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I2(RIOB33_X105Y101_IOB_X1Y101_I),
.I3(RIOB33_X105Y111_IOB_X1Y112_I),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y110_SLICE_X7Y110_AO5),
.O6(CLBLM_R_X5Y110_SLICE_X7Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6fffcfff06660ccc)
  ) CLBLM_R_X5Y111_SLICE_X6Y111_DLUT (
.I0(LIOB33_X0Y101_IOB_X0Y102_I),
.I1(CLBLM_R_X5Y110_SLICE_X6Y110_BO6),
.I2(LIOB33_X0Y113_IOB_X0Y114_I),
.I3(LIOB33_X0Y103_IOB_X0Y104_I),
.I4(LIOB33_X0Y115_IOB_X0Y116_I),
.I5(CLBLM_R_X5Y111_SLICE_X6Y111_BO6),
.O5(CLBLM_R_X5Y111_SLICE_X6Y111_DO5),
.O6(CLBLM_R_X5Y111_SLICE_X6Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6999699969aa5aaa)
  ) CLBLM_R_X5Y111_SLICE_X6Y111_CLUT (
.I0(CLBLM_R_X5Y113_SLICE_X6Y113_AO6),
.I1(CLBLM_R_X3Y111_SLICE_X3Y111_DO6),
.I2(LIOB33_X0Y115_IOB_X0Y116_I),
.I3(LIOB33_X0Y101_IOB_X0Y101_I),
.I4(LIOB33_X0Y113_IOB_X0Y114_I),
.I5(CLBLM_R_X3Y111_SLICE_X2Y111_AO6),
.O5(CLBLM_R_X5Y111_SLICE_X6Y111_CO5),
.O6(CLBLM_R_X5Y111_SLICE_X6Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'he8b2fcf3e8b2e8b2)
  ) CLBLM_R_X5Y111_SLICE_X6Y111_BLUT (
.I0(CLBLM_R_X3Y111_SLICE_X3Y111_DO6),
.I1(CLBLM_R_X5Y113_SLICE_X7Y113_AO6),
.I2(CLBLM_R_X7Y112_SLICE_X8Y112_AO6),
.I3(CLBLM_R_X5Y113_SLICE_X6Y113_AO6),
.I4(CLBLM_R_X3Y111_SLICE_X2Y111_AO6),
.I5(CLBLM_R_X3Y108_SLICE_X2Y108_AO5),
.O5(CLBLM_R_X5Y111_SLICE_X6Y111_BO5),
.O6(CLBLM_R_X5Y111_SLICE_X6Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h693c96c369699696)
  ) CLBLM_R_X5Y111_SLICE_X6Y111_ALUT (
.I0(CLBLM_R_X3Y111_SLICE_X3Y111_DO6),
.I1(CLBLM_R_X5Y113_SLICE_X7Y113_AO6),
.I2(CLBLM_R_X7Y112_SLICE_X8Y112_AO6),
.I3(CLBLM_R_X3Y111_SLICE_X2Y111_AO6),
.I4(CLBLM_R_X5Y113_SLICE_X6Y113_AO6),
.I5(CLBLM_R_X3Y108_SLICE_X2Y108_AO5),
.O5(CLBLM_R_X5Y111_SLICE_X6Y111_AO5),
.O6(CLBLM_R_X5Y111_SLICE_X6Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h69963cc3c33c6996)
  ) CLBLM_R_X5Y111_SLICE_X7Y111_DLUT (
.I0(CLBLM_R_X5Y111_SLICE_X7Y111_AO6),
.I1(CLBLM_R_X7Y110_SLICE_X9Y110_DO6),
.I2(CLBLM_R_X7Y111_SLICE_X8Y111_DO6),
.I3(CLBLM_R_X5Y111_SLICE_X7Y111_AO5),
.I4(CLBLM_R_X7Y111_SLICE_X8Y111_CO6),
.I5(CLBLM_R_X5Y112_SLICE_X7Y112_BO6),
.O5(CLBLM_R_X5Y111_SLICE_X7Y111_DO5),
.O6(CLBLM_R_X5Y111_SLICE_X7Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h65a69a599a5965a6)
  ) CLBLM_R_X5Y111_SLICE_X7Y111_CLUT (
.I0(CLBLM_R_X5Y111_SLICE_X7Y111_AO6),
.I1(CLBLL_L_X4Y111_SLICE_X5Y111_DO6),
.I2(CLBLM_R_X5Y112_SLICE_X7Y112_CO6),
.I3(CLBLM_R_X3Y111_SLICE_X3Y111_AO5),
.I4(CLBLM_R_X7Y111_SLICE_X8Y111_CO6),
.I5(CLBLM_R_X5Y112_SLICE_X7Y112_BO6),
.O5(CLBLM_R_X5Y111_SLICE_X7Y111_CO5),
.O6(CLBLM_R_X5Y111_SLICE_X7Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h134cb1ee66660000)
  ) CLBLM_R_X5Y111_SLICE_X7Y111_BLUT (
.I0(RIOB33_X105Y101_IOB_X1Y101_I),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(RIOB33_X105Y111_IOB_X1Y112_I),
.I3(RIOB33_X105Y101_IOB_X1Y102_I),
.I4(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I5(RIOB33_X105Y113_IOB_X1Y113_I),
.O5(CLBLM_R_X5Y111_SLICE_X7Y111_BO5),
.O6(CLBLM_R_X5Y111_SLICE_X7Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h7777777733ff33ff)
  ) CLBLM_R_X5Y111_SLICE_X7Y111_ALUT (
.I0(LIOB33_X0Y113_IOB_X0Y114_I),
.I1(LIOB33_X0Y107_IOB_X0Y107_I),
.I2(1'b1),
.I3(LIOB33_X0Y115_IOB_X0Y116_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y111_SLICE_X7Y111_AO5),
.O6(CLBLM_R_X5Y111_SLICE_X7Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fd5ffff15403fc0)
  ) CLBLM_R_X5Y112_SLICE_X6Y112_DLUT (
.I0(LIOB33_X0Y105_IOB_X0Y105_I),
.I1(LIOB33_X0Y115_IOB_X0Y116_I),
.I2(LIOB33_X0Y103_IOB_X0Y104_I),
.I3(CLBLM_R_X5Y112_SLICE_X6Y112_CO6),
.I4(LIOB33_X0Y113_IOB_X0Y114_I),
.I5(CLBLM_R_X5Y111_SLICE_X6Y111_DO6),
.O5(CLBLM_R_X5Y112_SLICE_X6Y112_DO5),
.O6(CLBLM_R_X5Y112_SLICE_X6Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h95a96a56ff0f00f0)
  ) CLBLM_R_X5Y112_SLICE_X6Y112_CLUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(LIOB33_X0Y115_IOB_X0Y116_I),
.I2(CLBLM_R_X7Y113_SLICE_X8Y113_AO6),
.I3(CLBLM_R_X5Y112_SLICE_X6Y112_AO5),
.I4(CLBLM_R_X7Y113_SLICE_X9Y113_CO6),
.I5(LIOB33_X0Y101_IOB_X0Y102_I),
.O5(CLBLM_R_X5Y112_SLICE_X6Y112_CO5),
.O6(CLBLM_R_X5Y112_SLICE_X6Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h693cc36996c33c96)
  ) CLBLM_R_X5Y112_SLICE_X6Y112_BLUT (
.I0(CLBLL_L_X4Y112_SLICE_X4Y112_AO5),
.I1(CLBLM_R_X7Y113_SLICE_X9Y113_BO6),
.I2(CLBLM_R_X7Y112_SLICE_X9Y112_AO6),
.I3(CLBLM_R_X5Y113_SLICE_X6Y113_BO6),
.I4(CLBLM_R_X5Y111_SLICE_X6Y111_BO6),
.I5(CLBLM_R_X5Y113_SLICE_X6Y113_CO6),
.O5(CLBLM_R_X5Y112_SLICE_X6Y112_BO5),
.O6(CLBLM_R_X5Y112_SLICE_X6Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc3c30f0f22bbaaff)
  ) CLBLM_R_X5Y112_SLICE_X6Y112_ALUT (
.I0(CLBLM_R_X5Y113_SLICE_X6Y113_DO6),
.I1(LIOB33_X0Y115_IOB_X0Y116_I),
.I2(CLBLM_R_X5Y113_SLICE_X6Y113_AO6),
.I3(CLBLM_R_X5Y110_SLICE_X7Y110_AO5),
.I4(LIOB33_X0Y101_IOB_X0Y101_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y112_SLICE_X6Y112_AO5),
.O6(CLBLM_R_X5Y112_SLICE_X6Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996c33c96963c3c)
  ) CLBLM_R_X5Y112_SLICE_X7Y112_DLUT (
.I0(LIOB33_X0Y103_IOB_X0Y104_I),
.I1(CLBLM_R_X5Y113_SLICE_X6Y113_CO6),
.I2(CLBLM_R_X7Y113_SLICE_X9Y113_CO6),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(LIOB33_X0Y115_IOB_X0Y116_I),
.I5(LIOB33_X0Y101_IOB_X0Y102_I),
.O5(CLBLM_R_X5Y112_SLICE_X7Y112_DO5),
.O6(CLBLM_R_X5Y112_SLICE_X7Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h78871ee18778e11e)
  ) CLBLM_R_X5Y112_SLICE_X7Y112_CLUT (
.I0(CLBLM_R_X5Y112_SLICE_X7Y112_AO6),
.I1(CLBLM_R_X5Y111_SLICE_X6Y111_DO6),
.I2(CLBLM_R_X5Y110_SLICE_X6Y110_AO5),
.I3(CLBLM_R_X5Y112_SLICE_X7Y112_AO5),
.I4(CLBLM_R_X5Y112_SLICE_X7Y112_DO6),
.I5(CLBLM_R_X7Y112_SLICE_X9Y112_DO6),
.O5(CLBLM_R_X5Y112_SLICE_X7Y112_CO5),
.O6(CLBLM_R_X5Y112_SLICE_X7Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdd0f440d0fd40f4)
  ) CLBLM_R_X5Y112_SLICE_X7Y112_BLUT (
.I0(CLBLM_R_X5Y112_SLICE_X7Y112_DO6),
.I1(CLBLM_R_X5Y111_SLICE_X6Y111_DO6),
.I2(CLBLM_R_X5Y110_SLICE_X6Y110_AO5),
.I3(CLBLM_R_X7Y112_SLICE_X9Y112_DO6),
.I4(CLBLM_R_X5Y112_SLICE_X7Y112_AO6),
.I5(CLBLM_R_X5Y112_SLICE_X7Y112_AO5),
.O5(CLBLM_R_X5Y112_SLICE_X7Y112_BO5),
.O6(CLBLM_R_X5Y112_SLICE_X7Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0fffff5555ffff)
  ) CLBLM_R_X5Y112_SLICE_X7Y112_ALUT (
.I0(LIOB33_X0Y115_IOB_X0Y116_I),
.I1(1'b1),
.I2(LIOB33_X0Y113_IOB_X0Y114_I),
.I3(1'b1),
.I4(LIOB33_X0Y105_IOB_X0Y105_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y112_SLICE_X7Y112_AO5),
.O6(CLBLM_R_X5Y112_SLICE_X7Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hd505d505ffffffff)
  ) CLBLM_R_X5Y113_SLICE_X6Y113_DLUT (
.I0(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I1(RIOB33_X105Y111_IOB_X1Y112_I),
.I2(RIOB33_X105Y113_IOB_X1Y113_I),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(1'b1),
.I5(LIOB33_X0Y115_IOB_X0Y116_I),
.O5(CLBLM_R_X5Y113_SLICE_X6Y113_DO5),
.O6(CLBLM_R_X5Y113_SLICE_X6Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'he8d48844eedde8d4)
  ) CLBLM_R_X5Y113_SLICE_X6Y113_CLUT (
.I0(CLBLM_R_X7Y113_SLICE_X9Y113_AO6),
.I1(CLBLM_R_X5Y113_SLICE_X7Y113_AO5),
.I2(CLBLM_R_X5Y113_SLICE_X7Y113_AO6),
.I3(CLBLM_R_X5Y111_SLICE_X7Y111_BO6),
.I4(CLBLM_R_X5Y113_SLICE_X6Y113_DO6),
.I5(CLBLM_R_X5Y110_SLICE_X7Y110_AO5),
.O5(CLBLM_R_X5Y113_SLICE_X6Y113_CO5),
.O6(CLBLM_R_X5Y113_SLICE_X6Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h4db2b24db24d4db2)
  ) CLBLM_R_X5Y113_SLICE_X6Y113_BLUT (
.I0(CLBLM_R_X5Y113_SLICE_X6Y113_DO6),
.I1(CLBLM_R_X5Y110_SLICE_X7Y110_AO5),
.I2(CLBLM_R_X5Y113_SLICE_X7Y113_AO6),
.I3(CLBLM_R_X5Y113_SLICE_X7Y113_AO5),
.I4(CLBLM_R_X7Y113_SLICE_X9Y113_AO6),
.I5(CLBLM_R_X5Y111_SLICE_X7Y111_BO6),
.O5(CLBLM_R_X5Y113_SLICE_X6Y113_BO5),
.O6(CLBLM_R_X5Y113_SLICE_X6Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h1d5500f02daaf000)
  ) CLBLM_R_X5Y113_SLICE_X6Y113_ALUT (
.I0(RIOB33_X105Y101_IOB_X1Y101_I),
.I1(RIOB33_X105Y111_IOB_X1Y112_I),
.I2(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(RIOB33_X105Y113_IOB_X1Y113_I),
.I5(LIOB33_X0Y115_IOB_X0Y116_I),
.O5(CLBLM_R_X5Y113_SLICE_X6Y113_AO5),
.O6(CLBLM_R_X5Y113_SLICE_X6Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y113_SLICE_X7Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y113_SLICE_X7Y113_DO5),
.O6(CLBLM_R_X5Y113_SLICE_X7Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y113_SLICE_X7Y113_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y113_SLICE_X7Y113_CO5),
.O6(CLBLM_R_X5Y113_SLICE_X7Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y113_SLICE_X7Y113_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y113_SLICE_X7Y113_BO5),
.O6(CLBLM_R_X5Y113_SLICE_X7Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f3f3f3f33ff33ff)
  ) CLBLM_R_X5Y113_SLICE_X7Y113_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y115_IOB_X0Y116_I),
.I2(LIOB33_X0Y101_IOB_X0Y101_I),
.I3(LIOB33_X0Y101_IOB_X0Y102_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y113_SLICE_X7Y113_AO5),
.O6(CLBLM_R_X5Y113_SLICE_X7Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y100_SLICE_X8Y100_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y100_SLICE_X8Y100_DO5),
.O6(CLBLM_R_X7Y100_SLICE_X8Y100_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y100_SLICE_X8Y100_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y100_SLICE_X8Y100_CO5),
.O6(CLBLM_R_X7Y100_SLICE_X8Y100_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y100_SLICE_X8Y100_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y100_SLICE_X8Y100_BO5),
.O6(CLBLM_R_X7Y100_SLICE_X8Y100_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f3f3f3f5f5f5f5f)
  ) CLBLM_R_X7Y100_SLICE_X8Y100_ALUT (
.I0(LIOB33_X0Y105_IOB_X0Y105_I),
.I1(LIOB33_X0Y105_IOB_X0Y106_I),
.I2(RIOB33_X105Y107_IOB_X1Y107_I),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y100_SLICE_X8Y100_AO5),
.O6(CLBLM_R_X7Y100_SLICE_X8Y100_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y100_SLICE_X9Y100_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y100_SLICE_X9Y100_DO5),
.O6(CLBLM_R_X7Y100_SLICE_X9Y100_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y100_SLICE_X9Y100_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y100_SLICE_X9Y100_CO5),
.O6(CLBLM_R_X7Y100_SLICE_X9Y100_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y100_SLICE_X9Y100_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y100_SLICE_X9Y100_BO5),
.O6(CLBLM_R_X7Y100_SLICE_X9Y100_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y100_SLICE_X9Y100_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y100_SLICE_X9Y100_AO5),
.O6(CLBLM_R_X7Y100_SLICE_X9Y100_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996696996966996)
  ) CLBLM_R_X7Y101_SLICE_X8Y101_DLUT (
.I0(CLBLM_L_X8Y101_SLICE_X11Y101_BO6),
.I1(CLBLL_L_X4Y100_SLICE_X4Y100_AO5),
.I2(CLBLM_R_X5Y100_SLICE_X6Y100_AO5),
.I3(CLBLM_L_X8Y103_SLICE_X11Y103_AO5),
.I4(CLBLM_L_X8Y101_SLICE_X11Y101_CO6),
.I5(CLBLM_L_X8Y100_SLICE_X10Y100_CO6),
.O5(CLBLM_R_X7Y101_SLICE_X8Y101_DO5),
.O6(CLBLM_R_X7Y101_SLICE_X8Y101_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h93ff6c00c95536aa)
  ) CLBLM_R_X7Y101_SLICE_X8Y101_CLUT (
.I0(CLBLM_L_X8Y101_SLICE_X10Y101_BO6),
.I1(RIOB33_X105Y107_IOB_X1Y108_I),
.I2(RIOB33_X105Y107_IOB_X1Y107_I),
.I3(LIOB33_X0Y105_IOB_X0Y105_I),
.I4(CLBLM_R_X7Y101_SLICE_X8Y101_DO6),
.I5(CLBLM_L_X8Y101_SLICE_X10Y101_CO6),
.O5(CLBLM_R_X7Y101_SLICE_X8Y101_CO5),
.O6(CLBLM_R_X7Y101_SLICE_X8Y101_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfab2f571b2a07150)
  ) CLBLM_R_X7Y101_SLICE_X8Y101_BLUT (
.I0(CLBLM_R_X7Y101_SLICE_X8Y101_DO6),
.I1(CLBLM_L_X8Y101_SLICE_X10Y101_BO6),
.I2(CLBLM_R_X7Y100_SLICE_X8Y100_AO6),
.I3(CLBLM_L_X8Y101_SLICE_X10Y101_CO6),
.I4(CLBLM_R_X7Y102_SLICE_X8Y102_AO6),
.I5(CLBLM_R_X7Y100_SLICE_X8Y100_AO5),
.O5(CLBLM_R_X7Y101_SLICE_X8Y101_BO5),
.O6(CLBLM_R_X7Y101_SLICE_X8Y101_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5a96a56996a5695a)
  ) CLBLM_R_X7Y101_SLICE_X8Y101_ALUT (
.I0(CLBLM_R_X7Y101_SLICE_X8Y101_DO6),
.I1(CLBLM_L_X8Y101_SLICE_X10Y101_BO6),
.I2(CLBLM_R_X7Y102_SLICE_X8Y102_AO6),
.I3(CLBLM_L_X8Y101_SLICE_X10Y101_CO6),
.I4(CLBLM_R_X7Y100_SLICE_X8Y100_AO6),
.I5(CLBLM_R_X7Y100_SLICE_X8Y100_AO5),
.O5(CLBLM_R_X7Y101_SLICE_X8Y101_AO5),
.O6(CLBLM_R_X7Y101_SLICE_X8Y101_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h55ff55ff55ff55ff)
  ) CLBLM_R_X7Y101_SLICE_X9Y101_DLUT (
.I0(LIOB33_X0Y107_IOB_X0Y107_I),
.I1(1'b1),
.I2(1'b1),
.I3(RIOB33_X105Y107_IOB_X1Y107_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y101_SLICE_X9Y101_DO5),
.O6(CLBLM_R_X7Y101_SLICE_X9Y101_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h054dcfcf4d5fffff)
  ) CLBLM_R_X7Y101_SLICE_X9Y101_CLUT (
.I0(LIOB33_X0Y103_IOB_X0Y104_I),
.I1(CLBLM_L_X8Y100_SLICE_X10Y100_AO5),
.I2(CLBLM_L_X8Y101_SLICE_X11Y101_CO6),
.I3(LIOB33_X0Y101_IOB_X0Y102_I),
.I4(RIOB33_X105Y107_IOB_X1Y108_I),
.I5(CLBLM_L_X8Y101_SLICE_X11Y101_AO6),
.O5(CLBLM_R_X7Y101_SLICE_X9Y101_CO5),
.O6(CLBLM_R_X7Y101_SLICE_X9Y101_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha5c369c369f05af0)
  ) CLBLM_R_X7Y101_SLICE_X9Y101_BLUT (
.I0(RIOB33_X105Y107_IOB_X1Y107_I),
.I1(CLBLM_L_X8Y102_SLICE_X10Y102_BO6),
.I2(CLBLM_R_X7Y101_SLICE_X8Y101_CO6),
.I3(LIOB33_X0Y105_IOB_X0Y106_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X7Y101_SLICE_X9Y101_AO5),
.O5(CLBLM_R_X7Y101_SLICE_X9Y101_BO5),
.O6(CLBLM_R_X7Y101_SLICE_X9Y101_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h44ccddff66cc9933)
  ) CLBLM_R_X7Y101_SLICE_X9Y101_ALUT (
.I0(RIOB33_X105Y107_IOB_X1Y107_I),
.I1(CLBLM_L_X8Y101_SLICE_X10Y101_CO6),
.I2(1'b1),
.I3(LIOB33_X0Y105_IOB_X0Y105_I),
.I4(CLBLM_L_X8Y101_SLICE_X10Y101_BO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y101_SLICE_X9Y101_AO5),
.O6(CLBLM_R_X7Y101_SLICE_X9Y101_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h9a956a956a9a6a6a)
  ) CLBLM_R_X7Y102_SLICE_X8Y102_DLUT (
.I0(CLBLM_R_X5Y101_SLICE_X7Y101_BO6),
.I1(LIOB33_X0Y105_IOB_X0Y106_I),
.I2(RIOB33_X105Y107_IOB_X1Y108_I),
.I3(CLBLM_R_X7Y101_SLICE_X9Y101_CO6),
.I4(LIOB33_X0Y105_IOB_X0Y105_I),
.I5(CLBLM_R_X5Y102_SLICE_X7Y102_BO6),
.O5(CLBLM_R_X7Y102_SLICE_X8Y102_DO5),
.O6(CLBLM_R_X7Y102_SLICE_X8Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h9f5f60a0a09f5f60)
  ) CLBLM_R_X7Y102_SLICE_X8Y102_CLUT (
.I0(LIOB33_X0Y107_IOB_X0Y107_I),
.I1(LIOB33_X0Y105_IOB_X0Y106_I),
.I2(RIOB33_X105Y107_IOB_X1Y107_I),
.I3(CLBLM_R_X7Y102_SLICE_X8Y102_AO5),
.I4(CLBLM_R_X7Y102_SLICE_X8Y102_DO6),
.I5(CLBLM_R_X7Y101_SLICE_X9Y101_AO6),
.O5(CLBLM_R_X7Y102_SLICE_X8Y102_CO5),
.O6(CLBLM_R_X7Y102_SLICE_X8Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h37157f157f377f7f)
  ) CLBLM_R_X7Y102_SLICE_X8Y102_BLUT (
.I0(CLBLM_R_X7Y102_SLICE_X8Y102_DO6),
.I1(RIOB33_X105Y107_IOB_X1Y107_I),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(CLBLM_R_X7Y101_SLICE_X9Y101_AO6),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(CLBLM_R_X7Y102_SLICE_X8Y102_AO5),
.O5(CLBLM_R_X7Y102_SLICE_X8Y102_BO5),
.O6(CLBLM_R_X7Y102_SLICE_X8Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ffffff66999999)
  ) CLBLM_R_X7Y102_SLICE_X8Y102_ALUT (
.I0(CLBLM_R_X7Y101_SLICE_X9Y101_CO6),
.I1(CLBLM_R_X5Y102_SLICE_X7Y102_BO6),
.I2(1'b1),
.I3(LIOB33_X0Y105_IOB_X0Y105_I),
.I4(RIOB33_X105Y107_IOB_X1Y108_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y102_SLICE_X8Y102_AO5),
.O6(CLBLM_R_X7Y102_SLICE_X8Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7888877787777888)
  ) CLBLM_R_X7Y102_SLICE_X9Y102_DLUT (
.I0(LIOB33_X0Y107_IOB_X0Y107_I),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(LIOB33_X0Y107_IOB_X0Y108_I),
.I3(RIOB33_X105Y103_IOB_X1Y104_I),
.I4(CLBLM_R_X7Y103_SLICE_X9Y103_DO6),
.I5(CLBLM_R_X7Y101_SLICE_X9Y101_BO6),
.O5(CLBLM_R_X7Y102_SLICE_X9Y102_DO5),
.O6(CLBLM_R_X7Y102_SLICE_X9Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fff07778fff0888)
  ) CLBLM_R_X7Y102_SLICE_X9Y102_CLUT (
.I0(LIOB33_X0Y107_IOB_X0Y107_I),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(LIOB33_X0Y107_IOB_X0Y108_I),
.I3(RIOB33_X105Y103_IOB_X1Y104_I),
.I4(CLBLM_R_X7Y103_SLICE_X9Y103_DO6),
.I5(CLBLM_R_X7Y101_SLICE_X9Y101_BO6),
.O5(CLBLM_R_X7Y102_SLICE_X9Y102_CO5),
.O6(CLBLM_R_X7Y102_SLICE_X9Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h69a55a69965aa596)
  ) CLBLM_R_X7Y102_SLICE_X9Y102_BLUT (
.I0(CLBLM_R_X7Y101_SLICE_X9Y101_DO6),
.I1(CLBLM_R_X7Y103_SLICE_X9Y103_AO6),
.I2(CLBLM_R_X7Y101_SLICE_X8Y101_BO6),
.I3(CLBLM_L_X8Y103_SLICE_X10Y103_DO6),
.I4(CLBLM_R_X7Y101_SLICE_X8Y101_AO6),
.I5(CLBLM_R_X7Y102_SLICE_X8Y102_DO6),
.O5(CLBLM_R_X7Y102_SLICE_X9Y102_BO5),
.O6(CLBLM_R_X7Y102_SLICE_X9Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5f5f5f5f7f7f1313)
  ) CLBLM_R_X7Y102_SLICE_X9Y102_ALUT (
.I0(LIOB33_X0Y109_IOB_X0Y109_I),
.I1(CLBLM_R_X7Y103_SLICE_X8Y103_AO5),
.I2(RIOB33_X105Y103_IOB_X1Y104_I),
.I3(1'b1),
.I4(CLBLM_R_X7Y102_SLICE_X9Y102_CO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y102_SLICE_X9Y102_AO5),
.O6(CLBLM_R_X7Y102_SLICE_X9Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h9a65a5a559a6aaaa)
  ) CLBLM_R_X7Y103_SLICE_X8Y103_DLUT (
.I0(CLBLM_R_X7Y102_SLICE_X9Y102_BO6),
.I1(RIOB33_X105Y103_IOB_X1Y104_I),
.I2(CLBLM_R_X7Y103_SLICE_X9Y103_DO6),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(LIOB33_X0Y107_IOB_X0Y108_I),
.I5(CLBLM_R_X7Y103_SLICE_X8Y103_BO6),
.O5(CLBLM_R_X7Y103_SLICE_X8Y103_DO5),
.O6(CLBLM_R_X7Y103_SLICE_X8Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h71f5b2fab2fab2fa)
  ) CLBLM_R_X7Y103_SLICE_X8Y103_CLUT (
.I0(CLBLM_R_X7Y101_SLICE_X8Y101_CO6),
.I1(LIOB33_X0Y107_IOB_X0Y107_I),
.I2(CLBLM_L_X8Y103_SLICE_X10Y103_DO6),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(RIOB33_X105Y107_IOB_X1Y107_I),
.O5(CLBLM_R_X7Y103_SLICE_X8Y103_CO5),
.O6(CLBLM_R_X7Y103_SLICE_X8Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h69c3963ca50f5af0)
  ) CLBLM_R_X7Y103_SLICE_X8Y103_BLUT (
.I0(LIOB33_X0Y107_IOB_X0Y107_I),
.I1(LIOB33_X0Y105_IOB_X0Y106_I),
.I2(CLBLM_R_X7Y101_SLICE_X8Y101_CO6),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_L_X8Y103_SLICE_X10Y103_DO6),
.I5(RIOB33_X105Y107_IOB_X1Y107_I),
.O5(CLBLM_R_X7Y103_SLICE_X8Y103_BO5),
.O6(CLBLM_R_X7Y103_SLICE_X8Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5fff050f5af0a50f)
  ) CLBLM_R_X7Y103_SLICE_X8Y103_ALUT (
.I0(LIOB33_X0Y107_IOB_X0Y108_I),
.I1(1'b1),
.I2(CLBLM_R_X7Y102_SLICE_X8Y102_CO6),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X7Y103_SLICE_X8Y103_CO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y103_SLICE_X8Y103_AO5),
.O6(CLBLM_R_X7Y103_SLICE_X8Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h1171f3ff7177f3ff)
  ) CLBLM_R_X7Y103_SLICE_X9Y103_DLUT (
.I0(LIOB33_X0Y107_IOB_X0Y107_I),
.I1(CLBLM_L_X8Y103_SLICE_X10Y103_BO6),
.I2(CLBLM_L_X10Y104_SLICE_X12Y104_DO6),
.I3(CLBLM_L_X8Y103_SLICE_X11Y103_CO6),
.I4(RIOB33_X105Y103_IOB_X1Y104_I),
.I5(LIOB33_X0Y105_IOB_X0Y106_I),
.O5(CLBLM_R_X7Y103_SLICE_X9Y103_DO5),
.O6(CLBLM_R_X7Y103_SLICE_X9Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h659aa6599a6559a6)
  ) CLBLM_R_X7Y103_SLICE_X9Y103_CLUT (
.I0(CLBLM_R_X7Y102_SLICE_X9Y102_AO6),
.I1(CLBLM_L_X8Y104_SLICE_X10Y104_AO5),
.I2(CLBLM_R_X7Y103_SLICE_X8Y103_BO6),
.I3(CLBLM_R_X7Y103_SLICE_X9Y103_AO5),
.I4(CLBLM_R_X7Y103_SLICE_X9Y103_DO6),
.I5(CLBLM_R_X7Y102_SLICE_X9Y102_BO6),
.O5(CLBLM_R_X7Y103_SLICE_X9Y103_CO5),
.O6(CLBLM_R_X7Y103_SLICE_X9Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6696996996996966)
  ) CLBLM_R_X7Y103_SLICE_X9Y103_BLUT (
.I0(CLBLM_L_X8Y103_SLICE_X10Y103_DO6),
.I1(CLBLM_R_X7Y101_SLICE_X8Y101_AO6),
.I2(CLBLM_L_X8Y103_SLICE_X10Y103_BO6),
.I3(CLBLM_L_X10Y103_SLICE_X12Y103_BO6),
.I4(CLBLM_R_X7Y103_SLICE_X9Y103_AO6),
.I5(CLBLM_R_X7Y105_SLICE_X9Y105_AO5),
.O5(CLBLM_R_X7Y103_SLICE_X9Y103_BO5),
.O6(CLBLM_R_X7Y103_SLICE_X9Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f3f3f3f77777777)
  ) CLBLM_R_X7Y103_SLICE_X9Y103_ALUT (
.I0(LIOB33_X0Y107_IOB_X0Y108_I),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y103_SLICE_X9Y103_AO5),
.O6(CLBLM_R_X7Y103_SLICE_X9Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h2a80bfeabfeabfea)
  ) CLBLM_R_X7Y104_SLICE_X8Y104_DLUT (
.I0(CLBLM_L_X8Y104_SLICE_X11Y104_BO6),
.I1(RIOB33_X105Y103_IOB_X1Y104_I),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(CLBLM_L_X8Y104_SLICE_X10Y104_BO6),
.I4(LIOB33_X0Y107_IOB_X0Y108_I),
.I5(RIOB33_X105Y103_IOB_X1Y103_I),
.O5(CLBLM_R_X7Y104_SLICE_X8Y104_DO5),
.O6(CLBLM_R_X7Y104_SLICE_X8Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h445d4cff55dfdfff)
  ) CLBLM_R_X7Y104_SLICE_X8Y104_CLUT (
.I0(RIOB33_X105Y101_IOB_X1Y102_I),
.I1(CLBLM_L_X8Y105_SLICE_X11Y105_DO6),
.I2(LIOB33_X0Y109_IOB_X0Y109_I),
.I3(CLBLM_R_X7Y105_SLICE_X8Y105_AO6),
.I4(LIOB33_X0Y109_IOB_X0Y110_I),
.I5(CLBLM_R_X7Y104_SLICE_X8Y104_BO6),
.O5(CLBLM_R_X7Y104_SLICE_X8Y104_CO5),
.O6(CLBLM_R_X7Y104_SLICE_X8Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7887877888777788)
  ) CLBLM_R_X7Y104_SLICE_X8Y104_BLUT (
.I0(LIOB33_X0Y107_IOB_X0Y108_I),
.I1(RIOB33_X105Y103_IOB_X1Y103_I),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(CLBLM_L_X8Y104_SLICE_X10Y104_BO6),
.I4(CLBLM_L_X8Y104_SLICE_X11Y104_BO6),
.I5(RIOB33_X105Y103_IOB_X1Y104_I),
.O5(CLBLM_R_X7Y104_SLICE_X8Y104_BO5),
.O6(CLBLM_R_X7Y104_SLICE_X8Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hda4f2abf25b0d540)
  ) CLBLM_R_X7Y104_SLICE_X8Y104_ALUT (
.I0(CLBLM_L_X8Y105_SLICE_X11Y105_DO6),
.I1(LIOB33_X0Y109_IOB_X0Y109_I),
.I2(RIOB33_X105Y101_IOB_X1Y102_I),
.I3(CLBLM_R_X7Y104_SLICE_X8Y104_BO6),
.I4(LIOB33_X0Y109_IOB_X0Y110_I),
.I5(CLBLM_R_X7Y105_SLICE_X8Y105_AO6),
.O5(CLBLM_R_X7Y104_SLICE_X8Y104_AO5),
.O6(CLBLM_R_X7Y104_SLICE_X8Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y104_SLICE_X9Y104_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y104_SLICE_X9Y104_DO5),
.O6(CLBLM_R_X7Y104_SLICE_X9Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y104_SLICE_X9Y104_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y104_SLICE_X9Y104_CO5),
.O6(CLBLM_R_X7Y104_SLICE_X9Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y104_SLICE_X9Y104_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y104_SLICE_X9Y104_BO5),
.O6(CLBLM_R_X7Y104_SLICE_X9Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hd42b2bd4bb44bb44)
  ) CLBLM_R_X7Y104_SLICE_X9Y104_ALUT (
.I0(CLBLM_L_X10Y104_SLICE_X12Y104_DO6),
.I1(CLBLM_L_X8Y103_SLICE_X11Y103_CO6),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(CLBLM_L_X8Y103_SLICE_X10Y103_BO6),
.I4(LIOB33_X0Y107_IOB_X0Y107_I),
.I5(RIOB33_X105Y103_IOB_X1Y104_I),
.O5(CLBLM_R_X7Y104_SLICE_X9Y104_AO5),
.O6(CLBLM_R_X7Y104_SLICE_X9Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hb478d21e3cf0965a)
  ) CLBLM_R_X7Y105_SLICE_X8Y105_DLUT (
.I0(CLBLM_R_X7Y104_SLICE_X9Y104_AO6),
.I1(LIOB33_X0Y107_IOB_X0Y108_I),
.I2(CLBLM_R_X7Y103_SLICE_X9Y103_BO6),
.I3(RIOB33_X105Y103_IOB_X1Y104_I),
.I4(CLBLM_L_X8Y104_SLICE_X11Y104_BO6),
.I5(RIOB33_X105Y103_IOB_X1Y103_I),
.O5(CLBLM_R_X7Y105_SLICE_X8Y105_DO5),
.O6(CLBLM_R_X7Y105_SLICE_X8Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfddff44fd00d4004)
  ) CLBLM_R_X7Y105_SLICE_X8Y105_CLUT (
.I0(CLBLM_R_X7Y104_SLICE_X9Y104_AO6),
.I1(CLBLM_L_X8Y106_SLICE_X11Y106_AO6),
.I2(CLBLM_R_X7Y103_SLICE_X9Y103_BO6),
.I3(CLBLM_L_X8Y104_SLICE_X10Y104_AO5),
.I4(CLBLM_L_X8Y104_SLICE_X11Y104_BO6),
.I5(CLBLM_R_X5Y105_SLICE_X7Y105_BO6),
.O5(CLBLM_R_X7Y105_SLICE_X8Y105_CO5),
.O6(CLBLM_R_X7Y105_SLICE_X8Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha69966a66a55aa6a)
  ) CLBLM_R_X7Y105_SLICE_X8Y105_BLUT (
.I0(CLBLM_R_X7Y105_SLICE_X8Y105_DO6),
.I1(LIOB33_X0Y109_IOB_X0Y109_I),
.I2(RIOB33_X105Y101_IOB_X1Y102_I),
.I3(CLBLM_L_X8Y105_SLICE_X11Y105_DO6),
.I4(CLBLM_R_X7Y104_SLICE_X8Y104_BO6),
.I5(RIOB33_X105Y103_IOB_X1Y103_I),
.O5(CLBLM_R_X7Y105_SLICE_X8Y105_BO5),
.O6(CLBLM_R_X7Y105_SLICE_X8Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6c9336c9936cc936)
  ) CLBLM_R_X7Y105_SLICE_X8Y105_ALUT (
.I0(CLBLM_L_X8Y104_SLICE_X11Y104_BO6),
.I1(CLBLM_R_X7Y103_SLICE_X9Y103_BO6),
.I2(CLBLM_L_X8Y106_SLICE_X11Y106_AO6),
.I3(CLBLM_R_X5Y105_SLICE_X7Y105_BO6),
.I4(CLBLM_R_X7Y104_SLICE_X9Y104_AO6),
.I5(CLBLM_L_X8Y104_SLICE_X10Y104_AO5),
.O5(CLBLM_R_X7Y105_SLICE_X8Y105_AO5),
.O6(CLBLM_R_X7Y105_SLICE_X8Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y105_SLICE_X9Y105_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y105_SLICE_X9Y105_DO5),
.O6(CLBLM_R_X7Y105_SLICE_X9Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y105_SLICE_X9Y105_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y105_SLICE_X9Y105_CO5),
.O6(CLBLM_R_X7Y105_SLICE_X9Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y105_SLICE_X9Y105_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y105_SLICE_X9Y105_BO5),
.O6(CLBLM_R_X7Y105_SLICE_X9Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0fffff0fff0fff)
  ) CLBLM_R_X7Y105_SLICE_X9Y105_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(RIOB33_X105Y103_IOB_X1Y104_I),
.I4(RIOB33_X105Y101_IOB_X1Y102_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y105_SLICE_X9Y105_AO5),
.O6(CLBLM_R_X7Y105_SLICE_X9Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hc6aa395563ff9c00)
  ) CLBLM_R_X7Y106_SLICE_X8Y106_DLUT (
.I0(CLBLM_R_X7Y106_SLICE_X8Y106_AO6),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(LIOB33_X0Y115_IOB_X0Y116_I),
.I3(LIOB33_X0Y109_IOB_X0Y109_I),
.I4(CLBLM_R_X7Y107_SLICE_X9Y107_CO6),
.I5(CLBLM_L_X8Y107_SLICE_X11Y107_BO6),
.O5(CLBLM_R_X7Y106_SLICE_X8Y106_DO5),
.O6(CLBLM_R_X7Y106_SLICE_X8Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h032bafaf2b3fffff)
  ) CLBLM_R_X7Y106_SLICE_X8Y106_CLUT (
.I0(CLBLM_R_X7Y106_SLICE_X8Y106_AO6),
.I1(LIOB33_X0Y109_IOB_X0Y110_I),
.I2(CLBLM_R_X7Y107_SLICE_X9Y107_BO6),
.I3(LIOB33_X0Y109_IOB_X0Y109_I),
.I4(LIOB33_X0Y115_IOB_X0Y116_I),
.I5(CLBLM_L_X8Y107_SLICE_X11Y107_BO6),
.O5(CLBLM_R_X7Y106_SLICE_X8Y106_CO5),
.O6(CLBLM_R_X7Y106_SLICE_X8Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc66c93c66c6c936c)
  ) CLBLM_R_X7Y106_SLICE_X8Y106_BLUT (
.I0(LIOB33_X0Y115_IOB_X0Y116_I),
.I1(CLBLM_R_X7Y107_SLICE_X9Y107_BO6),
.I2(LIOB33_X0Y109_IOB_X0Y110_I),
.I3(CLBLM_L_X8Y107_SLICE_X11Y107_BO6),
.I4(CLBLM_R_X7Y106_SLICE_X8Y106_AO6),
.I5(LIOB33_X0Y109_IOB_X0Y109_I),
.O5(CLBLM_R_X7Y106_SLICE_X8Y106_BO5),
.O6(CLBLM_R_X7Y106_SLICE_X8Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h7d14dd44ff3cffcc)
  ) CLBLM_R_X7Y106_SLICE_X8Y106_ALUT (
.I0(LIOB33_X0Y115_IOB_X0Y116_I),
.I1(CLBLM_L_X8Y108_SLICE_X11Y108_BO6),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(CLBLM_R_X7Y109_SLICE_X8Y109_BO6),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(LIOB33_X0Y107_IOB_X0Y108_I),
.O5(CLBLM_R_X7Y106_SLICE_X8Y106_AO5),
.O6(CLBLM_R_X7Y106_SLICE_X8Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y106_SLICE_X9Y106_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y106_SLICE_X9Y106_DO5),
.O6(CLBLM_R_X7Y106_SLICE_X9Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y106_SLICE_X9Y106_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y106_SLICE_X9Y106_CO5),
.O6(CLBLM_R_X7Y106_SLICE_X9Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y106_SLICE_X9Y106_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y106_SLICE_X9Y106_BO5),
.O6(CLBLM_R_X7Y106_SLICE_X9Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333ffff33ff33ff)
  ) CLBLM_R_X7Y106_SLICE_X9Y106_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y107_IOB_X0Y108_I),
.I2(1'b1),
.I3(RIOB33_X105Y101_IOB_X1Y101_I),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y106_SLICE_X9Y106_AO5),
.O6(CLBLM_R_X7Y106_SLICE_X9Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'heedd8e4d8e4d8844)
  ) CLBLM_R_X7Y107_SLICE_X8Y107_DLUT (
.I0(CLBLM_R_X7Y106_SLICE_X9Y106_AO6),
.I1(CLBLM_R_X7Y107_SLICE_X9Y107_AO6),
.I2(CLBLM_L_X8Y107_SLICE_X11Y107_AO6),
.I3(CLBLM_L_X8Y108_SLICE_X10Y108_BO6),
.I4(CLBLM_R_X7Y108_SLICE_X8Y108_AO5),
.I5(CLBLM_R_X7Y109_SLICE_X8Y109_BO6),
.O5(CLBLM_R_X7Y107_SLICE_X8Y107_DO5),
.O6(CLBLM_R_X7Y107_SLICE_X8Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hb74877888b748778)
  ) CLBLM_R_X7Y107_SLICE_X8Y107_CLUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(LIOB33_X0Y107_IOB_X0Y108_I),
.I2(CLBLM_L_X8Y107_SLICE_X11Y107_AO6),
.I3(CLBLM_L_X8Y108_SLICE_X10Y108_BO6),
.I4(LIOB33_X0Y115_IOB_X0Y116_I),
.I5(CLBLM_R_X7Y109_SLICE_X8Y109_BO6),
.O5(CLBLM_R_X7Y107_SLICE_X8Y107_CO5),
.O6(CLBLM_R_X7Y107_SLICE_X8Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6c93a05f936c5fa0)
  ) CLBLM_R_X7Y107_SLICE_X8Y107_BLUT (
.I0(LIOB33_X0Y115_IOB_X0Y116_I),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(LIOB33_X0Y107_IOB_X0Y108_I),
.I3(CLBLM_R_X7Y109_SLICE_X8Y109_BO6),
.I4(LIOB33_X0Y107_IOB_X0Y107_I),
.I5(CLBLM_L_X8Y108_SLICE_X11Y108_BO6),
.O5(CLBLM_R_X7Y107_SLICE_X8Y107_BO5),
.O6(CLBLM_R_X7Y107_SLICE_X8Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h4bb4b44bd22d2dd2)
  ) CLBLM_R_X7Y107_SLICE_X8Y107_ALUT (
.I0(CLBLM_R_X7Y108_SLICE_X8Y108_AO5),
.I1(CLBLM_L_X8Y107_SLICE_X11Y107_AO6),
.I2(CLBLM_R_X7Y107_SLICE_X9Y107_AO6),
.I3(CLBLM_L_X8Y108_SLICE_X10Y108_BO6),
.I4(CLBLM_R_X7Y106_SLICE_X9Y106_AO6),
.I5(CLBLM_R_X7Y109_SLICE_X8Y109_BO6),
.O5(CLBLM_R_X7Y107_SLICE_X8Y107_AO5),
.O6(CLBLM_R_X7Y107_SLICE_X8Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbb0f220bf0b2f02)
  ) CLBLM_R_X7Y107_SLICE_X9Y107_DLUT (
.I0(CLBLM_R_X7Y106_SLICE_X9Y106_AO6),
.I1(CLBLM_L_X8Y108_SLICE_X10Y108_CO6),
.I2(CLBLM_L_X8Y107_SLICE_X10Y107_AO6),
.I3(CLBLM_R_X7Y107_SLICE_X9Y107_AO5),
.I4(CLBLM_L_X8Y107_SLICE_X11Y107_CO6),
.I5(CLBLM_R_X7Y106_SLICE_X9Y106_AO5),
.O5(CLBLM_R_X7Y107_SLICE_X9Y107_DO5),
.O6(CLBLM_R_X7Y107_SLICE_X9Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h963cc396cccc33cc)
  ) CLBLM_R_X7Y107_SLICE_X9Y107_CLUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(CLBLM_L_X8Y107_SLICE_X10Y107_AO6),
.I2(RIOB33_X105Y101_IOB_X1Y101_I),
.I3(CLBLM_L_X8Y108_SLICE_X10Y108_CO6),
.I4(CLBLM_L_X8Y107_SLICE_X11Y107_CO6),
.I5(LIOB33_X0Y107_IOB_X0Y108_I),
.O5(CLBLM_R_X7Y107_SLICE_X9Y107_CO5),
.O6(CLBLM_R_X7Y107_SLICE_X9Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h399cc663c663399c)
  ) CLBLM_R_X7Y107_SLICE_X9Y107_BLUT (
.I0(CLBLM_L_X8Y108_SLICE_X10Y108_CO6),
.I1(CLBLM_L_X8Y107_SLICE_X10Y107_AO6),
.I2(CLBLM_R_X7Y106_SLICE_X9Y106_AO6),
.I3(CLBLM_L_X8Y107_SLICE_X11Y107_CO6),
.I4(CLBLM_R_X7Y106_SLICE_X9Y106_AO5),
.I5(CLBLM_R_X7Y107_SLICE_X9Y107_AO5),
.O5(CLBLM_R_X7Y107_SLICE_X9Y107_BO5),
.O6(CLBLM_R_X7Y107_SLICE_X9Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h7777777733ff33ff)
  ) CLBLM_R_X7Y107_SLICE_X9Y107_ALUT (
.I0(LIOB33_X0Y115_IOB_X0Y116_I),
.I1(LIOB33_X0Y109_IOB_X0Y109_I),
.I2(1'b1),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y107_SLICE_X9Y107_AO5),
.O6(CLBLM_R_X7Y107_SLICE_X9Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996c33c3cc36996)
  ) CLBLM_R_X7Y108_SLICE_X8Y108_DLUT (
.I0(CLBLM_R_X7Y108_SLICE_X8Y108_AO6),
.I1(CLBLM_R_X5Y108_SLICE_X6Y108_AO5),
.I2(CLBLM_R_X7Y108_SLICE_X9Y108_AO6),
.I3(CLBLM_R_X7Y108_SLICE_X8Y108_AO5),
.I4(CLBLM_R_X5Y110_SLICE_X7Y110_CO6),
.I5(CLBLM_R_X7Y109_SLICE_X8Y109_AO6),
.O5(CLBLM_R_X7Y108_SLICE_X8Y108_DO5),
.O6(CLBLM_R_X7Y108_SLICE_X8Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'he88ec00cfccfe88e)
  ) CLBLM_R_X7Y108_SLICE_X8Y108_CLUT (
.I0(CLBLM_R_X7Y108_SLICE_X8Y108_AO6),
.I1(CLBLM_R_X5Y108_SLICE_X6Y108_AO5),
.I2(CLBLM_R_X7Y108_SLICE_X9Y108_AO6),
.I3(CLBLM_R_X7Y108_SLICE_X8Y108_AO5),
.I4(CLBLM_R_X5Y110_SLICE_X7Y110_CO6),
.I5(CLBLM_R_X7Y109_SLICE_X8Y109_AO6),
.O5(CLBLM_R_X7Y108_SLICE_X8Y108_CO5),
.O6(CLBLM_R_X7Y108_SLICE_X8Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h96c3f00f3c96f0f0)
  ) CLBLM_R_X7Y108_SLICE_X8Y108_BLUT (
.I0(LIOB33_X0Y113_IOB_X0Y114_I),
.I1(LIOB33_X0Y115_IOB_X0Y116_I),
.I2(CLBLM_R_X7Y108_SLICE_X9Y108_AO6),
.I3(CLBLM_R_X5Y110_SLICE_X7Y110_CO6),
.I4(LIOB33_X0Y107_IOB_X0Y108_I),
.I5(CLBLM_R_X7Y109_SLICE_X8Y109_AO6),
.O5(CLBLM_R_X7Y108_SLICE_X8Y108_BO5),
.O6(CLBLM_R_X7Y108_SLICE_X8Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5f5f5f5f0fff0fff)
  ) CLBLM_R_X7Y108_SLICE_X8Y108_ALUT (
.I0(LIOB33_X0Y113_IOB_X0Y114_I),
.I1(1'b1),
.I2(LIOB33_X0Y107_IOB_X0Y108_I),
.I3(LIOB33_X0Y115_IOB_X0Y116_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y108_SLICE_X8Y108_AO5),
.O6(CLBLM_R_X7Y108_SLICE_X8Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y108_SLICE_X9Y108_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y108_SLICE_X9Y108_DO5),
.O6(CLBLM_R_X7Y108_SLICE_X9Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y108_SLICE_X9Y108_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y108_SLICE_X9Y108_CO5),
.O6(CLBLM_R_X7Y108_SLICE_X9Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y108_SLICE_X9Y108_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y108_SLICE_X9Y108_BO5),
.O6(CLBLM_R_X7Y108_SLICE_X9Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6c9336c9936cc936)
  ) CLBLM_R_X7Y108_SLICE_X9Y108_ALUT (
.I0(CLBLM_R_X7Y111_SLICE_X8Y111_DO6),
.I1(CLBLM_L_X10Y108_SLICE_X12Y108_BO6),
.I2(CLBLM_R_X5Y111_SLICE_X7Y111_AO5),
.I3(CLBLM_L_X8Y108_SLICE_X10Y108_AO6),
.I4(CLBLM_R_X7Y110_SLICE_X9Y110_DO6),
.I5(CLBLM_R_X7Y110_SLICE_X9Y110_CO6),
.O5(CLBLM_R_X7Y108_SLICE_X9Y108_AO5),
.O6(CLBLM_R_X7Y108_SLICE_X9Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y109_SLICE_X8Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y109_SLICE_X8Y109_DO5),
.O6(CLBLM_R_X7Y109_SLICE_X8Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y109_SLICE_X8Y109_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y109_SLICE_X8Y109_CO5),
.O6(CLBLM_R_X7Y109_SLICE_X8Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h2888beeebeeebeee)
  ) CLBLM_R_X7Y109_SLICE_X8Y109_BLUT (
.I0(CLBLM_R_X7Y111_SLICE_X8Y111_DO6),
.I1(CLBLM_R_X7Y110_SLICE_X9Y110_BO6),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(LIOB33_X0Y105_IOB_X0Y106_I),
.I4(LIOB33_X0Y107_IOB_X0Y107_I),
.I5(LIOB33_X0Y115_IOB_X0Y116_I),
.O5(CLBLM_R_X7Y109_SLICE_X8Y109_BO5),
.O6(CLBLM_R_X7Y109_SLICE_X8Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6999966696669666)
  ) CLBLM_R_X7Y109_SLICE_X8Y109_ALUT (
.I0(CLBLM_R_X7Y111_SLICE_X8Y111_DO6),
.I1(CLBLM_R_X7Y110_SLICE_X9Y110_BO6),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(LIOB33_X0Y105_IOB_X0Y106_I),
.I4(LIOB33_X0Y107_IOB_X0Y107_I),
.I5(LIOB33_X0Y115_IOB_X0Y116_I),
.O5(CLBLM_R_X7Y109_SLICE_X8Y109_AO5),
.O6(CLBLM_R_X7Y109_SLICE_X8Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y109_SLICE_X9Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y109_SLICE_X9Y109_DO5),
.O6(CLBLM_R_X7Y109_SLICE_X9Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y109_SLICE_X9Y109_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y109_SLICE_X9Y109_CO5),
.O6(CLBLM_R_X7Y109_SLICE_X9Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y109_SLICE_X9Y109_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y109_SLICE_X9Y109_BO5),
.O6(CLBLM_R_X7Y109_SLICE_X9Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y109_SLICE_X9Y109_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y109_SLICE_X9Y109_AO5),
.O6(CLBLM_R_X7Y109_SLICE_X9Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y110_SLICE_X8Y110_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y110_SLICE_X8Y110_DO5),
.O6(CLBLM_R_X7Y110_SLICE_X8Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y110_SLICE_X8Y110_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y110_SLICE_X8Y110_CO5),
.O6(CLBLM_R_X7Y110_SLICE_X8Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y110_SLICE_X8Y110_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y110_SLICE_X8Y110_BO5),
.O6(CLBLM_R_X7Y110_SLICE_X8Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y110_SLICE_X8Y110_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y110_SLICE_X8Y110_AO5),
.O6(CLBLM_R_X7Y110_SLICE_X8Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6c9336c9936cc936)
  ) CLBLM_R_X7Y110_SLICE_X9Y110_DLUT (
.I0(CLBLM_R_X7Y110_SLICE_X9Y110_AO6),
.I1(CLBLM_R_X7Y111_SLICE_X8Y111_AO5),
.I2(CLBLM_L_X8Y112_SLICE_X10Y112_DO6),
.I3(CLBLM_R_X7Y110_SLICE_X9Y110_AO5),
.I4(CLBLM_L_X8Y110_SLICE_X10Y110_AO6),
.I5(CLBLM_L_X8Y110_SLICE_X11Y110_CO6),
.O5(CLBLM_R_X7Y110_SLICE_X9Y110_DO5),
.O6(CLBLM_R_X7Y110_SLICE_X9Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hecb38020fefbc832)
  ) CLBLM_R_X7Y110_SLICE_X9Y110_CLUT (
.I0(CLBLM_R_X7Y110_SLICE_X9Y110_AO6),
.I1(CLBLM_L_X8Y110_SLICE_X11Y110_CO6),
.I2(CLBLM_L_X8Y112_SLICE_X10Y112_DO6),
.I3(CLBLM_R_X7Y110_SLICE_X9Y110_AO5),
.I4(CLBLM_R_X7Y111_SLICE_X8Y111_AO5),
.I5(CLBLM_L_X8Y110_SLICE_X10Y110_AO6),
.O5(CLBLM_R_X7Y110_SLICE_X9Y110_CO5),
.O6(CLBLM_R_X7Y110_SLICE_X9Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha659659acc33ff00)
  ) CLBLM_R_X7Y110_SLICE_X9Y110_BLUT (
.I0(RIOB33_X105Y101_IOB_X1Y101_I),
.I1(CLBLM_L_X8Y112_SLICE_X10Y112_DO6),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(CLBLM_L_X8Y110_SLICE_X11Y110_CO6),
.I4(CLBLM_L_X8Y110_SLICE_X10Y110_AO6),
.I5(LIOB33_X0Y105_IOB_X0Y105_I),
.O5(CLBLM_R_X7Y110_SLICE_X9Y110_BO5),
.O6(CLBLM_R_X7Y110_SLICE_X9Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555ffff5f5f5f5f)
  ) CLBLM_R_X7Y110_SLICE_X9Y110_ALUT (
.I0(LIOB33_X0Y105_IOB_X0Y105_I),
.I1(1'b1),
.I2(RIOB33_X105Y101_IOB_X1Y101_I),
.I3(1'b1),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y110_SLICE_X9Y110_AO5),
.O6(CLBLM_R_X7Y110_SLICE_X9Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'he8eed4dd88e844d4)
  ) CLBLM_R_X7Y111_SLICE_X8Y111_DLUT (
.I0(CLBLM_R_X7Y110_SLICE_X9Y110_AO6),
.I1(CLBLM_R_X7Y111_SLICE_X8Y111_AO6),
.I2(CLBLM_R_X7Y112_SLICE_X8Y112_BO6),
.I3(CLBLM_R_X7Y112_SLICE_X9Y112_CO6),
.I4(CLBLM_L_X8Y112_SLICE_X10Y112_CO6),
.I5(CLBLM_R_X5Y112_SLICE_X7Y112_AO5),
.O5(CLBLM_R_X7Y111_SLICE_X8Y111_DO5),
.O6(CLBLM_R_X7Y111_SLICE_X8Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6966969999696696)
  ) CLBLM_R_X7Y111_SLICE_X8Y111_CLUT (
.I0(CLBLM_R_X7Y110_SLICE_X9Y110_AO6),
.I1(CLBLM_R_X7Y111_SLICE_X8Y111_AO6),
.I2(CLBLM_R_X7Y112_SLICE_X8Y112_BO6),
.I3(CLBLM_R_X7Y112_SLICE_X9Y112_CO6),
.I4(CLBLM_L_X8Y112_SLICE_X10Y112_CO6),
.I5(CLBLM_R_X5Y112_SLICE_X7Y112_AO5),
.O5(CLBLM_R_X7Y111_SLICE_X8Y111_CO5),
.O6(CLBLM_R_X7Y111_SLICE_X8Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h69969696c33c3c3c)
  ) CLBLM_R_X7Y111_SLICE_X8Y111_BLUT (
.I0(LIOB33_X0Y115_IOB_X0Y116_I),
.I1(CLBLM_R_X7Y112_SLICE_X9Y112_BO6),
.I2(CLBLM_R_X7Y112_SLICE_X8Y112_BO6),
.I3(LIOB33_X0Y103_IOB_X0Y104_I),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(LIOB33_X0Y105_IOB_X0Y105_I),
.O5(CLBLM_R_X7Y111_SLICE_X8Y111_BO5),
.O6(CLBLM_R_X7Y111_SLICE_X8Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h777777773f3f3f3f)
  ) CLBLM_R_X7Y111_SLICE_X8Y111_ALUT (
.I0(LIOB33_X0Y115_IOB_X0Y116_I),
.I1(LIOB33_X0Y105_IOB_X0Y106_I),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y111_SLICE_X8Y111_AO5),
.O6(CLBLM_R_X7Y111_SLICE_X8Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y111_SLICE_X9Y111_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y111_SLICE_X9Y111_DO5),
.O6(CLBLM_R_X7Y111_SLICE_X9Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fff07778fff0888)
  ) CLBLM_R_X7Y111_SLICE_X9Y111_CLUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(LIOB33_X0Y103_IOB_X0Y104_I),
.I2(LIOB33_X0Y115_IOB_X0Y116_I),
.I3(LIOB33_X0Y105_IOB_X0Y105_I),
.I4(CLBLM_R_X7Y112_SLICE_X8Y112_BO6),
.I5(CLBLM_R_X7Y112_SLICE_X9Y112_BO6),
.O5(CLBLM_R_X7Y111_SLICE_X9Y111_CO5),
.O6(CLBLM_R_X7Y111_SLICE_X9Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h69a5965a995566aa)
  ) CLBLM_R_X7Y111_SLICE_X9Y111_BLUT (
.I0(CLBLM_L_X8Y112_SLICE_X10Y112_DO6),
.I1(LIOB33_X0Y103_IOB_X0Y104_I),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(RIOB33_X105Y101_IOB_X1Y101_I),
.I4(CLBLM_L_X8Y111_SLICE_X10Y111_AO6),
.I5(LIOB33_X0Y105_IOB_X0Y105_I),
.O5(CLBLM_R_X7Y111_SLICE_X9Y111_BO5),
.O6(CLBLM_R_X7Y111_SLICE_X9Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h9c3c6cccc39c336c)
  ) CLBLM_R_X7Y111_SLICE_X9Y111_ALUT (
.I0(LIOB33_X0Y115_IOB_X0Y116_I),
.I1(CLBLM_R_X7Y110_SLICE_X9Y110_BO6),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(CLBLM_R_X7Y111_SLICE_X9Y111_BO6),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(CLBLM_R_X7Y111_SLICE_X9Y111_CO6),
.O5(CLBLM_R_X7Y111_SLICE_X9Y111_AO5),
.O6(CLBLM_R_X7Y111_SLICE_X9Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y112_SLICE_X8Y112_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y112_SLICE_X8Y112_DO5),
.O6(CLBLM_R_X7Y112_SLICE_X8Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h96f05af0a53c963c)
  ) CLBLM_R_X7Y112_SLICE_X8Y112_CLUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(CLBLM_R_X7Y112_SLICE_X9Y112_CO6),
.I2(CLBLM_L_X8Y112_SLICE_X10Y112_CO6),
.I3(LIOB33_X0Y105_IOB_X0Y105_I),
.I4(LIOB33_X0Y115_IOB_X0Y116_I),
.I5(CLBLM_R_X7Y112_SLICE_X8Y112_BO6),
.O5(CLBLM_R_X7Y112_SLICE_X8Y112_CO5),
.O6(CLBLM_R_X7Y112_SLICE_X8Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7bffbbff125a22aa)
  ) CLBLM_R_X7Y112_SLICE_X8Y112_BLUT (
.I0(CLBLM_R_X7Y113_SLICE_X9Y113_CO6),
.I1(LIOB33_X0Y103_IOB_X0Y104_I),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(LIOB33_X0Y115_IOB_X0Y116_I),
.I4(LIOB33_X0Y101_IOB_X0Y102_I),
.I5(CLBLM_R_X5Y113_SLICE_X6Y113_CO6),
.O5(CLBLM_R_X7Y112_SLICE_X8Y112_BO5),
.O6(CLBLM_R_X7Y112_SLICE_X8Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ffffff0f0fffff)
  ) CLBLM_R_X7Y112_SLICE_X8Y112_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(LIOB33_X0Y113_IOB_X0Y114_I),
.I4(LIOB33_X0Y101_IOB_X0Y102_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y112_SLICE_X8Y112_AO5),
.O6(CLBLM_R_X7Y112_SLICE_X8Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h78871ee18778e11e)
  ) CLBLM_R_X7Y112_SLICE_X9Y112_DLUT (
.I0(CLBLM_R_X7Y112_SLICE_X9Y112_AO6),
.I1(CLBLM_R_X5Y113_SLICE_X6Y113_CO6),
.I2(CLBLM_R_X7Y113_SLICE_X9Y113_DO6),
.I3(CLBLM_L_X8Y112_SLICE_X11Y112_DO6),
.I4(CLBLM_R_X7Y113_SLICE_X9Y113_BO6),
.I5(CLBLM_R_X7Y113_SLICE_X9Y113_AO5),
.O5(CLBLM_R_X7Y112_SLICE_X9Y112_DO5),
.O6(CLBLM_R_X7Y112_SLICE_X9Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996a55ac33c0ff0)
  ) CLBLM_R_X7Y112_SLICE_X9Y112_CLUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(LIOB33_X0Y101_IOB_X0Y102_I),
.I2(CLBLM_R_X7Y113_SLICE_X9Y113_DO6),
.I3(CLBLM_L_X8Y112_SLICE_X10Y112_BO6),
.I4(RIOB33_X105Y101_IOB_X1Y101_I),
.I5(LIOB33_X0Y103_IOB_X0Y104_I),
.O5(CLBLM_R_X7Y112_SLICE_X9Y112_CO5),
.O6(CLBLM_R_X7Y112_SLICE_X9Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h9fa35f93605ca06c)
  ) CLBLM_R_X7Y112_SLICE_X9Y112_BLUT (
.I0(RIOB33_X105Y101_IOB_X1Y101_I),
.I1(CLBLM_L_X8Y112_SLICE_X10Y112_AO6),
.I2(LIOB33_X0Y101_IOB_X0Y102_I),
.I3(CLBLM_R_X7Y113_SLICE_X8Y113_AO5),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(CLBLM_L_X8Y112_SLICE_X10Y112_BO6),
.O5(CLBLM_R_X7Y112_SLICE_X9Y112_BO5),
.O6(CLBLM_R_X7Y112_SLICE_X9Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h55ff55ff0fff0fff)
  ) CLBLM_R_X7Y112_SLICE_X9Y112_ALUT (
.I0(LIOB33_X0Y115_IOB_X0Y116_I),
.I1(1'b1),
.I2(RIOB33_X105Y101_IOB_X1Y101_I),
.I3(LIOB33_X0Y103_IOB_X0Y104_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y112_SLICE_X9Y112_AO5),
.O6(CLBLM_R_X7Y112_SLICE_X9Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y113_SLICE_X8Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y113_SLICE_X8Y113_DO5),
.O6(CLBLM_R_X7Y113_SLICE_X8Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y113_SLICE_X8Y113_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y113_SLICE_X8Y113_CO5),
.O6(CLBLM_R_X7Y113_SLICE_X8Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h08086c280008e428)
  ) CLBLM_R_X7Y113_SLICE_X8Y113_BLUT (
.I0(RIOB33_X105Y101_IOB_X1Y101_I),
.I1(RIOB33_X105Y113_IOB_X1Y113_I),
.I2(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I3(RIOB33_X105Y101_IOB_X1Y102_I),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(RIOB33_X105Y111_IOB_X1Y112_I),
.O5(CLBLM_R_X7Y113_SLICE_X8Y113_BO5),
.O6(CLBLM_R_X7Y113_SLICE_X8Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h93939393ff13ff13)
  ) CLBLM_R_X7Y113_SLICE_X8Y113_ALUT (
.I0(LIOB33_X0Y101_IOB_X0Y101_I),
.I1(CLBLM_R_X5Y111_SLICE_X7Y111_BO6),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(CLBLM_R_X7Y113_SLICE_X8Y113_BO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y113_SLICE_X8Y113_AO5),
.O6(CLBLM_R_X7Y113_SLICE_X8Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfec0c8c0c8fcfe)
  ) CLBLM_R_X7Y113_SLICE_X9Y113_DLUT (
.I0(CLBLM_R_X7Y113_SLICE_X9Y113_AO6),
.I1(CLBLM_R_X7Y112_SLICE_X8Y112_AO5),
.I2(CLBLM_R_X7Y113_SLICE_X8Y113_BO6),
.I3(CLBLM_R_X5Y111_SLICE_X7Y111_BO6),
.I4(CLBLM_L_X8Y112_SLICE_X11Y112_AO6),
.I5(CLBLM_L_X8Y113_SLICE_X11Y113_AO6),
.O5(CLBLM_R_X7Y113_SLICE_X9Y113_DO5),
.O6(CLBLM_R_X7Y113_SLICE_X9Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3cf0c30f39ffc600)
  ) CLBLM_R_X7Y113_SLICE_X9Y113_CLUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(RIOB33_X105Y101_IOB_X1Y101_I),
.I2(CLBLM_R_X7Y113_SLICE_X8Y113_BO6),
.I3(LIOB33_X0Y101_IOB_X0Y101_I),
.I4(CLBLM_L_X8Y112_SLICE_X11Y112_AO6),
.I5(CLBLM_R_X5Y111_SLICE_X7Y111_BO6),
.O5(CLBLM_R_X7Y113_SLICE_X9Y113_CO5),
.O6(CLBLM_R_X7Y113_SLICE_X9Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h699669965aa56996)
  ) CLBLM_R_X7Y113_SLICE_X9Y113_BLUT (
.I0(CLBLM_R_X7Y112_SLICE_X8Y112_AO5),
.I1(CLBLM_R_X7Y113_SLICE_X8Y113_BO6),
.I2(CLBLM_L_X8Y112_SLICE_X11Y112_AO6),
.I3(CLBLM_L_X8Y113_SLICE_X11Y113_AO6),
.I4(CLBLM_R_X7Y113_SLICE_X9Y113_AO6),
.I5(CLBLM_R_X5Y111_SLICE_X7Y111_BO6),
.O5(CLBLM_R_X7Y113_SLICE_X9Y113_BO5),
.O6(CLBLM_R_X7Y113_SLICE_X9Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555ffff3333ffff)
  ) CLBLM_R_X7Y113_SLICE_X9Y113_ALUT (
.I0(LIOB33_X0Y101_IOB_X0Y101_I),
.I1(LIOB33_X0Y103_IOB_X0Y104_I),
.I2(1'b1),
.I3(1'b1),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y113_SLICE_X9Y113_AO5),
.O6(CLBLM_R_X7Y113_SLICE_X9Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5aa55a96aa55aaaa)
  ) CLBLM_R_X11Y106_SLICE_X14Y106_DLUT (
.I0(CLBLM_L_X10Y104_SLICE_X13Y104_AO6),
.I1(RIOB33_X105Y103_IOB_X1Y104_I),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_L_X10Y105_SLICE_X13Y105_AO6),
.I4(CLBLM_L_X10Y109_SLICE_X12Y109_BO6),
.I5(LIOB33_X0Y101_IOB_X0Y101_I),
.O5(CLBLM_R_X11Y106_SLICE_X14Y106_DO5),
.O6(CLBLM_R_X11Y106_SLICE_X14Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffc3ffc3c300eb82)
  ) CLBLM_R_X11Y106_SLICE_X14Y106_CLUT (
.I0(CLBLM_R_X11Y106_SLICE_X14Y106_AO6),
.I1(CLBLM_L_X10Y104_SLICE_X13Y104_AO6),
.I2(CLBLM_R_X5Y102_SLICE_X6Y102_AO6),
.I3(CLBLM_R_X11Y106_SLICE_X14Y106_AO5),
.I4(CLBLM_L_X10Y109_SLICE_X12Y109_BO6),
.I5(CLBLM_L_X10Y105_SLICE_X13Y105_AO6),
.O5(CLBLM_R_X11Y106_SLICE_X14Y106_CO5),
.O6(CLBLM_R_X11Y106_SLICE_X14Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3c963cc3c369c33c)
  ) CLBLM_R_X11Y106_SLICE_X14Y106_BLUT (
.I0(CLBLM_L_X10Y109_SLICE_X12Y109_BO6),
.I1(CLBLM_R_X5Y102_SLICE_X6Y102_AO6),
.I2(CLBLM_L_X10Y104_SLICE_X13Y104_AO6),
.I3(CLBLM_L_X10Y105_SLICE_X13Y105_AO6),
.I4(CLBLM_R_X11Y106_SLICE_X14Y106_AO6),
.I5(CLBLM_R_X11Y106_SLICE_X14Y106_AO5),
.O5(CLBLM_R_X11Y106_SLICE_X14Y106_BO5),
.O6(CLBLM_R_X11Y106_SLICE_X14Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ffffff0f0fffff)
  ) CLBLM_R_X11Y106_SLICE_X14Y106_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(LIOB33_X0Y101_IOB_X0Y102_I),
.I3(LIOB33_X0Y101_IOB_X0Y101_I),
.I4(RIOB33_X105Y103_IOB_X1Y104_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y106_SLICE_X14Y106_AO5),
.O6(CLBLM_R_X11Y106_SLICE_X14Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y106_SLICE_X15Y106_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y106_SLICE_X15Y106_DO5),
.O6(CLBLM_R_X11Y106_SLICE_X15Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y106_SLICE_X15Y106_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y106_SLICE_X15Y106_CO5),
.O6(CLBLM_R_X11Y106_SLICE_X15Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y106_SLICE_X15Y106_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y106_SLICE_X15Y106_BO5),
.O6(CLBLM_R_X11Y106_SLICE_X15Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y106_SLICE_X15Y106_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y106_SLICE_X15Y106_AO5),
.O6(CLBLM_R_X11Y106_SLICE_X15Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y101_IOB_X0Y101_IBUF (
.I(LIOB33_X0Y101_IOB_X0Y101_IPAD),
.O(LIOB33_X0Y101_IOB_X0Y101_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y101_IOB_X0Y102_IBUF (
.I(LIOB33_X0Y101_IOB_X0Y102_IPAD),
.O(LIOB33_X0Y101_IOB_X0Y102_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y103_IOB_X0Y103_IBUF (
.I(LIOB33_X0Y103_IOB_X0Y103_IPAD),
.O(LIOB33_X0Y103_IOB_X0Y103_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y103_IOB_X0Y104_IBUF (
.I(LIOB33_X0Y103_IOB_X0Y104_IPAD),
.O(LIOB33_X0Y103_IOB_X0Y104_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y105_IOB_X0Y105_IBUF (
.I(LIOB33_X0Y105_IOB_X0Y105_IPAD),
.O(LIOB33_X0Y105_IOB_X0Y105_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y105_IOB_X0Y106_IBUF (
.I(LIOB33_X0Y105_IOB_X0Y106_IPAD),
.O(LIOB33_X0Y105_IOB_X0Y106_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y107_IOB_X0Y107_IBUF (
.I(LIOB33_X0Y107_IOB_X0Y107_IPAD),
.O(LIOB33_X0Y107_IOB_X0Y107_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y107_IOB_X0Y108_IBUF (
.I(LIOB33_X0Y107_IOB_X0Y108_IPAD),
.O(LIOB33_X0Y107_IOB_X0Y108_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y109_IOB_X0Y109_IBUF (
.I(LIOB33_X0Y109_IOB_X0Y109_IPAD),
.O(LIOB33_X0Y109_IOB_X0Y109_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y109_IOB_X0Y110_IBUF (
.I(LIOB33_X0Y109_IOB_X0Y110_IPAD),
.O(LIOB33_X0Y109_IOB_X0Y110_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y111_IOB_X0Y111_IBUF (
.I(LIOB33_X0Y111_IOB_X0Y111_IPAD),
.O(LIOB33_X0Y111_IOB_X0Y111_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y111_IOB_X0Y112_IBUF (
.I(LIOB33_X0Y111_IOB_X0Y112_IPAD),
.O(LIOB33_X0Y111_IOB_X0Y112_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y113_IOB_X0Y113_IBUF (
.I(LIOB33_X0Y113_IOB_X0Y113_IPAD),
.O(LIOB33_X0Y113_IOB_X0Y113_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y113_IOB_X0Y114_IBUF (
.I(LIOB33_X0Y113_IOB_X0Y114_IPAD),
.O(LIOB33_X0Y113_IOB_X0Y114_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y115_IOB_X0Y115_IBUF (
.I(LIOB33_X0Y115_IOB_X0Y115_IPAD),
.O(LIOB33_X0Y115_IOB_X0Y115_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y115_IOB_X0Y116_IBUF (
.I(LIOB33_X0Y115_IOB_X0Y116_IPAD),
.O(LIOB33_X0Y115_IOB_X0Y116_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y117_IOB_X0Y117_IBUF (
.I(LIOB33_X0Y117_IOB_X0Y117_IPAD),
.O(LIOB33_X0Y117_IOB_X0Y117_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y117_IOB_X0Y118_OBUF (
.I(CLBLL_L_X2Y114_SLICE_X0Y114_AO5),
.O(LIOB33_X0Y117_IOB_X0Y118_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y119_IOB_X0Y119_OBUF (
.I(CLBLL_L_X2Y114_SLICE_X0Y114_AO6),
.O(LIOB33_X0Y119_IOB_X0Y119_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y119_IOB_X0Y120_OBUF (
.I(CLBLL_L_X2Y113_SLICE_X0Y113_AO5),
.O(LIOB33_X0Y119_IOB_X0Y120_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y121_IOB_X0Y121_OBUF (
.I(CLBLL_L_X2Y113_SLICE_X0Y113_BO5),
.O(LIOB33_X0Y121_IOB_X0Y121_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y121_IOB_X0Y122_OBUF (
.I(CLBLL_L_X2Y113_SLICE_X1Y113_AO6),
.O(LIOB33_X0Y121_IOB_X0Y122_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y123_IOB_X0Y123_OBUF (
.I(CLBLL_L_X2Y113_SLICE_X1Y113_CO6),
.O(LIOB33_X0Y123_IOB_X0Y123_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y123_IOB_X0Y124_OBUF (
.I(CLBLM_R_X3Y112_SLICE_X2Y112_AO6),
.O(LIOB33_X0Y123_IOB_X0Y124_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y125_IOB_X0Y125_OBUF (
.I(CLBLM_R_X3Y111_SLICE_X3Y111_AO6),
.O(LIOB33_X0Y125_IOB_X0Y125_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y125_IOB_X0Y126_OBUF (
.I(CLBLM_R_X3Y111_SLICE_X2Y111_BO6),
.O(LIOB33_X0Y125_IOB_X0Y126_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y127_IOB_X0Y127_OBUF (
.I(CLBLL_L_X4Y110_SLICE_X4Y110_AO5),
.O(LIOB33_X0Y127_IOB_X0Y127_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y127_IOB_X0Y128_OBUF (
.I(CLBLL_L_X4Y107_SLICE_X4Y107_AO6),
.O(LIOB33_X0Y127_IOB_X0Y128_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y129_IOB_X0Y129_OBUF (
.I(CLBLM_R_X3Y110_SLICE_X3Y110_BO6),
.O(LIOB33_X0Y129_IOB_X0Y129_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y129_IOB_X0Y130_OBUF (
.I(CLBLL_L_X2Y114_SLICE_X0Y114_BO5),
.O(LIOB33_X0Y129_IOB_X0Y130_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y131_IOB_X0Y131_OBUF (
.I(CLBLM_R_X3Y110_SLICE_X2Y110_AO5),
.O(LIOB33_X0Y131_IOB_X0Y131_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y131_IOB_X0Y132_OBUF (
.I(CLBLM_R_X3Y110_SLICE_X2Y110_BO6),
.O(LIOB33_X0Y131_IOB_X0Y132_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y133_IOB_X0Y133_OBUF (
.I(CLBLM_R_X3Y110_SLICE_X2Y110_CO6),
.O(LIOB33_X0Y133_IOB_X0Y133_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y133_IOB_X0Y134_OBUF (
.I(1'b0),
.O(LIOB33_X0Y133_IOB_X0Y134_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y135_IOB_X0Y135_OBUF (
.I(CLBLM_R_X3Y107_SLICE_X2Y107_AO5),
.O(LIOB33_X0Y135_IOB_X0Y135_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y135_IOB_X0Y136_OBUF (
.I(CLBLM_R_X3Y107_SLICE_X2Y107_AO6),
.O(LIOB33_X0Y135_IOB_X0Y136_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y137_IOB_X0Y137_OBUF (
.I(CLBLL_L_X2Y109_SLICE_X1Y109_AO6),
.O(LIOB33_X0Y137_IOB_X0Y137_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y137_IOB_X0Y138_OBUF (
.I(CLBLL_L_X2Y108_SLICE_X1Y108_DO6),
.O(LIOB33_X0Y137_IOB_X0Y138_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y139_IOB_X0Y139_OBUF (
.I(CLBLL_L_X2Y107_SLICE_X1Y107_CO6),
.O(LIOB33_X0Y139_IOB_X0Y139_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y139_IOB_X0Y140_OBUF (
.I(CLBLL_L_X2Y105_SLICE_X1Y105_DO6),
.O(LIOB33_X0Y139_IOB_X0Y140_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y141_IOB_X0Y141_OBUF (
.I(CLBLL_L_X2Y105_SLICE_X0Y105_AO6),
.O(LIOB33_X0Y141_IOB_X0Y141_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y141_IOB_X0Y142_OBUF (
.I(CLBLL_L_X2Y105_SLICE_X0Y105_AO5),
.O(LIOB33_X0Y141_IOB_X0Y142_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y143_IOB_X0Y143_OBUF (
.I(CLBLL_L_X2Y106_SLICE_X0Y106_BO6),
.O(LIOB33_X0Y143_IOB_X0Y143_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y145_IOB_X0Y145_OBUF (
.I(CLBLM_R_X3Y104_SLICE_X3Y104_DO6),
.O(LIOB33_X0Y145_IOB_X0Y145_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y145_IOB_X0Y146_OBUF (
.I(CLBLM_R_X3Y104_SLICE_X3Y104_BO6),
.O(LIOB33_X0Y145_IOB_X0Y146_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y147_IOB_X0Y147_OBUF (
.I(CLBLL_L_X2Y108_SLICE_X0Y108_DO6),
.O(LIOB33_X0Y147_IOB_X0Y147_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y147_IOB_X0Y148_OBUF (
.I(CLBLL_L_X2Y108_SLICE_X0Y108_BO6),
.O(LIOB33_X0Y147_IOB_X0Y148_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_SING_X0Y100_IOB_X0Y100_IBUF (
.I(LIOB33_SING_X0Y100_IOB_X0Y100_IPAD),
.O(LIOB33_SING_X0Y100_IOB_X0Y100_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y149_IOB_X0Y149_OBUF (
.I(CLBLL_L_X2Y108_SLICE_X0Y108_CO6),
.O(LIOB33_SING_X0Y149_IOB_X0Y149_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y101_IOB_X1Y101_IBUF (
.I(RIOB33_X105Y101_IOB_X1Y101_IPAD),
.O(RIOB33_X105Y101_IOB_X1Y101_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y101_IOB_X1Y102_IBUF (
.I(RIOB33_X105Y101_IOB_X1Y102_IPAD),
.O(RIOB33_X105Y101_IOB_X1Y102_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y103_IOB_X1Y103_IBUF (
.I(RIOB33_X105Y103_IOB_X1Y103_IPAD),
.O(RIOB33_X105Y103_IOB_X1Y103_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y103_IOB_X1Y104_IBUF (
.I(RIOB33_X105Y103_IOB_X1Y104_IPAD),
.O(RIOB33_X105Y103_IOB_X1Y104_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y105_IOB_X1Y105_IBUF (
.I(RIOB33_X105Y105_IOB_X1Y105_IPAD),
.O(RIOB33_X105Y105_IOB_X1Y105_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y105_IOB_X1Y106_IBUF (
.I(RIOB33_X105Y105_IOB_X1Y106_IPAD),
.O(RIOB33_X105Y105_IOB_X1Y106_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y107_IOB_X1Y107_IBUF (
.I(RIOB33_X105Y107_IOB_X1Y107_IPAD),
.O(RIOB33_X105Y107_IOB_X1Y107_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y107_IOB_X1Y108_IBUF (
.I(RIOB33_X105Y107_IOB_X1Y108_IPAD),
.O(RIOB33_X105Y107_IOB_X1Y108_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y109_IOB_X1Y109_IBUF (
.I(RIOB33_X105Y109_IOB_X1Y109_IPAD),
.O(RIOB33_X105Y109_IOB_X1Y109_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y109_IOB_X1Y110_IBUF (
.I(RIOB33_X105Y109_IOB_X1Y110_IPAD),
.O(RIOB33_X105Y109_IOB_X1Y110_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y111_IOB_X1Y111_IBUF (
.I(RIOB33_X105Y111_IOB_X1Y111_IPAD),
.O(RIOB33_X105Y111_IOB_X1Y111_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y111_IOB_X1Y112_IBUF (
.I(RIOB33_X105Y111_IOB_X1Y112_IPAD),
.O(RIOB33_X105Y111_IOB_X1Y112_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y113_IOB_X1Y113_IBUF (
.I(RIOB33_X105Y113_IOB_X1Y113_IPAD),
.O(RIOB33_X105Y113_IOB_X1Y113_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_SING_X105Y100_IOB_X1Y100_IBUF (
.I(RIOB33_SING_X105Y100_IOB_X1Y100_IPAD),
.O(RIOB33_SING_X105Y100_IOB_X1Y100_I)
  );
  assign CLBLL_L_X2Y102_SLICE_X0Y102_A = CLBLL_L_X2Y102_SLICE_X0Y102_AO6;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_B = CLBLL_L_X2Y102_SLICE_X0Y102_BO6;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_C = CLBLL_L_X2Y102_SLICE_X0Y102_CO6;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_D = CLBLL_L_X2Y102_SLICE_X0Y102_DO6;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_A = CLBLL_L_X2Y102_SLICE_X1Y102_AO6;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_B = CLBLL_L_X2Y102_SLICE_X1Y102_BO6;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_C = CLBLL_L_X2Y102_SLICE_X1Y102_CO6;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_D = CLBLL_L_X2Y102_SLICE_X1Y102_DO6;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_A = CLBLL_L_X2Y103_SLICE_X0Y103_AO6;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_B = CLBLL_L_X2Y103_SLICE_X0Y103_BO6;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_C = CLBLL_L_X2Y103_SLICE_X0Y103_CO6;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_D = CLBLL_L_X2Y103_SLICE_X0Y103_DO6;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_A = CLBLL_L_X2Y103_SLICE_X1Y103_AO6;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_B = CLBLL_L_X2Y103_SLICE_X1Y103_BO6;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_C = CLBLL_L_X2Y103_SLICE_X1Y103_CO6;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_D = CLBLL_L_X2Y103_SLICE_X1Y103_DO6;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_AMUX = CLBLL_L_X2Y103_SLICE_X1Y103_AO5;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_A = CLBLL_L_X2Y104_SLICE_X0Y104_AO6;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_B = CLBLL_L_X2Y104_SLICE_X0Y104_BO6;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_C = CLBLL_L_X2Y104_SLICE_X0Y104_CO6;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_D = CLBLL_L_X2Y104_SLICE_X0Y104_DO6;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_AMUX = CLBLL_L_X2Y104_SLICE_X0Y104_AO5;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_BMUX = CLBLL_L_X2Y104_SLICE_X0Y104_BO6;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_DMUX = CLBLL_L_X2Y104_SLICE_X0Y104_DO6;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_A = CLBLL_L_X2Y104_SLICE_X1Y104_AO6;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_B = CLBLL_L_X2Y104_SLICE_X1Y104_BO6;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_C = CLBLL_L_X2Y104_SLICE_X1Y104_CO6;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_D = CLBLL_L_X2Y104_SLICE_X1Y104_DO6;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_AMUX = CLBLL_L_X2Y104_SLICE_X1Y104_AO5;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_A = CLBLL_L_X2Y105_SLICE_X0Y105_AO6;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_B = CLBLL_L_X2Y105_SLICE_X0Y105_BO6;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_C = CLBLL_L_X2Y105_SLICE_X0Y105_CO6;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_D = CLBLL_L_X2Y105_SLICE_X0Y105_DO6;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_AMUX = CLBLL_L_X2Y105_SLICE_X0Y105_AO5;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_BMUX = CLBLL_L_X2Y105_SLICE_X0Y105_BO5;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_CMUX = CLBLL_L_X2Y105_SLICE_X0Y105_CO6;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_A = CLBLL_L_X2Y105_SLICE_X1Y105_AO6;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_B = CLBLL_L_X2Y105_SLICE_X1Y105_BO6;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_C = CLBLL_L_X2Y105_SLICE_X1Y105_CO6;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_D = CLBLL_L_X2Y105_SLICE_X1Y105_DO6;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_AMUX = CLBLL_L_X2Y105_SLICE_X1Y105_AO5;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_A = CLBLL_L_X2Y106_SLICE_X0Y106_AO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_B = CLBLL_L_X2Y106_SLICE_X0Y106_BO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_C = CLBLL_L_X2Y106_SLICE_X0Y106_CO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_D = CLBLL_L_X2Y106_SLICE_X0Y106_DO6;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_A = CLBLL_L_X2Y106_SLICE_X1Y106_AO6;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_B = CLBLL_L_X2Y106_SLICE_X1Y106_BO6;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_C = CLBLL_L_X2Y106_SLICE_X1Y106_CO6;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_D = CLBLL_L_X2Y106_SLICE_X1Y106_DO6;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_AMUX = CLBLL_L_X2Y106_SLICE_X1Y106_AO5;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_BMUX = CLBLL_L_X2Y106_SLICE_X1Y106_BO6;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_A = CLBLL_L_X2Y107_SLICE_X0Y107_AO6;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_B = CLBLL_L_X2Y107_SLICE_X0Y107_BO6;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_C = CLBLL_L_X2Y107_SLICE_X0Y107_CO6;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_D = CLBLL_L_X2Y107_SLICE_X0Y107_DO6;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_A = CLBLL_L_X2Y107_SLICE_X1Y107_AO6;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_B = CLBLL_L_X2Y107_SLICE_X1Y107_BO6;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_C = CLBLL_L_X2Y107_SLICE_X1Y107_CO6;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_D = CLBLL_L_X2Y107_SLICE_X1Y107_DO6;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_A = CLBLL_L_X2Y108_SLICE_X0Y108_AO6;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_B = CLBLL_L_X2Y108_SLICE_X0Y108_BO6;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_C = CLBLL_L_X2Y108_SLICE_X0Y108_CO6;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_D = CLBLL_L_X2Y108_SLICE_X0Y108_DO6;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_AMUX = CLBLL_L_X2Y108_SLICE_X0Y108_AO5;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_A = CLBLL_L_X2Y108_SLICE_X1Y108_AO6;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_B = CLBLL_L_X2Y108_SLICE_X1Y108_BO6;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_C = CLBLL_L_X2Y108_SLICE_X1Y108_CO6;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_D = CLBLL_L_X2Y108_SLICE_X1Y108_DO6;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_A = CLBLL_L_X2Y109_SLICE_X0Y109_AO6;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_B = CLBLL_L_X2Y109_SLICE_X0Y109_BO6;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_C = CLBLL_L_X2Y109_SLICE_X0Y109_CO6;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_D = CLBLL_L_X2Y109_SLICE_X0Y109_DO6;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_A = CLBLL_L_X2Y109_SLICE_X1Y109_AO6;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_B = CLBLL_L_X2Y109_SLICE_X1Y109_BO6;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_C = CLBLL_L_X2Y109_SLICE_X1Y109_CO6;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_D = CLBLL_L_X2Y109_SLICE_X1Y109_DO6;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_A = CLBLL_L_X2Y112_SLICE_X0Y112_AO6;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_B = CLBLL_L_X2Y112_SLICE_X0Y112_BO6;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_C = CLBLL_L_X2Y112_SLICE_X0Y112_CO6;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_D = CLBLL_L_X2Y112_SLICE_X0Y112_DO6;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_A = CLBLL_L_X2Y112_SLICE_X1Y112_AO6;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_B = CLBLL_L_X2Y112_SLICE_X1Y112_BO6;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_C = CLBLL_L_X2Y112_SLICE_X1Y112_CO6;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_D = CLBLL_L_X2Y112_SLICE_X1Y112_DO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_A = CLBLL_L_X2Y113_SLICE_X0Y113_AO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_B = CLBLL_L_X2Y113_SLICE_X0Y113_BO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_C = CLBLL_L_X2Y113_SLICE_X0Y113_CO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_D = CLBLL_L_X2Y113_SLICE_X0Y113_DO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_AMUX = CLBLL_L_X2Y113_SLICE_X0Y113_AO5;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_BMUX = CLBLL_L_X2Y113_SLICE_X0Y113_BO5;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_A = CLBLL_L_X2Y113_SLICE_X1Y113_AO6;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_B = CLBLL_L_X2Y113_SLICE_X1Y113_BO6;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_C = CLBLL_L_X2Y113_SLICE_X1Y113_CO6;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_D = CLBLL_L_X2Y113_SLICE_X1Y113_DO6;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_AMUX = CLBLL_L_X2Y113_SLICE_X1Y113_AO5;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_A = CLBLL_L_X2Y114_SLICE_X0Y114_AO6;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_B = CLBLL_L_X2Y114_SLICE_X0Y114_BO6;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_C = CLBLL_L_X2Y114_SLICE_X0Y114_CO6;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_D = CLBLL_L_X2Y114_SLICE_X0Y114_DO6;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_AMUX = CLBLL_L_X2Y114_SLICE_X0Y114_AO5;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_BMUX = CLBLL_L_X2Y114_SLICE_X0Y114_BO5;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_A = CLBLL_L_X2Y114_SLICE_X1Y114_AO6;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_B = CLBLL_L_X2Y114_SLICE_X1Y114_BO6;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_C = CLBLL_L_X2Y114_SLICE_X1Y114_CO6;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_D = CLBLL_L_X2Y114_SLICE_X1Y114_DO6;
  assign CLBLL_L_X4Y100_SLICE_X4Y100_A = CLBLL_L_X4Y100_SLICE_X4Y100_AO6;
  assign CLBLL_L_X4Y100_SLICE_X4Y100_B = CLBLL_L_X4Y100_SLICE_X4Y100_BO6;
  assign CLBLL_L_X4Y100_SLICE_X4Y100_C = CLBLL_L_X4Y100_SLICE_X4Y100_CO6;
  assign CLBLL_L_X4Y100_SLICE_X4Y100_D = CLBLL_L_X4Y100_SLICE_X4Y100_DO6;
  assign CLBLL_L_X4Y100_SLICE_X4Y100_AMUX = CLBLL_L_X4Y100_SLICE_X4Y100_AO5;
  assign CLBLL_L_X4Y100_SLICE_X4Y100_CMUX = CLBLL_L_X4Y100_SLICE_X4Y100_CO6;
  assign CLBLL_L_X4Y100_SLICE_X5Y100_A = CLBLL_L_X4Y100_SLICE_X5Y100_AO6;
  assign CLBLL_L_X4Y100_SLICE_X5Y100_B = CLBLL_L_X4Y100_SLICE_X5Y100_BO6;
  assign CLBLL_L_X4Y100_SLICE_X5Y100_C = CLBLL_L_X4Y100_SLICE_X5Y100_CO6;
  assign CLBLL_L_X4Y100_SLICE_X5Y100_D = CLBLL_L_X4Y100_SLICE_X5Y100_DO6;
  assign CLBLL_L_X4Y101_SLICE_X4Y101_A = CLBLL_L_X4Y101_SLICE_X4Y101_AO6;
  assign CLBLL_L_X4Y101_SLICE_X4Y101_B = CLBLL_L_X4Y101_SLICE_X4Y101_BO6;
  assign CLBLL_L_X4Y101_SLICE_X4Y101_C = CLBLL_L_X4Y101_SLICE_X4Y101_CO6;
  assign CLBLL_L_X4Y101_SLICE_X4Y101_D = CLBLL_L_X4Y101_SLICE_X4Y101_DO6;
  assign CLBLL_L_X4Y101_SLICE_X5Y101_A = CLBLL_L_X4Y101_SLICE_X5Y101_AO6;
  assign CLBLL_L_X4Y101_SLICE_X5Y101_B = CLBLL_L_X4Y101_SLICE_X5Y101_BO6;
  assign CLBLL_L_X4Y101_SLICE_X5Y101_C = CLBLL_L_X4Y101_SLICE_X5Y101_CO6;
  assign CLBLL_L_X4Y101_SLICE_X5Y101_D = CLBLL_L_X4Y101_SLICE_X5Y101_DO6;
  assign CLBLL_L_X4Y101_SLICE_X5Y101_AMUX = CLBLL_L_X4Y101_SLICE_X5Y101_AO5;
  assign CLBLL_L_X4Y101_SLICE_X5Y101_BMUX = CLBLL_L_X4Y101_SLICE_X5Y101_BO5;
  assign CLBLL_L_X4Y101_SLICE_X5Y101_CMUX = CLBLL_L_X4Y101_SLICE_X5Y101_CO5;
  assign CLBLL_L_X4Y102_SLICE_X4Y102_A = CLBLL_L_X4Y102_SLICE_X4Y102_AO6;
  assign CLBLL_L_X4Y102_SLICE_X4Y102_B = CLBLL_L_X4Y102_SLICE_X4Y102_BO6;
  assign CLBLL_L_X4Y102_SLICE_X4Y102_C = CLBLL_L_X4Y102_SLICE_X4Y102_CO6;
  assign CLBLL_L_X4Y102_SLICE_X4Y102_D = CLBLL_L_X4Y102_SLICE_X4Y102_DO6;
  assign CLBLL_L_X4Y102_SLICE_X4Y102_AMUX = CLBLL_L_X4Y102_SLICE_X4Y102_AO5;
  assign CLBLL_L_X4Y102_SLICE_X4Y102_BMUX = CLBLL_L_X4Y102_SLICE_X4Y102_BO5;
  assign CLBLL_L_X4Y102_SLICE_X5Y102_A = CLBLL_L_X4Y102_SLICE_X5Y102_AO6;
  assign CLBLL_L_X4Y102_SLICE_X5Y102_B = CLBLL_L_X4Y102_SLICE_X5Y102_BO6;
  assign CLBLL_L_X4Y102_SLICE_X5Y102_C = CLBLL_L_X4Y102_SLICE_X5Y102_CO6;
  assign CLBLL_L_X4Y102_SLICE_X5Y102_D = CLBLL_L_X4Y102_SLICE_X5Y102_DO6;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_A = CLBLL_L_X4Y103_SLICE_X4Y103_AO6;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_B = CLBLL_L_X4Y103_SLICE_X4Y103_BO6;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_C = CLBLL_L_X4Y103_SLICE_X4Y103_CO6;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_D = CLBLL_L_X4Y103_SLICE_X4Y103_DO6;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_A = CLBLL_L_X4Y103_SLICE_X5Y103_AO6;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_B = CLBLL_L_X4Y103_SLICE_X5Y103_BO6;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_C = CLBLL_L_X4Y103_SLICE_X5Y103_CO6;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_D = CLBLL_L_X4Y103_SLICE_X5Y103_DO6;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_AMUX = CLBLL_L_X4Y103_SLICE_X5Y103_AO5;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_BMUX = CLBLL_L_X4Y103_SLICE_X5Y103_BO5;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_CMUX = CLBLL_L_X4Y103_SLICE_X5Y103_CO6;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_A = CLBLL_L_X4Y104_SLICE_X4Y104_AO6;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_B = CLBLL_L_X4Y104_SLICE_X4Y104_BO6;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_C = CLBLL_L_X4Y104_SLICE_X4Y104_CO6;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_D = CLBLL_L_X4Y104_SLICE_X4Y104_DO6;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_AMUX = CLBLL_L_X4Y104_SLICE_X4Y104_AO5;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_BMUX = CLBLL_L_X4Y104_SLICE_X4Y104_BO5;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_CMUX = CLBLL_L_X4Y104_SLICE_X4Y104_CO5;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_A = CLBLL_L_X4Y104_SLICE_X5Y104_AO6;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_B = CLBLL_L_X4Y104_SLICE_X5Y104_BO6;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_C = CLBLL_L_X4Y104_SLICE_X5Y104_CO6;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_D = CLBLL_L_X4Y104_SLICE_X5Y104_DO6;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_AMUX = CLBLL_L_X4Y104_SLICE_X5Y104_AO5;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_BMUX = CLBLL_L_X4Y104_SLICE_X5Y104_BO5;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_A = CLBLL_L_X4Y105_SLICE_X4Y105_AO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_B = CLBLL_L_X4Y105_SLICE_X4Y105_BO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_C = CLBLL_L_X4Y105_SLICE_X4Y105_CO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_D = CLBLL_L_X4Y105_SLICE_X4Y105_DO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_AMUX = CLBLL_L_X4Y105_SLICE_X4Y105_AO5;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_A = CLBLL_L_X4Y105_SLICE_X5Y105_AO6;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_B = CLBLL_L_X4Y105_SLICE_X5Y105_BO6;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_C = CLBLL_L_X4Y105_SLICE_X5Y105_CO6;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_D = CLBLL_L_X4Y105_SLICE_X5Y105_DO6;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_BMUX = CLBLL_L_X4Y105_SLICE_X5Y105_BO6;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_CMUX = CLBLL_L_X4Y105_SLICE_X5Y105_CO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_A = CLBLL_L_X4Y106_SLICE_X4Y106_AO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_B = CLBLL_L_X4Y106_SLICE_X4Y106_BO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_C = CLBLL_L_X4Y106_SLICE_X4Y106_CO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_D = CLBLL_L_X4Y106_SLICE_X4Y106_DO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_AMUX = CLBLL_L_X4Y106_SLICE_X4Y106_AO5;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_A = CLBLL_L_X4Y106_SLICE_X5Y106_AO6;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_B = CLBLL_L_X4Y106_SLICE_X5Y106_BO6;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_C = CLBLL_L_X4Y106_SLICE_X5Y106_CO6;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_D = CLBLL_L_X4Y106_SLICE_X5Y106_DO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_A = CLBLL_L_X4Y107_SLICE_X4Y107_AO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_B = CLBLL_L_X4Y107_SLICE_X4Y107_BO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_C = CLBLL_L_X4Y107_SLICE_X4Y107_CO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_D = CLBLL_L_X4Y107_SLICE_X4Y107_DO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_AMUX = CLBLL_L_X4Y107_SLICE_X4Y107_AO5;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_A = CLBLL_L_X4Y107_SLICE_X5Y107_AO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_B = CLBLL_L_X4Y107_SLICE_X5Y107_BO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_C = CLBLL_L_X4Y107_SLICE_X5Y107_CO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_D = CLBLL_L_X4Y107_SLICE_X5Y107_DO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_AMUX = CLBLL_L_X4Y107_SLICE_X5Y107_AO5;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_A = CLBLL_L_X4Y108_SLICE_X4Y108_AO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_B = CLBLL_L_X4Y108_SLICE_X4Y108_BO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_C = CLBLL_L_X4Y108_SLICE_X4Y108_CO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_D = CLBLL_L_X4Y108_SLICE_X4Y108_DO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_A = CLBLL_L_X4Y108_SLICE_X5Y108_AO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_B = CLBLL_L_X4Y108_SLICE_X5Y108_BO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_C = CLBLL_L_X4Y108_SLICE_X5Y108_CO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_D = CLBLL_L_X4Y108_SLICE_X5Y108_DO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_BMUX = CLBLL_L_X4Y108_SLICE_X5Y108_BO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A = CLBLL_L_X4Y109_SLICE_X4Y109_AO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B = CLBLL_L_X4Y109_SLICE_X4Y109_BO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C = CLBLL_L_X4Y109_SLICE_X4Y109_CO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D = CLBLL_L_X4Y109_SLICE_X4Y109_DO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A = CLBLL_L_X4Y109_SLICE_X5Y109_AO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B = CLBLL_L_X4Y109_SLICE_X5Y109_BO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C = CLBLL_L_X4Y109_SLICE_X5Y109_CO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D = CLBLL_L_X4Y109_SLICE_X5Y109_DO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_AMUX = CLBLL_L_X4Y109_SLICE_X5Y109_AO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_DMUX = CLBLL_L_X4Y109_SLICE_X5Y109_DO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_A = CLBLL_L_X4Y110_SLICE_X4Y110_AO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_B = CLBLL_L_X4Y110_SLICE_X4Y110_BO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_C = CLBLL_L_X4Y110_SLICE_X4Y110_CO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_D = CLBLL_L_X4Y110_SLICE_X4Y110_DO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_AMUX = CLBLL_L_X4Y110_SLICE_X4Y110_AO5;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_A = CLBLL_L_X4Y110_SLICE_X5Y110_AO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_B = CLBLL_L_X4Y110_SLICE_X5Y110_BO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_C = CLBLL_L_X4Y110_SLICE_X5Y110_CO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_D = CLBLL_L_X4Y110_SLICE_X5Y110_DO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_AMUX = CLBLL_L_X4Y110_SLICE_X5Y110_AO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_CMUX = CLBLL_L_X4Y110_SLICE_X5Y110_CO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_A = CLBLL_L_X4Y111_SLICE_X4Y111_AO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_B = CLBLL_L_X4Y111_SLICE_X4Y111_BO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_C = CLBLL_L_X4Y111_SLICE_X4Y111_CO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_D = CLBLL_L_X4Y111_SLICE_X4Y111_DO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_A = CLBLL_L_X4Y111_SLICE_X5Y111_AO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_B = CLBLL_L_X4Y111_SLICE_X5Y111_BO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_C = CLBLL_L_X4Y111_SLICE_X5Y111_CO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_D = CLBLL_L_X4Y111_SLICE_X5Y111_DO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_BMUX = CLBLL_L_X4Y111_SLICE_X5Y111_BO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_A = CLBLL_L_X4Y112_SLICE_X4Y112_AO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_B = CLBLL_L_X4Y112_SLICE_X4Y112_BO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_C = CLBLL_L_X4Y112_SLICE_X4Y112_CO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_D = CLBLL_L_X4Y112_SLICE_X4Y112_DO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_AMUX = CLBLL_L_X4Y112_SLICE_X4Y112_AO5;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_A = CLBLL_L_X4Y112_SLICE_X5Y112_AO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_B = CLBLL_L_X4Y112_SLICE_X5Y112_BO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_C = CLBLL_L_X4Y112_SLICE_X5Y112_CO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_D = CLBLL_L_X4Y112_SLICE_X5Y112_DO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_DMUX = CLBLL_L_X4Y112_SLICE_X5Y112_DO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A = CLBLL_L_X4Y113_SLICE_X4Y113_AO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B = CLBLL_L_X4Y113_SLICE_X4Y113_BO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C = CLBLL_L_X4Y113_SLICE_X4Y113_CO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D = CLBLL_L_X4Y113_SLICE_X4Y113_DO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A = CLBLL_L_X4Y113_SLICE_X5Y113_AO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B = CLBLL_L_X4Y113_SLICE_X5Y113_BO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C = CLBLL_L_X4Y113_SLICE_X5Y113_CO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D = CLBLL_L_X4Y113_SLICE_X5Y113_DO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_AMUX = CLBLL_L_X4Y113_SLICE_X5Y113_AO5;
  assign CLBLM_L_X8Y100_SLICE_X10Y100_A = CLBLM_L_X8Y100_SLICE_X10Y100_AO6;
  assign CLBLM_L_X8Y100_SLICE_X10Y100_B = CLBLM_L_X8Y100_SLICE_X10Y100_BO6;
  assign CLBLM_L_X8Y100_SLICE_X10Y100_C = CLBLM_L_X8Y100_SLICE_X10Y100_CO6;
  assign CLBLM_L_X8Y100_SLICE_X10Y100_D = CLBLM_L_X8Y100_SLICE_X10Y100_DO6;
  assign CLBLM_L_X8Y100_SLICE_X10Y100_AMUX = CLBLM_L_X8Y100_SLICE_X10Y100_AO5;
  assign CLBLM_L_X8Y100_SLICE_X11Y100_A = CLBLM_L_X8Y100_SLICE_X11Y100_AO6;
  assign CLBLM_L_X8Y100_SLICE_X11Y100_B = CLBLM_L_X8Y100_SLICE_X11Y100_BO6;
  assign CLBLM_L_X8Y100_SLICE_X11Y100_C = CLBLM_L_X8Y100_SLICE_X11Y100_CO6;
  assign CLBLM_L_X8Y100_SLICE_X11Y100_D = CLBLM_L_X8Y100_SLICE_X11Y100_DO6;
  assign CLBLM_L_X8Y100_SLICE_X11Y100_DMUX = CLBLM_L_X8Y100_SLICE_X11Y100_DO6;
  assign CLBLM_L_X8Y101_SLICE_X10Y101_A = CLBLM_L_X8Y101_SLICE_X10Y101_AO6;
  assign CLBLM_L_X8Y101_SLICE_X10Y101_B = CLBLM_L_X8Y101_SLICE_X10Y101_BO6;
  assign CLBLM_L_X8Y101_SLICE_X10Y101_C = CLBLM_L_X8Y101_SLICE_X10Y101_CO6;
  assign CLBLM_L_X8Y101_SLICE_X10Y101_D = CLBLM_L_X8Y101_SLICE_X10Y101_DO6;
  assign CLBLM_L_X8Y101_SLICE_X11Y101_A = CLBLM_L_X8Y101_SLICE_X11Y101_AO6;
  assign CLBLM_L_X8Y101_SLICE_X11Y101_B = CLBLM_L_X8Y101_SLICE_X11Y101_BO6;
  assign CLBLM_L_X8Y101_SLICE_X11Y101_C = CLBLM_L_X8Y101_SLICE_X11Y101_CO6;
  assign CLBLM_L_X8Y101_SLICE_X11Y101_D = CLBLM_L_X8Y101_SLICE_X11Y101_DO6;
  assign CLBLM_L_X8Y101_SLICE_X11Y101_AMUX = CLBLM_L_X8Y101_SLICE_X11Y101_AO5;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_A = CLBLM_L_X8Y102_SLICE_X10Y102_AO6;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_B = CLBLM_L_X8Y102_SLICE_X10Y102_BO6;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_C = CLBLM_L_X8Y102_SLICE_X10Y102_CO6;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_D = CLBLM_L_X8Y102_SLICE_X10Y102_DO6;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_AMUX = CLBLM_L_X8Y102_SLICE_X10Y102_AO5;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_A = CLBLM_L_X8Y102_SLICE_X11Y102_AO6;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_B = CLBLM_L_X8Y102_SLICE_X11Y102_BO6;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_C = CLBLM_L_X8Y102_SLICE_X11Y102_CO6;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_D = CLBLM_L_X8Y102_SLICE_X11Y102_DO6;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_CMUX = CLBLM_L_X8Y102_SLICE_X11Y102_CO6;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_A = CLBLM_L_X8Y103_SLICE_X10Y103_AO6;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_B = CLBLM_L_X8Y103_SLICE_X10Y103_BO6;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_C = CLBLM_L_X8Y103_SLICE_X10Y103_CO6;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_D = CLBLM_L_X8Y103_SLICE_X10Y103_DO6;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_AMUX = CLBLM_L_X8Y103_SLICE_X10Y103_AO5;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_A = CLBLM_L_X8Y103_SLICE_X11Y103_AO6;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_B = CLBLM_L_X8Y103_SLICE_X11Y103_BO6;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_C = CLBLM_L_X8Y103_SLICE_X11Y103_CO6;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_D = CLBLM_L_X8Y103_SLICE_X11Y103_DO6;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_AMUX = CLBLM_L_X8Y103_SLICE_X11Y103_AO5;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_A = CLBLM_L_X8Y104_SLICE_X10Y104_AO6;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_B = CLBLM_L_X8Y104_SLICE_X10Y104_BO6;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_C = CLBLM_L_X8Y104_SLICE_X10Y104_CO6;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_D = CLBLM_L_X8Y104_SLICE_X10Y104_DO6;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_AMUX = CLBLM_L_X8Y104_SLICE_X10Y104_AO5;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_A = CLBLM_L_X8Y104_SLICE_X11Y104_AO6;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_B = CLBLM_L_X8Y104_SLICE_X11Y104_BO6;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_C = CLBLM_L_X8Y104_SLICE_X11Y104_CO6;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_D = CLBLM_L_X8Y104_SLICE_X11Y104_DO6;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_A = CLBLM_L_X8Y105_SLICE_X10Y105_AO6;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_B = CLBLM_L_X8Y105_SLICE_X10Y105_BO6;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_C = CLBLM_L_X8Y105_SLICE_X10Y105_CO6;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_D = CLBLM_L_X8Y105_SLICE_X10Y105_DO6;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_AMUX = CLBLM_L_X8Y105_SLICE_X10Y105_AO5;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_A = CLBLM_L_X8Y105_SLICE_X11Y105_AO6;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_B = CLBLM_L_X8Y105_SLICE_X11Y105_BO6;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_C = CLBLM_L_X8Y105_SLICE_X11Y105_CO6;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_D = CLBLM_L_X8Y105_SLICE_X11Y105_DO6;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_BMUX = CLBLM_L_X8Y105_SLICE_X11Y105_BO6;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_DMUX = CLBLM_L_X8Y105_SLICE_X11Y105_DO6;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_A = CLBLM_L_X8Y106_SLICE_X10Y106_AO6;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_B = CLBLM_L_X8Y106_SLICE_X10Y106_BO6;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_C = CLBLM_L_X8Y106_SLICE_X10Y106_CO6;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_D = CLBLM_L_X8Y106_SLICE_X10Y106_DO6;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_AMUX = CLBLM_L_X8Y106_SLICE_X10Y106_AO5;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_A = CLBLM_L_X8Y106_SLICE_X11Y106_AO6;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_B = CLBLM_L_X8Y106_SLICE_X11Y106_BO6;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_C = CLBLM_L_X8Y106_SLICE_X11Y106_CO6;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_D = CLBLM_L_X8Y106_SLICE_X11Y106_DO6;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_AMUX = CLBLM_L_X8Y106_SLICE_X11Y106_AO5;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_A = CLBLM_L_X8Y107_SLICE_X10Y107_AO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_B = CLBLM_L_X8Y107_SLICE_X10Y107_BO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_C = CLBLM_L_X8Y107_SLICE_X10Y107_CO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_D = CLBLM_L_X8Y107_SLICE_X10Y107_DO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_AMUX = CLBLM_L_X8Y107_SLICE_X10Y107_AO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_A = CLBLM_L_X8Y107_SLICE_X11Y107_AO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_B = CLBLM_L_X8Y107_SLICE_X11Y107_BO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_C = CLBLM_L_X8Y107_SLICE_X11Y107_CO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_D = CLBLM_L_X8Y107_SLICE_X11Y107_DO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_A = CLBLM_L_X8Y108_SLICE_X10Y108_AO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_B = CLBLM_L_X8Y108_SLICE_X10Y108_BO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_C = CLBLM_L_X8Y108_SLICE_X10Y108_CO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_D = CLBLM_L_X8Y108_SLICE_X10Y108_DO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_AMUX = CLBLM_L_X8Y108_SLICE_X10Y108_AO5;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_A = CLBLM_L_X8Y108_SLICE_X11Y108_AO6;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_B = CLBLM_L_X8Y108_SLICE_X11Y108_BO6;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_C = CLBLM_L_X8Y108_SLICE_X11Y108_CO6;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_D = CLBLM_L_X8Y108_SLICE_X11Y108_DO6;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_A = CLBLM_L_X8Y109_SLICE_X10Y109_AO6;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_B = CLBLM_L_X8Y109_SLICE_X10Y109_BO6;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_C = CLBLM_L_X8Y109_SLICE_X10Y109_CO6;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_D = CLBLM_L_X8Y109_SLICE_X10Y109_DO6;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_AMUX = CLBLM_L_X8Y109_SLICE_X10Y109_AO5;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_CMUX = CLBLM_L_X8Y109_SLICE_X10Y109_CO6;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_A = CLBLM_L_X8Y109_SLICE_X11Y109_AO6;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_B = CLBLM_L_X8Y109_SLICE_X11Y109_BO6;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_C = CLBLM_L_X8Y109_SLICE_X11Y109_CO6;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_D = CLBLM_L_X8Y109_SLICE_X11Y109_DO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_A = CLBLM_L_X8Y110_SLICE_X10Y110_AO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_B = CLBLM_L_X8Y110_SLICE_X10Y110_BO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_C = CLBLM_L_X8Y110_SLICE_X10Y110_CO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_D = CLBLM_L_X8Y110_SLICE_X10Y110_DO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_A = CLBLM_L_X8Y110_SLICE_X11Y110_AO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_B = CLBLM_L_X8Y110_SLICE_X11Y110_BO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_C = CLBLM_L_X8Y110_SLICE_X11Y110_CO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_D = CLBLM_L_X8Y110_SLICE_X11Y110_DO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_AMUX = CLBLM_L_X8Y110_SLICE_X11Y110_AO5;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_A = CLBLM_L_X8Y111_SLICE_X10Y111_AO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_B = CLBLM_L_X8Y111_SLICE_X10Y111_BO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_C = CLBLM_L_X8Y111_SLICE_X10Y111_CO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_D = CLBLM_L_X8Y111_SLICE_X10Y111_DO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_A = CLBLM_L_X8Y111_SLICE_X11Y111_AO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_B = CLBLM_L_X8Y111_SLICE_X11Y111_BO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_C = CLBLM_L_X8Y111_SLICE_X11Y111_CO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_D = CLBLM_L_X8Y111_SLICE_X11Y111_DO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_A = CLBLM_L_X8Y112_SLICE_X10Y112_AO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_B = CLBLM_L_X8Y112_SLICE_X10Y112_BO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_C = CLBLM_L_X8Y112_SLICE_X10Y112_CO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_D = CLBLM_L_X8Y112_SLICE_X10Y112_DO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_AMUX = CLBLM_L_X8Y112_SLICE_X10Y112_AO5;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_A = CLBLM_L_X8Y112_SLICE_X11Y112_AO6;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_B = CLBLM_L_X8Y112_SLICE_X11Y112_BO6;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_C = CLBLM_L_X8Y112_SLICE_X11Y112_CO6;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_D = CLBLM_L_X8Y112_SLICE_X11Y112_DO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_A = CLBLM_L_X8Y113_SLICE_X10Y113_AO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_B = CLBLM_L_X8Y113_SLICE_X10Y113_BO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_C = CLBLM_L_X8Y113_SLICE_X10Y113_CO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_D = CLBLM_L_X8Y113_SLICE_X10Y113_DO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_A = CLBLM_L_X8Y113_SLICE_X11Y113_AO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_B = CLBLM_L_X8Y113_SLICE_X11Y113_BO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_C = CLBLM_L_X8Y113_SLICE_X11Y113_CO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_D = CLBLM_L_X8Y113_SLICE_X11Y113_DO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_AMUX = CLBLM_L_X8Y113_SLICE_X11Y113_AO5;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_A = CLBLM_L_X10Y102_SLICE_X12Y102_AO6;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_B = CLBLM_L_X10Y102_SLICE_X12Y102_BO6;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_C = CLBLM_L_X10Y102_SLICE_X12Y102_CO6;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_D = CLBLM_L_X10Y102_SLICE_X12Y102_DO6;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_AMUX = CLBLM_L_X10Y102_SLICE_X12Y102_AO5;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_A = CLBLM_L_X10Y102_SLICE_X13Y102_AO6;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_B = CLBLM_L_X10Y102_SLICE_X13Y102_BO6;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_C = CLBLM_L_X10Y102_SLICE_X13Y102_CO6;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_D = CLBLM_L_X10Y102_SLICE_X13Y102_DO6;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_A = CLBLM_L_X10Y103_SLICE_X12Y103_AO6;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_B = CLBLM_L_X10Y103_SLICE_X12Y103_BO6;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_C = CLBLM_L_X10Y103_SLICE_X12Y103_CO6;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_D = CLBLM_L_X10Y103_SLICE_X12Y103_DO6;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_AMUX = CLBLM_L_X10Y103_SLICE_X12Y103_AO5;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_A = CLBLM_L_X10Y103_SLICE_X13Y103_AO6;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_B = CLBLM_L_X10Y103_SLICE_X13Y103_BO6;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_C = CLBLM_L_X10Y103_SLICE_X13Y103_CO6;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_D = CLBLM_L_X10Y103_SLICE_X13Y103_DO6;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_BMUX = CLBLM_L_X10Y103_SLICE_X13Y103_BO6;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_CMUX = CLBLM_L_X10Y103_SLICE_X13Y103_CO6;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_A = CLBLM_L_X10Y104_SLICE_X12Y104_AO6;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_B = CLBLM_L_X10Y104_SLICE_X12Y104_BO6;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_C = CLBLM_L_X10Y104_SLICE_X12Y104_CO6;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_D = CLBLM_L_X10Y104_SLICE_X12Y104_DO6;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_AMUX = CLBLM_L_X10Y104_SLICE_X12Y104_AO5;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_A = CLBLM_L_X10Y104_SLICE_X13Y104_AO6;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_B = CLBLM_L_X10Y104_SLICE_X13Y104_BO6;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_C = CLBLM_L_X10Y104_SLICE_X13Y104_CO6;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_D = CLBLM_L_X10Y104_SLICE_X13Y104_DO6;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_A = CLBLM_L_X10Y105_SLICE_X12Y105_AO6;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_B = CLBLM_L_X10Y105_SLICE_X12Y105_BO6;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_C = CLBLM_L_X10Y105_SLICE_X12Y105_CO6;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_D = CLBLM_L_X10Y105_SLICE_X12Y105_DO6;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_A = CLBLM_L_X10Y105_SLICE_X13Y105_AO6;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_B = CLBLM_L_X10Y105_SLICE_X13Y105_BO6;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_C = CLBLM_L_X10Y105_SLICE_X13Y105_CO6;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_D = CLBLM_L_X10Y105_SLICE_X13Y105_DO6;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_AMUX = CLBLM_L_X10Y105_SLICE_X13Y105_AO6;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_A = CLBLM_L_X10Y106_SLICE_X12Y106_AO6;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_B = CLBLM_L_X10Y106_SLICE_X12Y106_BO6;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_C = CLBLM_L_X10Y106_SLICE_X12Y106_CO6;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_D = CLBLM_L_X10Y106_SLICE_X12Y106_DO6;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_AMUX = CLBLM_L_X10Y106_SLICE_X12Y106_AO5;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_A = CLBLM_L_X10Y106_SLICE_X13Y106_AO6;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_B = CLBLM_L_X10Y106_SLICE_X13Y106_BO6;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_C = CLBLM_L_X10Y106_SLICE_X13Y106_CO6;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_D = CLBLM_L_X10Y106_SLICE_X13Y106_DO6;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_AMUX = CLBLM_L_X10Y106_SLICE_X13Y106_AO5;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_A = CLBLM_L_X10Y107_SLICE_X12Y107_AO6;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_B = CLBLM_L_X10Y107_SLICE_X12Y107_BO6;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_C = CLBLM_L_X10Y107_SLICE_X12Y107_CO6;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_D = CLBLM_L_X10Y107_SLICE_X12Y107_DO6;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_AMUX = CLBLM_L_X10Y107_SLICE_X12Y107_AO5;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_A = CLBLM_L_X10Y107_SLICE_X13Y107_AO6;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_B = CLBLM_L_X10Y107_SLICE_X13Y107_BO6;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_C = CLBLM_L_X10Y107_SLICE_X13Y107_CO6;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_D = CLBLM_L_X10Y107_SLICE_X13Y107_DO6;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_BMUX = CLBLM_L_X10Y107_SLICE_X13Y107_BO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_A = CLBLM_L_X10Y108_SLICE_X12Y108_AO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_B = CLBLM_L_X10Y108_SLICE_X12Y108_BO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_C = CLBLM_L_X10Y108_SLICE_X12Y108_CO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_D = CLBLM_L_X10Y108_SLICE_X12Y108_DO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_AMUX = CLBLM_L_X10Y108_SLICE_X12Y108_AO5;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_A = CLBLM_L_X10Y108_SLICE_X13Y108_AO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_B = CLBLM_L_X10Y108_SLICE_X13Y108_BO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_C = CLBLM_L_X10Y108_SLICE_X13Y108_CO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_D = CLBLM_L_X10Y108_SLICE_X13Y108_DO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_AMUX = CLBLM_L_X10Y108_SLICE_X13Y108_AO5;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_A = CLBLM_L_X10Y109_SLICE_X12Y109_AO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_B = CLBLM_L_X10Y109_SLICE_X12Y109_BO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_C = CLBLM_L_X10Y109_SLICE_X12Y109_CO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_D = CLBLM_L_X10Y109_SLICE_X12Y109_DO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_AMUX = CLBLM_L_X10Y109_SLICE_X12Y109_AO5;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_A = CLBLM_L_X10Y109_SLICE_X13Y109_AO6;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_B = CLBLM_L_X10Y109_SLICE_X13Y109_BO6;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_C = CLBLM_L_X10Y109_SLICE_X13Y109_CO6;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_D = CLBLM_L_X10Y109_SLICE_X13Y109_DO6;
  assign CLBLM_R_X3Y100_SLICE_X2Y100_A = CLBLM_R_X3Y100_SLICE_X2Y100_AO6;
  assign CLBLM_R_X3Y100_SLICE_X2Y100_B = CLBLM_R_X3Y100_SLICE_X2Y100_BO6;
  assign CLBLM_R_X3Y100_SLICE_X2Y100_C = CLBLM_R_X3Y100_SLICE_X2Y100_CO6;
  assign CLBLM_R_X3Y100_SLICE_X2Y100_D = CLBLM_R_X3Y100_SLICE_X2Y100_DO6;
  assign CLBLM_R_X3Y100_SLICE_X3Y100_A = CLBLM_R_X3Y100_SLICE_X3Y100_AO6;
  assign CLBLM_R_X3Y100_SLICE_X3Y100_B = CLBLM_R_X3Y100_SLICE_X3Y100_BO6;
  assign CLBLM_R_X3Y100_SLICE_X3Y100_C = CLBLM_R_X3Y100_SLICE_X3Y100_CO6;
  assign CLBLM_R_X3Y100_SLICE_X3Y100_D = CLBLM_R_X3Y100_SLICE_X3Y100_DO6;
  assign CLBLM_R_X3Y100_SLICE_X3Y100_AMUX = CLBLM_R_X3Y100_SLICE_X3Y100_AO5;
  assign CLBLM_R_X3Y101_SLICE_X2Y101_A = CLBLM_R_X3Y101_SLICE_X2Y101_AO6;
  assign CLBLM_R_X3Y101_SLICE_X2Y101_B = CLBLM_R_X3Y101_SLICE_X2Y101_BO6;
  assign CLBLM_R_X3Y101_SLICE_X2Y101_C = CLBLM_R_X3Y101_SLICE_X2Y101_CO6;
  assign CLBLM_R_X3Y101_SLICE_X2Y101_D = CLBLM_R_X3Y101_SLICE_X2Y101_DO6;
  assign CLBLM_R_X3Y101_SLICE_X3Y101_A = CLBLM_R_X3Y101_SLICE_X3Y101_AO6;
  assign CLBLM_R_X3Y101_SLICE_X3Y101_B = CLBLM_R_X3Y101_SLICE_X3Y101_BO6;
  assign CLBLM_R_X3Y101_SLICE_X3Y101_C = CLBLM_R_X3Y101_SLICE_X3Y101_CO6;
  assign CLBLM_R_X3Y101_SLICE_X3Y101_D = CLBLM_R_X3Y101_SLICE_X3Y101_DO6;
  assign CLBLM_R_X3Y101_SLICE_X3Y101_AMUX = CLBLM_R_X3Y101_SLICE_X3Y101_AO5;
  assign CLBLM_R_X3Y102_SLICE_X2Y102_A = CLBLM_R_X3Y102_SLICE_X2Y102_AO6;
  assign CLBLM_R_X3Y102_SLICE_X2Y102_B = CLBLM_R_X3Y102_SLICE_X2Y102_BO6;
  assign CLBLM_R_X3Y102_SLICE_X2Y102_C = CLBLM_R_X3Y102_SLICE_X2Y102_CO6;
  assign CLBLM_R_X3Y102_SLICE_X2Y102_D = CLBLM_R_X3Y102_SLICE_X2Y102_DO6;
  assign CLBLM_R_X3Y102_SLICE_X3Y102_A = CLBLM_R_X3Y102_SLICE_X3Y102_AO6;
  assign CLBLM_R_X3Y102_SLICE_X3Y102_B = CLBLM_R_X3Y102_SLICE_X3Y102_BO6;
  assign CLBLM_R_X3Y102_SLICE_X3Y102_C = CLBLM_R_X3Y102_SLICE_X3Y102_CO6;
  assign CLBLM_R_X3Y102_SLICE_X3Y102_D = CLBLM_R_X3Y102_SLICE_X3Y102_DO6;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_A = CLBLM_R_X3Y103_SLICE_X2Y103_AO6;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_B = CLBLM_R_X3Y103_SLICE_X2Y103_BO6;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_C = CLBLM_R_X3Y103_SLICE_X2Y103_CO6;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_D = CLBLM_R_X3Y103_SLICE_X2Y103_DO6;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_AMUX = CLBLM_R_X3Y103_SLICE_X2Y103_AO5;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_A = CLBLM_R_X3Y103_SLICE_X3Y103_AO6;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_B = CLBLM_R_X3Y103_SLICE_X3Y103_BO6;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_C = CLBLM_R_X3Y103_SLICE_X3Y103_CO6;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_D = CLBLM_R_X3Y103_SLICE_X3Y103_DO6;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_AMUX = CLBLM_R_X3Y103_SLICE_X3Y103_AO5;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_CMUX = CLBLM_R_X3Y103_SLICE_X3Y103_CO6;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_A = CLBLM_R_X3Y104_SLICE_X2Y104_AO6;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_B = CLBLM_R_X3Y104_SLICE_X2Y104_BO6;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_C = CLBLM_R_X3Y104_SLICE_X2Y104_CO6;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_D = CLBLM_R_X3Y104_SLICE_X2Y104_DO6;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_A = CLBLM_R_X3Y104_SLICE_X3Y104_AO6;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_B = CLBLM_R_X3Y104_SLICE_X3Y104_BO6;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_C = CLBLM_R_X3Y104_SLICE_X3Y104_CO6;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_D = CLBLM_R_X3Y104_SLICE_X3Y104_DO6;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_AMUX = CLBLM_R_X3Y104_SLICE_X3Y104_AO5;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_A = CLBLM_R_X3Y105_SLICE_X2Y105_AO6;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_B = CLBLM_R_X3Y105_SLICE_X2Y105_BO6;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_C = CLBLM_R_X3Y105_SLICE_X2Y105_CO6;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_D = CLBLM_R_X3Y105_SLICE_X2Y105_DO6;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_AMUX = CLBLM_R_X3Y105_SLICE_X2Y105_AO5;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_A = CLBLM_R_X3Y105_SLICE_X3Y105_AO6;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_B = CLBLM_R_X3Y105_SLICE_X3Y105_BO6;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_C = CLBLM_R_X3Y105_SLICE_X3Y105_CO6;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_D = CLBLM_R_X3Y105_SLICE_X3Y105_DO6;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_A = CLBLM_R_X3Y106_SLICE_X2Y106_AO6;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_B = CLBLM_R_X3Y106_SLICE_X2Y106_BO6;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_C = CLBLM_R_X3Y106_SLICE_X2Y106_CO6;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_D = CLBLM_R_X3Y106_SLICE_X2Y106_DO6;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_AMUX = CLBLM_R_X3Y106_SLICE_X2Y106_AO5;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_A = CLBLM_R_X3Y106_SLICE_X3Y106_AO6;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_B = CLBLM_R_X3Y106_SLICE_X3Y106_BO6;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_C = CLBLM_R_X3Y106_SLICE_X3Y106_CO6;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_D = CLBLM_R_X3Y106_SLICE_X3Y106_DO6;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_AMUX = CLBLM_R_X3Y106_SLICE_X3Y106_AO5;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_A = CLBLM_R_X3Y107_SLICE_X2Y107_AO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_B = CLBLM_R_X3Y107_SLICE_X2Y107_BO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_C = CLBLM_R_X3Y107_SLICE_X2Y107_CO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_D = CLBLM_R_X3Y107_SLICE_X2Y107_DO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_AMUX = CLBLM_R_X3Y107_SLICE_X2Y107_AO5;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_CMUX = CLBLM_R_X3Y107_SLICE_X2Y107_CO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_A = CLBLM_R_X3Y107_SLICE_X3Y107_AO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_B = CLBLM_R_X3Y107_SLICE_X3Y107_BO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_C = CLBLM_R_X3Y107_SLICE_X3Y107_CO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_D = CLBLM_R_X3Y107_SLICE_X3Y107_DO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_AMUX = CLBLM_R_X3Y107_SLICE_X3Y107_AO5;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_A = CLBLM_R_X3Y108_SLICE_X2Y108_AO6;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_B = CLBLM_R_X3Y108_SLICE_X2Y108_BO6;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_C = CLBLM_R_X3Y108_SLICE_X2Y108_CO6;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_D = CLBLM_R_X3Y108_SLICE_X2Y108_DO6;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_AMUX = CLBLM_R_X3Y108_SLICE_X2Y108_AO5;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_A = CLBLM_R_X3Y108_SLICE_X3Y108_AO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_B = CLBLM_R_X3Y108_SLICE_X3Y108_BO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_C = CLBLM_R_X3Y108_SLICE_X3Y108_CO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_D = CLBLM_R_X3Y108_SLICE_X3Y108_DO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_BMUX = CLBLM_R_X3Y108_SLICE_X3Y108_BO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_DMUX = CLBLM_R_X3Y108_SLICE_X3Y108_DO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_A = CLBLM_R_X3Y109_SLICE_X2Y109_AO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_B = CLBLM_R_X3Y109_SLICE_X2Y109_BO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_C = CLBLM_R_X3Y109_SLICE_X2Y109_CO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_D = CLBLM_R_X3Y109_SLICE_X2Y109_DO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_A = CLBLM_R_X3Y109_SLICE_X3Y109_AO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_B = CLBLM_R_X3Y109_SLICE_X3Y109_BO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_C = CLBLM_R_X3Y109_SLICE_X3Y109_CO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_D = CLBLM_R_X3Y109_SLICE_X3Y109_DO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_A = CLBLM_R_X3Y110_SLICE_X2Y110_AO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_B = CLBLM_R_X3Y110_SLICE_X2Y110_BO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_C = CLBLM_R_X3Y110_SLICE_X2Y110_CO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_D = CLBLM_R_X3Y110_SLICE_X2Y110_DO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_AMUX = CLBLM_R_X3Y110_SLICE_X2Y110_AO5;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_BMUX = CLBLM_R_X3Y110_SLICE_X2Y110_BO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_A = CLBLM_R_X3Y110_SLICE_X3Y110_AO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_B = CLBLM_R_X3Y110_SLICE_X3Y110_BO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_C = CLBLM_R_X3Y110_SLICE_X3Y110_CO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_D = CLBLM_R_X3Y110_SLICE_X3Y110_DO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_A = CLBLM_R_X3Y111_SLICE_X2Y111_AO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_B = CLBLM_R_X3Y111_SLICE_X2Y111_BO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_C = CLBLM_R_X3Y111_SLICE_X2Y111_CO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_D = CLBLM_R_X3Y111_SLICE_X2Y111_DO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_A = CLBLM_R_X3Y111_SLICE_X3Y111_AO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_B = CLBLM_R_X3Y111_SLICE_X3Y111_BO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_C = CLBLM_R_X3Y111_SLICE_X3Y111_CO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_D = CLBLM_R_X3Y111_SLICE_X3Y111_DO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_AMUX = CLBLM_R_X3Y111_SLICE_X3Y111_AO5;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_BMUX = CLBLM_R_X3Y111_SLICE_X3Y111_BO5;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_CMUX = CLBLM_R_X3Y111_SLICE_X3Y111_CO5;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_A = CLBLM_R_X3Y112_SLICE_X2Y112_AO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_B = CLBLM_R_X3Y112_SLICE_X2Y112_BO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_C = CLBLM_R_X3Y112_SLICE_X2Y112_CO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_D = CLBLM_R_X3Y112_SLICE_X2Y112_DO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_AMUX = CLBLM_R_X3Y112_SLICE_X2Y112_AO5;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_CMUX = CLBLM_R_X3Y112_SLICE_X2Y112_CO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_A = CLBLM_R_X3Y112_SLICE_X3Y112_AO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_B = CLBLM_R_X3Y112_SLICE_X3Y112_BO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_C = CLBLM_R_X3Y112_SLICE_X3Y112_CO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_D = CLBLM_R_X3Y112_SLICE_X3Y112_DO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_AMUX = CLBLM_R_X3Y112_SLICE_X3Y112_AO5;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_BMUX = CLBLM_R_X3Y112_SLICE_X3Y112_BO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_A = CLBLM_R_X3Y113_SLICE_X2Y113_AO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_B = CLBLM_R_X3Y113_SLICE_X2Y113_BO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_C = CLBLM_R_X3Y113_SLICE_X2Y113_CO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_D = CLBLM_R_X3Y113_SLICE_X2Y113_DO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_AMUX = CLBLM_R_X3Y113_SLICE_X2Y113_AO5;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_BMUX = CLBLM_R_X3Y113_SLICE_X2Y113_BO5;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_A = CLBLM_R_X3Y113_SLICE_X3Y113_AO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_B = CLBLM_R_X3Y113_SLICE_X3Y113_BO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_C = CLBLM_R_X3Y113_SLICE_X3Y113_CO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_D = CLBLM_R_X3Y113_SLICE_X3Y113_DO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_AMUX = CLBLM_R_X3Y113_SLICE_X3Y113_AO5;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_DMUX = CLBLM_R_X3Y113_SLICE_X3Y113_DO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_A = CLBLM_R_X3Y114_SLICE_X2Y114_AO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_B = CLBLM_R_X3Y114_SLICE_X2Y114_BO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_C = CLBLM_R_X3Y114_SLICE_X2Y114_CO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_D = CLBLM_R_X3Y114_SLICE_X2Y114_DO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_AMUX = CLBLM_R_X3Y114_SLICE_X2Y114_AO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_A = CLBLM_R_X3Y114_SLICE_X3Y114_AO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_B = CLBLM_R_X3Y114_SLICE_X3Y114_BO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_C = CLBLM_R_X3Y114_SLICE_X3Y114_CO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_D = CLBLM_R_X3Y114_SLICE_X3Y114_DO6;
  assign CLBLM_R_X5Y100_SLICE_X6Y100_A = CLBLM_R_X5Y100_SLICE_X6Y100_AO6;
  assign CLBLM_R_X5Y100_SLICE_X6Y100_B = CLBLM_R_X5Y100_SLICE_X6Y100_BO6;
  assign CLBLM_R_X5Y100_SLICE_X6Y100_C = CLBLM_R_X5Y100_SLICE_X6Y100_CO6;
  assign CLBLM_R_X5Y100_SLICE_X6Y100_D = CLBLM_R_X5Y100_SLICE_X6Y100_DO6;
  assign CLBLM_R_X5Y100_SLICE_X6Y100_AMUX = CLBLM_R_X5Y100_SLICE_X6Y100_AO5;
  assign CLBLM_R_X5Y100_SLICE_X7Y100_A = CLBLM_R_X5Y100_SLICE_X7Y100_AO6;
  assign CLBLM_R_X5Y100_SLICE_X7Y100_B = CLBLM_R_X5Y100_SLICE_X7Y100_BO6;
  assign CLBLM_R_X5Y100_SLICE_X7Y100_C = CLBLM_R_X5Y100_SLICE_X7Y100_CO6;
  assign CLBLM_R_X5Y100_SLICE_X7Y100_D = CLBLM_R_X5Y100_SLICE_X7Y100_DO6;
  assign CLBLM_R_X5Y101_SLICE_X6Y101_A = CLBLM_R_X5Y101_SLICE_X6Y101_AO6;
  assign CLBLM_R_X5Y101_SLICE_X6Y101_B = CLBLM_R_X5Y101_SLICE_X6Y101_BO6;
  assign CLBLM_R_X5Y101_SLICE_X6Y101_C = CLBLM_R_X5Y101_SLICE_X6Y101_CO6;
  assign CLBLM_R_X5Y101_SLICE_X6Y101_D = CLBLM_R_X5Y101_SLICE_X6Y101_DO6;
  assign CLBLM_R_X5Y101_SLICE_X6Y101_AMUX = CLBLM_R_X5Y101_SLICE_X6Y101_AO5;
  assign CLBLM_R_X5Y101_SLICE_X6Y101_CMUX = CLBLM_R_X5Y101_SLICE_X6Y101_CO6;
  assign CLBLM_R_X5Y101_SLICE_X7Y101_A = CLBLM_R_X5Y101_SLICE_X7Y101_AO6;
  assign CLBLM_R_X5Y101_SLICE_X7Y101_B = CLBLM_R_X5Y101_SLICE_X7Y101_BO6;
  assign CLBLM_R_X5Y101_SLICE_X7Y101_C = CLBLM_R_X5Y101_SLICE_X7Y101_CO6;
  assign CLBLM_R_X5Y101_SLICE_X7Y101_D = CLBLM_R_X5Y101_SLICE_X7Y101_DO6;
  assign CLBLM_R_X5Y101_SLICE_X7Y101_AMUX = CLBLM_R_X5Y101_SLICE_X7Y101_AO5;
  assign CLBLM_R_X5Y102_SLICE_X6Y102_A = CLBLM_R_X5Y102_SLICE_X6Y102_AO6;
  assign CLBLM_R_X5Y102_SLICE_X6Y102_B = CLBLM_R_X5Y102_SLICE_X6Y102_BO6;
  assign CLBLM_R_X5Y102_SLICE_X6Y102_C = CLBLM_R_X5Y102_SLICE_X6Y102_CO6;
  assign CLBLM_R_X5Y102_SLICE_X6Y102_D = CLBLM_R_X5Y102_SLICE_X6Y102_DO6;
  assign CLBLM_R_X5Y102_SLICE_X6Y102_AMUX = CLBLM_R_X5Y102_SLICE_X6Y102_AO5;
  assign CLBLM_R_X5Y102_SLICE_X6Y102_BMUX = CLBLM_R_X5Y102_SLICE_X6Y102_BO5;
  assign CLBLM_R_X5Y102_SLICE_X6Y102_DMUX = CLBLM_R_X5Y102_SLICE_X6Y102_DO6;
  assign CLBLM_R_X5Y102_SLICE_X7Y102_A = CLBLM_R_X5Y102_SLICE_X7Y102_AO6;
  assign CLBLM_R_X5Y102_SLICE_X7Y102_B = CLBLM_R_X5Y102_SLICE_X7Y102_BO6;
  assign CLBLM_R_X5Y102_SLICE_X7Y102_C = CLBLM_R_X5Y102_SLICE_X7Y102_CO6;
  assign CLBLM_R_X5Y102_SLICE_X7Y102_D = CLBLM_R_X5Y102_SLICE_X7Y102_DO6;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_A = CLBLM_R_X5Y103_SLICE_X6Y103_AO6;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_B = CLBLM_R_X5Y103_SLICE_X6Y103_BO6;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_C = CLBLM_R_X5Y103_SLICE_X6Y103_CO6;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_D = CLBLM_R_X5Y103_SLICE_X6Y103_DO6;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_AMUX = CLBLM_R_X5Y103_SLICE_X6Y103_AO6;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_A = CLBLM_R_X5Y103_SLICE_X7Y103_AO6;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_B = CLBLM_R_X5Y103_SLICE_X7Y103_BO6;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_C = CLBLM_R_X5Y103_SLICE_X7Y103_CO6;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_D = CLBLM_R_X5Y103_SLICE_X7Y103_DO6;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_A = CLBLM_R_X5Y104_SLICE_X6Y104_AO6;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_B = CLBLM_R_X5Y104_SLICE_X6Y104_BO6;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_C = CLBLM_R_X5Y104_SLICE_X6Y104_CO6;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_D = CLBLM_R_X5Y104_SLICE_X6Y104_DO6;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_A = CLBLM_R_X5Y104_SLICE_X7Y104_AO6;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_B = CLBLM_R_X5Y104_SLICE_X7Y104_BO6;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_C = CLBLM_R_X5Y104_SLICE_X7Y104_CO6;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_D = CLBLM_R_X5Y104_SLICE_X7Y104_DO6;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_A = CLBLM_R_X5Y105_SLICE_X6Y105_AO6;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_B = CLBLM_R_X5Y105_SLICE_X6Y105_BO6;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_C = CLBLM_R_X5Y105_SLICE_X6Y105_CO6;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_D = CLBLM_R_X5Y105_SLICE_X6Y105_DO6;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_A = CLBLM_R_X5Y105_SLICE_X7Y105_AO6;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_B = CLBLM_R_X5Y105_SLICE_X7Y105_BO6;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_C = CLBLM_R_X5Y105_SLICE_X7Y105_CO6;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_D = CLBLM_R_X5Y105_SLICE_X7Y105_DO6;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_AMUX = CLBLM_R_X5Y105_SLICE_X7Y105_AO5;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_BMUX = CLBLM_R_X5Y105_SLICE_X7Y105_BO5;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_A = CLBLM_R_X5Y106_SLICE_X6Y106_AO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_B = CLBLM_R_X5Y106_SLICE_X6Y106_BO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_C = CLBLM_R_X5Y106_SLICE_X6Y106_CO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_D = CLBLM_R_X5Y106_SLICE_X6Y106_DO6;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_A = CLBLM_R_X5Y106_SLICE_X7Y106_AO6;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_B = CLBLM_R_X5Y106_SLICE_X7Y106_BO6;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_C = CLBLM_R_X5Y106_SLICE_X7Y106_CO6;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_D = CLBLM_R_X5Y106_SLICE_X7Y106_DO6;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_AMUX = CLBLM_R_X5Y106_SLICE_X7Y106_AO5;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_A = CLBLM_R_X5Y107_SLICE_X6Y107_AO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_B = CLBLM_R_X5Y107_SLICE_X6Y107_BO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_C = CLBLM_R_X5Y107_SLICE_X6Y107_CO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_D = CLBLM_R_X5Y107_SLICE_X6Y107_DO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_AMUX = CLBLM_R_X5Y107_SLICE_X6Y107_AO5;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_A = CLBLM_R_X5Y107_SLICE_X7Y107_AO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_B = CLBLM_R_X5Y107_SLICE_X7Y107_BO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_C = CLBLM_R_X5Y107_SLICE_X7Y107_CO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_D = CLBLM_R_X5Y107_SLICE_X7Y107_DO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_A = CLBLM_R_X5Y108_SLICE_X6Y108_AO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_B = CLBLM_R_X5Y108_SLICE_X6Y108_BO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_C = CLBLM_R_X5Y108_SLICE_X6Y108_CO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_D = CLBLM_R_X5Y108_SLICE_X6Y108_DO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_AMUX = CLBLM_R_X5Y108_SLICE_X6Y108_AO5;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_A = CLBLM_R_X5Y108_SLICE_X7Y108_AO6;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_B = CLBLM_R_X5Y108_SLICE_X7Y108_BO6;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_C = CLBLM_R_X5Y108_SLICE_X7Y108_CO6;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_D = CLBLM_R_X5Y108_SLICE_X7Y108_DO6;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_AMUX = CLBLM_R_X5Y108_SLICE_X7Y108_AO5;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_A = CLBLM_R_X5Y109_SLICE_X6Y109_AO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_B = CLBLM_R_X5Y109_SLICE_X6Y109_BO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_C = CLBLM_R_X5Y109_SLICE_X6Y109_CO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_D = CLBLM_R_X5Y109_SLICE_X6Y109_DO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_AMUX = CLBLM_R_X5Y109_SLICE_X6Y109_AO5;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_A = CLBLM_R_X5Y109_SLICE_X7Y109_AO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_B = CLBLM_R_X5Y109_SLICE_X7Y109_BO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_C = CLBLM_R_X5Y109_SLICE_X7Y109_CO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_D = CLBLM_R_X5Y109_SLICE_X7Y109_DO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_A = CLBLM_R_X5Y110_SLICE_X6Y110_AO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_B = CLBLM_R_X5Y110_SLICE_X6Y110_BO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_C = CLBLM_R_X5Y110_SLICE_X6Y110_CO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_D = CLBLM_R_X5Y110_SLICE_X6Y110_DO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_AMUX = CLBLM_R_X5Y110_SLICE_X6Y110_AO5;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_A = CLBLM_R_X5Y110_SLICE_X7Y110_AO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_B = CLBLM_R_X5Y110_SLICE_X7Y110_BO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_C = CLBLM_R_X5Y110_SLICE_X7Y110_CO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_D = CLBLM_R_X5Y110_SLICE_X7Y110_DO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_AMUX = CLBLM_R_X5Y110_SLICE_X7Y110_AO5;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_A = CLBLM_R_X5Y111_SLICE_X6Y111_AO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_B = CLBLM_R_X5Y111_SLICE_X6Y111_BO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_C = CLBLM_R_X5Y111_SLICE_X6Y111_CO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_D = CLBLM_R_X5Y111_SLICE_X6Y111_DO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_A = CLBLM_R_X5Y111_SLICE_X7Y111_AO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_B = CLBLM_R_X5Y111_SLICE_X7Y111_BO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_C = CLBLM_R_X5Y111_SLICE_X7Y111_CO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_D = CLBLM_R_X5Y111_SLICE_X7Y111_DO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_AMUX = CLBLM_R_X5Y111_SLICE_X7Y111_AO5;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_A = CLBLM_R_X5Y112_SLICE_X6Y112_AO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_B = CLBLM_R_X5Y112_SLICE_X6Y112_BO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_C = CLBLM_R_X5Y112_SLICE_X6Y112_CO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_D = CLBLM_R_X5Y112_SLICE_X6Y112_DO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_AMUX = CLBLM_R_X5Y112_SLICE_X6Y112_AO5;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_DMUX = CLBLM_R_X5Y112_SLICE_X6Y112_DO6;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_A = CLBLM_R_X5Y112_SLICE_X7Y112_AO6;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_B = CLBLM_R_X5Y112_SLICE_X7Y112_BO6;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_C = CLBLM_R_X5Y112_SLICE_X7Y112_CO6;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_D = CLBLM_R_X5Y112_SLICE_X7Y112_DO6;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_AMUX = CLBLM_R_X5Y112_SLICE_X7Y112_AO5;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_A = CLBLM_R_X5Y113_SLICE_X6Y113_AO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_B = CLBLM_R_X5Y113_SLICE_X6Y113_BO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_C = CLBLM_R_X5Y113_SLICE_X6Y113_CO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_D = CLBLM_R_X5Y113_SLICE_X6Y113_DO6;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_A = CLBLM_R_X5Y113_SLICE_X7Y113_AO6;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_B = CLBLM_R_X5Y113_SLICE_X7Y113_BO6;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_C = CLBLM_R_X5Y113_SLICE_X7Y113_CO6;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_D = CLBLM_R_X5Y113_SLICE_X7Y113_DO6;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_AMUX = CLBLM_R_X5Y113_SLICE_X7Y113_AO5;
  assign CLBLM_R_X7Y100_SLICE_X8Y100_A = CLBLM_R_X7Y100_SLICE_X8Y100_AO6;
  assign CLBLM_R_X7Y100_SLICE_X8Y100_B = CLBLM_R_X7Y100_SLICE_X8Y100_BO6;
  assign CLBLM_R_X7Y100_SLICE_X8Y100_C = CLBLM_R_X7Y100_SLICE_X8Y100_CO6;
  assign CLBLM_R_X7Y100_SLICE_X8Y100_D = CLBLM_R_X7Y100_SLICE_X8Y100_DO6;
  assign CLBLM_R_X7Y100_SLICE_X8Y100_AMUX = CLBLM_R_X7Y100_SLICE_X8Y100_AO5;
  assign CLBLM_R_X7Y100_SLICE_X9Y100_A = CLBLM_R_X7Y100_SLICE_X9Y100_AO6;
  assign CLBLM_R_X7Y100_SLICE_X9Y100_B = CLBLM_R_X7Y100_SLICE_X9Y100_BO6;
  assign CLBLM_R_X7Y100_SLICE_X9Y100_C = CLBLM_R_X7Y100_SLICE_X9Y100_CO6;
  assign CLBLM_R_X7Y100_SLICE_X9Y100_D = CLBLM_R_X7Y100_SLICE_X9Y100_DO6;
  assign CLBLM_R_X7Y101_SLICE_X8Y101_A = CLBLM_R_X7Y101_SLICE_X8Y101_AO6;
  assign CLBLM_R_X7Y101_SLICE_X8Y101_B = CLBLM_R_X7Y101_SLICE_X8Y101_BO6;
  assign CLBLM_R_X7Y101_SLICE_X8Y101_C = CLBLM_R_X7Y101_SLICE_X8Y101_CO6;
  assign CLBLM_R_X7Y101_SLICE_X8Y101_D = CLBLM_R_X7Y101_SLICE_X8Y101_DO6;
  assign CLBLM_R_X7Y101_SLICE_X8Y101_CMUX = CLBLM_R_X7Y101_SLICE_X8Y101_CO6;
  assign CLBLM_R_X7Y101_SLICE_X9Y101_A = CLBLM_R_X7Y101_SLICE_X9Y101_AO6;
  assign CLBLM_R_X7Y101_SLICE_X9Y101_B = CLBLM_R_X7Y101_SLICE_X9Y101_BO6;
  assign CLBLM_R_X7Y101_SLICE_X9Y101_C = CLBLM_R_X7Y101_SLICE_X9Y101_CO6;
  assign CLBLM_R_X7Y101_SLICE_X9Y101_D = CLBLM_R_X7Y101_SLICE_X9Y101_DO6;
  assign CLBLM_R_X7Y101_SLICE_X9Y101_AMUX = CLBLM_R_X7Y101_SLICE_X9Y101_AO5;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_A = CLBLM_R_X7Y102_SLICE_X8Y102_AO6;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_B = CLBLM_R_X7Y102_SLICE_X8Y102_BO6;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_C = CLBLM_R_X7Y102_SLICE_X8Y102_CO6;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_D = CLBLM_R_X7Y102_SLICE_X8Y102_DO6;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_AMUX = CLBLM_R_X7Y102_SLICE_X8Y102_AO5;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_A = CLBLM_R_X7Y102_SLICE_X9Y102_AO6;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_B = CLBLM_R_X7Y102_SLICE_X9Y102_BO6;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_C = CLBLM_R_X7Y102_SLICE_X9Y102_CO6;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_D = CLBLM_R_X7Y102_SLICE_X9Y102_DO6;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_AMUX = CLBLM_R_X7Y102_SLICE_X9Y102_AO5;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_CMUX = CLBLM_R_X7Y102_SLICE_X9Y102_CO6;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_A = CLBLM_R_X7Y103_SLICE_X8Y103_AO6;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_B = CLBLM_R_X7Y103_SLICE_X8Y103_BO6;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_C = CLBLM_R_X7Y103_SLICE_X8Y103_CO6;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_D = CLBLM_R_X7Y103_SLICE_X8Y103_DO6;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_AMUX = CLBLM_R_X7Y103_SLICE_X8Y103_AO5;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_BMUX = CLBLM_R_X7Y103_SLICE_X8Y103_BO6;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_CMUX = CLBLM_R_X7Y103_SLICE_X8Y103_CO6;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_A = CLBLM_R_X7Y103_SLICE_X9Y103_AO6;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_B = CLBLM_R_X7Y103_SLICE_X9Y103_BO6;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_C = CLBLM_R_X7Y103_SLICE_X9Y103_CO6;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_D = CLBLM_R_X7Y103_SLICE_X9Y103_DO6;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_AMUX = CLBLM_R_X7Y103_SLICE_X9Y103_AO5;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_A = CLBLM_R_X7Y104_SLICE_X8Y104_AO6;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_B = CLBLM_R_X7Y104_SLICE_X8Y104_BO6;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_C = CLBLM_R_X7Y104_SLICE_X8Y104_CO6;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_D = CLBLM_R_X7Y104_SLICE_X8Y104_DO6;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_A = CLBLM_R_X7Y104_SLICE_X9Y104_AO6;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_B = CLBLM_R_X7Y104_SLICE_X9Y104_BO6;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_C = CLBLM_R_X7Y104_SLICE_X9Y104_CO6;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_D = CLBLM_R_X7Y104_SLICE_X9Y104_DO6;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_A = CLBLM_R_X7Y105_SLICE_X8Y105_AO6;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_B = CLBLM_R_X7Y105_SLICE_X8Y105_BO6;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_C = CLBLM_R_X7Y105_SLICE_X8Y105_CO6;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_D = CLBLM_R_X7Y105_SLICE_X8Y105_DO6;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_A = CLBLM_R_X7Y105_SLICE_X9Y105_AO6;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_B = CLBLM_R_X7Y105_SLICE_X9Y105_BO6;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_C = CLBLM_R_X7Y105_SLICE_X9Y105_CO6;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_D = CLBLM_R_X7Y105_SLICE_X9Y105_DO6;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_AMUX = CLBLM_R_X7Y105_SLICE_X9Y105_AO5;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_A = CLBLM_R_X7Y106_SLICE_X8Y106_AO6;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_B = CLBLM_R_X7Y106_SLICE_X8Y106_BO6;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_C = CLBLM_R_X7Y106_SLICE_X8Y106_CO6;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_D = CLBLM_R_X7Y106_SLICE_X8Y106_DO6;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_A = CLBLM_R_X7Y106_SLICE_X9Y106_AO6;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_B = CLBLM_R_X7Y106_SLICE_X9Y106_BO6;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_C = CLBLM_R_X7Y106_SLICE_X9Y106_CO6;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_D = CLBLM_R_X7Y106_SLICE_X9Y106_DO6;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_AMUX = CLBLM_R_X7Y106_SLICE_X9Y106_AO5;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_A = CLBLM_R_X7Y107_SLICE_X8Y107_AO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_B = CLBLM_R_X7Y107_SLICE_X8Y107_BO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_C = CLBLM_R_X7Y107_SLICE_X8Y107_CO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_D = CLBLM_R_X7Y107_SLICE_X8Y107_DO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_A = CLBLM_R_X7Y107_SLICE_X9Y107_AO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_B = CLBLM_R_X7Y107_SLICE_X9Y107_BO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_C = CLBLM_R_X7Y107_SLICE_X9Y107_CO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_D = CLBLM_R_X7Y107_SLICE_X9Y107_DO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_AMUX = CLBLM_R_X7Y107_SLICE_X9Y107_AO5;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_A = CLBLM_R_X7Y108_SLICE_X8Y108_AO6;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_B = CLBLM_R_X7Y108_SLICE_X8Y108_BO6;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_C = CLBLM_R_X7Y108_SLICE_X8Y108_CO6;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_D = CLBLM_R_X7Y108_SLICE_X8Y108_DO6;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_AMUX = CLBLM_R_X7Y108_SLICE_X8Y108_AO5;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_A = CLBLM_R_X7Y108_SLICE_X9Y108_AO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_B = CLBLM_R_X7Y108_SLICE_X9Y108_BO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_C = CLBLM_R_X7Y108_SLICE_X9Y108_CO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_D = CLBLM_R_X7Y108_SLICE_X9Y108_DO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_A = CLBLM_R_X7Y109_SLICE_X8Y109_AO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_B = CLBLM_R_X7Y109_SLICE_X8Y109_BO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_C = CLBLM_R_X7Y109_SLICE_X8Y109_CO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_D = CLBLM_R_X7Y109_SLICE_X8Y109_DO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_A = CLBLM_R_X7Y109_SLICE_X9Y109_AO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_B = CLBLM_R_X7Y109_SLICE_X9Y109_BO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_C = CLBLM_R_X7Y109_SLICE_X9Y109_CO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_D = CLBLM_R_X7Y109_SLICE_X9Y109_DO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_A = CLBLM_R_X7Y110_SLICE_X8Y110_AO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_B = CLBLM_R_X7Y110_SLICE_X8Y110_BO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_C = CLBLM_R_X7Y110_SLICE_X8Y110_CO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_D = CLBLM_R_X7Y110_SLICE_X8Y110_DO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_A = CLBLM_R_X7Y110_SLICE_X9Y110_AO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_B = CLBLM_R_X7Y110_SLICE_X9Y110_BO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_C = CLBLM_R_X7Y110_SLICE_X9Y110_CO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_D = CLBLM_R_X7Y110_SLICE_X9Y110_DO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_AMUX = CLBLM_R_X7Y110_SLICE_X9Y110_AO5;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_A = CLBLM_R_X7Y111_SLICE_X8Y111_AO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_B = CLBLM_R_X7Y111_SLICE_X8Y111_BO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_C = CLBLM_R_X7Y111_SLICE_X8Y111_CO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_D = CLBLM_R_X7Y111_SLICE_X8Y111_DO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_AMUX = CLBLM_R_X7Y111_SLICE_X8Y111_AO5;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_A = CLBLM_R_X7Y111_SLICE_X9Y111_AO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_B = CLBLM_R_X7Y111_SLICE_X9Y111_BO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_C = CLBLM_R_X7Y111_SLICE_X9Y111_CO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_D = CLBLM_R_X7Y111_SLICE_X9Y111_DO6;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_A = CLBLM_R_X7Y112_SLICE_X8Y112_AO6;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_B = CLBLM_R_X7Y112_SLICE_X8Y112_BO6;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_C = CLBLM_R_X7Y112_SLICE_X8Y112_CO6;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_D = CLBLM_R_X7Y112_SLICE_X8Y112_DO6;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_AMUX = CLBLM_R_X7Y112_SLICE_X8Y112_AO5;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_A = CLBLM_R_X7Y112_SLICE_X9Y112_AO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_B = CLBLM_R_X7Y112_SLICE_X9Y112_BO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_C = CLBLM_R_X7Y112_SLICE_X9Y112_CO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_D = CLBLM_R_X7Y112_SLICE_X9Y112_DO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_AMUX = CLBLM_R_X7Y112_SLICE_X9Y112_AO5;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_A = CLBLM_R_X7Y113_SLICE_X8Y113_AO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_B = CLBLM_R_X7Y113_SLICE_X8Y113_BO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_C = CLBLM_R_X7Y113_SLICE_X8Y113_CO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_D = CLBLM_R_X7Y113_SLICE_X8Y113_DO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_AMUX = CLBLM_R_X7Y113_SLICE_X8Y113_AO5;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_BMUX = CLBLM_R_X7Y113_SLICE_X8Y113_BO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_A = CLBLM_R_X7Y113_SLICE_X9Y113_AO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_B = CLBLM_R_X7Y113_SLICE_X9Y113_BO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_C = CLBLM_R_X7Y113_SLICE_X9Y113_CO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_D = CLBLM_R_X7Y113_SLICE_X9Y113_DO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_AMUX = CLBLM_R_X7Y113_SLICE_X9Y113_AO5;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_A = CLBLM_R_X11Y106_SLICE_X14Y106_AO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_B = CLBLM_R_X11Y106_SLICE_X14Y106_BO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_C = CLBLM_R_X11Y106_SLICE_X14Y106_CO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_D = CLBLM_R_X11Y106_SLICE_X14Y106_DO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_AMUX = CLBLM_R_X11Y106_SLICE_X14Y106_AO5;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_A = CLBLM_R_X11Y106_SLICE_X15Y106_AO6;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_B = CLBLM_R_X11Y106_SLICE_X15Y106_BO6;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_C = CLBLM_R_X11Y106_SLICE_X15Y106_CO6;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_D = CLBLM_R_X11Y106_SLICE_X15Y106_DO6;
  assign LIOI3_X0Y101_ILOGIC_X0Y102_O = LIOB33_X0Y101_IOB_X0Y102_I;
  assign LIOI3_X0Y101_ILOGIC_X0Y101_O = LIOB33_X0Y101_IOB_X0Y101_I;
  assign LIOI3_X0Y103_ILOGIC_X0Y104_O = LIOB33_X0Y103_IOB_X0Y104_I;
  assign LIOI3_X0Y103_ILOGIC_X0Y103_O = LIOB33_X0Y103_IOB_X0Y103_I;
  assign LIOI3_X0Y105_ILOGIC_X0Y106_O = LIOB33_X0Y105_IOB_X0Y106_I;
  assign LIOI3_X0Y105_ILOGIC_X0Y105_O = LIOB33_X0Y105_IOB_X0Y105_I;
  assign LIOI3_X0Y109_ILOGIC_X0Y110_O = LIOB33_X0Y109_IOB_X0Y110_I;
  assign LIOI3_X0Y109_ILOGIC_X0Y109_O = LIOB33_X0Y109_IOB_X0Y109_I;
  assign LIOI3_X0Y111_ILOGIC_X0Y112_O = LIOB33_X0Y111_IOB_X0Y112_I;
  assign LIOI3_X0Y111_ILOGIC_X0Y111_O = LIOB33_X0Y111_IOB_X0Y111_I;
  assign LIOI3_X0Y115_ILOGIC_X0Y116_O = LIOB33_X0Y115_IOB_X0Y116_I;
  assign LIOI3_X0Y115_ILOGIC_X0Y115_O = LIOB33_X0Y115_IOB_X0Y115_I;
  assign LIOI3_X0Y117_ILOGIC_X0Y117_O = LIOB33_X0Y117_IOB_X0Y117_I;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_OQ = CLBLL_L_X2Y114_SLICE_X0Y114_AO5;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_TQ = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_OQ = CLBLL_L_X2Y113_SLICE_X1Y113_AO6;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_TQ = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_OQ = CLBLL_L_X2Y113_SLICE_X0Y113_BO5;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_TQ = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_OQ = CLBLM_R_X3Y112_SLICE_X2Y112_AO6;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_TQ = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_OQ = CLBLL_L_X2Y113_SLICE_X1Y113_CO6;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_TQ = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_OQ = CLBLM_R_X3Y111_SLICE_X2Y111_BO6;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_TQ = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_OQ = CLBLM_R_X3Y111_SLICE_X3Y111_AO6;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_TQ = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_OQ = CLBLL_L_X4Y107_SLICE_X4Y107_AO6;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_TQ = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_OQ = CLBLL_L_X4Y110_SLICE_X4Y110_AO5;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_TQ = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_OQ = CLBLL_L_X2Y114_SLICE_X0Y114_BO5;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_TQ = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_OQ = CLBLM_R_X3Y110_SLICE_X3Y110_BO6;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_TQ = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_OQ = 1'b0;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_TQ = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_OQ = CLBLM_R_X3Y110_SLICE_X2Y110_CO6;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_TQ = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_OQ = CLBLM_R_X3Y107_SLICE_X2Y107_AO6;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_TQ = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_OQ = CLBLM_R_X3Y107_SLICE_X2Y107_AO5;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_TQ = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_OQ = CLBLL_L_X2Y105_SLICE_X1Y105_DO6;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_TQ = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_OQ = CLBLL_L_X2Y107_SLICE_X1Y107_CO6;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_TQ = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_OQ = CLBLL_L_X2Y105_SLICE_X0Y105_AO5;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_TQ = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_OQ = CLBLL_L_X2Y105_SLICE_X0Y105_AO6;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_TQ = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_OQ = CLBLM_R_X3Y104_SLICE_X3Y104_BO6;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_TQ = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_OQ = CLBLM_R_X3Y104_SLICE_X3Y104_DO6;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_TQ = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_OQ = CLBLL_L_X2Y108_SLICE_X0Y108_BO6;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_TQ = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_OQ = CLBLL_L_X2Y108_SLICE_X0Y108_DO6;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_TQ = 1'b1;
  assign LIOI3_SING_X0Y100_ILOGIC_X0Y100_O = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_OQ = CLBLL_L_X2Y108_SLICE_X0Y108_CO6;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y108_O = LIOB33_X0Y107_IOB_X0Y108_I;
  assign LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y107_O = LIOB33_X0Y107_IOB_X0Y107_I;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_OQ = CLBLL_L_X2Y113_SLICE_X0Y113_AO5;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_OQ = CLBLL_L_X2Y114_SLICE_X0Y114_AO6;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_OQ = CLBLM_R_X3Y110_SLICE_X2Y110_BO6;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_OQ = CLBLM_R_X3Y110_SLICE_X2Y110_AO5;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_OQ = CLBLL_L_X2Y104_SLICE_X1Y104_CO6;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_OQ = CLBLL_L_X2Y106_SLICE_X0Y106_BO6;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y114_O = LIOB33_X0Y113_IOB_X0Y114_I;
  assign LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y113_O = LIOB33_X0Y113_IOB_X0Y113_I;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_OQ = CLBLL_L_X2Y108_SLICE_X1Y108_DO6;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_OQ = CLBLL_L_X2Y109_SLICE_X1Y109_AO6;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_TQ = 1'b1;
  assign RIOI3_X105Y101_ILOGIC_X1Y102_O = RIOB33_X105Y101_IOB_X1Y102_I;
  assign RIOI3_X105Y101_ILOGIC_X1Y101_O = RIOB33_X105Y101_IOB_X1Y101_I;
  assign RIOI3_X105Y103_ILOGIC_X1Y104_O = RIOB33_X105Y103_IOB_X1Y104_I;
  assign RIOI3_X105Y103_ILOGIC_X1Y103_O = RIOB33_X105Y103_IOB_X1Y103_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y106_O = RIOB33_X105Y105_IOB_X1Y106_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y105_O = RIOB33_X105Y105_IOB_X1Y105_I;
  assign RIOI3_X105Y109_ILOGIC_X1Y110_O = RIOB33_X105Y109_IOB_X1Y110_I;
  assign RIOI3_X105Y109_ILOGIC_X1Y109_O = RIOB33_X105Y109_IOB_X1Y109_I;
  assign RIOI3_X105Y111_ILOGIC_X1Y112_O = RIOB33_X105Y111_IOB_X1Y112_I;
  assign RIOI3_X105Y111_ILOGIC_X1Y111_O = RIOB33_X105Y111_IOB_X1Y111_I;
  assign RIOI3_SING_X105Y100_ILOGIC_X1Y100_O = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_O = RIOB33_X105Y107_IOB_X1Y108_I;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_O = RIOB33_X105Y107_IOB_X1Y107_I;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_O = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_C6 = CLBLM_L_X8Y104_SLICE_X10Y104_AO6;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_D1 = CLBLM_L_X8Y102_SLICE_X11Y102_AO6;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_D2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_D3 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_D4 = CLBLM_L_X10Y102_SLICE_X12Y102_CO6;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_D5 = CLBLM_L_X10Y104_SLICE_X13Y104_CO6;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_D6 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_A4 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_A5 = 1'b1;
  assign LIOB33_X0Y147_IOB_X0Y147_O = CLBLL_L_X2Y108_SLICE_X0Y108_DO6;
  assign LIOB33_X0Y147_IOB_X0Y148_O = CLBLL_L_X2Y108_SLICE_X0Y108_BO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_A6 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_B6 = CLBLM_R_X3Y103_SLICE_X2Y103_CO6;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_A1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_A2 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_A3 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_A4 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_A5 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_A6 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_B2 = CLBLM_L_X10Y103_SLICE_X13Y103_DO6;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_B3 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_B4 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_B5 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_B6 = CLBLM_R_X11Y106_SLICE_X14Y106_CO6;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_C1 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_C2 = CLBLM_L_X10Y103_SLICE_X13Y103_DO6;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_C4 = CLBLM_R_X11Y106_SLICE_X14Y106_CO6;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_C5 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_C6 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_C1 = CLBLM_R_X5Y111_SLICE_X7Y111_AO6;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_D1 = 1'b1;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_D2 = 1'b1;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_D3 = 1'b1;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_D4 = 1'b1;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_D5 = 1'b1;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_D6 = 1'b1;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_C2 = CLBLL_L_X4Y111_SLICE_X5Y111_DO6;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_A1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_A2 = 1'b1;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_A3 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_A4 = 1'b1;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_A5 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_A6 = 1'b1;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_B1 = CLBLM_L_X10Y103_SLICE_X13Y103_AO6;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_B2 = CLBLM_L_X10Y102_SLICE_X12Y102_BO6;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_B3 = CLBLM_L_X10Y103_SLICE_X13Y103_CO6;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_B4 = CLBLM_R_X11Y106_SLICE_X14Y106_CO6;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_B5 = CLBLM_L_X10Y104_SLICE_X12Y104_AO6;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_B6 = CLBLM_L_X10Y103_SLICE_X12Y103_AO5;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_C1 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_C2 = CLBLM_L_X10Y104_SLICE_X13Y104_CO6;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_C4 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_C5 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_C6 = CLBLM_L_X8Y102_SLICE_X11Y102_BO6;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_D1 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_D2 = CLBLM_L_X10Y104_SLICE_X13Y104_CO6;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_D3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_D4 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_D5 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_D6 = CLBLM_L_X8Y102_SLICE_X11Y102_BO6;
  assign CLBLL_L_X4Y100_SLICE_X4Y100_A1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X4Y100_SLICE_X4Y100_A2 = CLBLL_L_X4Y100_SLICE_X5Y100_BO6;
  assign CLBLL_L_X4Y100_SLICE_X4Y100_A3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X4Y100_SLICE_X4Y100_A4 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLL_L_X4Y100_SLICE_X4Y100_A5 = CLBLL_L_X4Y100_SLICE_X4Y100_CO6;
  assign CLBLL_L_X4Y100_SLICE_X4Y100_A6 = 1'b1;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_D3 = CLBLM_R_X7Y111_SLICE_X8Y111_DO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_D4 = CLBLM_R_X5Y111_SLICE_X7Y111_AO5;
  assign CLBLL_L_X4Y100_SLICE_X4Y100_B1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X4Y100_SLICE_X4Y100_B2 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLL_L_X4Y100_SLICE_X4Y100_B3 = CLBLL_L_X4Y100_SLICE_X5Y100_AO6;
  assign CLBLL_L_X4Y100_SLICE_X4Y100_B4 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLL_L_X4Y100_SLICE_X4Y100_B5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y100_SLICE_X4Y100_B6 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLL_L_X4Y100_SLICE_X4Y100_C1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y100_SLICE_X4Y100_C2 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLL_L_X4Y100_SLICE_X4Y100_C3 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLL_L_X4Y100_SLICE_X4Y100_C4 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLL_L_X4Y100_SLICE_X4Y100_C5 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X4Y100_SLICE_X4Y100_C6 = CLBLL_L_X4Y100_SLICE_X5Y100_AO6;
  assign CLBLL_L_X4Y100_SLICE_X4Y100_D1 = 1'b1;
  assign CLBLL_L_X4Y100_SLICE_X4Y100_D2 = 1'b1;
  assign CLBLL_L_X4Y100_SLICE_X4Y100_D3 = 1'b1;
  assign CLBLL_L_X4Y100_SLICE_X4Y100_D4 = 1'b1;
  assign CLBLL_L_X4Y100_SLICE_X4Y100_D5 = 1'b1;
  assign CLBLL_L_X4Y100_SLICE_X4Y100_D6 = 1'b1;
  assign CLBLL_L_X4Y100_SLICE_X5Y100_A1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X4Y100_SLICE_X5Y100_A2 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X4Y100_SLICE_X5Y100_A3 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLL_L_X4Y100_SLICE_X5Y100_A4 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLL_L_X4Y100_SLICE_X5Y100_A5 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLL_L_X4Y100_SLICE_X5Y100_A6 = CLBLM_R_X5Y103_SLICE_X6Y103_CO6;
  assign CLBLL_L_X4Y100_SLICE_X5Y100_B1 = CLBLL_L_X4Y100_SLICE_X5Y100_DO6;
  assign CLBLL_L_X4Y100_SLICE_X5Y100_B2 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLL_L_X4Y100_SLICE_X5Y100_B3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y100_SLICE_X5Y100_B4 = CLBLM_R_X5Y101_SLICE_X7Y101_AO6;
  assign CLBLL_L_X4Y100_SLICE_X5Y100_B5 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLL_L_X4Y100_SLICE_X5Y100_B6 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLL_L_X4Y100_SLICE_X5Y100_C1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y100_SLICE_X5Y100_C2 = CLBLL_L_X4Y100_SLICE_X4Y100_CO6;
  assign CLBLL_L_X4Y100_SLICE_X5Y100_C3 = CLBLM_R_X5Y101_SLICE_X7Y101_AO6;
  assign CLBLL_L_X4Y100_SLICE_X5Y100_C4 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X4Y100_SLICE_X5Y100_C5 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLL_L_X4Y100_SLICE_X5Y100_C6 = CLBLM_R_X5Y100_SLICE_X6Y100_AO6;
  assign CLBLL_L_X4Y100_SLICE_X5Y100_D1 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLL_L_X4Y100_SLICE_X5Y100_D2 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLL_L_X4Y100_SLICE_X5Y100_D3 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X4Y100_SLICE_X5Y100_D4 = CLBLM_R_X5Y103_SLICE_X6Y103_CO6;
  assign CLBLL_L_X4Y100_SLICE_X5Y100_D5 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLL_L_X4Y100_SLICE_X5Y100_D6 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_A1 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_A2 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_A3 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_A4 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_A6 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_B1 = CLBLM_L_X10Y105_SLICE_X13Y105_DO6;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_B2 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_B3 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_B4 = CLBLM_L_X10Y106_SLICE_X13Y106_BO6;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_B5 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_B6 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_C1 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_C2 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_C3 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_C4 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_C5 = CLBLM_L_X10Y105_SLICE_X13Y105_DO6;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_C6 = CLBLM_L_X10Y106_SLICE_X13Y106_BO6;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_D1 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_D2 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_D3 = CLBLM_L_X10Y106_SLICE_X13Y106_AO5;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_D4 = CLBLM_L_X10Y103_SLICE_X13Y103_DO6;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_D5 = CLBLM_L_X8Y101_SLICE_X11Y101_AO5;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_D6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_A1 = CLBLM_L_X8Y105_SLICE_X10Y105_AO6;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_A2 = CLBLM_L_X10Y106_SLICE_X13Y106_BO6;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_A3 = CLBLM_L_X10Y104_SLICE_X12Y104_AO5;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_A4 = CLBLM_L_X10Y104_SLICE_X12Y104_BO6;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_A5 = CLBLM_L_X10Y104_SLICE_X13Y104_BO6;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_A6 = CLBLM_L_X10Y106_SLICE_X12Y106_AO5;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_B1 = CLBLM_L_X8Y105_SLICE_X10Y105_AO6;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_B2 = CLBLM_L_X10Y104_SLICE_X12Y104_BO6;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_B3 = CLBLM_L_X10Y104_SLICE_X12Y104_AO5;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_B4 = CLBLM_L_X10Y106_SLICE_X13Y106_BO6;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_B5 = CLBLM_L_X10Y104_SLICE_X13Y104_BO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_D4 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_B6 = CLBLM_L_X10Y106_SLICE_X12Y106_AO5;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_C1 = CLBLM_L_X10Y104_SLICE_X13Y104_BO6;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_C2 = CLBLM_L_X10Y104_SLICE_X12Y104_BO6;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_C3 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_C4 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_C5 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_C6 = CLBLM_L_X10Y106_SLICE_X13Y106_BO6;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_D1 = 1'b1;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_D2 = 1'b1;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_D3 = 1'b1;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_D4 = 1'b1;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_D5 = 1'b1;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_D6 = 1'b1;
  assign CLBLL_L_X4Y101_SLICE_X4Y101_A1 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLL_L_X4Y101_SLICE_X4Y101_A2 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLL_L_X4Y101_SLICE_X4Y101_A3 = CLBLL_L_X4Y100_SLICE_X4Y100_AO6;
  assign CLBLL_L_X4Y101_SLICE_X4Y101_A4 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X4Y101_SLICE_X4Y101_A5 = CLBLL_L_X4Y100_SLICE_X4Y100_BO6;
  assign CLBLL_L_X4Y101_SLICE_X4Y101_A6 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLL_L_X4Y101_SLICE_X4Y101_B1 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X4Y101_SLICE_X4Y101_B2 = CLBLL_L_X4Y101_SLICE_X5Y101_BO5;
  assign CLBLL_L_X4Y101_SLICE_X4Y101_B3 = CLBLL_L_X4Y101_SLICE_X5Y101_CO5;
  assign CLBLL_L_X4Y101_SLICE_X4Y101_B4 = CLBLL_L_X4Y102_SLICE_X5Y102_BO6;
  assign CLBLL_L_X4Y101_SLICE_X4Y101_B5 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X4Y101_SLICE_X4Y101_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y101_SLICE_X4Y101_C1 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X4Y101_SLICE_X4Y101_C2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y101_SLICE_X4Y101_C3 = CLBLL_L_X4Y101_SLICE_X5Y101_BO5;
  assign CLBLL_L_X4Y101_SLICE_X4Y101_C4 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X4Y101_SLICE_X4Y101_C5 = CLBLL_L_X4Y101_SLICE_X5Y101_CO5;
  assign CLBLL_L_X4Y101_SLICE_X4Y101_C6 = CLBLL_L_X4Y102_SLICE_X5Y102_BO6;
  assign CLBLL_L_X4Y101_SLICE_X4Y101_D1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y101_SLICE_X4Y101_D2 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLL_L_X4Y101_SLICE_X4Y101_D3 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X4Y101_SLICE_X4Y101_D4 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLL_L_X4Y101_SLICE_X4Y101_D5 = CLBLL_L_X4Y100_SLICE_X5Y100_AO6;
  assign CLBLL_L_X4Y101_SLICE_X4Y101_D6 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X5Y101_SLICE_X7Y101_A3 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLL_L_X4Y101_SLICE_X5Y101_A1 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLL_L_X4Y101_SLICE_X5Y101_A2 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLL_L_X4Y101_SLICE_X5Y101_A3 = CLBLL_L_X4Y101_SLICE_X4Y101_AO6;
  assign CLBLL_L_X4Y101_SLICE_X5Y101_A4 = CLBLM_R_X5Y100_SLICE_X6Y100_BO6;
  assign CLBLL_L_X4Y101_SLICE_X5Y101_A5 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLL_L_X4Y101_SLICE_X5Y101_A6 = 1'b1;
  assign CLBLL_L_X4Y101_SLICE_X5Y101_B1 = CLBLM_R_X5Y101_SLICE_X6Y101_DO6;
  assign CLBLL_L_X4Y101_SLICE_X5Y101_B2 = CLBLL_L_X4Y101_SLICE_X5Y101_AO5;
  assign CLBLL_L_X4Y101_SLICE_X5Y101_B3 = 1'b1;
  assign CLBLL_L_X4Y101_SLICE_X5Y101_B4 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLL_L_X4Y101_SLICE_X5Y101_B5 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLL_L_X4Y101_SLICE_X5Y101_B6 = 1'b1;
  assign CLBLL_L_X4Y101_SLICE_X5Y101_C1 = CLBLM_R_X5Y101_SLICE_X6Y101_BO6;
  assign CLBLL_L_X4Y101_SLICE_X5Y101_C2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y101_SLICE_X5Y101_C3 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLL_L_X4Y101_SLICE_X5Y101_C4 = CLBLM_R_X5Y102_SLICE_X6Y102_AO5;
  assign CLBLL_L_X4Y101_SLICE_X5Y101_C5 = 1'b1;
  assign CLBLL_L_X4Y101_SLICE_X5Y101_C6 = 1'b1;
  assign CLBLL_L_X4Y101_SLICE_X5Y101_D1 = CLBLM_R_X5Y101_SLICE_X6Y101_BO6;
  assign CLBLL_L_X4Y101_SLICE_X5Y101_D2 = CLBLM_R_X5Y102_SLICE_X6Y102_AO5;
  assign CLBLL_L_X4Y101_SLICE_X5Y101_D3 = CLBLL_L_X4Y101_SLICE_X5Y101_AO5;
  assign CLBLL_L_X4Y101_SLICE_X5Y101_D4 = CLBLL_L_X4Y101_SLICE_X5Y101_CO6;
  assign CLBLL_L_X4Y101_SLICE_X5Y101_D5 = CLBLM_R_X5Y101_SLICE_X6Y101_DO6;
  assign CLBLL_L_X4Y101_SLICE_X5Y101_D6 = CLBLL_L_X4Y101_SLICE_X5Y101_BO6;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_A1 = CLBLM_L_X10Y109_SLICE_X12Y109_BO6;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_A2 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_A3 = 1'b1;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_A4 = CLBLM_L_X10Y105_SLICE_X13Y105_AO6;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_A5 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_A6 = 1'b1;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_B1 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_B2 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_B3 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_B4 = CLBLM_L_X10Y108_SLICE_X13Y108_DO6;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_B5 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_B6 = CLBLM_R_X11Y106_SLICE_X14Y106_DO6;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_C1 = CLBLM_L_X10Y106_SLICE_X13Y106_AO6;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_C2 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_C3 = CLBLM_L_X10Y109_SLICE_X12Y109_AO5;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_C4 = CLBLM_R_X11Y106_SLICE_X14Y106_DO6;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_C5 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_C6 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_D1 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_D2 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_D3 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_D4 = CLBLM_L_X10Y106_SLICE_X13Y106_CO6;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_D5 = CLBLM_L_X10Y107_SLICE_X12Y107_DO6;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_D6 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_A1 = 1'b1;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_A2 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_A3 = 1'b1;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_A4 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_A5 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_A6 = 1'b1;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_B1 = CLBLM_L_X10Y103_SLICE_X13Y103_AO6;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_B2 = CLBLM_R_X11Y106_SLICE_X14Y106_BO6;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_B3 = CLBLM_L_X10Y104_SLICE_X12Y104_AO6;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_B4 = CLBLM_L_X10Y108_SLICE_X13Y108_DO6;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_B5 = CLBLM_L_X10Y106_SLICE_X12Y106_AO6;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_B6 = CLBLM_R_X11Y106_SLICE_X14Y106_CO6;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_C1 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_C2 = CLBLM_L_X10Y106_SLICE_X13Y106_CO6;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_C3 = CLBLM_L_X10Y107_SLICE_X12Y107_DO6;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_C4 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_C5 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_C6 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_D1 = CLBLM_L_X10Y105_SLICE_X12Y105_CO6;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_D2 = CLBLM_L_X10Y105_SLICE_X13Y105_CO6;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_D3 = CLBLM_L_X10Y106_SLICE_X13Y106_DO6;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_D4 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_D5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_D6 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLL_L_X4Y102_SLICE_X4Y102_A1 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLL_L_X4Y102_SLICE_X4Y102_A2 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLL_L_X4Y102_SLICE_X4Y102_A3 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X4Y102_SLICE_X4Y102_A4 = 1'b1;
  assign CLBLL_L_X4Y102_SLICE_X4Y102_A5 = 1'b1;
  assign CLBLL_L_X4Y102_SLICE_X4Y102_A6 = 1'b1;
  assign CLBLL_L_X4Y102_SLICE_X4Y102_B1 = CLBLM_R_X5Y103_SLICE_X6Y103_DO6;
  assign CLBLL_L_X4Y102_SLICE_X4Y102_B2 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLL_L_X4Y102_SLICE_X4Y102_B3 = CLBLM_R_X5Y102_SLICE_X6Y102_DO6;
  assign CLBLL_L_X4Y102_SLICE_X4Y102_B4 = CLBLM_R_X7Y102_SLICE_X9Y102_AO5;
  assign CLBLL_L_X4Y102_SLICE_X4Y102_B5 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLL_L_X4Y102_SLICE_X4Y102_B6 = 1'b1;
  assign CLBLL_L_X4Y102_SLICE_X4Y102_C1 = CLBLL_L_X4Y102_SLICE_X4Y102_AO6;
  assign CLBLL_L_X4Y102_SLICE_X4Y102_C2 = CLBLM_R_X5Y102_SLICE_X6Y102_CO6;
  assign CLBLL_L_X4Y102_SLICE_X4Y102_C3 = CLBLL_L_X4Y106_SLICE_X4Y106_AO5;
  assign CLBLL_L_X4Y102_SLICE_X4Y102_C4 = CLBLL_L_X4Y102_SLICE_X4Y102_AO5;
  assign CLBLL_L_X4Y102_SLICE_X4Y102_C5 = CLBLM_R_X5Y103_SLICE_X6Y103_DO6;
  assign CLBLL_L_X4Y102_SLICE_X4Y102_C6 = CLBLL_L_X4Y102_SLICE_X4Y102_BO6;
  assign CLBLL_L_X4Y102_SLICE_X4Y102_D1 = CLBLM_R_X3Y102_SLICE_X3Y102_BO6;
  assign CLBLL_L_X4Y102_SLICE_X4Y102_D2 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X4Y102_SLICE_X4Y102_D3 = CLBLL_L_X4Y102_SLICE_X5Y102_DO6;
  assign CLBLL_L_X4Y102_SLICE_X4Y102_D4 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X4Y102_SLICE_X4Y102_D5 = CLBLM_R_X3Y102_SLICE_X3Y102_CO6;
  assign CLBLL_L_X4Y102_SLICE_X4Y102_D6 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B1 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B3 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_C4 = CLBLM_R_X5Y110_SLICE_X6Y110_DO6;
  assign CLBLL_L_X4Y102_SLICE_X5Y102_A1 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLL_L_X4Y102_SLICE_X5Y102_A2 = CLBLM_R_X5Y101_SLICE_X6Y101_DO6;
  assign CLBLL_L_X4Y102_SLICE_X5Y102_A3 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X4Y102_SLICE_X5Y102_A4 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLL_L_X4Y102_SLICE_X5Y102_A5 = CLBLL_L_X4Y101_SLICE_X5Y101_AO5;
  assign CLBLL_L_X4Y102_SLICE_X5Y102_A6 = CLBLL_L_X4Y102_SLICE_X5Y102_CO6;
  assign CLBLL_L_X4Y102_SLICE_X5Y102_B1 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLL_L_X4Y102_SLICE_X5Y102_B2 = CLBLM_R_X5Y101_SLICE_X6Y101_DO6;
  assign CLBLL_L_X4Y102_SLICE_X5Y102_B3 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X4Y102_SLICE_X5Y102_B4 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLL_L_X4Y102_SLICE_X5Y102_B5 = CLBLL_L_X4Y101_SLICE_X5Y101_AO5;
  assign CLBLL_L_X4Y102_SLICE_X5Y102_B6 = CLBLL_L_X4Y102_SLICE_X5Y102_CO6;
  assign CLBLL_L_X4Y102_SLICE_X5Y102_C1 = CLBLL_L_X4Y101_SLICE_X4Y101_AO6;
  assign CLBLL_L_X4Y102_SLICE_X5Y102_C2 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLL_L_X4Y102_SLICE_X5Y102_C3 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLL_L_X4Y102_SLICE_X5Y102_C4 = CLBLM_R_X3Y101_SLICE_X3Y101_CO6;
  assign CLBLL_L_X4Y102_SLICE_X5Y102_C5 = CLBLM_R_X5Y100_SLICE_X6Y100_BO6;
  assign CLBLL_L_X4Y102_SLICE_X5Y102_C6 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLL_L_X4Y102_SLICE_X5Y102_D1 = CLBLL_L_X4Y101_SLICE_X4Y101_AO6;
  assign CLBLL_L_X4Y102_SLICE_X5Y102_D2 = CLBLM_R_X3Y101_SLICE_X3Y101_CO6;
  assign CLBLL_L_X4Y102_SLICE_X5Y102_D3 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLL_L_X4Y102_SLICE_X5Y102_D4 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLL_L_X4Y102_SLICE_X5Y102_D5 = CLBLM_R_X5Y100_SLICE_X6Y100_BO6;
  assign CLBLL_L_X4Y102_SLICE_X5Y102_D6 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C1 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_A1 = CLBLM_L_X10Y107_SLICE_X13Y107_BO6;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_A2 = CLBLM_L_X10Y108_SLICE_X12Y108_AO5;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_A3 = CLBLM_L_X10Y106_SLICE_X12Y106_BO6;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_A4 = CLBLM_L_X10Y107_SLICE_X12Y107_AO5;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_A5 = CLBLM_L_X10Y107_SLICE_X12Y107_DO6;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_A6 = CLBLM_L_X10Y106_SLICE_X12Y106_AO5;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_B1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_B2 = CLBLM_L_X10Y108_SLICE_X13Y108_DO6;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_B3 = CLBLM_R_X11Y106_SLICE_X14Y106_DO6;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_B4 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_B5 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_B6 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_C1 = CLBLM_L_X10Y107_SLICE_X12Y107_AO5;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_C2 = CLBLM_L_X10Y106_SLICE_X12Y106_AO5;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_C3 = CLBLM_L_X10Y107_SLICE_X12Y107_DO6;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_C4 = CLBLM_L_X10Y108_SLICE_X12Y108_AO5;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_C5 = CLBLM_L_X10Y106_SLICE_X12Y106_BO6;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_C6 = CLBLM_L_X10Y107_SLICE_X13Y107_BO6;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_D1 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_D2 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_D3 = CLBLM_L_X10Y107_SLICE_X12Y107_DO6;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_D4 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_D5 = CLBLM_L_X10Y106_SLICE_X12Y106_BO6;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_D6 = CLBLM_L_X10Y107_SLICE_X13Y107_BO6;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_A1 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_A2 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_A3 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_A4 = 1'b1;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_A5 = 1'b1;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_A6 = 1'b1;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_B1 = CLBLM_L_X8Y110_SLICE_X11Y110_DO6;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_B2 = CLBLM_R_X11Y106_SLICE_X14Y106_BO6;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_B3 = CLBLM_L_X10Y106_SLICE_X12Y106_AO6;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_B4 = CLBLM_L_X10Y108_SLICE_X13Y108_BO6;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_B5 = CLBLM_L_X10Y107_SLICE_X12Y107_AO6;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_B6 = CLBLM_L_X10Y108_SLICE_X13Y108_DO6;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_C1 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_C2 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_C3 = CLBLM_L_X8Y110_SLICE_X11Y110_DO6;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_C4 = CLBLM_L_X10Y109_SLICE_X12Y109_CO6;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_C5 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_C6 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_D1 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_D2 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_D3 = CLBLM_L_X8Y110_SLICE_X11Y110_DO6;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_D4 = CLBLM_L_X10Y109_SLICE_X12Y109_CO6;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_D5 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_D6 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_A1 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_A3 = CLBLL_L_X4Y103_SLICE_X5Y103_AO5;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_A4 = CLBLL_L_X4Y103_SLICE_X4Y103_BO6;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_A5 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_A6 = CLBLL_L_X4Y101_SLICE_X4Y101_CO6;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_B1 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_B2 = CLBLL_L_X4Y103_SLICE_X5Y103_BO5;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_B3 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_B4 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_B5 = CLBLL_L_X4Y102_SLICE_X5Y102_AO6;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_B6 = CLBLL_L_X4Y102_SLICE_X4Y102_DO6;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_C1 = CLBLL_L_X4Y102_SLICE_X5Y102_AO6;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_C2 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_C3 = CLBLL_L_X4Y103_SLICE_X5Y103_BO5;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_C4 = CLBLL_L_X4Y102_SLICE_X4Y102_DO6;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_C5 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_C6 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_D1 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_D2 = CLBLL_L_X4Y103_SLICE_X5Y103_AO5;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_D3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_D4 = CLBLL_L_X4Y101_SLICE_X4Y101_CO6;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_D5 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_D6 = CLBLL_L_X4Y103_SLICE_X4Y103_BO6;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_A1 = CLBLL_L_X4Y103_SLICE_X5Y103_BO5;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_A2 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_A3 = CLBLL_L_X4Y102_SLICE_X5Y102_AO6;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_A4 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_A5 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_A6 = 1'b1;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_B1 = CLBLL_L_X4Y102_SLICE_X5Y102_DO6;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_B2 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_B3 = CLBLM_R_X3Y102_SLICE_X3Y102_CO6;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_B4 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_B5 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_B6 = 1'b1;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_C1 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_C2 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_C3 = CLBLL_L_X4Y102_SLICE_X4Y102_BO5;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_C4 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_C5 = CLBLM_R_X5Y103_SLICE_X6Y103_AO6;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_C6 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_D1 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_D2 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_D3 = CLBLL_L_X4Y102_SLICE_X4Y102_BO5;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_D4 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_D5 = CLBLM_R_X5Y103_SLICE_X6Y103_AO6;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_D6 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_A1 = 1'b1;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_A2 = 1'b1;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_A3 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_A4 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_A5 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_A6 = 1'b1;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_B1 = CLBLM_L_X10Y109_SLICE_X12Y109_BO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_B2 = CLBLM_L_X10Y108_SLICE_X13Y108_CO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_B3 = CLBLM_R_X11Y106_SLICE_X14Y106_AO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_B4 = CLBLM_L_X10Y109_SLICE_X12Y109_DO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_B5 = CLBLM_L_X10Y108_SLICE_X13Y108_AO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_B6 = CLBLM_L_X10Y108_SLICE_X13Y108_AO5;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_C1 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_C2 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_C4 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_C5 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_C6 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_D1 = CLBLM_L_X10Y108_SLICE_X13Y108_AO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_D2 = CLBLM_R_X11Y106_SLICE_X14Y106_AO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_D3 = CLBLM_L_X10Y109_SLICE_X12Y109_DO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_D4 = CLBLM_L_X10Y108_SLICE_X13Y108_AO5;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_D5 = CLBLM_L_X10Y108_SLICE_X13Y108_CO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_D6 = CLBLM_L_X10Y109_SLICE_X12Y109_BO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_A1 = 1'b1;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_A2 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_A3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_A4 = 1'b1;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_A5 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_A6 = 1'b1;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_B1 = CLBLM_R_X7Y110_SLICE_X9Y110_AO5;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_B2 = CLBLM_L_X10Y107_SLICE_X12Y107_BO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_B3 = CLBLM_L_X10Y107_SLICE_X12Y107_AO5;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_B4 = CLBLM_L_X8Y110_SLICE_X10Y110_BO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_B5 = CLBLM_L_X10Y108_SLICE_X12Y108_AO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_B6 = CLBLM_L_X10Y107_SLICE_X12Y107_CO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_C1 = CLBLM_L_X10Y107_SLICE_X12Y107_AO5;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_C2 = CLBLM_L_X10Y107_SLICE_X12Y107_BO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_C3 = CLBLM_L_X10Y108_SLICE_X12Y108_AO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_C4 = CLBLM_L_X10Y107_SLICE_X12Y107_CO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_C5 = CLBLM_R_X7Y110_SLICE_X9Y110_AO5;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_C6 = CLBLM_L_X8Y110_SLICE_X10Y110_BO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_D1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_D2 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_D3 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_D4 = CLBLM_L_X10Y107_SLICE_X12Y107_CO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_D5 = CLBLM_L_X10Y107_SLICE_X12Y107_BO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_D6 = CLBLM_L_X8Y110_SLICE_X10Y110_BO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_A3 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_A1 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_A2 = CLBLL_L_X4Y104_SLICE_X5Y104_BO6;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_A3 = 1'b1;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_A4 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_A5 = CLBLL_L_X4Y103_SLICE_X5Y103_CO6;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_A6 = 1'b1;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_B1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_B2 = CLBLL_L_X4Y103_SLICE_X5Y103_AO5;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_B3 = CLBLL_L_X4Y101_SLICE_X4Y101_CO6;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_B4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_B5 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_B6 = 1'b1;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_C1 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_C2 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_C3 = CLBLL_L_X4Y103_SLICE_X4Y103_CO6;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_C4 = CLBLM_R_X3Y103_SLICE_X3Y103_AO5;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_C5 = CLBLL_L_X4Y103_SLICE_X4Y103_DO6;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_C6 = 1'b1;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_D1 = CLBLL_L_X4Y103_SLICE_X5Y103_CO6;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_D2 = CLBLL_L_X4Y104_SLICE_X5Y104_CO6;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_D3 = CLBLL_L_X4Y104_SLICE_X5Y104_BO6;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_D4 = CLBLL_L_X4Y105_SLICE_X4Y105_AO5;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_D5 = CLBLM_R_X3Y103_SLICE_X3Y103_AO6;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_D6 = CLBLL_L_X4Y104_SLICE_X4Y104_BO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_B1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_B2 = CLBLM_L_X8Y112_SLICE_X10Y112_DO6;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_A1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_A2 = 1'b1;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_A3 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_A4 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_A5 = 1'b1;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_A6 = 1'b1;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_B1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_B2 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_B3 = 1'b1;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_B4 = CLBLM_R_X5Y104_SLICE_X6Y104_AO6;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_B5 = CLBLM_R_X5Y104_SLICE_X6Y104_BO6;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_B6 = 1'b1;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_C1 = CLBLL_L_X4Y104_SLICE_X5Y104_AO6;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_C2 = CLBLM_R_X5Y105_SLICE_X6Y105_AO6;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_C3 = CLBLM_R_X7Y104_SLICE_X8Y104_AO6;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_C4 = CLBLL_L_X4Y104_SLICE_X5Y104_AO5;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_C5 = CLBLL_L_X4Y104_SLICE_X5Y104_BO5;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_C6 = CLBLM_R_X5Y105_SLICE_X7Y105_CO6;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_D1 = 1'b1;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_D2 = 1'b1;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_D3 = 1'b1;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_D4 = 1'b1;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_D5 = 1'b1;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_D6 = 1'b1;
  assign LIOI3_X0Y101_ILOGIC_X0Y102_D = LIOB33_X0Y101_IOB_X0Y102_I;
  assign LIOI3_X0Y101_ILOGIC_X0Y101_D = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_A1 = 1'b1;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_A2 = 1'b1;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_A3 = 1'b1;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_A4 = 1'b1;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_A5 = 1'b1;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_A6 = 1'b1;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_B1 = 1'b1;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_B2 = 1'b1;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_B3 = 1'b1;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_B4 = 1'b1;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_B5 = 1'b1;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_B6 = 1'b1;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_C1 = 1'b1;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_C2 = 1'b1;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_C3 = 1'b1;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_C4 = 1'b1;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_C5 = 1'b1;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_C6 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_A6 = 1'b1;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_D1 = 1'b1;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_D2 = 1'b1;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_D3 = 1'b1;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_D4 = 1'b1;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_D5 = 1'b1;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_D6 = 1'b1;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_A1 = CLBLM_L_X10Y109_SLICE_X12Y109_DO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_A2 = CLBLM_L_X10Y108_SLICE_X13Y108_CO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_A3 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_A4 = 1'b1;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_A5 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_A6 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_C3 = CLBLM_R_X5Y110_SLICE_X6Y110_AO5;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_B2 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_B3 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_B4 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_B5 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_B6 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_C1 = CLBLM_L_X10Y108_SLICE_X13Y108_CO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_C2 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_C3 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_C4 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_C5 = CLBLM_L_X10Y109_SLICE_X12Y109_DO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_C6 = CLBLM_L_X10Y109_SLICE_X12Y109_BO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_D1 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_D2 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_D3 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_D4 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_D5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_A1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_A2 = CLBLL_L_X4Y105_SLICE_X5Y105_BO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_A3 = 1'b1;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_A4 = CLBLM_R_X5Y105_SLICE_X6Y105_CO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_A5 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_A6 = 1'b1;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_D6 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_B1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_B2 = CLBLL_L_X4Y105_SLICE_X5Y105_BO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_B3 = CLBLL_L_X4Y105_SLICE_X5Y105_CO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_B4 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_B5 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_B6 = CLBLM_R_X5Y105_SLICE_X6Y105_CO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_C1 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_C2 = CLBLL_L_X4Y105_SLICE_X5Y105_CO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_C3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_C4 = CLBLL_L_X4Y105_SLICE_X4Y105_AO5;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_C5 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_C6 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_C1 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_C2 = 1'b1;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_D1 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_D2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_D3 = CLBLL_L_X4Y105_SLICE_X5Y105_BO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_D4 = CLBLL_L_X4Y104_SLICE_X5Y104_CO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_D5 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_D6 = CLBLM_R_X5Y105_SLICE_X6Y105_CO6;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_D3 = CLBLM_R_X7Y113_SLICE_X9Y113_CO6;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_D4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_C3 = 1'b1;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_A1 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_A2 = CLBLM_R_X5Y106_SLICE_X6Y106_BO6;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_A3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_A4 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_A5 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_A6 = CLBLM_R_X5Y106_SLICE_X6Y106_CO6;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_B1 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_B2 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_B3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_B4 = CLBLM_R_X5Y106_SLICE_X6Y106_BO6;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_B5 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_B6 = CLBLM_R_X5Y106_SLICE_X6Y106_CO6;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_C1 = CLBLM_R_X5Y105_SLICE_X6Y105_AO6;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_C2 = CLBLM_R_X7Y104_SLICE_X8Y104_AO6;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_C3 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_C4 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_C5 = CLBLM_R_X5Y105_SLICE_X7Y105_CO6;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_C6 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_D1 = 1'b1;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_D2 = 1'b1;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_D3 = 1'b1;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_D4 = 1'b1;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_D5 = 1'b1;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_D6 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_D4 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_C1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_C2 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_C3 = CLBLM_R_X7Y113_SLICE_X8Y113_AO6;
  assign CLBLM_L_X8Y100_SLICE_X11Y100_A1 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_L_X8Y100_SLICE_X11Y100_A2 = CLBLM_L_X8Y102_SLICE_X10Y102_DO6;
  assign CLBLM_L_X8Y100_SLICE_X11Y100_A3 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X8Y100_SLICE_X11Y100_A4 = CLBLM_L_X8Y100_SLICE_X11Y100_DO6;
  assign CLBLM_L_X8Y100_SLICE_X11Y100_A5 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_L_X8Y100_SLICE_X11Y100_A6 = CLBLM_L_X8Y100_SLICE_X11Y100_CO6;
  assign CLBLM_L_X8Y100_SLICE_X11Y100_B1 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_L_X8Y100_SLICE_X11Y100_B2 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_L_X8Y100_SLICE_X11Y100_B3 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X8Y100_SLICE_X11Y100_B4 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_L_X8Y100_SLICE_X11Y100_B5 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_L_X8Y100_SLICE_X11Y100_B6 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_L_X8Y100_SLICE_X11Y100_C1 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X8Y100_SLICE_X11Y100_C2 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_L_X8Y100_SLICE_X11Y100_C3 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_L_X8Y100_SLICE_X11Y100_C4 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_L_X8Y100_SLICE_X11Y100_C5 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_L_X8Y100_SLICE_X11Y100_C6 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_L_X8Y100_SLICE_X11Y100_D1 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X8Y100_SLICE_X11Y100_D2 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_L_X8Y100_SLICE_X11Y100_D3 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_L_X8Y100_SLICE_X11Y100_D4 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_L_X8Y100_SLICE_X11Y100_D5 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_L_X8Y100_SLICE_X11Y100_D6 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_L_X8Y100_SLICE_X10Y100_A1 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_L_X8Y100_SLICE_X10Y100_A2 = CLBLM_L_X8Y100_SLICE_X11Y100_DO6;
  assign CLBLM_L_X8Y100_SLICE_X10Y100_A3 = 1'b1;
  assign CLBLM_L_X8Y100_SLICE_X10Y100_A4 = CLBLM_L_X8Y102_SLICE_X10Y102_DO6;
  assign CLBLM_L_X8Y100_SLICE_X10Y100_A5 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X8Y100_SLICE_X10Y100_A6 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_D4 = CLBLM_R_X5Y112_SLICE_X6Y112_CO6;
  assign CLBLM_L_X8Y100_SLICE_X10Y100_B1 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_L_X8Y100_SLICE_X10Y100_B2 = CLBLM_L_X8Y102_SLICE_X10Y102_AO5;
  assign CLBLM_L_X8Y100_SLICE_X10Y100_B3 = CLBLM_L_X8Y100_SLICE_X11Y100_AO6;
  assign CLBLM_L_X8Y100_SLICE_X10Y100_B4 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X8Y100_SLICE_X10Y100_B5 = CLBLM_L_X8Y100_SLICE_X10Y100_AO6;
  assign CLBLM_L_X8Y100_SLICE_X10Y100_B6 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_A1 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_A2 = CLBLM_R_X5Y102_SLICE_X6Y102_DO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_A3 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_A4 = CLBLM_R_X7Y102_SLICE_X9Y102_AO5;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_A5 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_A6 = 1'b1;
  assign CLBLM_L_X8Y100_SLICE_X10Y100_C1 = CLBLL_L_X4Y103_SLICE_X5Y103_BO6;
  assign CLBLM_L_X8Y100_SLICE_X10Y100_C2 = CLBLM_L_X8Y100_SLICE_X11Y100_CO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_B1 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_B2 = CLBLM_R_X5Y106_SLICE_X7Y106_BO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_B3 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_B4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_B5 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_B6 = CLBLM_R_X7Y106_SLICE_X8Y106_CO6;
  assign CLBLM_L_X8Y100_SLICE_X10Y100_C4 = CLBLL_L_X4Y101_SLICE_X5Y101_AO6;
  assign CLBLM_L_X8Y100_SLICE_X10Y100_C5 = CLBLM_L_X8Y102_SLICE_X10Y102_DO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_C1 = CLBLM_R_X5Y106_SLICE_X7Y106_BO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_C2 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_C3 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_L_X8Y100_SLICE_X10Y100_D4 = CLBLL_L_X4Y101_SLICE_X5Y101_AO6;
  assign CLBLM_L_X8Y100_SLICE_X10Y100_D5 = CLBLM_L_X8Y102_SLICE_X10Y102_DO6;
  assign CLBLM_L_X8Y100_SLICE_X10Y100_D6 = CLBLM_R_X3Y100_SLICE_X3Y100_AO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_C4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_C6 = CLBLM_R_X7Y106_SLICE_X8Y106_CO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_C5 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_L_X8Y100_SLICE_X10Y100_D2 = CLBLM_L_X8Y100_SLICE_X11Y100_CO6;
  assign CLBLM_L_X8Y100_SLICE_X10Y100_D3 = CLBLM_L_X8Y100_SLICE_X11Y100_DO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_D1 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_D2 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_D3 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_D4 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_D5 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_D6 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_A1 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_A2 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_A3 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_A4 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_A5 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_A6 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_B1 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_B2 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_B3 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_B4 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_B5 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_B6 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_C1 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_C2 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_C3 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_C4 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_C5 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_C6 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_D1 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_D2 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_D3 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_D4 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_D5 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_D6 = 1'b1;
  assign CLBLM_L_X8Y101_SLICE_X11Y101_A1 = CLBLM_L_X10Y104_SLICE_X13Y104_AO6;
  assign CLBLM_L_X8Y101_SLICE_X11Y101_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y101_SLICE_X11Y101_A3 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X8Y101_SLICE_X11Y101_A4 = CLBLM_L_X8Y100_SLICE_X11Y100_CO6;
  assign CLBLM_L_X8Y101_SLICE_X11Y101_A5 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_L_X8Y101_SLICE_X11Y101_A6 = 1'b1;
  assign CLBLM_L_X8Y101_SLICE_X11Y101_B1 = CLBLM_L_X8Y101_SLICE_X11Y101_DO6;
  assign CLBLM_L_X8Y101_SLICE_X11Y101_B2 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X8Y101_SLICE_X11Y101_B3 = CLBLM_L_X8Y100_SLICE_X11Y100_BO6;
  assign CLBLM_L_X8Y101_SLICE_X11Y101_B4 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_L_X8Y101_SLICE_X11Y101_B5 = CLBLM_L_X8Y100_SLICE_X11Y100_CO6;
  assign CLBLM_L_X8Y101_SLICE_X11Y101_B6 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X8Y101_SLICE_X11Y101_C1 = CLBLM_L_X8Y100_SLICE_X11Y100_CO6;
  assign CLBLM_L_X8Y101_SLICE_X11Y101_C2 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X8Y101_SLICE_X11Y101_C3 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X8Y101_SLICE_X11Y101_C4 = CLBLM_L_X8Y100_SLICE_X11Y100_BO6;
  assign CLBLM_L_X8Y101_SLICE_X11Y101_C5 = CLBLM_L_X8Y101_SLICE_X11Y101_DO6;
  assign CLBLM_L_X8Y101_SLICE_X11Y101_C6 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_L_X8Y101_SLICE_X11Y101_D1 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X8Y101_SLICE_X11Y101_D2 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_L_X8Y101_SLICE_X11Y101_D3 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_L_X8Y101_SLICE_X11Y101_D4 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X8Y101_SLICE_X11Y101_D5 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_L_X8Y101_SLICE_X11Y101_D6 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_L_X8Y101_SLICE_X10Y101_A1 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_L_X8Y101_SLICE_X10Y101_A2 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X8Y101_SLICE_X10Y101_A3 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_L_X8Y101_SLICE_X10Y101_A4 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_L_X8Y101_SLICE_X10Y101_A5 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_L_X8Y101_SLICE_X10Y101_A6 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X8Y101_SLICE_X10Y101_B1 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_L_X8Y101_SLICE_X10Y101_B2 = CLBLM_L_X8Y100_SLICE_X10Y100_AO5;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_A1 = CLBLL_L_X4Y110_SLICE_X4Y110_BO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_A2 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_L_X8Y101_SLICE_X10Y101_B5 = CLBLM_L_X8Y101_SLICE_X11Y101_CO6;
  assign CLBLM_L_X8Y101_SLICE_X10Y101_B6 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_A3 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_A4 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_A5 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_A6 = 1'b1;
  assign CLBLM_L_X8Y101_SLICE_X10Y101_C1 = CLBLM_L_X8Y100_SLICE_X11Y100_AO6;
  assign CLBLM_L_X8Y101_SLICE_X10Y101_C2 = CLBLM_L_X10Y102_SLICE_X12Y102_DO6;
  assign CLBLM_L_X8Y101_SLICE_X10Y101_C3 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_L_X8Y101_SLICE_X10Y101_C4 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X8Y101_SLICE_X10Y101_C5 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X8Y101_SLICE_X10Y101_C6 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_B5 = CLBLL_L_X4Y108_SLICE_X4Y108_AO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_B6 = CLBLL_L_X4Y109_SLICE_X4Y109_CO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_B1 = CLBLL_L_X2Y105_SLICE_X1Y105_AO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_B2 = CLBLL_L_X4Y107_SLICE_X5Y107_BO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_B3 = CLBLM_R_X3Y106_SLICE_X3Y106_AO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_B4 = CLBLL_L_X4Y107_SLICE_X5Y107_AO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_C3 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_C5 = CLBLM_R_X5Y108_SLICE_X6Y108_DO6;
  assign CLBLM_L_X8Y101_SLICE_X10Y101_D1 = CLBLM_L_X8Y100_SLICE_X11Y100_AO6;
  assign CLBLM_L_X8Y101_SLICE_X10Y101_D2 = CLBLM_L_X10Y102_SLICE_X12Y102_DO6;
  assign CLBLM_L_X8Y101_SLICE_X10Y101_D3 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X8Y101_SLICE_X10Y101_D4 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X8Y101_SLICE_X10Y101_D5 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_L_X8Y101_SLICE_X10Y101_D6 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_C4 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_C6 = CLBLL_L_X4Y108_SLICE_X5Y108_BO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_D1 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_D2 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_D3 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_D4 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_D5 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_D6 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_A1 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_A2 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_A3 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_A4 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_A5 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_A6 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_B2 = CLBLL_L_X4Y110_SLICE_X5Y110_BO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_B3 = CLBLL_L_X4Y110_SLICE_X5Y110_AO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_B1 = CLBLM_R_X7Y108_SLICE_X8Y108_DO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_B2 = CLBLL_L_X4Y109_SLICE_X5Y109_BO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_B3 = CLBLM_R_X7Y107_SLICE_X8Y107_AO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_B4 = CLBLL_L_X4Y107_SLICE_X4Y107_AO5;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_B5 = CLBLL_L_X4Y106_SLICE_X4Y106_AO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_B6 = CLBLM_R_X7Y108_SLICE_X8Y108_CO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_B5 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_C1 = CLBLM_R_X5Y107_SLICE_X6Y107_BO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_C2 = CLBLL_L_X4Y107_SLICE_X5Y107_AO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_C3 = CLBLM_R_X7Y106_SLICE_X8Y106_BO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_C4 = CLBLL_L_X4Y107_SLICE_X5Y107_AO5;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_C5 = CLBLL_L_X4Y108_SLICE_X4Y108_BO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_C6 = CLBLM_R_X5Y107_SLICE_X7Y107_BO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_D1 = CLBLM_R_X5Y107_SLICE_X6Y107_BO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_D2 = CLBLM_R_X5Y107_SLICE_X7Y107_DO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_D3 = CLBLL_L_X4Y107_SLICE_X5Y107_AO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_D4 = CLBLL_L_X4Y107_SLICE_X5Y107_AO5;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_D5 = CLBLL_L_X4Y108_SLICE_X4Y108_BO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_D6 = CLBLL_L_X4Y103_SLICE_X5Y103_AO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_C4 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_C5 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_D5 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_A1 = CLBLM_L_X8Y102_SLICE_X11Y102_DO6;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_A2 = CLBLM_L_X10Y103_SLICE_X13Y103_CO6;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_A3 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_A4 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_A6 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_B1 = CLBLM_L_X8Y102_SLICE_X11Y102_DO6;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_B2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_B3 = CLBLM_L_X8Y102_SLICE_X10Y102_AO6;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_B4 = CLBLM_L_X8Y103_SLICE_X11Y103_BO6;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_B5 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_B6 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_C2 = CLBLM_L_X10Y103_SLICE_X13Y103_CO6;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_C3 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_C4 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_C5 = CLBLM_L_X8Y102_SLICE_X11Y102_DO6;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_C6 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_D1 = CLBLM_L_X8Y101_SLICE_X10Y101_AO6;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_D2 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_D3 = CLBLM_L_X8Y102_SLICE_X10Y102_DO6;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_D4 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_D5 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_D6 = CLBLM_L_X10Y102_SLICE_X13Y102_AO6;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_A1 = 1'b1;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_A2 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_A3 = CLBLM_L_X10Y102_SLICE_X13Y102_AO6;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_A4 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_A5 = CLBLM_L_X8Y101_SLICE_X10Y101_AO6;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_A6 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_A1 = CLBLM_R_X7Y108_SLICE_X8Y108_DO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_A2 = CLBLM_R_X5Y108_SLICE_X7Y108_BO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_A3 = CLBLM_R_X5Y109_SLICE_X6Y109_DO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_A4 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_A5 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_A6 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_B1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_B2 = CLBLM_L_X8Y100_SLICE_X10Y100_BO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_B1 = CLBLM_R_X7Y108_SLICE_X8Y108_DO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_B2 = CLBLM_R_X5Y108_SLICE_X7Y108_BO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_B3 = CLBLM_R_X5Y109_SLICE_X6Y109_DO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_B4 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_B5 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_B6 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_B5 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_B6 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_C1 = CLBLM_L_X10Y102_SLICE_X12Y102_AO5;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_C2 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_C3 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_C2 = CLBLM_L_X8Y101_SLICE_X11Y101_CO6;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_C3 = CLBLM_L_X8Y100_SLICE_X10Y100_DO6;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_C4 = CLBLM_L_X8Y103_SLICE_X11Y103_AO5;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_C5 = CLBLM_L_X10Y102_SLICE_X12Y102_DO6;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_C6 = CLBLM_L_X8Y100_SLICE_X10Y100_CO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_C1 = CLBLM_R_X5Y107_SLICE_X7Y107_AO6;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_D1 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_D2 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_D3 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_D4 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_D5 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_D6 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_D1 = CLBLL_L_X4Y106_SLICE_X4Y106_BO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_D2 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_D3 = CLBLL_L_X4Y108_SLICE_X5Y108_BO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_D4 = CLBLM_R_X5Y107_SLICE_X6Y107_CO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_D5 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_D6 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_A1 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_A2 = CLBLL_L_X4Y108_SLICE_X4Y108_BO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_A3 = CLBLM_R_X5Y107_SLICE_X7Y107_AO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_A4 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_A5 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_A6 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_A1 = 1'b1;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_A2 = 1'b1;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_A3 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_B1 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_B2 = CLBLM_R_X7Y106_SLICE_X8Y106_DO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_B3 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_B4 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_B5 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_B6 = CLBLM_R_X5Y107_SLICE_X7Y107_BO6;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_B1 = 1'b1;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_B2 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_C1 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_C2 = CLBLM_R_X5Y107_SLICE_X7Y107_BO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_C3 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_C4 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_C5 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_C6 = CLBLM_R_X7Y106_SLICE_X8Y106_DO6;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_C1 = 1'b1;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_C2 = 1'b1;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_C3 = 1'b1;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_C4 = 1'b1;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_C5 = 1'b1;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_C6 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_D1 = CLBLL_L_X4Y108_SLICE_X5Y108_AO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_D2 = CLBLL_L_X4Y107_SLICE_X5Y107_DO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_D3 = CLBLL_L_X4Y109_SLICE_X5Y109_CO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_D4 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_D5 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_D6 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_D4 = 1'b1;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_D5 = 1'b1;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_D6 = 1'b1;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_D3 = 1'b1;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_A1 = 1'b1;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_A2 = 1'b1;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_A3 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_A4 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_A5 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_A6 = 1'b1;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_B1 = CLBLM_L_X10Y109_SLICE_X12Y109_BO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_B2 = CLBLM_R_X5Y102_SLICE_X6Y102_AO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_B3 = CLBLM_L_X10Y104_SLICE_X13Y104_AO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_B4 = CLBLM_L_X10Y105_SLICE_X13Y105_AO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_B5 = CLBLM_R_X11Y106_SLICE_X14Y106_AO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_B6 = CLBLM_R_X11Y106_SLICE_X14Y106_AO5;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_C1 = CLBLM_R_X11Y106_SLICE_X14Y106_AO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_C2 = CLBLM_L_X10Y104_SLICE_X13Y104_AO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_C3 = CLBLM_R_X5Y102_SLICE_X6Y102_AO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_C4 = CLBLM_R_X11Y106_SLICE_X14Y106_AO5;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_C5 = CLBLM_L_X10Y109_SLICE_X12Y109_BO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_C6 = CLBLM_L_X10Y105_SLICE_X13Y105_AO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_D1 = CLBLM_L_X10Y104_SLICE_X13Y104_AO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_D2 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_D3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_D4 = CLBLM_L_X10Y105_SLICE_X13Y105_AO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_D5 = CLBLM_L_X10Y109_SLICE_X12Y109_BO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_D6 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_A1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_A2 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_A3 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_A4 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_A5 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_A6 = 1'b1;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_B1 = CLBLM_L_X8Y103_SLICE_X11Y103_DO6;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_B2 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_B3 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_B4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_B5 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_B6 = CLBLM_L_X8Y103_SLICE_X11Y103_AO6;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_C1 = CLBLM_L_X8Y102_SLICE_X11Y102_CO6;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_C2 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_C3 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_C5 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_C6 = CLBLM_L_X8Y100_SLICE_X10Y100_BO6;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_D1 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_D2 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_D3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_D4 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_D5 = 1'b1;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_D6 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_A1 = 1'b1;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_A3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_A4 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_A5 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A1 = CLBLL_L_X4Y110_SLICE_X4Y110_DO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_A6 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A3 = CLBLM_R_X5Y109_SLICE_X6Y109_BO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A4 = CLBLM_R_X5Y109_SLICE_X6Y109_CO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A5 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A6 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_B1 = CLBLM_L_X8Y101_SLICE_X10Y101_DO6;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_B2 = CLBLM_R_X7Y100_SLICE_X8Y100_AO5;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_B3 = CLBLM_L_X8Y102_SLICE_X11Y102_CO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B4 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B5 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B6 = CLBLL_L_X4Y109_SLICE_X4Y109_CO6;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_B4 = CLBLM_L_X8Y102_SLICE_X10Y102_CO6;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_B5 = CLBLM_L_X8Y103_SLICE_X10Y103_AO6;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_B6 = CLBLM_L_X8Y103_SLICE_X10Y103_AO5;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B2 = CLBLM_R_X5Y108_SLICE_X6Y108_BO6;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_C1 = CLBLM_L_X8Y102_SLICE_X11Y102_CO6;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_C2 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_C3 = CLBLM_L_X8Y101_SLICE_X10Y101_DO6;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_C4 = CLBLM_L_X8Y102_SLICE_X10Y102_CO6;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_C5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_C6 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C2 = CLBLL_L_X4Y109_SLICE_X5Y109_AO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C3 = CLBLL_L_X4Y110_SLICE_X4Y110_DO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C5 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C4 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C6 = CLBLM_R_X5Y109_SLICE_X6Y109_CO6;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_D1 = CLBLM_L_X8Y103_SLICE_X10Y103_AO6;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_D2 = CLBLM_L_X8Y102_SLICE_X10Y102_CO6;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_D3 = CLBLM_L_X8Y101_SLICE_X10Y101_DO6;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_D4 = CLBLM_L_X8Y103_SLICE_X10Y103_AO5;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_D5 = CLBLM_L_X8Y102_SLICE_X11Y102_CO6;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_D6 = CLBLM_R_X7Y100_SLICE_X8Y100_AO5;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D1 = CLBLL_L_X4Y108_SLICE_X5Y108_AO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D2 = CLBLL_L_X4Y109_SLICE_X5Y109_CO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D3 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D4 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D5 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D6 = CLBLL_L_X4Y107_SLICE_X5Y107_CO6;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_C5 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_C6 = CLBLM_R_X3Y110_SLICE_X2Y110_AO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A1 = CLBLM_R_X5Y110_SLICE_X6Y110_CO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A2 = CLBLM_R_X5Y110_SLICE_X7Y110_BO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A3 = CLBLM_R_X7Y108_SLICE_X8Y108_AO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A4 = CLBLM_R_X5Y109_SLICE_X6Y109_AO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A5 = CLBLM_R_X5Y108_SLICE_X6Y108_AO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A6 = CLBLM_R_X5Y111_SLICE_X7Y111_DO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B1 = CLBLM_R_X5Y110_SLICE_X6Y110_CO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B2 = CLBLM_R_X5Y110_SLICE_X7Y110_BO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B3 = CLBLM_R_X5Y108_SLICE_X6Y108_AO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B4 = CLBLM_R_X5Y109_SLICE_X6Y109_AO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B5 = CLBLM_R_X7Y108_SLICE_X8Y108_AO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B6 = CLBLM_R_X5Y111_SLICE_X7Y111_DO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C1 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C2 = CLBLL_L_X4Y109_SLICE_X4Y109_CO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C3 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C4 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C5 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C6 = CLBLM_R_X5Y108_SLICE_X6Y108_BO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_B5 = CLBLM_L_X8Y111_SLICE_X10Y111_AO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_B6 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D1 = CLBLL_L_X4Y108_SLICE_X5Y108_AO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D2 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D3 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D4 = CLBLL_L_X4Y109_SLICE_X5Y109_CO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D5 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D6 = CLBLL_L_X4Y107_SLICE_X5Y107_DO6;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_D4 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_D5 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_C1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_D6 = CLBLM_R_X3Y106_SLICE_X2Y106_CO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_C2 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_C3 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign LIOI3_X0Y105_ILOGIC_X0Y106_D = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_C4 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign LIOI3_X0Y105_ILOGIC_X0Y105_D = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_C5 = CLBLM_R_X7Y112_SLICE_X8Y112_BO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_C6 = CLBLM_R_X7Y112_SLICE_X9Y112_BO6;
  assign LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y114_D = LIOB33_X0Y113_IOB_X0Y114_I;
  assign LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y113_D = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_D1 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_D2 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_D5 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_D6 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_A1 = CLBLM_L_X10Y104_SLICE_X12Y104_CO6;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_A2 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_A3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_A4 = CLBLM_L_X10Y103_SLICE_X12Y103_DO6;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_A5 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_A6 = CLBLM_L_X10Y105_SLICE_X13Y105_BO6;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_B1 = CLBLM_L_X10Y105_SLICE_X13Y105_BO6;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_B2 = CLBLM_L_X10Y103_SLICE_X12Y103_CO6;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_B3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_B4 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_B5 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_B6 = CLBLM_L_X10Y104_SLICE_X12Y104_CO6;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_C1 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_C2 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_C3 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_C4 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_C5 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_C6 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_D1 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_D2 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_D3 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_D4 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_D5 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_D6 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_A1 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_A2 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_A3 = CLBLL_L_X4Y110_SLICE_X5Y110_AO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_A4 = CLBLM_R_X3Y110_SLICE_X3Y110_AO6;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_A3 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_A5 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_A4 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_A5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_A6 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_A6 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_B1 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_A1 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_A2 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_B4 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_B6 = CLBLM_R_X3Y110_SLICE_X3Y110_AO6;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_B1 = CLBLM_L_X10Y104_SLICE_X12Y104_DO6;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_B2 = CLBLM_L_X8Y103_SLICE_X10Y103_CO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_C1 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_C2 = CLBLL_L_X4Y110_SLICE_X5Y110_AO6;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_B3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_B4 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_B6 = CLBLM_L_X8Y103_SLICE_X11Y103_CO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_C3 = CLBLL_L_X4Y110_SLICE_X5Y110_DO6;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_C1 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_C2 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_C3 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_C4 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_C5 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_C6 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_C6 = CLBLM_R_X3Y110_SLICE_X3Y110_AO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_D1 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_D2 = CLBLM_R_X5Y110_SLICE_X6Y110_AO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_D3 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_D4 = CLBLL_L_X4Y111_SLICE_X4Y111_CO6;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_D1 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_D2 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_D3 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_D4 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_D5 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_D6 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_D6 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_A1 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_A2 = CLBLM_R_X5Y110_SLICE_X6Y110_AO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_A3 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_A4 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_A5 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_A6 = CLBLL_L_X4Y111_SLICE_X4Y111_CO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_B1 = CLBLM_R_X5Y110_SLICE_X6Y110_CO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_B2 = CLBLM_R_X5Y109_SLICE_X6Y109_AO5;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_B3 = CLBLM_R_X5Y109_SLICE_X6Y109_AO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_B4 = CLBLM_R_X5Y110_SLICE_X7Y110_BO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_B5 = CLBLL_L_X4Y110_SLICE_X5Y110_CO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_B6 = CLBLL_L_X4Y111_SLICE_X4Y111_CO6;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_D5 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_D6 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_C1 = CLBLM_R_X5Y112_SLICE_X6Y112_DO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_C2 = CLBLM_R_X3Y111_SLICE_X3Y111_AO5;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_C3 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_C4 = CLBLM_R_X7Y111_SLICE_X8Y111_BO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_C5 = CLBLL_L_X4Y111_SLICE_X5Y111_DO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_C6 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_D1 = CLBLL_L_X4Y110_SLICE_X5Y110_CO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_D2 = CLBLM_R_X5Y111_SLICE_X7Y111_CO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_D3 = CLBLM_R_X5Y109_SLICE_X6Y109_AO5;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_D4 = CLBLL_L_X4Y111_SLICE_X4Y111_CO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_D5 = CLBLM_R_X5Y109_SLICE_X6Y109_AO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_D6 = CLBLL_L_X4Y110_SLICE_X4Y110_AO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_D2 = CLBLM_R_X7Y111_SLICE_X8Y111_AO6;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_A3 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_B6 = CLBLM_R_X5Y111_SLICE_X7Y111_BO6;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_B1 = CLBLM_R_X7Y105_SLICE_X9Y105_AO5;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_B2 = CLBLM_L_X8Y103_SLICE_X10Y103_BO6;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_B6 = CLBLM_L_X8Y105_SLICE_X10Y105_AO5;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_C5 = CLBLM_R_X5Y113_SLICE_X6Y113_DO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_C6 = CLBLM_R_X5Y110_SLICE_X7Y110_AO5;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_A1 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_A2 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_A3 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_A4 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_A5 = CLBLM_L_X8Y104_SLICE_X11Y104_AO6;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_A6 = CLBLM_L_X8Y105_SLICE_X11Y105_CO6;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_B1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_B2 = CLBLM_L_X10Y105_SLICE_X13Y105_BO6;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_B3 = CLBLM_L_X10Y104_SLICE_X12Y104_CO6;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_B4 = CLBLM_L_X10Y103_SLICE_X12Y103_CO6;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_B5 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_B6 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_C1 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_C2 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_C3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_C4 = CLBLM_L_X10Y105_SLICE_X12Y105_CO6;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_C5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_C6 = CLBLM_L_X10Y107_SLICE_X13Y107_CO6;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_D1 = CLBLM_L_X8Y104_SLICE_X11Y104_AO6;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_D2 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_D3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_D4 = CLBLM_L_X8Y105_SLICE_X11Y105_CO6;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_D5 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_D6 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_A1 = CLBLL_L_X4Y112_SLICE_X4Y112_DO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_A2 = CLBLL_L_X4Y111_SLICE_X5Y111_BO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_A3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_A4 = CLBLL_L_X4Y111_SLICE_X4Y111_BO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_A5 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_A6 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_A1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_A2 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_B1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_A5 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_B2 = CLBLL_L_X4Y112_SLICE_X5Y112_DO6;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_A6 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_B3 = CLBLL_L_X4Y111_SLICE_X5Y111_AO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_B4 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_B5 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_B6 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_A4 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_B4 = CLBLM_L_X10Y103_SLICE_X12Y103_BO6;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_B5 = CLBLM_L_X10Y105_SLICE_X12Y105_BO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_C1 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_C2 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_C3 = CLBLL_L_X4Y111_SLICE_X5Y111_BO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_C4 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_C5 = CLBLL_L_X4Y111_SLICE_X4Y111_DO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_C6 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_B3 = CLBLM_L_X10Y103_SLICE_X12Y103_CO6;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_C2 = CLBLM_L_X10Y103_SLICE_X12Y103_CO6;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_C3 = CLBLM_L_X10Y105_SLICE_X12Y105_AO6;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_C4 = CLBLM_L_X8Y105_SLICE_X10Y105_AO5;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_C5 = CLBLM_L_X10Y107_SLICE_X13Y107_CO6;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_C6 = CLBLM_R_X7Y105_SLICE_X9Y105_AO6;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_C1 = CLBLM_L_X10Y105_SLICE_X12Y105_BO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_D1 = CLBLM_R_X3Y112_SLICE_X3Y112_DO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_D2 = CLBLM_R_X3Y111_SLICE_X3Y111_BO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_D3 = CLBLL_L_X4Y112_SLICE_X5Y112_BO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_D4 = CLBLL_L_X4Y112_SLICE_X5Y112_AO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_D5 = CLBLM_R_X3Y111_SLICE_X3Y111_BO5;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_D6 = CLBLM_R_X3Y111_SLICE_X3Y111_CO5;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_D1 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_D2 = CLBLM_L_X10Y105_SLICE_X12Y105_CO6;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_D3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_D4 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_D5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_D6 = CLBLM_L_X10Y107_SLICE_X13Y107_CO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_A1 = CLBLL_L_X4Y113_SLICE_X5Y113_AO5;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_A2 = CLBLM_R_X5Y110_SLICE_X6Y110_BO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_A3 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_A4 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_A5 = CLBLM_R_X5Y112_SLICE_X6Y112_AO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_A6 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_B1 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_B2 = CLBLM_R_X5Y112_SLICE_X6Y112_BO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_B3 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_B4 = CLBLL_L_X4Y112_SLICE_X5Y112_DO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_B5 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_B6 = CLBLL_L_X4Y111_SLICE_X5Y111_CO6;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_D1 = CLBLL_L_X2Y108_SLICE_X1Y108_DO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_C1 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_C2 = CLBLM_R_X5Y111_SLICE_X6Y111_BO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_C3 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_C4 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_C5 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_C6 = CLBLM_R_X5Y110_SLICE_X6Y110_BO6;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_T1 = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_D1 = CLBLM_R_X3Y110_SLICE_X2Y110_CO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_D1 = CLBLM_R_X3Y111_SLICE_X3Y111_CO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_D2 = CLBLL_L_X4Y112_SLICE_X5Y112_DO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_D3 = CLBLM_R_X3Y111_SLICE_X3Y111_BO5;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_D4 = CLBLL_L_X4Y111_SLICE_X5Y111_CO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_D5 = CLBLM_R_X5Y112_SLICE_X7Y112_AO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_D6 = CLBLM_R_X5Y112_SLICE_X6Y112_BO6;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_D1 = CLBLL_L_X2Y109_SLICE_X1Y109_AO6;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_T1 = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_T1 = 1'b1;
  assign LIOI3_X0Y109_ILOGIC_X0Y110_D = LIOB33_X0Y109_IOB_X0Y110_I;
  assign LIOI3_X0Y109_ILOGIC_X0Y109_D = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_A1 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_A2 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_A3 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_A4 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_A5 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_A6 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_B1 = CLBLM_L_X8Y105_SLICE_X11Y105_BO6;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_B2 = CLBLM_L_X8Y106_SLICE_X11Y106_AO5;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_B3 = CLBLM_L_X8Y106_SLICE_X10Y106_AO6;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_B4 = CLBLM_L_X8Y105_SLICE_X10Y105_BO6;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_B5 = CLBLM_L_X8Y106_SLICE_X11Y106_AO6;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_B6 = CLBLM_L_X8Y105_SLICE_X11Y105_CO6;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_C1 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_C2 = CLBLM_L_X8Y105_SLICE_X10Y105_BO6;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_C3 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_C4 = CLBLM_L_X8Y105_SLICE_X11Y105_CO6;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_C5 = CLBLM_L_X8Y105_SLICE_X11Y105_BO6;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_C6 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_D1 = CLBLM_L_X8Y106_SLICE_X11Y106_AO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_A1 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_A2 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_D4 = CLBLM_L_X8Y105_SLICE_X11Y105_CO6;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_D5 = CLBLM_L_X8Y106_SLICE_X10Y106_AO6;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_D6 = CLBLM_L_X8Y106_SLICE_X11Y106_AO5;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_A3 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_A4 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_A5 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_A6 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_B1 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_A1 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_A2 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_A3 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_A4 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_A5 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_B2 = CLBLL_L_X4Y112_SLICE_X5Y112_BO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_B3 = CLBLL_L_X4Y112_SLICE_X5Y112_AO6;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_A6 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_C1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_C2 = CLBLL_L_X4Y112_SLICE_X5Y112_CO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_C3 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_C4 = CLBLM_R_X3Y112_SLICE_X3Y112_DO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_C5 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_C6 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_B1 = CLBLM_R_X7Y106_SLICE_X9Y106_AO5;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_B2 = CLBLM_L_X8Y107_SLICE_X10Y107_DO6;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_B3 = CLBLM_L_X8Y106_SLICE_X11Y106_AO5;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_B4 = CLBLM_L_X8Y105_SLICE_X10Y105_DO6;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_B5 = CLBLM_L_X8Y105_SLICE_X10Y105_CO6;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_C1 = CLBLM_L_X8Y105_SLICE_X10Y105_CO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_D1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_D2 = CLBLL_L_X4Y112_SLICE_X5Y112_CO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_D3 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_D4 = CLBLM_R_X3Y112_SLICE_X3Y112_DO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_D5 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_D6 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_C2 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_C3 = CLBLM_L_X8Y107_SLICE_X10Y107_DO6;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_C4 = CLBLM_L_X8Y105_SLICE_X10Y105_DO6;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_C5 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_C6 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_D1 = CLBLM_L_X8Y105_SLICE_X10Y105_CO6;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_D2 = CLBLM_L_X8Y106_SLICE_X11Y106_AO5;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_D3 = CLBLM_L_X8Y107_SLICE_X10Y107_DO6;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_D4 = CLBLM_L_X8Y106_SLICE_X10Y106_AO5;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_D5 = CLBLM_R_X7Y106_SLICE_X9Y106_AO5;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_D6 = CLBLM_L_X8Y105_SLICE_X10Y105_DO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_A1 = CLBLL_L_X4Y112_SLICE_X4Y112_AO5;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_A2 = CLBLM_R_X5Y113_SLICE_X6Y113_BO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_A3 = CLBLL_L_X4Y112_SLICE_X4Y112_AO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_A4 = CLBLM_R_X5Y111_SLICE_X6Y111_AO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_A5 = CLBLM_R_X5Y111_SLICE_X6Y111_BO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_A6 = CLBLM_R_X3Y113_SLICE_X3Y113_CO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_B1 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_B2 = CLBLM_R_X5Y111_SLICE_X6Y111_CO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_B3 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_B4 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_B5 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_B6 = CLBLM_R_X3Y113_SLICE_X3Y113_CO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_C1 = CLBLL_L_X4Y113_SLICE_X5Y113_AO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_C2 = CLBLM_R_X5Y111_SLICE_X6Y111_CO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_C3 = CLBLM_R_X3Y113_SLICE_X2Y113_BO5;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_C4 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_C5 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_C6 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_D1 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_D2 = CLBLM_R_X5Y111_SLICE_X6Y111_CO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_D3 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_D4 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_D5 = CLBLM_R_X3Y113_SLICE_X3Y113_CO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_D6 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X7Y100_SLICE_X9Y100_A1 = 1'b1;
  assign CLBLM_R_X7Y100_SLICE_X9Y100_A2 = 1'b1;
  assign CLBLM_R_X7Y100_SLICE_X9Y100_A3 = 1'b1;
  assign CLBLM_R_X7Y100_SLICE_X9Y100_A4 = 1'b1;
  assign CLBLM_R_X7Y100_SLICE_X9Y100_A5 = 1'b1;
  assign CLBLM_R_X7Y100_SLICE_X9Y100_A6 = 1'b1;
  assign CLBLM_R_X7Y100_SLICE_X9Y100_B1 = 1'b1;
  assign CLBLM_R_X7Y100_SLICE_X9Y100_B2 = 1'b1;
  assign CLBLM_R_X7Y100_SLICE_X9Y100_B3 = 1'b1;
  assign CLBLM_R_X7Y100_SLICE_X9Y100_B4 = 1'b1;
  assign CLBLM_R_X7Y100_SLICE_X9Y100_B5 = 1'b1;
  assign CLBLM_R_X7Y100_SLICE_X9Y100_B6 = 1'b1;
  assign CLBLM_R_X7Y100_SLICE_X9Y100_C1 = 1'b1;
  assign CLBLM_R_X7Y100_SLICE_X9Y100_C2 = 1'b1;
  assign CLBLM_R_X7Y100_SLICE_X9Y100_C3 = 1'b1;
  assign CLBLM_R_X7Y100_SLICE_X9Y100_C4 = 1'b1;
  assign CLBLM_R_X7Y100_SLICE_X9Y100_C5 = 1'b1;
  assign CLBLM_R_X7Y100_SLICE_X9Y100_C6 = 1'b1;
  assign CLBLM_R_X7Y100_SLICE_X9Y100_D1 = 1'b1;
  assign CLBLM_R_X7Y100_SLICE_X9Y100_D2 = 1'b1;
  assign CLBLM_R_X7Y100_SLICE_X9Y100_D3 = 1'b1;
  assign CLBLM_R_X7Y100_SLICE_X9Y100_D4 = 1'b1;
  assign CLBLM_R_X7Y100_SLICE_X9Y100_D5 = 1'b1;
  assign CLBLM_R_X7Y100_SLICE_X9Y100_D6 = 1'b1;
  assign CLBLM_R_X7Y100_SLICE_X8Y100_A1 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X7Y100_SLICE_X8Y100_A2 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X7Y100_SLICE_X8Y100_A3 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X7Y100_SLICE_X8Y100_A4 = 1'b1;
  assign CLBLM_R_X7Y100_SLICE_X8Y100_A5 = 1'b1;
  assign CLBLM_R_X7Y100_SLICE_X8Y100_A6 = 1'b1;
  assign CLBLM_R_X7Y100_SLICE_X8Y100_B1 = 1'b1;
  assign CLBLM_R_X7Y100_SLICE_X8Y100_B2 = 1'b1;
  assign CLBLM_R_X7Y100_SLICE_X8Y100_B3 = 1'b1;
  assign CLBLM_R_X7Y100_SLICE_X8Y100_B4 = 1'b1;
  assign CLBLM_R_X7Y100_SLICE_X8Y100_B5 = 1'b1;
  assign CLBLM_R_X7Y100_SLICE_X8Y100_B6 = 1'b1;
  assign CLBLM_R_X7Y100_SLICE_X8Y100_C1 = 1'b1;
  assign CLBLM_R_X7Y100_SLICE_X8Y100_C2 = 1'b1;
  assign CLBLM_R_X7Y100_SLICE_X8Y100_C3 = 1'b1;
  assign CLBLM_R_X7Y100_SLICE_X8Y100_C4 = 1'b1;
  assign CLBLM_R_X7Y100_SLICE_X8Y100_C5 = 1'b1;
  assign CLBLM_R_X7Y100_SLICE_X8Y100_C6 = 1'b1;
  assign CLBLM_R_X7Y100_SLICE_X8Y100_D1 = 1'b1;
  assign CLBLM_R_X7Y100_SLICE_X8Y100_D2 = 1'b1;
  assign CLBLM_R_X7Y100_SLICE_X8Y100_D3 = 1'b1;
  assign CLBLM_R_X7Y100_SLICE_X8Y100_D4 = 1'b1;
  assign CLBLM_R_X7Y100_SLICE_X8Y100_D5 = 1'b1;
  assign CLBLM_R_X7Y100_SLICE_X8Y100_D6 = 1'b1;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_A1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_A2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_A3 = CLBLM_L_X10Y108_SLICE_X12Y108_DO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_A4 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_A5 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_A6 = CLBLM_R_X7Y110_SLICE_X9Y110_CO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_B1 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_B2 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_B3 = CLBLM_L_X8Y108_SLICE_X11Y108_AO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_B4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_B5 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_B6 = CLBLM_L_X8Y107_SLICE_X11Y107_CO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_C1 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_C2 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_C3 = CLBLM_L_X10Y108_SLICE_X12Y108_DO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_C4 = CLBLM_R_X7Y110_SLICE_X9Y110_CO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_C5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_C6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A1 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A2 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A3 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A4 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A5 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A6 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_D1 = CLBLM_L_X8Y108_SLICE_X11Y108_AO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_D2 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B1 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B2 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B3 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B4 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B5 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B6 = 1'b1;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_D4 = CLBLM_L_X8Y107_SLICE_X11Y107_CO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_D5 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_A1 = CLBLM_R_X7Y105_SLICE_X9Y105_AO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C2 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C3 = 1'b1;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_A2 = CLBLM_L_X10Y107_SLICE_X13Y107_CO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C5 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C6 = 1'b1;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_A3 = CLBLM_L_X10Y107_SLICE_X13Y107_AO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_A4 = CLBLM_L_X10Y108_SLICE_X12Y108_CO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_A5 = CLBLM_L_X10Y105_SLICE_X12Y105_AO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_A6 = CLBLM_L_X8Y108_SLICE_X10Y108_AO5;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_B1 = CLBLM_L_X8Y107_SLICE_X10Y107_DO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_B2 = CLBLM_L_X10Y106_SLICE_X12Y106_DO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_B3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D1 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D2 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D3 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D4 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D5 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D6 = 1'b1;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_B5 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_B6 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_C1 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_C2 = CLBLM_L_X10Y106_SLICE_X12Y106_DO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_C3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_C4 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_C5 = CLBLM_L_X8Y107_SLICE_X10Y107_DO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_C6 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_D1 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_D2 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_D3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_D4 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_D5 = CLBLM_L_X10Y107_SLICE_X13Y107_DO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_D6 = CLBLM_L_X10Y108_SLICE_X12Y108_CO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A1 = CLBLM_R_X3Y111_SLICE_X2Y111_AO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A2 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A3 = CLBLM_R_X3Y111_SLICE_X3Y111_DO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A4 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A5 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A6 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B1 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B2 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B3 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B4 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B5 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B6 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C1 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C2 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C3 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C4 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C5 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C6 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D1 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D2 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D3 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D4 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D5 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D6 = 1'b1;
  assign CLBLM_R_X7Y101_SLICE_X9Y101_A1 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X7Y101_SLICE_X9Y101_A2 = CLBLM_L_X8Y101_SLICE_X10Y101_CO6;
  assign CLBLM_R_X7Y101_SLICE_X9Y101_A3 = 1'b1;
  assign CLBLM_R_X7Y101_SLICE_X9Y101_A4 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X7Y101_SLICE_X9Y101_A5 = CLBLM_L_X8Y101_SLICE_X10Y101_BO6;
  assign CLBLM_R_X7Y101_SLICE_X9Y101_A6 = 1'b1;
  assign CLBLM_R_X7Y101_SLICE_X9Y101_B1 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X7Y101_SLICE_X9Y101_B2 = CLBLM_L_X8Y102_SLICE_X10Y102_BO6;
  assign CLBLM_R_X7Y101_SLICE_X9Y101_B3 = CLBLM_R_X7Y101_SLICE_X8Y101_CO6;
  assign CLBLM_R_X7Y101_SLICE_X9Y101_B4 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X7Y101_SLICE_X9Y101_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y101_SLICE_X9Y101_B6 = CLBLM_R_X7Y101_SLICE_X9Y101_AO5;
  assign CLBLM_R_X7Y101_SLICE_X9Y101_C1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X7Y101_SLICE_X9Y101_C2 = CLBLM_L_X8Y100_SLICE_X10Y100_AO5;
  assign CLBLM_R_X7Y101_SLICE_X9Y101_C3 = CLBLM_L_X8Y101_SLICE_X11Y101_CO6;
  assign CLBLM_R_X7Y101_SLICE_X9Y101_C4 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X7Y101_SLICE_X9Y101_C5 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X7Y101_SLICE_X9Y101_C6 = CLBLM_L_X8Y101_SLICE_X11Y101_AO6;
  assign CLBLM_R_X7Y101_SLICE_X9Y101_D1 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X7Y101_SLICE_X9Y101_D2 = 1'b1;
  assign CLBLM_R_X7Y101_SLICE_X9Y101_D3 = 1'b1;
  assign CLBLM_R_X7Y101_SLICE_X9Y101_D4 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X7Y101_SLICE_X9Y101_D5 = 1'b1;
  assign CLBLM_R_X7Y101_SLICE_X9Y101_D6 = 1'b1;
  assign CLBLM_R_X7Y101_SLICE_X8Y101_A1 = CLBLM_R_X7Y101_SLICE_X8Y101_DO6;
  assign CLBLM_R_X7Y101_SLICE_X8Y101_A2 = CLBLM_L_X8Y101_SLICE_X10Y101_BO6;
  assign CLBLM_R_X7Y101_SLICE_X8Y101_A3 = CLBLM_R_X7Y102_SLICE_X8Y102_AO6;
  assign CLBLM_R_X7Y101_SLICE_X8Y101_A4 = CLBLM_L_X8Y101_SLICE_X10Y101_CO6;
  assign CLBLM_R_X7Y101_SLICE_X8Y101_A5 = CLBLM_R_X7Y100_SLICE_X8Y100_AO6;
  assign CLBLM_R_X7Y101_SLICE_X8Y101_A6 = CLBLM_R_X7Y100_SLICE_X8Y100_AO5;
  assign CLBLM_R_X7Y101_SLICE_X8Y101_B1 = CLBLM_R_X7Y101_SLICE_X8Y101_DO6;
  assign CLBLM_R_X7Y101_SLICE_X8Y101_B2 = CLBLM_L_X8Y101_SLICE_X10Y101_BO6;
  assign CLBLM_R_X7Y101_SLICE_X8Y101_B3 = CLBLM_R_X7Y100_SLICE_X8Y100_AO6;
  assign CLBLM_R_X7Y101_SLICE_X8Y101_B4 = CLBLM_L_X8Y101_SLICE_X10Y101_CO6;
  assign CLBLM_R_X7Y101_SLICE_X8Y101_B5 = CLBLM_R_X7Y102_SLICE_X8Y102_AO6;
  assign CLBLM_R_X7Y101_SLICE_X8Y101_B6 = CLBLM_R_X7Y100_SLICE_X8Y100_AO5;
  assign CLBLM_R_X7Y101_SLICE_X8Y101_C1 = CLBLM_L_X8Y101_SLICE_X10Y101_BO6;
  assign CLBLM_R_X7Y101_SLICE_X8Y101_C2 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X7Y101_SLICE_X8Y101_C3 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X7Y101_SLICE_X8Y101_C4 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X7Y101_SLICE_X8Y101_C5 = CLBLM_R_X7Y101_SLICE_X8Y101_DO6;
  assign CLBLM_R_X7Y101_SLICE_X8Y101_C6 = CLBLM_L_X8Y101_SLICE_X10Y101_CO6;
  assign CLBLM_R_X7Y101_SLICE_X8Y101_D1 = CLBLM_L_X8Y101_SLICE_X11Y101_BO6;
  assign CLBLM_R_X7Y101_SLICE_X8Y101_D2 = CLBLL_L_X4Y100_SLICE_X4Y100_AO5;
  assign CLBLM_R_X7Y101_SLICE_X8Y101_D3 = CLBLM_R_X5Y100_SLICE_X6Y100_AO5;
  assign CLBLM_R_X7Y101_SLICE_X8Y101_D4 = CLBLM_L_X8Y103_SLICE_X11Y103_AO5;
  assign CLBLM_R_X7Y101_SLICE_X8Y101_D5 = CLBLM_L_X8Y101_SLICE_X11Y101_CO6;
  assign CLBLM_R_X7Y101_SLICE_X8Y101_D6 = CLBLM_L_X8Y100_SLICE_X10Y100_CO6;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_A1 = CLBLM_L_X10Y106_SLICE_X12Y106_CO6;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_A2 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_A3 = CLBLM_L_X10Y107_SLICE_X13Y107_DO6;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_A4 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_A5 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_A6 = CLBLM_L_X8Y108_SLICE_X11Y108_CO6;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_B1 = CLBLM_L_X8Y108_SLICE_X11Y108_DO6;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_B2 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_B3 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_B4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_B5 = CLBLM_L_X10Y108_SLICE_X12Y108_DO6;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_B6 = CLBLM_L_X8Y111_SLICE_X10Y111_BO6;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_C1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_C2 = CLBLM_L_X8Y109_SLICE_X11Y109_AO6;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_C3 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_C4 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_C5 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_C6 = CLBLM_L_X8Y110_SLICE_X10Y110_BO6;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_D1 = CLBLM_L_X8Y109_SLICE_X11Y109_AO6;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_D2 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_D3 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_D4 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_D5 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_D6 = CLBLM_L_X8Y110_SLICE_X10Y110_BO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_A1 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_A2 = 1'b1;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_A3 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_A4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_A5 = 1'b1;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_A6 = 1'b1;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_B1 = CLBLM_R_X7Y110_SLICE_X9Y110_CO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_B2 = CLBLM_L_X10Y107_SLICE_X13Y107_AO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_B3 = CLBLM_L_X10Y108_SLICE_X12Y108_CO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_B4 = CLBLM_L_X10Y108_SLICE_X12Y108_BO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_B5 = CLBLM_L_X8Y108_SLICE_X10Y108_AO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_B6 = CLBLM_L_X8Y108_SLICE_X10Y108_AO5;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_C1 = CLBLM_L_X10Y107_SLICE_X13Y107_DO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_C2 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_C3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_C4 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_C5 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_C6 = CLBLM_L_X10Y108_SLICE_X12Y108_CO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_D1 = 1'b1;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_D2 = 1'b1;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_D3 = 1'b1;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_D4 = 1'b1;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_D5 = 1'b1;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_D6 = 1'b1;
  assign LIOI3_X0Y111_ILOGIC_X0Y112_D = LIOB33_X0Y111_IOB_X0Y112_I;
  assign LIOI3_X0Y111_ILOGIC_X0Y111_D = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_A1 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_A2 = CLBLM_R_X7Y103_SLICE_X8Y103_AO5;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_A3 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_A4 = 1'b1;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_A5 = CLBLM_R_X7Y102_SLICE_X9Y102_CO6;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_A6 = 1'b1;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_B1 = CLBLM_R_X7Y101_SLICE_X9Y101_DO6;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_B2 = CLBLM_R_X7Y103_SLICE_X9Y103_AO6;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_B3 = CLBLM_R_X7Y101_SLICE_X8Y101_BO6;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_B4 = CLBLM_L_X8Y103_SLICE_X10Y103_DO6;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_B5 = CLBLM_R_X7Y101_SLICE_X8Y101_AO6;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_B6 = CLBLM_R_X7Y102_SLICE_X8Y102_DO6;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_C1 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_C2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_C3 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_C4 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_C5 = CLBLM_R_X7Y103_SLICE_X9Y103_DO6;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_C6 = CLBLM_R_X7Y101_SLICE_X9Y101_BO6;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_D1 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_D2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_D3 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_D4 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_D5 = CLBLM_R_X7Y103_SLICE_X9Y103_DO6;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_D6 = CLBLM_R_X7Y101_SLICE_X9Y101_BO6;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_A1 = CLBLM_R_X7Y101_SLICE_X9Y101_CO6;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_A2 = CLBLM_R_X5Y102_SLICE_X7Y102_BO6;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_A3 = 1'b1;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_A4 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_A5 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_A6 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_C4 = CLBLM_L_X8Y112_SLICE_X10Y112_BO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_C5 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_B1 = CLBLM_R_X7Y102_SLICE_X8Y102_DO6;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_B2 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_B3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_B4 = CLBLM_R_X7Y101_SLICE_X9Y101_AO6;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_B5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_B6 = CLBLM_R_X7Y102_SLICE_X8Y102_AO5;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_C6 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_C1 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_C2 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_C3 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_C4 = CLBLM_R_X7Y102_SLICE_X8Y102_AO5;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_C5 = CLBLM_R_X7Y102_SLICE_X8Y102_DO6;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_C6 = CLBLM_R_X7Y101_SLICE_X9Y101_AO6;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_D1 = CLBLM_R_X5Y101_SLICE_X7Y101_BO6;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_D2 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_D3 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_D4 = CLBLM_R_X7Y101_SLICE_X9Y101_CO6;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_D5 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_D6 = CLBLM_R_X5Y102_SLICE_X7Y102_BO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_D5 = CLBLM_R_X7Y113_SLICE_X9Y113_BO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_D6 = CLBLM_R_X7Y113_SLICE_X9Y113_AO5;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_A1 = CLBLM_L_X10Y109_SLICE_X12Y109_CO6;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_A2 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_A3 = CLBLM_L_X8Y109_SLICE_X10Y109_AO6;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_A4 = CLBLM_L_X10Y109_SLICE_X12Y109_AO6;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_A5 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_A6 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_B1 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_B2 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_B3 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_B4 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_B5 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_B6 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_C1 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_C2 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_C3 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_C4 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_C5 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_C6 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_D1 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_D2 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_D3 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_D4 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_D5 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_D6 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_A1 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_A2 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_A3 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_A4 = CLBLM_L_X8Y109_SLICE_X10Y109_BO6;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_A5 = CLBLM_L_X8Y109_SLICE_X10Y109_CO6;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_A6 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_B1 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_B2 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_B3 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_B4 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_B5 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_B6 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_C1 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_C2 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_C3 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_C4 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_C5 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_C6 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_D1 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_D2 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_D3 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_D4 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_D5 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_D6 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_B6 = CLBLM_R_X5Y113_SLICE_X6Y113_CO6;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_C4 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_C5 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_C6 = CLBLM_R_X7Y112_SLICE_X8Y112_BO6;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_A1 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_A3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_A4 = 1'b1;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_A5 = 1'b1;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_A6 = 1'b1;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_B1 = CLBLM_L_X8Y103_SLICE_X10Y103_DO6;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_B2 = CLBLM_R_X7Y101_SLICE_X8Y101_AO6;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_B3 = CLBLM_L_X8Y103_SLICE_X10Y103_BO6;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_B4 = CLBLM_L_X10Y103_SLICE_X12Y103_BO6;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_B5 = CLBLM_R_X7Y103_SLICE_X9Y103_AO6;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_B6 = CLBLM_R_X7Y105_SLICE_X9Y105_AO5;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_D2 = CLBLM_L_X8Y105_SLICE_X10Y105_BO6;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_C1 = CLBLM_R_X7Y102_SLICE_X9Y102_AO6;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_C2 = CLBLM_L_X8Y104_SLICE_X10Y104_AO5;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_D3 = CLBLM_L_X8Y105_SLICE_X11Y105_BO6;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_C3 = CLBLM_R_X7Y103_SLICE_X8Y103_BO6;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_C4 = CLBLM_R_X7Y103_SLICE_X9Y103_AO5;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_C5 = CLBLM_R_X7Y103_SLICE_X9Y103_DO6;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_C6 = CLBLM_R_X7Y102_SLICE_X9Y102_BO6;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_D1 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_D2 = CLBLM_L_X8Y103_SLICE_X10Y103_BO6;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_D3 = CLBLM_L_X10Y104_SLICE_X12Y104_DO6;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_D4 = CLBLM_L_X8Y103_SLICE_X11Y103_CO6;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_D5 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_D6 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_A1 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_A2 = 1'b1;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_A3 = CLBLM_R_X7Y102_SLICE_X8Y102_CO6;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_A5 = CLBLM_R_X7Y103_SLICE_X8Y103_CO6;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_A6 = 1'b1;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_B1 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_B2 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_B3 = CLBLM_R_X7Y101_SLICE_X8Y101_CO6;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_B4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_B5 = CLBLM_L_X8Y103_SLICE_X10Y103_DO6;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_B6 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_C1 = CLBLM_R_X7Y101_SLICE_X8Y101_CO6;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_C2 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_C3 = CLBLM_L_X8Y103_SLICE_X10Y103_DO6;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_C5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_C6 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_D1 = CLBLM_R_X7Y102_SLICE_X9Y102_BO6;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_D2 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_D3 = CLBLM_R_X7Y103_SLICE_X9Y103_DO6;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_D4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_D5 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_D6 = CLBLM_R_X7Y103_SLICE_X8Y103_BO6;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_B6 = CLBLM_L_X8Y106_SLICE_X10Y106_AO5;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_A1 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_A2 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_A3 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_A4 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_A5 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_A6 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_B1 = CLBLM_L_X10Y109_SLICE_X12Y109_DO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_B2 = CLBLM_L_X8Y109_SLICE_X10Y109_BO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_B3 = CLBLM_L_X10Y108_SLICE_X13Y108_AO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_B4 = CLBLM_L_X8Y109_SLICE_X10Y109_CO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_B5 = CLBLM_L_X8Y110_SLICE_X11Y110_AO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_B6 = CLBLM_L_X8Y110_SLICE_X11Y110_AO5;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_C1 = CLBLM_L_X10Y108_SLICE_X13Y108_BO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_C2 = CLBLM_L_X10Y107_SLICE_X12Y107_AO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_C3 = CLBLM_R_X7Y112_SLICE_X9Y112_AO5;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_C4 = CLBLM_L_X8Y112_SLICE_X11Y112_CO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_C5 = CLBLM_L_X8Y110_SLICE_X11Y110_DO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_C6 = CLBLM_L_X8Y110_SLICE_X11Y110_BO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_D1 = CLBLM_L_X8Y110_SLICE_X11Y110_AO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_D2 = CLBLM_L_X8Y109_SLICE_X10Y109_CO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_D3 = CLBLM_L_X10Y109_SLICE_X12Y109_DO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_D4 = CLBLM_L_X8Y110_SLICE_X11Y110_AO5;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_D5 = CLBLM_L_X10Y108_SLICE_X13Y108_AO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_D6 = CLBLM_L_X8Y109_SLICE_X10Y109_BO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_A1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_A2 = CLBLM_L_X8Y112_SLICE_X11Y112_CO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_A3 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_A4 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_A5 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_A6 = CLBLM_L_X8Y110_SLICE_X10Y110_CO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_B1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_B2 = CLBLM_L_X8Y112_SLICE_X11Y112_CO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_B3 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_B4 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_B5 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_B6 = CLBLM_L_X8Y110_SLICE_X10Y110_CO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_C1 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_C2 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_C3 = CLBLM_L_X10Y109_SLICE_X12Y109_DO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_C4 = CLBLM_L_X8Y109_SLICE_X10Y109_CO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_C5 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_C6 = CLBLM_L_X8Y109_SLICE_X10Y109_BO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_D1 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_D2 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_D3 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_D4 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_D5 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_D6 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_A1 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_A2 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_A3 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_A4 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_A5 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_A6 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_B1 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_B2 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_B3 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_B4 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_B5 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_B6 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_C1 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_C2 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_C3 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_C4 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_C5 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_C6 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_D1 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_D2 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_D3 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_D4 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_D5 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X0Y102_D6 = 1'b1;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_A1 = CLBLM_L_X10Y104_SLICE_X12Y104_DO6;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_A2 = CLBLM_L_X8Y103_SLICE_X11Y103_CO6;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_A3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_A4 = CLBLM_L_X8Y103_SLICE_X10Y103_BO6;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_A5 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_A6 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_B1 = 1'b1;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_B2 = 1'b1;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_B3 = 1'b1;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_B4 = 1'b1;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_B5 = 1'b1;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_B6 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_A1 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_A2 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_A3 = CLBLL_L_X4Y101_SLICE_X4Y101_DO6;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_A4 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_A5 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_A6 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_C1 = 1'b1;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_C2 = 1'b1;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_C3 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_B1 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_B2 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_B3 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_B4 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_B5 = CLBLL_L_X2Y102_SLICE_X1Y102_AO6;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_B6 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_D1 = 1'b1;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_D2 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_C1 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_C2 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_C3 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_C4 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_C5 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_C6 = 1'b1;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_D4 = 1'b1;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_A1 = CLBLM_L_X8Y105_SLICE_X11Y105_DO6;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_A2 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_A3 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_A4 = CLBLM_R_X7Y104_SLICE_X8Y104_BO6;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_A5 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_A6 = CLBLM_R_X7Y105_SLICE_X8Y105_AO6;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_D1 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_D2 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_D3 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_D4 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_D5 = 1'b1;
  assign CLBLL_L_X2Y102_SLICE_X1Y102_D6 = 1'b1;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_B4 = CLBLM_L_X8Y104_SLICE_X10Y104_BO6;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_B6 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_B1 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_B2 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_B3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_B5 = CLBLM_L_X8Y104_SLICE_X11Y104_BO6;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_C1 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_C2 = CLBLM_L_X8Y105_SLICE_X11Y105_DO6;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_C3 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_C4 = CLBLM_R_X7Y105_SLICE_X8Y105_AO6;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_C5 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_C6 = CLBLM_R_X7Y104_SLICE_X8Y104_BO6;
  assign LIOI3_X0Y115_ILOGIC_X0Y115_D = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_D1 = CLBLM_L_X8Y104_SLICE_X11Y104_BO6;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_D2 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_D3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_D4 = CLBLM_L_X8Y104_SLICE_X10Y104_BO6;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_D5 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_D6 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_A1 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_A2 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_A3 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_A4 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_A5 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_A6 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_B1 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_B2 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_B3 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_B4 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_B5 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_B6 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_C1 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_C2 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_C3 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_C4 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_C5 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_C6 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_D1 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_D2 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_D3 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_D4 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_D5 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_D6 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_A1 = CLBLM_L_X8Y112_SLICE_X10Y112_AO5;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_A2 = CLBLM_L_X8Y110_SLICE_X10Y110_CO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_A3 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_A4 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_A5 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_A6 = CLBLM_L_X8Y109_SLICE_X10Y109_AO5;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_B1 = CLBLM_L_X8Y112_SLICE_X10Y112_DO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_B2 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_B3 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_B4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_B5 = CLBLM_L_X8Y111_SLICE_X10Y111_AO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_B6 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_C1 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_C2 = CLBLM_L_X8Y110_SLICE_X10Y110_CO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_C3 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_C4 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_C5 = CLBLM_L_X8Y112_SLICE_X10Y112_AO5;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_C6 = CLBLM_L_X8Y109_SLICE_X10Y109_AO5;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_D1 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_D2 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_D3 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_D4 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_D5 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_D6 = 1'b1;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_A1 = 1'b1;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_A2 = CLBLM_R_X5Y102_SLICE_X6Y102_CO6;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_A3 = CLBLL_L_X2Y103_SLICE_X1Y103_AO6;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_A4 = CLBLL_L_X4Y106_SLICE_X4Y106_AO5;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_A5 = 1'b1;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_A6 = 1'b1;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_B1 = 1'b1;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_B2 = 1'b1;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_B3 = 1'b1;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_B4 = 1'b1;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_B5 = 1'b1;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_B6 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_B4 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_C1 = 1'b1;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_C2 = 1'b1;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_C3 = 1'b1;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_C4 = 1'b1;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_C5 = 1'b1;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_C6 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_B5 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_B6 = CLBLM_R_X3Y112_SLICE_X3Y112_DO6;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_D1 = 1'b1;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_D2 = 1'b1;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_D3 = 1'b1;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_D4 = 1'b1;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_D5 = 1'b1;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_D6 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_A1 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_A2 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_A3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_A4 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_A5 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_A6 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_B1 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_B2 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_B3 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_B4 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_B5 = 1'b1;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_A1 = 1'b1;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_A2 = CLBLL_L_X4Y106_SLICE_X4Y106_AO5;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_A3 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_A4 = CLBLM_R_X5Y102_SLICE_X6Y102_CO6;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_A5 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_A6 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_C2 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_B6 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_C5 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_C1 = 1'b1;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_B1 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_B2 = CLBLL_L_X4Y106_SLICE_X4Y106_AO5;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_B3 = CLBLL_L_X4Y101_SLICE_X5Y101_DO6;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_B4 = CLBLM_R_X5Y102_SLICE_X6Y102_CO6;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_B5 = CLBLL_L_X2Y103_SLICE_X1Y103_AO6;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_C6 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_D1 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_D2 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_D3 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_D4 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_D5 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_D6 = 1'b1;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_C1 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_C2 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_C3 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_C4 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_C5 = CLBLL_L_X2Y103_SLICE_X1Y103_DO6;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_C6 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_A1 = CLBLM_L_X8Y104_SLICE_X11Y104_BO6;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_A2 = CLBLM_R_X7Y103_SLICE_X9Y103_BO6;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_A3 = CLBLM_L_X8Y106_SLICE_X11Y106_AO6;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_A4 = CLBLM_R_X5Y105_SLICE_X7Y105_BO6;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_A5 = CLBLM_R_X7Y104_SLICE_X9Y104_AO6;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_A6 = CLBLM_L_X8Y104_SLICE_X10Y104_AO5;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_D1 = CLBLL_L_X2Y102_SLICE_X1Y102_AO6;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_D2 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_D3 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_B1 = CLBLM_R_X7Y105_SLICE_X8Y105_DO6;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_D4 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_D5 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_B4 = CLBLM_L_X8Y105_SLICE_X11Y105_DO6;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_D6 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_B6 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_B2 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_B3 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_B5 = CLBLM_R_X7Y104_SLICE_X8Y104_BO6;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_C1 = CLBLM_R_X7Y104_SLICE_X9Y104_AO6;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_C2 = CLBLM_L_X8Y106_SLICE_X11Y106_AO6;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_C3 = CLBLM_R_X7Y103_SLICE_X9Y103_BO6;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_C4 = CLBLM_L_X8Y104_SLICE_X10Y104_AO5;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_C5 = CLBLM_L_X8Y104_SLICE_X11Y104_BO6;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_C6 = CLBLM_R_X5Y105_SLICE_X7Y105_BO6;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_D1 = CLBLM_R_X7Y104_SLICE_X9Y104_AO6;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_D2 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_D3 = CLBLM_R_X7Y103_SLICE_X9Y103_BO6;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_D4 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_D5 = CLBLM_L_X8Y104_SLICE_X11Y104_BO6;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_D6 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_C6 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_C4 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_C5 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_C6 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_A1 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_A2 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_A3 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_A4 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_A5 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_A6 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_B1 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_B2 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_B3 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_B4 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_B5 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_B6 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_C1 = CLBLM_L_X8Y113_SLICE_X11Y113_AO6;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_C2 = CLBLM_L_X8Y109_SLICE_X10Y109_BO6;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_C3 = CLBLM_L_X8Y113_SLICE_X11Y113_AO5;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_C4 = CLBLM_L_X8Y110_SLICE_X11Y110_AO5;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_C5 = CLBLM_L_X8Y112_SLICE_X11Y112_AO6;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_C6 = CLBLM_L_X8Y112_SLICE_X11Y112_BO6;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_D1 = CLBLM_L_X8Y113_SLICE_X11Y113_AO6;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_D2 = CLBLM_L_X8Y110_SLICE_X11Y110_AO5;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_D3 = CLBLM_L_X8Y113_SLICE_X11Y113_AO5;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_D4 = CLBLM_L_X8Y112_SLICE_X11Y112_AO6;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_D5 = CLBLM_L_X8Y109_SLICE_X10Y109_BO6;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_D6 = CLBLM_L_X8Y112_SLICE_X11Y112_BO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_A1 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_A2 = CLBLM_L_X8Y112_SLICE_X11Y112_BO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_A3 = CLBLM_L_X8Y112_SLICE_X11Y112_AO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_A4 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_A5 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_A6 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_B1 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_B2 = CLBLM_L_X8Y112_SLICE_X11Y112_BO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_B3 = CLBLM_L_X8Y112_SLICE_X11Y112_AO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_B4 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_B5 = CLBLM_L_X8Y109_SLICE_X10Y109_BO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_B6 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_C1 = CLBLM_R_X7Y113_SLICE_X9Y113_DO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_C2 = CLBLM_L_X8Y112_SLICE_X11Y112_CO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_C3 = CLBLM_L_X8Y112_SLICE_X11Y112_DO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_C4 = CLBLM_R_X7Y113_SLICE_X9Y113_AO5;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_C5 = CLBLM_R_X7Y112_SLICE_X9Y112_AO5;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_C6 = CLBLM_L_X8Y110_SLICE_X11Y110_BO6;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_A1 = CLBLL_L_X4Y104_SLICE_X4Y104_BO5;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_A2 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_A3 = CLBLL_L_X2Y105_SLICE_X0Y105_DO6;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_A4 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_A5 = 1'b1;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_A6 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_D6 = CLBLM_L_X8Y112_SLICE_X10Y112_BO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_D1 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_B1 = CLBLL_L_X2Y105_SLICE_X0Y105_BO5;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_B2 = CLBLL_L_X4Y103_SLICE_X4Y103_AO6;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_B3 = CLBLL_L_X4Y104_SLICE_X4Y104_BO5;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_B4 = CLBLL_L_X2Y104_SLICE_X0Y104_DO6;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_B5 = CLBLL_L_X2Y105_SLICE_X0Y105_DO6;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_B6 = CLBLL_L_X2Y105_SLICE_X1Y105_CO6;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_C1 = CLBLL_L_X2Y104_SLICE_X0Y104_AO6;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_C2 = CLBLL_L_X2Y105_SLICE_X1Y105_CO6;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_C3 = CLBLL_L_X2Y105_SLICE_X0Y105_BO5;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_C4 = CLBLL_L_X2Y104_SLICE_X0Y104_AO5;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_C5 = CLBLL_L_X4Y103_SLICE_X4Y103_AO6;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_C6 = CLBLL_L_X4Y104_SLICE_X4Y104_CO5;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_D1 = CLBLL_L_X2Y114_SLICE_X0Y114_AO5;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_D1 = 1'b1;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_D2 = 1'b1;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_D3 = 1'b1;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_D4 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_D5 = 1'b1;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_D6 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_T1 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_A1 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_A2 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_A3 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_A4 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_A5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_A6 = 1'b1;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_A1 = CLBLM_R_X3Y103_SLICE_X2Y103_BO6;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_A2 = CLBLL_L_X4Y104_SLICE_X4Y104_AO5;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_A3 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_B4 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_B5 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_B6 = 1'b1;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_A4 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_A5 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_A6 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_B1 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_B2 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_C3 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_C4 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_C5 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_C6 = 1'b1;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_B1 = CLBLL_L_X2Y103_SLICE_X1Y103_DO6;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_B2 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_B3 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_B4 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_B5 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_B6 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_C1 = CLBLL_L_X4Y104_SLICE_X4Y104_CO5;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_C2 = 1'b1;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_C3 = CLBLL_L_X2Y104_SLICE_X0Y104_BO6;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_D2 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_D3 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_D4 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_D5 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_D6 = 1'b1;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_C4 = 1'b1;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_C5 = 1'b1;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_C6 = 1'b1;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_D1 = 1'b1;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_D2 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_A1 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_A2 = CLBLM_L_X8Y108_SLICE_X11Y108_BO6;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_A3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_A4 = CLBLM_R_X7Y109_SLICE_X8Y109_BO6;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_A5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_A6 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_D3 = 1'b1;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_D4 = 1'b1;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_D5 = 1'b1;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_D6 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_B2 = CLBLM_R_X7Y107_SLICE_X9Y107_BO6;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_B3 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_B4 = CLBLM_L_X8Y107_SLICE_X11Y107_BO6;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_B5 = CLBLM_R_X7Y106_SLICE_X8Y106_AO6;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_B6 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_B1 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_C1 = CLBLM_R_X7Y106_SLICE_X8Y106_AO6;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_C2 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_C3 = CLBLM_R_X7Y107_SLICE_X9Y107_BO6;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_C4 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_C5 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_C6 = CLBLM_L_X8Y107_SLICE_X11Y107_BO6;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_D1 = CLBLM_R_X7Y106_SLICE_X8Y106_AO6;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_D2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_D3 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_D4 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_D5 = CLBLM_R_X7Y107_SLICE_X9Y107_CO6;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_D6 = CLBLM_L_X8Y107_SLICE_X11Y107_BO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_A1 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_A2 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_A3 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_A4 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_A5 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_A6 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_B1 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_B2 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_B3 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_B4 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_B5 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_B6 = 1'b1;
  assign LIOI3_X0Y117_ILOGIC_X0Y117_D = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_C1 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_C2 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_C3 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_C4 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_C5 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_C6 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_D1 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_D2 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_D3 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_D4 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_D5 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_D6 = 1'b1;
  assign RIOI3_X105Y101_ILOGIC_X1Y102_D = RIOB33_X105Y101_IOB_X1Y102_I;
  assign RIOI3_X105Y101_ILOGIC_X1Y101_D = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_A1 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_A2 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_A3 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_A4 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_A5 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_A6 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_B1 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_B2 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_B3 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_B4 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_B5 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_B6 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_C1 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_C2 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_C3 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_C4 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_C5 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_C6 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_A1 = CLBLL_L_X2Y105_SLICE_X0Y105_BO5;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_A2 = CLBLL_L_X2Y105_SLICE_X1Y105_BO6;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_A3 = CLBLM_R_X3Y106_SLICE_X3Y106_CO6;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_A4 = CLBLL_L_X2Y105_SLICE_X0Y105_BO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_D1 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_D2 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_D3 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_D4 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_D5 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_D6 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_A5 = CLBLL_L_X2Y104_SLICE_X0Y104_AO6;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_A6 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_B1 = CLBLL_L_X2Y106_SLICE_X1Y106_BO6;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_B2 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_B3 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_B4 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_B5 = CLBLL_L_X2Y105_SLICE_X0Y105_CO6;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_B6 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_C1 = CLBLL_L_X2Y103_SLICE_X0Y103_AO6;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_C2 = CLBLL_L_X2Y105_SLICE_X1Y105_AO5;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_C3 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_C4 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_C5 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_C6 = CLBLL_L_X4Y101_SLICE_X4Y101_BO6;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_D1 = CLBLL_L_X2Y103_SLICE_X0Y103_AO6;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_D2 = CLBLL_L_X2Y105_SLICE_X1Y105_AO5;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_D3 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_D4 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_D5 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_D6 = CLBLL_L_X4Y101_SLICE_X4Y101_BO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_A1 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_A2 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_A3 = 1'b1;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_A4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_A5 = 1'b1;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_A6 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_A1 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_A3 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_A4 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_A5 = CLBLL_L_X4Y101_SLICE_X5Y101_DO6;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_A6 = 1'b1;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_B1 = CLBLM_L_X8Y108_SLICE_X10Y108_CO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_B2 = CLBLM_L_X8Y107_SLICE_X10Y107_AO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_B3 = CLBLM_R_X7Y106_SLICE_X9Y106_AO6;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_B1 = CLBLL_L_X4Y104_SLICE_X4Y104_AO5;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_B2 = CLBLM_R_X3Y106_SLICE_X3Y106_BO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_C1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_C2 = CLBLM_L_X8Y107_SLICE_X10Y107_AO6;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_B3 = CLBLL_L_X2Y106_SLICE_X1Y106_AO6;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_B4 = CLBLM_R_X3Y105_SLICE_X2Y105_AO5;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_B5 = CLBLL_L_X2Y107_SLICE_X1Y107_AO6;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_B6 = CLBLM_R_X3Y103_SLICE_X2Y103_BO6;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_C1 = CLBLL_L_X2Y105_SLICE_X0Y105_BO6;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_C2 = CLBLM_R_X3Y105_SLICE_X2Y105_CO6;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_C3 = CLBLM_R_X3Y106_SLICE_X2Y106_DO6;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_C4 = CLBLM_R_X3Y106_SLICE_X3Y106_CO6;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_C5 = CLBLL_L_X2Y104_SLICE_X1Y104_AO6;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_C6 = CLBLM_R_X3Y106_SLICE_X3Y106_BO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_C5 = CLBLM_L_X8Y107_SLICE_X11Y107_CO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_C6 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_D1 = CLBLM_R_X7Y106_SLICE_X9Y106_AO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_D2 = CLBLM_L_X8Y108_SLICE_X10Y108_CO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_D3 = CLBLM_L_X8Y107_SLICE_X10Y107_AO6;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_D1 = CLBLL_L_X2Y107_SLICE_X1Y107_AO6;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_D2 = CLBLL_L_X2Y104_SLICE_X1Y104_AO5;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_D3 = CLBLL_L_X2Y104_SLICE_X1Y104_AO6;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_D4 = CLBLM_R_X3Y105_SLICE_X2Y105_AO5;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_D5 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_D6 = CLBLM_R_X3Y106_SLICE_X3Y106_BO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_D4 = CLBLM_R_X7Y107_SLICE_X9Y107_AO5;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_A1 = CLBLM_R_X7Y108_SLICE_X8Y108_AO5;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_A2 = CLBLM_L_X8Y107_SLICE_X11Y107_AO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_A3 = CLBLM_R_X7Y107_SLICE_X9Y107_AO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_A4 = CLBLM_L_X8Y108_SLICE_X10Y108_BO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_A5 = CLBLM_R_X7Y106_SLICE_X9Y106_AO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_A6 = CLBLM_R_X7Y109_SLICE_X8Y109_BO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_B1 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_B2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_B3 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_B4 = CLBLM_R_X7Y109_SLICE_X8Y109_BO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_B5 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_B6 = CLBLM_L_X8Y108_SLICE_X11Y108_BO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_C4 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_C5 = CLBLM_L_X8Y112_SLICE_X11Y112_AO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_C1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_C2 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_C3 = CLBLM_L_X8Y107_SLICE_X11Y107_AO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_C4 = CLBLM_L_X8Y108_SLICE_X10Y108_BO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_C5 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_C6 = CLBLM_R_X7Y109_SLICE_X8Y109_BO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_C6 = CLBLM_R_X5Y111_SLICE_X7Y111_BO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_D1 = CLBLM_R_X7Y106_SLICE_X9Y106_AO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_D2 = CLBLM_R_X7Y107_SLICE_X9Y107_AO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_D3 = CLBLM_L_X8Y107_SLICE_X11Y107_AO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_D4 = CLBLM_L_X8Y108_SLICE_X10Y108_BO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_D5 = CLBLM_R_X7Y108_SLICE_X8Y108_AO5;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_D6 = CLBLM_R_X7Y109_SLICE_X8Y109_BO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_D2 = CLBLM_R_X7Y112_SLICE_X8Y112_AO5;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_D3 = CLBLM_R_X7Y113_SLICE_X8Y113_BO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_D4 = CLBLM_R_X5Y111_SLICE_X7Y111_BO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_A1 = CLBLM_R_X3Y106_SLICE_X3Y106_CO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_A2 = CLBLL_L_X2Y106_SLICE_X1Y106_BO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_A3 = CLBLL_L_X2Y106_SLICE_X1Y106_AO5;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_A4 = CLBLL_L_X2Y105_SLICE_X1Y105_BO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_A5 = CLBLL_L_X2Y104_SLICE_X0Y104_AO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_A6 = CLBLL_L_X2Y105_SLICE_X0Y105_CO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_B1 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_B2 = CLBLL_L_X4Y103_SLICE_X4Y103_AO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_B3 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_B4 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_B5 = CLBLL_L_X2Y106_SLICE_X0Y106_AO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_B6 = CLBLL_L_X2Y104_SLICE_X0Y104_AO5;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_C1 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_C2 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_C3 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_C4 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_C5 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_C6 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_B6 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_D1 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_D2 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_D3 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_D4 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_D5 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_D6 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_C4 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_A1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_A2 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_A3 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_A4 = CLBLM_L_X8Y108_SLICE_X10Y108_AO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_A5 = CLBLM_R_X7Y110_SLICE_X9Y110_DO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_A6 = CLBLM_R_X7Y110_SLICE_X9Y110_CO6;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_A4 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_A5 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_A6 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_A2 = CLBLM_L_X10Y108_SLICE_X12Y108_BO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_B2 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_B3 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_B4 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_B5 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_B6 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_B1 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_B2 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_B3 = CLBLL_L_X2Y103_SLICE_X1Y103_BO6;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_B4 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_B5 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_C4 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_C5 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_C1 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_C2 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_C3 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_C4 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_C5 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_C6 = 1'b1;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_D3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_D1 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_D1 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_D3 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_D4 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_D5 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_D2 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_D3 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_D4 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_D5 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_D6 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_D6 = 1'b1;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_D6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_A1 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_A2 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_A3 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_A4 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_A5 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_A6 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_B1 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_B2 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_B3 = CLBLM_R_X7Y108_SLICE_X9Y108_AO6;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_B4 = CLBLM_R_X5Y110_SLICE_X7Y110_CO6;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_B5 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_B6 = CLBLM_R_X7Y109_SLICE_X8Y109_AO6;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_C1 = CLBLM_R_X7Y108_SLICE_X8Y108_AO6;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_C2 = CLBLM_R_X5Y108_SLICE_X6Y108_AO5;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_C3 = CLBLM_R_X7Y108_SLICE_X9Y108_AO6;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_C4 = CLBLM_R_X7Y108_SLICE_X8Y108_AO5;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_C5 = CLBLM_R_X5Y110_SLICE_X7Y110_CO6;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_C6 = CLBLM_R_X7Y109_SLICE_X8Y109_AO6;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_D1 = CLBLM_R_X7Y108_SLICE_X8Y108_AO6;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_D2 = CLBLM_R_X5Y108_SLICE_X6Y108_AO5;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_D3 = CLBLM_R_X7Y108_SLICE_X9Y108_AO6;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_D4 = CLBLM_R_X7Y108_SLICE_X8Y108_AO5;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_D5 = CLBLM_R_X5Y110_SLICE_X7Y110_CO6;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_D6 = CLBLM_R_X7Y109_SLICE_X8Y109_AO6;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_D1 = CLBLL_L_X2Y113_SLICE_X1Y113_AO6;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_T1 = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_D1 = CLBLL_L_X2Y113_SLICE_X0Y113_BO5;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_T1 = 1'b1;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_B4 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_A1 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_A2 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_A3 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_A4 = CLBLL_L_X2Y104_SLICE_X1Y104_BO6;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_A5 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_A6 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_B1 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_B2 = CLBLL_L_X2Y104_SLICE_X1Y104_BO6;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_B3 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_B4 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_B5 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_B6 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_C1 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_C2 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_C3 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_C4 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_C5 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_C6 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_D1 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_D2 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_D3 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_D4 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_D5 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_D6 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_A1 = CLBLM_R_X3Y109_SLICE_X2Y109_AO6;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_A2 = CLBLM_R_X3Y106_SLICE_X2Y106_BO6;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_A3 = CLBLM_R_X3Y105_SLICE_X2Y105_AO6;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_A4 = CLBLL_L_X2Y107_SLICE_X1Y107_BO6;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_A5 = CLBLM_R_X3Y108_SLICE_X2Y108_DO6;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_A6 = CLBLM_R_X3Y106_SLICE_X2Y106_CO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_A1 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_A2 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_A3 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_B1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_B2 = CLBLL_L_X2Y107_SLICE_X0Y107_BO6;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_B3 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_B4 = CLBLL_L_X4Y104_SLICE_X4Y104_DO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_B1 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_B2 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_B3 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_B4 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_B5 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_B6 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_B5 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_B6 = CLBLL_L_X2Y108_SLICE_X1Y108_CO6;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_C1 = CLBLL_L_X2Y107_SLICE_X1Y107_AO6;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_C2 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_C3 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_C4 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_C5 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_C6 = CLBLM_R_X3Y105_SLICE_X2Y105_BO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_C1 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_C2 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_C3 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_C4 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_C5 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_C6 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_D1 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_D2 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_D3 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_D4 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_D5 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_D6 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_D1 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_D2 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_D3 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_D4 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_D5 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_D6 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_A1 = CLBLM_R_X7Y111_SLICE_X8Y111_DO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_A2 = CLBLM_R_X7Y110_SLICE_X9Y110_BO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_A3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_A4 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_A5 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_A6 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_B1 = CLBLM_R_X7Y111_SLICE_X8Y111_DO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_B2 = CLBLM_R_X7Y110_SLICE_X9Y110_BO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_B3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_B4 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_B5 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_B6 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_C1 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_C2 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_C3 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_C4 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_C5 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_C6 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_D1 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_D2 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_D3 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_D4 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_D5 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_D6 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_A1 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_A2 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_A3 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_A4 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_A5 = CLBLL_L_X2Y107_SLICE_X0Y107_BO6;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_A6 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_B1 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_B2 = CLBLM_R_X3Y104_SLICE_X2Y104_CO6;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_B3 = CLBLL_L_X2Y107_SLICE_X0Y107_AO6;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_B4 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_B5 = CLBLL_L_X2Y107_SLICE_X0Y107_BO6;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_B6 = CLBLM_R_X3Y104_SLICE_X3Y104_CO6;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_C1 = CLBLM_R_X3Y104_SLICE_X2Y104_CO6;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_C2 = CLBLL_L_X2Y107_SLICE_X0Y107_AO6;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_C3 = CLBLM_R_X3Y104_SLICE_X3Y104_CO6;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_C4 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_C5 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_C6 = CLBLL_L_X2Y107_SLICE_X0Y107_BO6;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_D1 = CLBLM_R_X3Y104_SLICE_X2Y104_CO6;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_D2 = CLBLL_L_X2Y107_SLICE_X0Y107_AO6;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_D3 = CLBLM_R_X3Y104_SLICE_X3Y104_CO6;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_D4 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_D5 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_D6 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C1 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_A1 = CLBLL_L_X2Y108_SLICE_X0Y108_AO5;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_A2 = CLBLM_R_X3Y105_SLICE_X2Y105_AO6;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_A3 = CLBLM_R_X3Y106_SLICE_X2Y106_BO6;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_A4 = CLBLL_L_X2Y108_SLICE_X1Y108_BO6;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_A5 = CLBLM_R_X3Y109_SLICE_X2Y109_AO6;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_A6 = CLBLM_R_X3Y108_SLICE_X2Y108_DO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C4 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_B1 = CLBLM_R_X5Y110_SLICE_X6Y110_DO6;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_B2 = CLBLL_L_X4Y106_SLICE_X4Y106_AO5;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_B3 = CLBLL_L_X2Y107_SLICE_X0Y107_BO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_A4 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_A5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_A6 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_B4 = CLBLM_R_X3Y110_SLICE_X2Y110_AO6;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_B5 = CLBLM_R_X5Y102_SLICE_X6Y102_CO6;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_B6 = CLBLL_L_X4Y107_SLICE_X4Y107_BO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_A1 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_A2 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_B3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_B4 = CLBLM_L_X8Y110_SLICE_X11Y110_CO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_B5 = CLBLM_L_X8Y110_SLICE_X10Y110_AO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_B6 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_C1 = CLBLM_R_X5Y102_SLICE_X6Y102_CO6;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_C2 = CLBLL_L_X4Y106_SLICE_X4Y106_AO5;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_C3 = CLBLL_L_X4Y107_SLICE_X4Y107_BO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_C1 = CLBLM_R_X7Y110_SLICE_X9Y110_AO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_C2 = CLBLM_L_X8Y110_SLICE_X11Y110_CO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_C3 = CLBLM_L_X8Y112_SLICE_X10Y112_DO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_C4 = CLBLM_R_X7Y110_SLICE_X9Y110_AO5;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_C5 = CLBLM_R_X7Y111_SLICE_X8Y111_AO5;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_C6 = CLBLM_L_X8Y110_SLICE_X10Y110_AO6;
  assign CLBLM_R_X5Y100_SLICE_X7Y100_A1 = 1'b1;
  assign CLBLM_R_X5Y100_SLICE_X7Y100_A2 = 1'b1;
  assign CLBLM_R_X5Y100_SLICE_X7Y100_A3 = 1'b1;
  assign CLBLM_R_X5Y100_SLICE_X7Y100_A4 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_D1 = CLBLL_L_X2Y108_SLICE_X1Y108_AO6;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_D2 = CLBLM_R_X3Y105_SLICE_X2Y105_AO6;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_D3 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_D1 = CLBLM_R_X7Y110_SLICE_X9Y110_AO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_D2 = CLBLM_R_X7Y111_SLICE_X8Y111_AO5;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_D3 = CLBLM_L_X8Y112_SLICE_X10Y112_DO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_D4 = CLBLM_R_X7Y110_SLICE_X9Y110_AO5;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_D5 = CLBLM_L_X8Y110_SLICE_X10Y110_AO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_D6 = CLBLM_L_X8Y110_SLICE_X11Y110_CO6;
  assign CLBLM_R_X5Y100_SLICE_X7Y100_B4 = 1'b1;
  assign CLBLM_R_X5Y100_SLICE_X7Y100_B6 = 1'b1;
  assign CLBLM_R_X5Y100_SLICE_X7Y100_C1 = 1'b1;
  assign CLBLM_R_X5Y100_SLICE_X7Y100_C2 = 1'b1;
  assign CLBLM_R_X5Y100_SLICE_X7Y100_C3 = 1'b1;
  assign CLBLM_R_X5Y100_SLICE_X7Y100_C4 = 1'b1;
  assign CLBLM_R_X5Y100_SLICE_X7Y100_C5 = 1'b1;
  assign CLBLM_R_X5Y100_SLICE_X7Y100_C6 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_A1 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_A2 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_A3 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_A4 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_A5 = 1'b1;
  assign CLBLM_R_X5Y100_SLICE_X7Y100_D1 = 1'b1;
  assign CLBLM_R_X5Y100_SLICE_X7Y100_D2 = 1'b1;
  assign CLBLM_R_X5Y100_SLICE_X7Y100_D3 = 1'b1;
  assign CLBLM_R_X5Y100_SLICE_X7Y100_D4 = 1'b1;
  assign CLBLM_R_X5Y100_SLICE_X7Y100_D5 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_B5 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_B6 = 1'b1;
  assign CLBLM_R_X5Y100_SLICE_X7Y100_D6 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_B1 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_B2 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_B3 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_B4 = 1'b1;
  assign CLBLM_R_X5Y100_SLICE_X6Y100_A1 = CLBLM_R_X5Y100_SLICE_X6Y100_DO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_C4 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_C5 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_C6 = 1'b1;
  assign CLBLM_R_X5Y100_SLICE_X6Y100_A2 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X5Y100_SLICE_X6Y100_A3 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X5Y100_SLICE_X6Y100_A4 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X5Y100_SLICE_X6Y100_A5 = CLBLL_L_X4Y100_SLICE_X5Y100_DO6;
  assign CLBLM_R_X5Y100_SLICE_X6Y100_A6 = 1'b1;
  assign CLBLM_R_X5Y100_SLICE_X6Y100_B1 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X5Y100_SLICE_X6Y100_B2 = CLBLL_L_X4Y100_SLICE_X5Y100_CO6;
  assign CLBLM_R_X5Y100_SLICE_X6Y100_B3 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X5Y100_SLICE_X6Y100_B4 = CLBLM_R_X5Y102_SLICE_X7Y102_AO6;
  assign CLBLM_R_X5Y100_SLICE_X6Y100_B5 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X5Y100_SLICE_X6Y100_B6 = CLBLM_R_X5Y100_SLICE_X6Y100_CO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_D1 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_D2 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_D3 = 1'b1;
  assign CLBLM_R_X5Y100_SLICE_X6Y100_C1 = CLBLM_R_X5Y101_SLICE_X7Y101_AO6;
  assign CLBLM_R_X5Y100_SLICE_X6Y100_C2 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X5Y100_SLICE_X6Y100_C3 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X5Y100_SLICE_X6Y100_C4 = CLBLL_L_X4Y100_SLICE_X5Y100_DO6;
  assign CLBLM_R_X5Y100_SLICE_X6Y100_C5 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X5Y100_SLICE_X6Y100_C6 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_D5 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_D6 = 1'b1;
  assign CLBLM_R_X5Y100_SLICE_X6Y100_D1 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X5Y100_SLICE_X6Y100_D2 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X5Y100_SLICE_X6Y100_D3 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X5Y100_SLICE_X6Y100_D4 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X5Y100_SLICE_X6Y100_D5 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X5Y100_SLICE_X6Y100_D6 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_D1 = CLBLM_R_X3Y112_SLICE_X2Y112_AO6;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_T1 = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_D1 = CLBLL_L_X2Y113_SLICE_X1Y113_CO6;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_A1 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_A2 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_A3 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_A4 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_A5 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_A6 = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_T1 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_B1 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_B2 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_B3 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_B4 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_B5 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_B6 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_C1 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_C2 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_C3 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_C4 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_C5 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_C6 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_D1 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_D2 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_D3 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_D4 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_D5 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_D6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_D1 = CLBLL_L_X2Y113_SLICE_X0Y113_AO5;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_A1 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_A2 = CLBLM_R_X3Y109_SLICE_X2Y109_AO6;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_A3 = CLBLM_R_X3Y108_SLICE_X2Y108_DO6;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_A4 = CLBLM_R_X3Y106_SLICE_X2Y106_BO6;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_A5 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_A6 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_B1 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_B2 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_B3 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_B4 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_B5 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_B6 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_A1 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_A2 = CLBLM_R_X7Y110_SLICE_X9Y110_BO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_A3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_C1 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_C2 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_C3 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_C4 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_C5 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_C6 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_A4 = CLBLM_R_X7Y111_SLICE_X9Y111_BO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_A5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_A6 = CLBLM_R_X7Y111_SLICE_X9Y111_CO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_B1 = CLBLM_L_X8Y112_SLICE_X10Y112_DO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_B2 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_B3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_B4 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_D1 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_D2 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_D3 = 1'b1;
  assign CLBLM_R_X5Y101_SLICE_X7Y101_A4 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X5Y101_SLICE_X7Y101_A5 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X5Y101_SLICE_X7Y101_A6 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_D4 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_D5 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_D6 = 1'b1;
  assign CLBLM_R_X5Y101_SLICE_X7Y101_A1 = CLBLM_R_X5Y101_SLICE_X7Y101_DO6;
  assign CLBLM_R_X5Y101_SLICE_X7Y101_A2 = CLBLM_R_X5Y101_SLICE_X7Y101_CO6;
  assign CLBLM_R_X5Y101_SLICE_X7Y101_B1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X5Y101_SLICE_X7Y101_B2 = CLBLM_R_X5Y101_SLICE_X7Y101_CO6;
  assign CLBLM_R_X5Y101_SLICE_X7Y101_B3 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X5Y101_SLICE_X7Y101_B4 = CLBLM_R_X5Y100_SLICE_X6Y100_AO5;
  assign CLBLM_R_X5Y101_SLICE_X7Y101_B5 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X5Y101_SLICE_X7Y101_B6 = CLBLM_L_X8Y101_SLICE_X11Y101_BO6;
  assign CLBLM_R_X5Y101_SLICE_X7Y101_C1 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X5Y101_SLICE_X7Y101_C2 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X5Y101_SLICE_X7Y101_C3 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X5Y101_SLICE_X7Y101_C4 = CLBLM_R_X5Y103_SLICE_X6Y103_CO6;
  assign CLBLM_R_X5Y101_SLICE_X7Y101_C5 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X5Y101_SLICE_X7Y101_C6 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_D3 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_D4 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_A1 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_A2 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_A3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_A4 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_A5 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_A6 = 1'b1;
  assign CLBLM_R_X5Y101_SLICE_X7Y101_D1 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X5Y101_SLICE_X7Y101_D2 = CLBLM_L_X8Y101_SLICE_X11Y101_BO6;
  assign CLBLM_R_X5Y101_SLICE_X7Y101_D3 = CLBLM_R_X5Y100_SLICE_X6Y100_DO6;
  assign CLBLM_R_X5Y101_SLICE_X7Y101_D4 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X5Y101_SLICE_X7Y101_D5 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X5Y101_SLICE_X7Y101_D6 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_B1 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_B6 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_B2 = CLBLM_R_X7Y112_SLICE_X9Y112_BO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_B3 = CLBLM_R_X7Y112_SLICE_X8Y112_BO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_B4 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_B5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y101_SLICE_X6Y101_A1 = CLBLM_R_X7Y102_SLICE_X8Y102_BO6;
  assign CLBLM_R_X5Y101_SLICE_X6Y101_A2 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X5Y101_SLICE_X6Y101_A3 = CLBLM_R_X5Y100_SLICE_X6Y100_CO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_C3 = CLBLM_R_X7Y112_SLICE_X8Y112_BO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_C4 = CLBLM_R_X7Y112_SLICE_X9Y112_CO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_C5 = CLBLM_L_X8Y112_SLICE_X10Y112_CO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_C6 = CLBLM_R_X5Y112_SLICE_X7Y112_AO5;
  assign CLBLM_R_X5Y101_SLICE_X6Y101_A4 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X5Y101_SLICE_X6Y101_A5 = CLBLM_R_X5Y102_SLICE_X7Y102_AO6;
  assign CLBLM_R_X5Y101_SLICE_X6Y101_A6 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_C1 = CLBLM_R_X7Y110_SLICE_X9Y110_AO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_C2 = CLBLM_R_X7Y111_SLICE_X8Y111_AO6;
  assign CLBLM_R_X5Y101_SLICE_X6Y101_B1 = CLBLM_R_X7Y102_SLICE_X8Y102_BO6;
  assign CLBLM_R_X5Y101_SLICE_X6Y101_B2 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X5Y101_SLICE_X6Y101_B3 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X5Y101_SLICE_X6Y101_B4 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X5Y101_SLICE_X6Y101_B5 = CLBLM_R_X5Y101_SLICE_X6Y101_CO6;
  assign CLBLM_R_X5Y101_SLICE_X6Y101_B6 = CLBLM_R_X5Y101_SLICE_X6Y101_AO5;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_D1 = CLBLM_R_X7Y110_SLICE_X9Y110_AO6;
  assign CLBLM_R_X5Y101_SLICE_X6Y101_C1 = CLBLM_R_X5Y102_SLICE_X7Y102_AO6;
  assign CLBLM_R_X5Y101_SLICE_X6Y101_C2 = CLBLM_R_X5Y100_SLICE_X6Y100_CO6;
  assign CLBLM_R_X5Y101_SLICE_X6Y101_C3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X5Y101_SLICE_X6Y101_C4 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X5Y101_SLICE_X6Y101_C5 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X5Y101_SLICE_X6Y101_C6 = CLBLL_L_X4Y100_SLICE_X5Y100_CO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_D3 = CLBLM_R_X7Y112_SLICE_X8Y112_BO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_D4 = CLBLM_R_X7Y112_SLICE_X9Y112_CO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_D5 = CLBLM_L_X8Y112_SLICE_X10Y112_CO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_D6 = CLBLM_R_X5Y112_SLICE_X7Y112_AO5;
  assign CLBLM_R_X5Y101_SLICE_X6Y101_D1 = CLBLM_R_X5Y101_SLICE_X6Y101_CO6;
  assign CLBLM_R_X5Y101_SLICE_X6Y101_D2 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X5Y101_SLICE_X6Y101_D3 = CLBLM_R_X7Y102_SLICE_X8Y102_BO6;
  assign CLBLM_R_X5Y101_SLICE_X6Y101_D4 = CLBLM_R_X5Y101_SLICE_X6Y101_AO5;
  assign CLBLM_R_X5Y101_SLICE_X6Y101_D5 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X5Y101_SLICE_X6Y101_D6 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y106_D = RIOB33_X105Y105_IOB_X1Y106_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y105_D = RIOB33_X105Y105_IOB_X1Y105_I;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y108_D = LIOB33_X0Y107_IOB_X0Y108_I;
  assign LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y107_D = LIOB33_X0Y107_IOB_X0Y107_I;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_D = RIOB33_X105Y113_IOB_X1Y113_I;
  assign RIOI3_SING_X105Y100_ILOGIC_X1Y100_D = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_A1 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_A2 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_A3 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_A4 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_A5 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_A6 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_B1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_B2 = CLBLM_L_X8Y112_SLICE_X10Y112_AO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_B3 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_B4 = CLBLM_R_X7Y113_SLICE_X8Y113_AO5;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_B5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_B6 = CLBLM_L_X8Y112_SLICE_X10Y112_BO6;
  assign CLBLM_R_X5Y102_SLICE_X7Y102_A1 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X5Y102_SLICE_X7Y102_A2 = CLBLM_R_X7Y101_SLICE_X9Y101_CO6;
  assign CLBLM_R_X5Y102_SLICE_X7Y102_A3 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X5Y102_SLICE_X7Y102_A4 = CLBLM_R_X5Y102_SLICE_X7Y102_BO6;
  assign CLBLM_R_X5Y102_SLICE_X7Y102_A5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y102_SLICE_X7Y102_A6 = CLBLM_R_X5Y101_SLICE_X7Y101_BO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_C1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_C2 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_C3 = CLBLM_R_X7Y113_SLICE_X9Y113_DO6;
  assign CLBLM_R_X5Y102_SLICE_X7Y102_B1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X5Y102_SLICE_X7Y102_B2 = CLBLM_R_X5Y100_SLICE_X6Y100_DO6;
  assign CLBLM_R_X5Y102_SLICE_X7Y102_B3 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X5Y102_SLICE_X7Y102_B4 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X5Y102_SLICE_X7Y102_B5 = CLBLM_L_X8Y101_SLICE_X11Y101_BO6;
  assign CLBLM_R_X5Y102_SLICE_X7Y102_B6 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_D1 = CLBLM_R_X7Y112_SLICE_X9Y112_AO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_D2 = CLBLM_R_X5Y113_SLICE_X6Y113_CO6;
  assign CLBLM_R_X5Y102_SLICE_X7Y102_C1 = 1'b1;
  assign CLBLM_R_X5Y102_SLICE_X7Y102_C2 = 1'b1;
  assign CLBLM_R_X5Y102_SLICE_X7Y102_C3 = 1'b1;
  assign CLBLM_R_X5Y102_SLICE_X7Y102_C4 = 1'b1;
  assign CLBLM_R_X5Y102_SLICE_X7Y102_C5 = 1'b1;
  assign CLBLM_R_X5Y102_SLICE_X7Y102_C6 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_D3 = CLBLM_R_X7Y113_SLICE_X9Y113_DO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_D4 = CLBLM_L_X8Y112_SLICE_X11Y112_DO6;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_A1 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_A2 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_A3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_A4 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_A5 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_A6 = 1'b1;
  assign CLBLM_R_X5Y102_SLICE_X7Y102_D1 = 1'b1;
  assign CLBLM_R_X5Y102_SLICE_X7Y102_D2 = 1'b1;
  assign CLBLM_R_X5Y102_SLICE_X7Y102_D3 = 1'b1;
  assign CLBLM_R_X5Y102_SLICE_X7Y102_D4 = 1'b1;
  assign CLBLM_R_X5Y102_SLICE_X7Y102_D5 = 1'b1;
  assign CLBLM_R_X5Y102_SLICE_X7Y102_D6 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_B1 = CLBLM_R_X7Y113_SLICE_X9Y113_CO6;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_B2 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_B3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_B4 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_B5 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X5Y102_SLICE_X6Y102_A1 = CLBLM_R_X5Y102_SLICE_X6Y102_BO5;
  assign CLBLM_R_X5Y102_SLICE_X6Y102_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y102_SLICE_X6Y102_A3 = CLBLM_R_X7Y103_SLICE_X8Y103_AO6;
  assign CLBLM_R_X5Y102_SLICE_X6Y102_A4 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X5Y102_SLICE_X6Y102_A5 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X5Y102_SLICE_X6Y102_A6 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_C1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_C2 = CLBLM_R_X7Y112_SLICE_X9Y112_CO6;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_C3 = CLBLM_L_X8Y112_SLICE_X10Y112_CO6;
  assign CLBLM_R_X5Y102_SLICE_X6Y102_B1 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X5Y102_SLICE_X6Y102_B2 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X5Y102_SLICE_X6Y102_B3 = CLBLM_R_X5Y101_SLICE_X6Y101_AO6;
  assign CLBLM_R_X5Y102_SLICE_X6Y102_B4 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X5Y102_SLICE_X6Y102_B5 = 1'b1;
  assign CLBLM_R_X5Y102_SLICE_X6Y102_B6 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_D1 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_D2 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_D3 = 1'b1;
  assign CLBLM_R_X5Y102_SLICE_X6Y102_C1 = CLBLM_R_X5Y101_SLICE_X6Y101_BO6;
  assign CLBLM_R_X5Y102_SLICE_X6Y102_C2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y102_SLICE_X6Y102_C3 = CLBLM_R_X7Y103_SLICE_X8Y103_AO6;
  assign CLBLM_R_X5Y102_SLICE_X6Y102_C4 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X5Y102_SLICE_X6Y102_C5 = CLBLM_R_X5Y102_SLICE_X6Y102_BO5;
  assign CLBLM_R_X5Y102_SLICE_X6Y102_C6 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_D4 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_D5 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_D6 = 1'b1;
  assign CLBLM_R_X5Y102_SLICE_X6Y102_D1 = CLBLM_R_X5Y101_SLICE_X6Y101_AO6;
  assign CLBLM_R_X5Y102_SLICE_X6Y102_D2 = CLBLM_R_X7Y103_SLICE_X8Y103_AO6;
  assign CLBLM_R_X5Y102_SLICE_X6Y102_D3 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X5Y102_SLICE_X6Y102_D4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y102_SLICE_X6Y102_D5 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X5Y102_SLICE_X6Y102_D6 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_A1 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_A2 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_A3 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_A4 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_A5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_A6 = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_D1 = CLBLM_R_X3Y111_SLICE_X2Y111_BO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_B1 = CLBLM_R_X7Y112_SLICE_X8Y112_AO5;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_B2 = CLBLM_R_X7Y113_SLICE_X8Y113_BO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_B3 = CLBLM_L_X8Y112_SLICE_X11Y112_AO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_B4 = CLBLM_L_X8Y113_SLICE_X11Y113_AO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_B5 = CLBLM_R_X7Y113_SLICE_X9Y113_AO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_B6 = CLBLM_R_X5Y111_SLICE_X7Y111_BO6;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_T1 = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_T1 = 1'b1;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_A1 = 1'b1;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_A2 = 1'b1;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_A3 = 1'b1;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_A4 = 1'b1;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_A5 = 1'b1;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_A6 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_C1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_C2 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_C3 = CLBLM_R_X7Y113_SLICE_X8Y113_BO6;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_B1 = 1'b1;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_B2 = 1'b1;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_B3 = 1'b1;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_B4 = 1'b1;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_B5 = 1'b1;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_B6 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_D1 = CLBLM_R_X7Y113_SLICE_X9Y113_AO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_D5 = CLBLM_L_X8Y112_SLICE_X11Y112_AO6;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_C1 = 1'b1;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_C2 = 1'b1;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_C3 = 1'b1;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_C4 = 1'b1;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_C5 = 1'b1;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_C6 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_D6 = CLBLM_L_X8Y113_SLICE_X11Y113_AO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_A1 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_A2 = CLBLM_R_X5Y111_SLICE_X7Y111_BO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_A3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_A4 = CLBLM_R_X7Y113_SLICE_X8Y113_BO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_A5 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_A6 = 1'b1;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_D1 = 1'b1;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_D2 = 1'b1;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_D3 = 1'b1;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_D4 = 1'b1;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_D5 = 1'b1;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_D6 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_B1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_B2 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_B3 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_B4 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_B5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_A1 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_A2 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_A3 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_A4 = CLBLM_R_X5Y103_SLICE_X6Y103_BO6;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_A5 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_A6 = CLBLM_R_X7Y104_SLICE_X8Y104_CO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_C1 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_C2 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_C3 = 1'b1;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_B1 = CLBLM_R_X7Y103_SLICE_X8Y103_DO6;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_B2 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_B3 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_B4 = CLBLM_R_X7Y104_SLICE_X8Y104_DO6;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_B5 = CLBLM_R_X7Y102_SLICE_X9Y102_DO6;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_B6 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_D1 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_D2 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_D3 = 1'b1;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_C1 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_C2 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_C3 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_C4 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_C5 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_C6 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_D4 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_D5 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_D6 = 1'b1;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_D1 = CLBLM_R_X7Y102_SLICE_X9Y102_DO6;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_D2 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_D3 = CLBLM_R_X7Y103_SLICE_X9Y103_CO6;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_D4 = CLBLM_R_X7Y104_SLICE_X8Y104_DO6;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_D5 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_D6 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_A1 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_A2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_A3 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_A4 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_A5 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_A6 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_B1 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_B2 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_B3 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_B4 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_B5 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_B6 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_C1 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_C2 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_C3 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_C4 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_C5 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_C6 = 1'b1;
  assign RIOI3_X105Y109_ILOGIC_X1Y110_D = RIOB33_X105Y109_IOB_X1Y110_I;
  assign RIOI3_X105Y109_ILOGIC_X1Y109_D = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_D1 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_D2 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_D3 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_D4 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_D5 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_D6 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_A1 = CLBLM_R_X3Y113_SLICE_X2Y113_CO6;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_A2 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_A3 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_A4 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_A5 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_A6 = CLBLL_L_X2Y113_SLICE_X1Y113_DO6;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_C4 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_B1 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_B2 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_B3 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_B4 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_B5 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_B6 = 1'b1;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_C5 = 1'b1;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_C6 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_C1 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_C2 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_C3 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_C4 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_C5 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_C6 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_D1 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_D2 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_D3 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_D4 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_D5 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_D6 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_A1 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_A2 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_A3 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_A4 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_A5 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_A6 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_B1 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_B2 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_B3 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_B4 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_B5 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_B6 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_C1 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_C2 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_C3 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_C4 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_C5 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_C6 = 1'b1;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_D3 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_D1 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_D2 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_D3 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_D4 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_D5 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_D6 = 1'b1;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_D5 = 1'b1;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_D6 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_A1 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_A2 = CLBLM_R_X7Y104_SLICE_X8Y104_CO6;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_A3 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_A4 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_A5 = CLBLM_R_X5Y103_SLICE_X6Y103_BO6;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_A6 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_B1 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_B2 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_B3 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_B4 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_B5 = CLBLM_R_X5Y105_SLICE_X6Y105_AO6;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_B6 = CLBLM_R_X7Y105_SLICE_X8Y105_BO6;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_C1 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_C2 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_C3 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_C4 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_C5 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_C6 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_D1 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_D2 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_D3 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_D4 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_D5 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_D6 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_A1 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_A2 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_A3 = CLBLL_L_X2Y112_SLICE_X0Y112_AO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_A4 = CLBLL_L_X2Y112_SLICE_X0Y112_BO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_A5 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_A6 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_B1 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_B2 = CLBLL_L_X2Y113_SLICE_X0Y113_CO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_B3 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_B4 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_B5 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_B6 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_C1 = CLBLL_L_X2Y112_SLICE_X0Y112_AO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_C2 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_C3 = CLBLM_R_X3Y114_SLICE_X2Y114_AO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_C4 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_C5 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_C6 = CLBLL_L_X2Y112_SLICE_X0Y112_BO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_D1 = CLBLL_L_X2Y112_SLICE_X0Y112_AO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_D2 = CLBLM_R_X3Y113_SLICE_X3Y113_AO5;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_D3 = CLBLL_L_X2Y114_SLICE_X0Y114_BO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_D4 = CLBLM_R_X3Y114_SLICE_X2Y114_AO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_D5 = CLBLL_L_X2Y112_SLICE_X0Y112_BO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_D6 = CLBLL_L_X2Y113_SLICE_X0Y113_BO6;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_A1 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_A2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_A3 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_A4 = CLBLL_L_X2Y113_SLICE_X1Y113_BO6;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_A5 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_A6 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_B1 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_B2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_B3 = CLBLL_L_X2Y113_SLICE_X0Y113_AO6;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_B4 = CLBLM_R_X3Y114_SLICE_X2Y114_BO6;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_B5 = CLBLM_R_X3Y113_SLICE_X2Y113_AO6;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_B6 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_C1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_C2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_C3 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_C4 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_C5 = CLBLL_L_X2Y113_SLICE_X1Y113_DO6;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_C6 = CLBLM_R_X3Y113_SLICE_X2Y113_CO6;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_D1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_D2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_D3 = CLBLL_L_X2Y113_SLICE_X0Y113_DO6;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_D4 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_D5 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_D6 = CLBLM_R_X3Y114_SLICE_X2Y114_BO6;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_A1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_A2 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_A3 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_A4 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_A5 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_A6 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_B1 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_B2 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_B3 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_B4 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_B5 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_B6 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_C1 = CLBLM_R_X7Y105_SLICE_X8Y105_AO6;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_C2 = CLBLM_R_X7Y105_SLICE_X8Y105_CO6;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_C3 = CLBLM_L_X8Y106_SLICE_X11Y106_DO6;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_C4 = CLBLM_R_X5Y105_SLICE_X7Y105_AO5;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_C5 = CLBLM_R_X7Y103_SLICE_X9Y103_CO6;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_C6 = CLBLM_R_X5Y105_SLICE_X7Y105_BO5;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_D1 = CLBLM_R_X5Y105_SLICE_X7Y105_AO6;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_D2 = CLBLM_R_X7Y105_SLICE_X8Y105_AO6;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_D3 = CLBLM_L_X8Y106_SLICE_X10Y106_DO6;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_D4 = CLBLM_R_X5Y105_SLICE_X7Y105_AO5;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_D5 = CLBLM_L_X8Y106_SLICE_X11Y106_DO6;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_D6 = CLBLM_L_X8Y106_SLICE_X11Y106_BO6;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_A1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_A2 = CLBLM_L_X8Y105_SLICE_X11Y105_AO6;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_A3 = CLBLM_L_X8Y107_SLICE_X10Y107_BO6;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_A4 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_A5 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_A6 = CLBLM_L_X8Y106_SLICE_X11Y106_BO6;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_B1 = CLBLM_R_X5Y107_SLICE_X6Y107_AO6;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_B2 = CLBLM_R_X7Y104_SLICE_X8Y104_AO6;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_B3 = CLBLL_L_X4Y104_SLICE_X5Y104_AO6;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_B4 = CLBLM_R_X5Y106_SLICE_X6Y106_AO6;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_B5 = CLBLM_R_X5Y105_SLICE_X6Y105_AO6;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_B6 = CLBLM_R_X5Y106_SLICE_X6Y106_BO6;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_C1 = CLBLM_R_X5Y105_SLICE_X6Y105_AO6;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_C2 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_C3 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_C4 = CLBLM_R_X7Y105_SLICE_X8Y105_BO6;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_C5 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_C6 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_D1 = CLBLL_L_X4Y104_SLICE_X5Y104_AO6;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_D2 = CLBLM_R_X5Y106_SLICE_X6Y106_BO6;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_D3 = CLBLM_R_X5Y105_SLICE_X7Y105_DO6;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_D4 = CLBLM_R_X5Y106_SLICE_X6Y106_AO6;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_D5 = CLBLM_R_X5Y107_SLICE_X6Y107_AO6;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_D6 = CLBLL_L_X4Y105_SLICE_X4Y105_AO6;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_D1 = CLBLM_R_X3Y111_SLICE_X3Y111_AO6;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_D1 = CLBLL_L_X4Y107_SLICE_X4Y107_AO6;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_T1 = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_D1 = CLBLL_L_X4Y110_SLICE_X4Y110_AO5;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_D1 = CLBLM_R_X3Y110_SLICE_X2Y110_BO6;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_D1 = CLBLM_R_X3Y110_SLICE_X2Y110_AO5;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_T1 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_A1 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_A2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_A3 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_A4 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_A5 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_A6 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_B1 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_B2 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_B3 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_B4 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_B5 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_B6 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_C1 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_C2 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_C3 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_C4 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_C5 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_C6 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_D1 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_D2 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_D3 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_D4 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_D5 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_D6 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_A1 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_A2 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_A3 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_A4 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_A5 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_A6 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_B1 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_B2 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_B3 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_B4 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_B5 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_B6 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_C1 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_C2 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_C3 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_C4 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_C5 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_C6 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_D1 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_D2 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_D3 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_D4 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_D5 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_D6 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_A1 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_A2 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_A3 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_A4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_A5 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_A6 = 1'b1;
  assign RIOI3_X105Y103_ILOGIC_X1Y104_D = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_B1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_B2 = CLBLM_L_X8Y106_SLICE_X10Y106_CO6;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_B3 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_B4 = CLBLM_L_X8Y107_SLICE_X11Y107_DO6;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_B5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_B6 = CLBLM_L_X8Y107_SLICE_X10Y107_CO6;
  assign RIOI3_X105Y111_ILOGIC_X1Y112_D = RIOB33_X105Y111_IOB_X1Y112_I;
  assign RIOI3_X105Y111_ILOGIC_X1Y111_D = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_C1 = CLBLM_R_X5Y106_SLICE_X7Y106_AO6;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_C2 = CLBLM_L_X8Y106_SLICE_X10Y106_BO6;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_C3 = CLBLM_R_X7Y107_SLICE_X9Y107_DO6;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_C4 = CLBLM_L_X8Y106_SLICE_X10Y106_DO6;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_C5 = CLBLM_R_X5Y105_SLICE_X7Y105_AO6;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_C6 = CLBLM_L_X8Y106_SLICE_X11Y106_BO6;
  assign RIOI3_X105Y103_ILOGIC_X1Y103_D = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_D1 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_D2 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_D3 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_D4 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_D5 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_D6 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_A1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_A2 = CLBLM_L_X8Y105_SLICE_X11Y105_AO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_A3 = CLBLM_L_X8Y106_SLICE_X11Y106_BO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_A4 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_A5 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_A6 = CLBLM_L_X8Y107_SLICE_X10Y107_BO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_B1 = CLBLM_L_X8Y107_SLICE_X11Y107_DO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_B2 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_B3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_B4 = CLBLM_L_X8Y106_SLICE_X10Y106_BO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_B5 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_B6 = CLBLM_L_X8Y107_SLICE_X10Y107_CO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_C1 = CLBLM_L_X8Y105_SLICE_X11Y105_AO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_C2 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_C3 = CLBLM_L_X8Y106_SLICE_X11Y106_CO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_C4 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_C5 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_C6 = CLBLM_L_X8Y107_SLICE_X10Y107_BO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_D1 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_D2 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_D3 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_D4 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_D5 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_D6 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_A1 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_A2 = CLBLM_R_X7Y107_SLICE_X8Y107_BO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_A3 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_A4 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_A5 = CLBLM_R_X7Y107_SLICE_X8Y107_CO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_A6 = CLBLM_R_X5Y108_SLICE_X7Y108_CO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_B1 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_B2 = CLBLM_R_X7Y107_SLICE_X8Y107_BO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_B3 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_B4 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_B5 = CLBLM_R_X7Y107_SLICE_X8Y107_AO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_B6 = CLBLM_R_X5Y108_SLICE_X7Y108_CO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_C1 = CLBLM_R_X5Y106_SLICE_X7Y106_AO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_C2 = CLBLM_R_X5Y106_SLICE_X7Y106_AO5;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_C3 = CLBLM_R_X7Y107_SLICE_X9Y107_DO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_C4 = CLBLM_R_X7Y107_SLICE_X8Y107_DO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_C5 = CLBLM_R_X7Y107_SLICE_X9Y107_BO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_C6 = CLBLM_L_X8Y106_SLICE_X10Y106_BO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_D1 = CLBLM_R_X7Y107_SLICE_X8Y107_AO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_D2 = CLBLM_R_X7Y107_SLICE_X8Y107_DO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_D3 = CLBLL_L_X4Y107_SLICE_X4Y107_AO5;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_D4 = CLBLM_R_X5Y106_SLICE_X7Y106_AO5;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_D5 = CLBLM_R_X7Y107_SLICE_X9Y107_BO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_D6 = CLBLM_R_X7Y108_SLICE_X8Y108_CO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_A1 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_A2 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_A3 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_A4 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_A5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_A6 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_B1 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_B2 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_B3 = CLBLM_R_X7Y107_SLICE_X8Y107_AO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_B4 = CLBLM_R_X7Y107_SLICE_X8Y107_BO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_B5 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_B6 = CLBLM_R_X5Y108_SLICE_X7Y108_CO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_C1 = CLBLM_R_X5Y107_SLICE_X6Y107_AO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_C2 = CLBLM_R_X7Y106_SLICE_X8Y106_CO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_C3 = CLBLM_R_X5Y106_SLICE_X6Y106_AO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_C4 = CLBLM_R_X5Y107_SLICE_X6Y107_AO5;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_C5 = CLBLM_R_X5Y107_SLICE_X6Y107_DO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_C6 = CLBLM_R_X5Y106_SLICE_X6Y106_BO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_D1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_D2 = CLBLM_L_X8Y106_SLICE_X10Y106_BO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_D3 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_D4 = CLBLM_L_X8Y107_SLICE_X11Y107_DO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_D5 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_D6 = CLBLM_L_X8Y107_SLICE_X10Y107_CO6;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_D1 = CLBLL_L_X2Y114_SLICE_X0Y114_BO5;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_T1 = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_D1 = CLBLM_R_X3Y110_SLICE_X3Y110_BO6;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_D1 = CLBLL_L_X2Y104_SLICE_X1Y104_CO6;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_D1 = CLBLL_L_X2Y106_SLICE_X0Y106_BO6;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_T1 = 1'b1;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_A1 = 1'b1;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_A2 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_A3 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_A4 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_A5 = 1'b1;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_A6 = 1'b1;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_B1 = CLBLM_R_X5Y110_SLICE_X7Y110_CO6;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_B2 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_B3 = CLBLM_R_X7Y111_SLICE_X9Y111_AO6;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_B4 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_B5 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_B6 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_C1 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_C2 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_C3 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_C4 = CLBLM_R_X5Y110_SLICE_X7Y110_CO6;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_C5 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_C6 = CLBLM_R_X7Y111_SLICE_X9Y111_AO6;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_D1 = CLBLM_R_X5Y108_SLICE_X7Y108_AO6;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_D2 = CLBLL_L_X4Y107_SLICE_X5Y107_AO5;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_D3 = CLBLM_R_X5Y107_SLICE_X7Y107_BO6;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_D4 = CLBLM_R_X5Y107_SLICE_X6Y107_AO5;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_D5 = CLBLM_R_X7Y106_SLICE_X8Y106_BO6;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_D6 = CLBLM_R_X5Y107_SLICE_X7Y107_CO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_A1 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_A2 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_A3 = 1'b1;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_A4 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_A5 = 1'b1;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_A6 = 1'b1;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_B1 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_B2 = CLBLM_R_X5Y108_SLICE_X7Y108_BO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_B3 = CLBLM_R_X5Y109_SLICE_X6Y109_DO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_B4 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_B5 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_B6 = CLBLM_R_X7Y108_SLICE_X8Y108_BO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_C1 = CLBLM_R_X7Y106_SLICE_X8Y106_BO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_C2 = CLBLM_R_X5Y107_SLICE_X6Y107_AO5;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_C3 = CLBLM_R_X7Y106_SLICE_X8Y106_CO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_C4 = CLBLL_L_X4Y107_SLICE_X5Y107_AO5;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_C5 = CLBLM_R_X5Y107_SLICE_X6Y107_DO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_C6 = CLBLM_R_X5Y107_SLICE_X7Y107_BO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_D1 = CLBLM_R_X5Y107_SLICE_X6Y107_AO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_D2 = CLBLM_R_X5Y108_SLICE_X7Y108_AO5;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_D3 = CLBLM_R_X7Y106_SLICE_X8Y106_CO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_D4 = CLBLM_R_X5Y107_SLICE_X6Y107_AO5;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_D5 = CLBLM_R_X5Y107_SLICE_X6Y107_DO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_D6 = CLBLM_R_X5Y106_SLICE_X7Y106_CO6;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_C3 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_C4 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_A1 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_A2 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_A3 = CLBLM_R_X5Y110_SLICE_X7Y110_AO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_A4 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_A5 = CLBLM_L_X8Y103_SLICE_X11Y103_AO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_A6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_B1 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_B2 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_B3 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_B4 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_B5 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_B6 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_C1 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_C2 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_C3 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_C4 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_C5 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_C6 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_D1 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_D2 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_D3 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_D4 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_D5 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_D6 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_A1 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_A2 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_A3 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_A4 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_A5 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_A6 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_B1 = CLBLM_R_X5Y110_SLICE_X7Y110_CO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_B2 = CLBLM_R_X7Y108_SLICE_X8Y108_AO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_B3 = CLBLM_R_X7Y109_SLICE_X8Y109_AO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_B4 = CLBLM_R_X5Y110_SLICE_X7Y110_BO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_B5 = CLBLM_R_X5Y109_SLICE_X6Y109_AO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_B6 = CLBLM_R_X5Y110_SLICE_X6Y110_CO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_C1 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_C2 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_C3 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_C4 = CLBLM_R_X5Y110_SLICE_X6Y110_CO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_C5 = CLBLM_R_X5Y110_SLICE_X7Y110_DO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_C6 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_D1 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_D2 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_D3 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_D4 = CLBLM_R_X5Y110_SLICE_X6Y110_CO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_D5 = CLBLM_R_X5Y110_SLICE_X7Y110_DO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_D6 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_A1 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_A2 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_A3 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_A4 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_A5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_A6 = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_D1 = 1'b0;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_B1 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_B2 = CLBLM_R_X5Y112_SLICE_X6Y112_DO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_B3 = CLBLM_R_X7Y111_SLICE_X8Y111_BO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_B4 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_B5 = CLBLM_R_X7Y111_SLICE_X8Y111_CO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_B6 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y100_SLICE_X3Y100_A1 = CLBLM_R_X3Y101_SLICE_X3Y101_DO6;
  assign CLBLM_R_X3Y100_SLICE_X3Y100_A2 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X3Y100_SLICE_X3Y100_A3 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X3Y100_SLICE_X3Y100_A4 = CLBLM_R_X3Y100_SLICE_X3Y100_BO6;
  assign CLBLM_R_X3Y100_SLICE_X3Y100_A5 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X3Y100_SLICE_X3Y100_A6 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_C1 = CLBLM_R_X7Y111_SLICE_X8Y111_BO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_C2 = CLBLM_R_X5Y112_SLICE_X6Y112_DO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_C3 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X3Y100_SLICE_X3Y100_B1 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X3Y100_SLICE_X3Y100_B2 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X3Y100_SLICE_X3Y100_B3 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X3Y100_SLICE_X3Y100_B4 = CLBLL_L_X4Y100_SLICE_X4Y100_AO6;
  assign CLBLM_R_X3Y100_SLICE_X3Y100_B5 = CLBLL_L_X4Y100_SLICE_X4Y100_BO6;
  assign CLBLM_R_X3Y100_SLICE_X3Y100_B6 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_D1 = CLBLM_R_X7Y111_SLICE_X8Y111_BO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_D2 = CLBLM_R_X7Y112_SLICE_X8Y112_CO6;
  assign CLBLM_R_X3Y100_SLICE_X3Y100_C1 = 1'b1;
  assign CLBLM_R_X3Y100_SLICE_X3Y100_C2 = 1'b1;
  assign CLBLM_R_X3Y100_SLICE_X3Y100_C3 = 1'b1;
  assign CLBLM_R_X3Y100_SLICE_X3Y100_C4 = 1'b1;
  assign CLBLM_R_X3Y100_SLICE_X3Y100_C5 = 1'b1;
  assign CLBLM_R_X3Y100_SLICE_X3Y100_C6 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_D3 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_D4 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_A1 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_A2 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_A3 = CLBLM_R_X7Y111_SLICE_X8Y111_BO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_A4 = CLBLM_R_X5Y112_SLICE_X6Y112_DO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_A5 = CLBLL_L_X4Y111_SLICE_X5Y111_DO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_A6 = 1'b1;
  assign CLBLM_R_X3Y100_SLICE_X3Y100_D1 = 1'b1;
  assign CLBLM_R_X3Y100_SLICE_X3Y100_D2 = 1'b1;
  assign CLBLM_R_X3Y100_SLICE_X3Y100_D3 = 1'b1;
  assign CLBLM_R_X3Y100_SLICE_X3Y100_D4 = 1'b1;
  assign CLBLM_R_X3Y100_SLICE_X3Y100_D5 = 1'b1;
  assign CLBLM_R_X3Y100_SLICE_X3Y100_D6 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_B1 = CLBLM_R_X5Y113_SLICE_X6Y113_DO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_B2 = CLBLM_R_X5Y111_SLICE_X7Y111_BO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_B3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_B4 = CLBLM_R_X5Y110_SLICE_X7Y110_AO5;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_B5 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X3Y100_SLICE_X2Y100_A1 = 1'b1;
  assign CLBLM_R_X3Y100_SLICE_X2Y100_A2 = 1'b1;
  assign CLBLM_R_X3Y100_SLICE_X2Y100_A3 = 1'b1;
  assign CLBLM_R_X3Y100_SLICE_X2Y100_A4 = 1'b1;
  assign CLBLM_R_X3Y100_SLICE_X2Y100_A5 = 1'b1;
  assign CLBLM_R_X3Y100_SLICE_X2Y100_A6 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_C1 = CLBLM_R_X7Y111_SLICE_X8Y111_BO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_C2 = CLBLL_L_X4Y111_SLICE_X5Y111_DO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_C3 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y100_SLICE_X2Y100_B1 = 1'b1;
  assign CLBLM_R_X3Y100_SLICE_X2Y100_B2 = 1'b1;
  assign CLBLM_R_X3Y100_SLICE_X2Y100_B3 = 1'b1;
  assign CLBLM_R_X3Y100_SLICE_X2Y100_B4 = 1'b1;
  assign CLBLM_R_X3Y100_SLICE_X2Y100_B5 = 1'b1;
  assign CLBLM_R_X3Y100_SLICE_X2Y100_B6 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_D1 = CLBLM_R_X5Y109_SLICE_X7Y109_AO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_D2 = CLBLL_L_X4Y101_SLICE_X4Y101_AO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_D3 = CLBLM_R_X5Y113_SLICE_X6Y113_DO6;
  assign CLBLM_R_X3Y100_SLICE_X2Y100_C1 = 1'b1;
  assign CLBLM_R_X3Y100_SLICE_X2Y100_C2 = 1'b1;
  assign CLBLM_R_X3Y100_SLICE_X2Y100_C3 = 1'b1;
  assign CLBLM_R_X3Y100_SLICE_X2Y100_C4 = 1'b1;
  assign CLBLM_R_X3Y100_SLICE_X2Y100_C5 = 1'b1;
  assign CLBLM_R_X3Y100_SLICE_X2Y100_C6 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_D4 = CLBLM_L_X8Y111_SLICE_X10Y111_CO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_D5 = CLBLM_R_X3Y110_SLICE_X3Y110_DO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_D6 = CLBLM_R_X5Y112_SLICE_X6Y112_DO6;
  assign CLBLM_R_X3Y100_SLICE_X2Y100_D1 = 1'b1;
  assign CLBLM_R_X3Y100_SLICE_X2Y100_D2 = 1'b1;
  assign CLBLM_R_X3Y100_SLICE_X2Y100_D3 = 1'b1;
  assign CLBLM_R_X3Y100_SLICE_X2Y100_D4 = 1'b1;
  assign CLBLM_R_X3Y100_SLICE_X2Y100_D5 = 1'b1;
  assign CLBLM_R_X3Y100_SLICE_X2Y100_D6 = 1'b1;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_A1 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_A2 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_A3 = 1'b1;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_A4 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_A5 = 1'b1;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_A6 = 1'b1;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_B1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_B2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_B3 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_B4 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_B5 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_B6 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X3Y101_SLICE_X3Y101_A1 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X3Y101_SLICE_X3Y101_A2 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_C3 = CLBLM_R_X5Y112_SLICE_X7Y112_CO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_C4 = CLBLM_R_X3Y111_SLICE_X3Y111_AO5;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_C5 = CLBLM_R_X7Y111_SLICE_X8Y111_CO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_C6 = CLBLM_R_X5Y112_SLICE_X7Y112_BO6;
  assign CLBLM_R_X3Y101_SLICE_X3Y101_A3 = CLBLL_L_X4Y100_SLICE_X4Y100_BO6;
  assign CLBLM_R_X3Y101_SLICE_X3Y101_A4 = CLBLM_R_X3Y101_SLICE_X3Y101_BO6;
  assign CLBLM_R_X3Y101_SLICE_X3Y101_A5 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X3Y101_SLICE_X3Y101_A6 = 1'b1;
  assign CLBLM_R_X3Y101_SLICE_X3Y101_B1 = CLBLL_L_X4Y101_SLICE_X4Y101_DO6;
  assign CLBLM_R_X3Y101_SLICE_X3Y101_B2 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X3Y101_SLICE_X3Y101_B3 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X3Y101_SLICE_X3Y101_B4 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y101_SLICE_X3Y101_B5 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X3Y101_SLICE_X3Y101_B6 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_D1 = CLBLM_R_X5Y111_SLICE_X7Y111_AO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_D5 = CLBLM_R_X7Y111_SLICE_X8Y111_CO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_D6 = CLBLM_R_X5Y112_SLICE_X7Y112_BO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_D2 = CLBLM_R_X7Y110_SLICE_X9Y110_DO6;
  assign CLBLM_R_X3Y101_SLICE_X3Y101_C1 = CLBLL_L_X4Y100_SLICE_X4Y100_AO6;
  assign CLBLM_R_X3Y101_SLICE_X3Y101_C2 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X3Y101_SLICE_X3Y101_C3 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X3Y101_SLICE_X3Y101_C4 = CLBLM_R_X3Y101_SLICE_X3Y101_AO5;
  assign CLBLM_R_X3Y101_SLICE_X3Y101_C5 = CLBLM_R_X3Y101_SLICE_X3Y101_DO6;
  assign CLBLM_R_X3Y101_SLICE_X3Y101_C6 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_A1 = CLBLM_R_X3Y111_SLICE_X3Y111_DO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_A2 = CLBLM_R_X5Y113_SLICE_X7Y113_AO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_A3 = CLBLM_R_X7Y112_SLICE_X8Y112_AO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_A4 = CLBLM_R_X3Y111_SLICE_X2Y111_AO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_A5 = CLBLM_R_X5Y113_SLICE_X6Y113_AO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_A6 = CLBLM_R_X3Y108_SLICE_X2Y108_AO5;
  assign CLBLM_R_X3Y101_SLICE_X3Y101_D1 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X3Y101_SLICE_X3Y101_D2 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X3Y101_SLICE_X3Y101_D3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X3Y101_SLICE_X3Y101_D4 = CLBLL_L_X4Y101_SLICE_X4Y101_DO6;
  assign CLBLM_R_X3Y101_SLICE_X3Y101_D5 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X3Y101_SLICE_X3Y101_D6 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_B1 = CLBLM_R_X3Y111_SLICE_X3Y111_DO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_B2 = CLBLM_R_X5Y113_SLICE_X7Y113_AO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_B3 = CLBLM_R_X7Y112_SLICE_X8Y112_AO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_B4 = CLBLM_R_X5Y113_SLICE_X6Y113_AO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_B5 = CLBLM_R_X3Y111_SLICE_X2Y111_AO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_B6 = CLBLM_R_X3Y108_SLICE_X2Y108_AO5;
  assign CLBLM_R_X3Y101_SLICE_X2Y101_A1 = 1'b1;
  assign CLBLM_R_X3Y101_SLICE_X2Y101_A2 = 1'b1;
  assign CLBLM_R_X3Y101_SLICE_X2Y101_A3 = 1'b1;
  assign CLBLM_R_X3Y101_SLICE_X2Y101_A4 = 1'b1;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_C4 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_C5 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_C6 = CLBLM_R_X3Y111_SLICE_X2Y111_AO6;
  assign CLBLM_R_X3Y101_SLICE_X2Y101_A5 = 1'b1;
  assign CLBLM_R_X3Y101_SLICE_X2Y101_A6 = 1'b1;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_C1 = CLBLM_R_X5Y113_SLICE_X6Y113_AO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_C2 = CLBLM_R_X3Y111_SLICE_X3Y111_DO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_C3 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X3Y101_SLICE_X2Y101_B1 = 1'b1;
  assign CLBLM_R_X3Y101_SLICE_X2Y101_B2 = 1'b1;
  assign CLBLM_R_X3Y101_SLICE_X2Y101_B3 = 1'b1;
  assign CLBLM_R_X3Y101_SLICE_X2Y101_B4 = 1'b1;
  assign CLBLM_R_X3Y101_SLICE_X2Y101_B5 = 1'b1;
  assign CLBLM_R_X3Y101_SLICE_X2Y101_B6 = 1'b1;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_D1 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_D2 = CLBLM_R_X5Y110_SLICE_X6Y110_BO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_D3 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X3Y101_SLICE_X2Y101_C1 = 1'b1;
  assign CLBLM_R_X3Y101_SLICE_X2Y101_C2 = 1'b1;
  assign CLBLM_R_X3Y101_SLICE_X2Y101_C3 = 1'b1;
  assign CLBLM_R_X3Y101_SLICE_X2Y101_C4 = 1'b1;
  assign CLBLM_R_X3Y101_SLICE_X2Y101_C5 = 1'b1;
  assign CLBLM_R_X3Y101_SLICE_X2Y101_C6 = 1'b1;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_D5 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_D6 = CLBLM_R_X5Y111_SLICE_X6Y111_BO6;
  assign CLBLM_R_X3Y101_SLICE_X2Y101_D1 = 1'b1;
  assign CLBLM_R_X3Y101_SLICE_X2Y101_D2 = 1'b1;
  assign CLBLM_R_X3Y101_SLICE_X2Y101_D3 = 1'b1;
  assign CLBLM_R_X3Y101_SLICE_X2Y101_D4 = 1'b1;
  assign CLBLM_R_X3Y101_SLICE_X2Y101_D5 = 1'b1;
  assign CLBLM_R_X3Y101_SLICE_X2Y101_D6 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_A1 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_A2 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_A3 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_A4 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_A5 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_A6 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_B1 = CLBLM_R_X5Y112_SLICE_X7Y112_DO6;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_B2 = CLBLM_R_X5Y111_SLICE_X6Y111_DO6;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_B3 = CLBLM_R_X5Y110_SLICE_X6Y110_AO5;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_B4 = CLBLM_R_X7Y112_SLICE_X9Y112_DO6;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_B5 = CLBLM_R_X5Y112_SLICE_X7Y112_AO6;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_B6 = CLBLM_R_X5Y112_SLICE_X7Y112_AO5;
  assign CLBLM_R_X3Y102_SLICE_X3Y102_A1 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X3Y102_SLICE_X3Y102_A2 = CLBLM_R_X3Y102_SLICE_X2Y102_BO6;
  assign CLBLM_R_X3Y102_SLICE_X3Y102_A3 = CLBLM_R_X3Y101_SLICE_X3Y101_AO6;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_C4 = CLBLM_R_X5Y112_SLICE_X7Y112_AO5;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_C5 = CLBLM_R_X5Y112_SLICE_X7Y112_DO6;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_C6 = CLBLM_R_X7Y112_SLICE_X9Y112_DO6;
  assign CLBLM_R_X3Y102_SLICE_X3Y102_A4 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X3Y102_SLICE_X3Y102_A5 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X3Y102_SLICE_X3Y102_A6 = CLBLM_R_X3Y100_SLICE_X3Y100_AO5;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_C1 = CLBLM_R_X5Y112_SLICE_X7Y112_AO6;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_C2 = CLBLM_R_X5Y111_SLICE_X6Y111_DO6;
  assign CLBLM_R_X3Y102_SLICE_X3Y102_B1 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X3Y102_SLICE_X3Y102_B2 = CLBLM_R_X3Y102_SLICE_X2Y102_BO6;
  assign CLBLM_R_X3Y102_SLICE_X3Y102_B3 = CLBLM_R_X3Y101_SLICE_X3Y101_AO6;
  assign CLBLM_R_X3Y102_SLICE_X3Y102_B4 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X3Y102_SLICE_X3Y102_B5 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X3Y102_SLICE_X3Y102_B6 = CLBLM_R_X3Y100_SLICE_X3Y100_AO5;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_D5 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_D6 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_D1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_D2 = CLBLM_R_X5Y113_SLICE_X6Y113_CO6;
  assign CLBLM_R_X3Y102_SLICE_X3Y102_C1 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X3Y102_SLICE_X3Y102_C2 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X3Y102_SLICE_X3Y102_C3 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X3Y102_SLICE_X3Y102_C4 = CLBLM_R_X3Y100_SLICE_X3Y100_AO5;
  assign CLBLM_R_X3Y102_SLICE_X3Y102_C5 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X3Y102_SLICE_X3Y102_C6 = CLBLM_R_X3Y101_SLICE_X3Y101_BO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_A1 = CLBLM_R_X5Y113_SLICE_X6Y113_DO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_A2 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_A3 = CLBLM_R_X5Y113_SLICE_X6Y113_AO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_A4 = CLBLM_R_X5Y110_SLICE_X7Y110_AO5;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_A5 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_A6 = 1'b1;
  assign CLBLM_R_X3Y102_SLICE_X3Y102_D1 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X3Y102_SLICE_X3Y102_D2 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X3Y102_SLICE_X3Y102_D3 = CLBLL_L_X4Y102_SLICE_X5Y102_DO6;
  assign CLBLM_R_X3Y102_SLICE_X3Y102_D4 = CLBLM_R_X3Y102_SLICE_X3Y102_CO6;
  assign CLBLM_R_X3Y102_SLICE_X3Y102_D5 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X3Y102_SLICE_X3Y102_D6 = CLBLM_R_X3Y102_SLICE_X3Y102_BO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_B6 = CLBLM_R_X5Y113_SLICE_X6Y113_CO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_B1 = CLBLL_L_X4Y112_SLICE_X4Y112_AO5;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_B2 = CLBLM_R_X7Y113_SLICE_X9Y113_BO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_B3 = CLBLM_R_X7Y112_SLICE_X9Y112_AO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_B4 = CLBLM_R_X5Y113_SLICE_X6Y113_BO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_B5 = CLBLM_R_X5Y111_SLICE_X6Y111_BO6;
  assign CLBLM_R_X3Y102_SLICE_X2Y102_A1 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_C4 = CLBLM_R_X5Y112_SLICE_X6Y112_AO5;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_C5 = CLBLM_R_X7Y113_SLICE_X9Y113_CO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_C6 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X3Y102_SLICE_X2Y102_A2 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X3Y102_SLICE_X2Y102_A3 = CLBLM_R_X3Y102_SLICE_X3Y102_AO6;
  assign CLBLM_R_X3Y102_SLICE_X2Y102_A4 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X3Y102_SLICE_X2Y102_A5 = CLBLL_L_X2Y102_SLICE_X1Y102_BO6;
  assign CLBLM_R_X3Y102_SLICE_X2Y102_A6 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X3Y102_SLICE_X2Y102_B1 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X3Y102_SLICE_X2Y102_B2 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X3Y102_SLICE_X2Y102_B3 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X3Y102_SLICE_X2Y102_B4 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X3Y102_SLICE_X2Y102_B5 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X3Y102_SLICE_X2Y102_B6 = CLBLL_L_X2Y102_SLICE_X1Y102_AO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_D1 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_D2 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_D3 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X3Y102_SLICE_X2Y102_C1 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X3Y102_SLICE_X2Y102_C2 = CLBLM_R_X3Y102_SLICE_X3Y102_AO6;
  assign CLBLM_R_X3Y102_SLICE_X2Y102_C3 = CLBLL_L_X2Y102_SLICE_X1Y102_BO6;
  assign CLBLM_R_X3Y102_SLICE_X2Y102_C4 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X3Y102_SLICE_X2Y102_C5 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X3Y102_SLICE_X2Y102_C6 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_D5 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_D6 = CLBLM_R_X5Y111_SLICE_X6Y111_DO6;
  assign CLBLM_R_X3Y102_SLICE_X2Y102_D1 = 1'b1;
  assign CLBLM_R_X3Y102_SLICE_X2Y102_D2 = 1'b1;
  assign CLBLM_R_X3Y102_SLICE_X2Y102_D3 = 1'b1;
  assign CLBLM_R_X3Y102_SLICE_X2Y102_D4 = 1'b1;
  assign CLBLM_R_X3Y102_SLICE_X2Y102_D5 = 1'b1;
  assign CLBLM_R_X3Y102_SLICE_X2Y102_D6 = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_D1 = CLBLM_R_X3Y107_SLICE_X2Y107_AO6;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_T1 = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_D1 = CLBLM_R_X3Y107_SLICE_X2Y107_AO5;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_T1 = 1'b1;
  assign LIOI3_X0Y115_ILOGIC_X0Y116_D = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_A1 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_A2 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_A3 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_A4 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_A5 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_A6 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_B1 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_B2 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_B3 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_B4 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_B5 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_B6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_D1 = CLBLL_L_X2Y114_SLICE_X0Y114_AO6;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_A1 = CLBLM_R_X3Y102_SLICE_X3Y102_DO6;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_A2 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_A3 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_A4 = CLBLM_R_X3Y102_SLICE_X2Y102_CO6;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_A5 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_A6 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_C1 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_C2 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_C3 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_B1 = CLBLL_L_X4Y103_SLICE_X5Y103_DO6;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_B2 = CLBLL_L_X4Y102_SLICE_X4Y102_CO6;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_B3 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_B4 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_B5 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_B6 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_D1 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_D2 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_C1 = CLBLM_R_X3Y102_SLICE_X2Y102_CO6;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_C2 = CLBLM_R_X3Y102_SLICE_X3Y102_DO6;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_C3 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_C4 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_C5 = CLBLM_R_X3Y103_SLICE_X2Y103_AO6;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_C6 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_D3 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_D4 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_A1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_A2 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_A3 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_A4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_A5 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_A6 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_D1 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_D2 = CLBLM_R_X3Y102_SLICE_X2Y102_CO6;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_D3 = CLBLM_R_X3Y102_SLICE_X3Y102_DO6;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_D4 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_D5 = CLBLM_R_X3Y103_SLICE_X2Y103_AO6;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_D6 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_B1 = CLBLM_R_X5Y113_SLICE_X6Y113_DO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_B2 = CLBLM_R_X5Y110_SLICE_X7Y110_AO5;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_B3 = CLBLM_R_X5Y113_SLICE_X7Y113_AO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_B4 = CLBLM_R_X5Y113_SLICE_X7Y113_AO5;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_B5 = CLBLM_R_X7Y113_SLICE_X9Y113_AO6;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_A1 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_A2 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_A3 = CLBLM_R_X3Y102_SLICE_X2Y102_AO6;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_A4 = CLBLL_L_X2Y103_SLICE_X1Y103_CO6;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_A5 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_A6 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_C1 = CLBLM_R_X7Y113_SLICE_X9Y113_AO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_C2 = CLBLM_R_X5Y113_SLICE_X7Y113_AO5;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_C3 = CLBLM_R_X5Y113_SLICE_X7Y113_AO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_C4 = CLBLM_R_X5Y111_SLICE_X7Y111_BO6;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_B1 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_B2 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_B3 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_B4 = CLBLL_L_X4Y102_SLICE_X4Y102_CO6;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_B5 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_B6 = CLBLL_L_X4Y103_SLICE_X5Y103_DO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_D1 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_D2 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_D3 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_C1 = CLBLL_L_X2Y103_SLICE_X1Y103_AO5;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_C2 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_C3 = CLBLL_L_X4Y102_SLICE_X4Y102_BO6;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_C4 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_C5 = CLBLM_R_X5Y103_SLICE_X6Y103_DO6;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_C6 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_D4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_D5 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_D6 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_D1 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_D2 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_D3 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_D4 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_D5 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_D6 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_B3 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_C1 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_C2 = 1'b1;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_A1 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_A2 = CLBLL_L_X4Y103_SLICE_X4Y103_CO6;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_A3 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_A4 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_A5 = CLBLM_R_X3Y103_SLICE_X3Y103_AO5;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_A6 = 1'b1;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_B1 = CLBLL_L_X4Y104_SLICE_X4Y104_CO6;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_B2 = CLBLM_R_X3Y103_SLICE_X3Y103_DO6;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_B3 = CLBLM_R_X3Y104_SLICE_X2Y104_AO6;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_B4 = CLBLL_L_X2Y104_SLICE_X0Y104_CO6;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_B5 = CLBLM_R_X3Y103_SLICE_X3Y103_CO6;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_B6 = CLBLM_R_X3Y104_SLICE_X3Y104_AO5;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_D1 = 1'b1;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_C1 = CLBLM_R_X3Y103_SLICE_X3Y103_CO6;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_C2 = CLBLM_R_X3Y103_SLICE_X3Y103_DO6;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_C3 = CLBLL_L_X4Y104_SLICE_X4Y104_CO6;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_C4 = CLBLM_R_X3Y104_SLICE_X3Y104_AO5;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_C5 = CLBLM_R_X3Y104_SLICE_X2Y104_AO6;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_C6 = CLBLL_L_X2Y104_SLICE_X0Y104_CO6;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_D1 = CLBLM_R_X3Y103_SLICE_X3Y103_CO6;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_D2 = 1'b1;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_D3 = 1'b1;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_D4 = CLBLM_R_X3Y104_SLICE_X3Y104_AO5;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_D5 = CLBLL_L_X4Y104_SLICE_X4Y104_CO6;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_D6 = CLBLL_L_X2Y104_SLICE_X0Y104_CO6;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_A1 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_A2 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_A3 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_A4 = CLBLM_R_X3Y104_SLICE_X2Y104_BO6;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_A5 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_A6 = CLBLM_R_X3Y103_SLICE_X2Y103_AO5;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_B1 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_B2 = CLBLL_L_X2Y103_SLICE_X1Y103_DO6;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_B3 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_B4 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_B5 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_B6 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_C1 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_C2 = CLBLM_R_X3Y103_SLICE_X2Y103_AO5;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_C3 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_C4 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_C5 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_C6 = CLBLM_R_X3Y104_SLICE_X2Y104_BO6;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_D1 = 1'b1;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_D2 = 1'b1;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_D3 = 1'b1;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_D4 = 1'b1;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_D5 = 1'b1;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_D6 = 1'b1;
  assign LIOB33_SING_X0Y149_IOB_X0Y149_O = CLBLL_L_X2Y108_SLICE_X0Y108_CO6;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_D1 = CLBLL_L_X2Y105_SLICE_X1Y105_DO6;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_T1 = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_D1 = CLBLL_L_X2Y107_SLICE_X1Y107_CO6;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_T1 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_A1 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_A2 = CLBLM_R_X5Y105_SLICE_X6Y105_BO6;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_A3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_A4 = CLBLL_L_X4Y105_SLICE_X5Y105_AO6;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_A5 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_A6 = CLBLL_L_X4Y106_SLICE_X4Y106_CO6;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_B1 = CLBLL_L_X4Y106_SLICE_X4Y106_CO6;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_B2 = CLBLL_L_X4Y105_SLICE_X5Y105_AO6;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_B3 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_B4 = CLBLM_R_X5Y105_SLICE_X6Y105_DO6;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_B5 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_B6 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_C1 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_C2 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_C3 = CLBLM_R_X5Y105_SLICE_X6Y105_DO6;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_C4 = CLBLL_L_X4Y106_SLICE_X4Y106_CO6;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_C5 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_C6 = CLBLL_L_X4Y105_SLICE_X5Y105_AO6;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_D1 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_D2 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_D3 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_D4 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_D5 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_D6 = 1'b1;
  assign LIOB33_X0Y117_IOB_X0Y118_O = CLBLL_L_X2Y114_SLICE_X0Y114_AO5;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_A1 = CLBLL_L_X4Y105_SLICE_X4Y105_CO6;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_A2 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_A3 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_A4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_A5 = CLBLL_L_X4Y104_SLICE_X4Y104_AO6;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_A6 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_B1 = CLBLL_L_X4Y105_SLICE_X4Y105_CO6;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_B2 = CLBLM_R_X3Y103_SLICE_X2Y103_BO6;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_B3 = CLBLL_L_X4Y104_SLICE_X4Y104_AO5;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_B4 = CLBLM_R_X3Y106_SLICE_X2Y106_AO6;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_B5 = CLBLL_L_X4Y104_SLICE_X4Y104_AO6;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_B6 = CLBLL_L_X2Y106_SLICE_X1Y106_AO6;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_C1 = CLBLL_L_X4Y104_SLICE_X4Y104_AO6;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_C2 = CLBLM_R_X3Y103_SLICE_X2Y103_BO6;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_C3 = CLBLL_L_X4Y105_SLICE_X4Y105_CO6;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_C4 = CLBLM_R_X3Y106_SLICE_X2Y106_AO6;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_C5 = CLBLL_L_X4Y104_SLICE_X4Y104_AO5;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_C6 = CLBLL_L_X2Y106_SLICE_X1Y106_AO6;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_D1 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_D2 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_D3 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_D4 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_D5 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_D6 = 1'b1;
  assign CLBLM_L_X8Y100_SLICE_X10Y100_C3 = CLBLM_L_X8Y100_SLICE_X11Y100_DO6;
  assign CLBLM_L_X8Y100_SLICE_X10Y100_C6 = CLBLM_R_X3Y100_SLICE_X3Y100_AO6;
  assign CLBLM_L_X8Y100_SLICE_X10Y100_D1 = CLBLL_L_X4Y103_SLICE_X5Y103_BO6;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_D = RIOB33_X105Y107_IOB_X1Y108_I;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_D = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_A1 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_A2 = CLBLL_L_X2Y103_SLICE_X1Y103_BO6;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_A3 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_A4 = CLBLM_R_X3Y103_SLICE_X2Y103_CO6;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_A5 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_A6 = 1'b1;
  assign LIOB33_X0Y119_IOB_X0Y119_O = CLBLL_L_X2Y114_SLICE_X0Y114_AO6;
  assign LIOB33_X0Y119_IOB_X0Y120_O = CLBLL_L_X2Y113_SLICE_X0Y113_AO5;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_B1 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_B2 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_B3 = CLBLM_R_X3Y103_SLICE_X3Y103_BO6;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_B4 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_B5 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_B6 = CLBLM_R_X3Y106_SLICE_X3Y106_AO5;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_C1 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_C2 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_C3 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_C4 = CLBLM_R_X3Y106_SLICE_X3Y106_AO5;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_C5 = CLBLM_R_X3Y103_SLICE_X3Y103_BO6;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_C6 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_D1 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_D2 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_D3 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_D4 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_D5 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_D6 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_A1 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_A2 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_A3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_A4 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_A5 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_A6 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_B1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_B2 = CLBLL_L_X4Y105_SLICE_X4Y105_BO6;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_B3 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_B4 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_B5 = CLBLM_R_X3Y105_SLICE_X3Y105_BO6;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_B6 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_C1 = CLBLM_R_X3Y105_SLICE_X3Y105_BO6;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_C2 = CLBLL_L_X4Y105_SLICE_X4Y105_BO6;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_C3 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_C4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_C5 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_C6 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_D1 = CLBLM_R_X3Y105_SLICE_X2Y105_AO6;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_D2 = CLBLM_R_X3Y107_SLICE_X3Y107_BO6;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_D3 = CLBLM_R_X3Y107_SLICE_X2Y107_DO6;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_D4 = CLBLM_R_X3Y106_SLICE_X2Y106_CO6;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_D5 = CLBLL_L_X2Y107_SLICE_X1Y107_BO6;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_D6 = CLBLM_R_X3Y105_SLICE_X2Y105_BO6;
  assign LIOB33_X0Y121_IOB_X0Y122_O = CLBLL_L_X2Y113_SLICE_X1Y113_AO6;
  assign LIOB33_X0Y121_IOB_X0Y121_O = CLBLL_L_X2Y113_SLICE_X0Y113_BO5;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_A1 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_A2 = 1'b1;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_A3 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_A4 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_A5 = 1'b1;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_A6 = 1'b1;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_B1 = CLBLM_R_X3Y106_SLICE_X2Y106_AO5;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_B2 = CLBLL_L_X4Y105_SLICE_X4Y105_DO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_B3 = CLBLL_L_X4Y107_SLICE_X4Y107_CO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_B4 = CLBLM_R_X3Y105_SLICE_X3Y105_CO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_B5 = CLBLM_R_X3Y105_SLICE_X3Y105_BO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_B6 = CLBLM_R_X3Y107_SLICE_X3Y107_AO5;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_D1 = CLBLL_L_X2Y105_SLICE_X0Y105_AO5;
  assign LIOI3_X0Y103_ILOGIC_X0Y104_D = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_C1 = CLBLM_R_X3Y105_SLICE_X3Y105_BO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_C2 = CLBLL_L_X4Y105_SLICE_X4Y105_DO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_C3 = CLBLL_L_X4Y107_SLICE_X4Y107_CO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_C4 = CLBLM_R_X3Y107_SLICE_X3Y107_AO5;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_C5 = CLBLM_R_X3Y106_SLICE_X2Y106_AO5;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_C6 = CLBLM_R_X3Y105_SLICE_X3Y105_CO6;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_T1 = 1'b1;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_D1 = 1'b1;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_D2 = 1'b1;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_D3 = 1'b1;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_D4 = 1'b1;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_D5 = 1'b1;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_D6 = 1'b1;
  assign LIOI3_X0Y103_ILOGIC_X0Y103_D = LIOB33_X0Y103_IOB_X0Y103_I;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_D1 = CLBLL_L_X2Y105_SLICE_X0Y105_AO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_A1 = CLBLM_R_X3Y108_SLICE_X3Y108_BO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_A2 = CLBLM_R_X3Y108_SLICE_X2Y108_BO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_A3 = CLBLM_R_X3Y108_SLICE_X2Y108_CO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_A4 = CLBLM_R_X3Y107_SLICE_X2Y107_BO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_A5 = CLBLM_R_X3Y107_SLICE_X2Y107_CO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_A6 = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_T1 = 1'b1;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_B1 = CLBLL_L_X4Y108_SLICE_X4Y108_DO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_B2 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_B3 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_B4 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_B5 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_B6 = CLBLM_R_X3Y108_SLICE_X3Y108_CO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_C1 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_C2 = CLBLM_R_X3Y108_SLICE_X3Y108_CO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_C3 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_C4 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_C5 = CLBLL_L_X4Y108_SLICE_X4Y108_DO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_C6 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_D1 = CLBLM_R_X3Y108_SLICE_X2Y108_BO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_D2 = CLBLM_R_X3Y107_SLICE_X3Y107_CO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_D3 = CLBLM_R_X3Y108_SLICE_X3Y108_BO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_D4 = CLBLM_R_X3Y107_SLICE_X2Y107_CO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_D5 = CLBLM_R_X3Y108_SLICE_X2Y108_CO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_D6 = CLBLM_R_X3Y107_SLICE_X2Y107_BO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_C5 = 1'b1;
  assign LIOB33_X0Y123_IOB_X0Y124_O = CLBLM_R_X3Y112_SLICE_X2Y112_AO6;
  assign LIOB33_X0Y123_IOB_X0Y123_O = CLBLL_L_X2Y113_SLICE_X1Y113_CO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_A1 = CLBLL_L_X4Y108_SLICE_X5Y108_CO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_A2 = CLBLL_L_X4Y108_SLICE_X4Y108_CO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_A3 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_A4 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_A5 = CLBLM_R_X5Y108_SLICE_X7Y108_DO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_A6 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_B1 = CLBLM_R_X3Y110_SLICE_X2Y110_DO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_B2 = CLBLL_L_X2Y108_SLICE_X0Y108_AO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_B3 = CLBLM_R_X3Y104_SLICE_X3Y104_AO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_B4 = CLBLL_L_X4Y109_SLICE_X5Y109_DO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_B5 = CLBLM_R_X3Y108_SLICE_X3Y108_AO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_B6 = CLBLL_L_X4Y108_SLICE_X5Y108_DO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_C1 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_C2 = CLBLL_L_X4Y108_SLICE_X4Y108_CO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_C3 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_C4 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_C5 = CLBLL_L_X4Y108_SLICE_X5Y108_CO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_C6 = CLBLM_R_X5Y108_SLICE_X7Y108_DO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_D1 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_D2 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_D3 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_D4 = CLBLM_R_X5Y108_SLICE_X6Y108_CO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_D5 = CLBLL_L_X4Y108_SLICE_X5Y108_CO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_D6 = CLBLL_L_X4Y108_SLICE_X4Y108_CO6;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_A1 = CLBLL_L_X4Y108_SLICE_X4Y108_DO6;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_A2 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_A3 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_A4 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_A5 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_A6 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_B1 = CLBLL_L_X4Y109_SLICE_X5Y109_DO6;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_B2 = CLBLM_R_X3Y108_SLICE_X3Y108_DO6;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_B3 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_B4 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_B5 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_B6 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_C1 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_C2 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_C3 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_C4 = CLBLL_L_X4Y107_SLICE_X4Y107_CO6;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_C5 = CLBLM_R_X3Y105_SLICE_X3Y105_AO6;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_C6 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_D1 = CLBLM_R_X3Y108_SLICE_X2Y108_AO6;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_D2 = CLBLM_R_X3Y108_SLICE_X3Y108_CO6;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_D3 = CLBLM_R_X3Y108_SLICE_X3Y108_BO6;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_D4 = CLBLM_R_X3Y108_SLICE_X2Y108_CO6;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_D5 = CLBLM_R_X3Y107_SLICE_X3Y107_AO6;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_D6 = CLBLM_R_X3Y108_SLICE_X2Y108_BO6;
  assign LIOB33_X0Y125_IOB_X0Y126_O = CLBLM_R_X3Y111_SLICE_X2Y111_BO6;
  assign LIOB33_X0Y125_IOB_X0Y125_O = CLBLM_R_X3Y111_SLICE_X3Y111_AO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_B4 = CLBLM_L_X8Y107_SLICE_X11Y107_CO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_B5 = CLBLM_R_X7Y106_SLICE_X9Y106_AO5;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_B6 = CLBLM_R_X7Y107_SLICE_X9Y107_AO5;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_C3 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_C4 = CLBLM_L_X8Y108_SLICE_X10Y108_CO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_A1 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_A2 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_A3 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_A4 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_A5 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_A6 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_B1 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_B2 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_B3 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_B4 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_B5 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_B6 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_C1 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_C2 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_C3 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_C4 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_C5 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_C6 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_D1 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_D2 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_D3 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_D4 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_D5 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_D6 = 1'b1;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_D5 = CLBLM_L_X8Y107_SLICE_X11Y107_CO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_A1 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_A2 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_A3 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_A4 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_A5 = CLBLM_R_X3Y105_SLICE_X3Y105_AO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_A6 = CLBLL_L_X4Y107_SLICE_X4Y107_CO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_D6 = CLBLM_R_X7Y106_SLICE_X9Y106_AO5;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_B1 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_B2 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_B3 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_B4 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_B5 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_B6 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_C1 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_C2 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_C3 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_C4 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_C5 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_C6 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_D1 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_D2 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_D3 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_D4 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_D5 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_D6 = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_D1 = CLBLM_R_X3Y104_SLICE_X3Y104_BO6;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_T1 = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_D1 = CLBLM_R_X3Y104_SLICE_X3Y104_DO6;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_T1 = 1'b1;
  assign LIOB33_X0Y127_IOB_X0Y128_O = CLBLL_L_X4Y107_SLICE_X4Y107_AO6;
  assign LIOB33_X0Y127_IOB_X0Y127_O = CLBLL_L_X4Y110_SLICE_X4Y110_AO5;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_A1 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_A2 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_A3 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_A4 = CLBLM_R_X3Y111_SLICE_X2Y111_CO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_A5 = CLBLL_L_X4Y111_SLICE_X4Y111_AO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_A6 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_B1 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_B2 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_B3 = CLBLL_L_X4Y109_SLICE_X4Y109_AO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_B4 = CLBLL_L_X4Y110_SLICE_X4Y110_CO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_B5 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_B6 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_C1 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_C2 = CLBLL_L_X4Y109_SLICE_X4Y109_AO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_C3 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_C4 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_C5 = CLBLL_L_X4Y110_SLICE_X4Y110_CO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_C6 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_D1 = CLBLL_L_X4Y111_SLICE_X4Y111_AO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_D2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_D3 = CLBLM_R_X3Y111_SLICE_X2Y111_CO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_D4 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_D5 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_D6 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_A1 = CLBLM_R_X3Y110_SLICE_X3Y110_CO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_A2 = CLBLL_L_X4Y109_SLICE_X4Y109_BO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_A3 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_A4 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_A5 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_A6 = 1'b1;
  assign CLBLM_L_X8Y101_SLICE_X10Y101_B3 = CLBLM_L_X8Y101_SLICE_X11Y101_AO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_B1 = CLBLM_R_X3Y110_SLICE_X3Y110_CO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_B2 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_B3 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_L_X8Y101_SLICE_X10Y101_B4 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_B4 = CLBLL_L_X4Y107_SLICE_X4Y107_BO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_B5 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_B6 = CLBLL_L_X4Y109_SLICE_X4Y109_BO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_C1 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_C2 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_C3 = CLBLL_L_X4Y109_SLICE_X4Y109_DO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_C4 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_C5 = CLBLM_R_X3Y110_SLICE_X2Y110_DO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_C6 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_D1 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_D2 = CLBLM_R_X3Y110_SLICE_X3Y110_CO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_D3 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_D4 = CLBLL_L_X4Y109_SLICE_X4Y109_BO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_D5 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_D6 = CLBLL_L_X4Y107_SLICE_X4Y107_BO6;
  assign LIOB33_X0Y129_IOB_X0Y130_O = CLBLL_L_X2Y114_SLICE_X0Y114_BO5;
  assign LIOB33_X0Y129_IOB_X0Y129_O = CLBLM_R_X3Y110_SLICE_X3Y110_BO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_A1 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_A2 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_A3 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_A4 = CLBLM_R_X3Y112_SLICE_X3Y112_CO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_A5 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_A6 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_B1 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_B2 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_B3 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_B4 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_B5 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_B6 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_C1 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_C2 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_C3 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_C4 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_C5 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_C6 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_D1 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_D2 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_D3 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_D4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_D5 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_D6 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_A1 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_A2 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_A3 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_A4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_A5 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_A6 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_B1 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_B2 = CLBLL_L_X4Y111_SLICE_X4Y111_AO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_B3 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_B4 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_B5 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_B6 = CLBLM_R_X3Y111_SLICE_X2Y111_CO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_C1 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_C2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_C3 = CLBLM_R_X3Y112_SLICE_X2Y112_DO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_C4 = CLBLL_L_X4Y112_SLICE_X4Y112_BO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_C5 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_C6 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_D1 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_D2 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_D3 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_D4 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_D5 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_D6 = 1'b1;
  assign LIOB33_X0Y131_IOB_X0Y132_O = CLBLM_R_X3Y110_SLICE_X2Y110_BO6;
  assign LIOB33_X0Y131_IOB_X0Y131_O = CLBLM_R_X3Y110_SLICE_X2Y110_AO5;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_D1 = CLBLL_L_X2Y108_SLICE_X0Y108_BO6;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_T1 = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_D1 = CLBLL_L_X2Y108_SLICE_X0Y108_DO6;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_T1 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_A1 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_A2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_A3 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_A4 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_A5 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_A6 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_B1 = CLBLM_R_X3Y113_SLICE_X3Y113_DO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_B2 = CLBLM_R_X3Y113_SLICE_X3Y113_BO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_B3 = CLBLL_L_X4Y112_SLICE_X4Y112_AO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_B4 = CLBLL_L_X2Y113_SLICE_X1Y113_AO5;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_B5 = CLBLM_R_X5Y111_SLICE_X6Y111_AO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_B6 = CLBLM_R_X3Y113_SLICE_X3Y113_CO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_C1 = CLBLL_L_X4Y112_SLICE_X4Y112_BO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_C2 = CLBLL_L_X4Y112_SLICE_X4Y112_CO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_C3 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_C4 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_C5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_C6 = CLBLL_L_X2Y112_SLICE_X1Y112_AO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_D1 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_D2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_D3 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_D4 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_D5 = CLBLM_R_X3Y113_SLICE_X2Y113_DO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_C1 = CLBLL_L_X4Y106_SLICE_X4Y106_BO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_D6 = CLBLM_R_X3Y113_SLICE_X3Y113_BO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_C2 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_A1 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_A2 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_A3 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_A4 = CLBLM_R_X3Y112_SLICE_X2Y112_BO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_A5 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_A6 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_B1 = CLBLL_L_X2Y113_SLICE_X1Y113_DO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_B2 = CLBLM_R_X3Y112_SLICE_X3Y112_BO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_B3 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_B4 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_B5 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_B6 = CLBLM_R_X3Y112_SLICE_X2Y112_CO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_C1 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_C2 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_C3 = CLBLM_R_X3Y113_SLICE_X2Y113_DO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_C4 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_C5 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_C6 = CLBLM_R_X3Y113_SLICE_X3Y113_BO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_D1 = CLBLM_R_X3Y112_SLICE_X2Y112_CO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_D2 = CLBLM_R_X5Y101_SLICE_X7Y101_AO5;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_D3 = CLBLM_R_X3Y112_SLICE_X3Y112_BO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_D4 = CLBLM_R_X3Y112_SLICE_X2Y112_AO5;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_D5 = CLBLL_L_X2Y113_SLICE_X1Y113_DO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_D6 = CLBLM_R_X3Y111_SLICE_X3Y111_BO6;
  assign LIOB33_X0Y133_IOB_X0Y134_O = 1'b0;
  assign LIOB33_X0Y133_IOB_X0Y133_O = CLBLM_R_X3Y110_SLICE_X2Y110_CO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_A1 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_A2 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_A3 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_A4 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_A5 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_A6 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_B1 = CLBLM_R_X3Y114_SLICE_X2Y114_DO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_B2 = CLBLM_R_X3Y113_SLICE_X3Y113_AO5;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_B3 = CLBLM_R_X3Y114_SLICE_X2Y114_AO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_B4 = CLBLM_R_X3Y114_SLICE_X2Y114_CO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_B5 = CLBLM_R_X3Y113_SLICE_X3Y113_AO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_B6 = CLBLM_R_X3Y112_SLICE_X3Y112_AO5;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_A4 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_C1 = CLBLM_R_X3Y113_SLICE_X3Y113_AO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_C2 = CLBLL_L_X4Y113_SLICE_X4Y113_AO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_C3 = CLBLM_R_X3Y112_SLICE_X3Y112_AO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_C4 = CLBLM_R_X3Y108_SLICE_X2Y108_AO5;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_C5 = CLBLM_R_X3Y111_SLICE_X2Y111_AO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_C6 = CLBLM_R_X3Y114_SLICE_X2Y114_CO6;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_A5 = 1'b1;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_A6 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_D1 = CLBLM_R_X3Y113_SLICE_X3Y113_AO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_D2 = CLBLL_L_X4Y113_SLICE_X4Y113_AO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_D3 = CLBLM_R_X3Y112_SLICE_X3Y112_AO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_D4 = CLBLM_R_X3Y108_SLICE_X2Y108_AO5;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_D5 = CLBLM_R_X3Y111_SLICE_X2Y111_AO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_D6 = CLBLM_R_X3Y114_SLICE_X2Y114_CO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_A1 = CLBLM_R_X3Y114_SLICE_X2Y114_DO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_A2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_A3 = CLBLM_R_X3Y114_SLICE_X2Y114_AO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_A4 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_A5 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_A6 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_B1 = CLBLM_R_X3Y114_SLICE_X2Y114_CO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_B2 = CLBLL_L_X4Y113_SLICE_X4Y113_AO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_B3 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_B4 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_B5 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_B6 = 1'b1;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_B3 = 1'b1;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_B4 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_C1 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_C2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_C3 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_C4 = CLBLM_R_X3Y113_SLICE_X2Y113_AO5;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_C5 = CLBLM_R_X3Y113_SLICE_X2Y113_DO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_C6 = CLBLM_R_X3Y113_SLICE_X2Y113_BO6;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_B5 = 1'b1;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_B6 = 1'b1;
  assign LIOB33_X0Y135_IOB_X0Y135_O = CLBLM_R_X3Y107_SLICE_X2Y107_AO5;
  assign LIOB33_X0Y135_IOB_X0Y136_O = CLBLM_R_X3Y107_SLICE_X2Y107_AO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_D1 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_D2 = CLBLM_R_X3Y111_SLICE_X2Y111_AO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_D3 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_D4 = CLBLL_L_X4Y113_SLICE_X4Y113_AO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_D5 = CLBLM_R_X3Y114_SLICE_X2Y114_CO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_D6 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_A1 = CLBLM_R_X7Y111_SLICE_X8Y111_DO6;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_D1 = 1'b1;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_D2 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_A3 = CLBLM_R_X5Y111_SLICE_X7Y111_AO5;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_B1 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_C1 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_C2 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_C3 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_D2 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_D3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_C6 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_D4 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_D5 = CLBLM_R_X7Y113_SLICE_X9Y113_DO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_A1 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_A2 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_A3 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_A4 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_A5 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_A6 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_B1 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_B2 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_B3 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_B4 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_B5 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_B6 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_C1 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_C2 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_C3 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_C4 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_C5 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_C6 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_D1 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_D2 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_D3 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_D4 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_D5 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_D6 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_D2 = 1'b1;
  assign LIOB33_X0Y137_IOB_X0Y137_O = CLBLL_L_X2Y109_SLICE_X1Y109_AO6;
  assign LIOB33_X0Y137_IOB_X0Y138_O = CLBLL_L_X2Y108_SLICE_X1Y108_DO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_A1 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_A2 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_A3 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_A4 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_A5 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_A6 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_B1 = CLBLM_R_X3Y114_SLICE_X2Y114_DO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_B2 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_B3 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_B4 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_B5 = CLBLM_R_X3Y114_SLICE_X2Y114_AO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_B6 = CLBLM_R_X3Y114_SLICE_X2Y114_CO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_C1 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_C2 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_C3 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_C4 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_C5 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_C6 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_D1 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_D2 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_D3 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_D4 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_D5 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_D6 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_C4 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_C5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_C6 = CLBLM_R_X7Y111_SLICE_X8Y111_CO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_D5 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_D6 = CLBLM_R_X5Y112_SLICE_X6Y112_DO6;
  assign LIOB33_X0Y139_IOB_X0Y140_O = CLBLL_L_X2Y105_SLICE_X1Y105_DO6;
  assign LIOB33_X0Y139_IOB_X0Y139_O = CLBLL_L_X2Y107_SLICE_X1Y107_CO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_B6 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_B3 = CLBLM_L_X8Y102_SLICE_X11Y102_CO6;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_B4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_C4 = CLBLM_R_X5Y110_SLICE_X6Y110_AO5;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_C5 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_C6 = CLBLM_R_X5Y112_SLICE_X6Y112_DO6;
  assign CLBLM_R_X5Y100_SLICE_X7Y100_A5 = 1'b1;
  assign CLBLM_R_X5Y100_SLICE_X7Y100_A6 = 1'b1;
  assign LIOB33_X0Y141_IOB_X0Y142_O = CLBLL_L_X2Y105_SLICE_X0Y105_AO5;
  assign LIOB33_X0Y141_IOB_X0Y141_O = CLBLL_L_X2Y105_SLICE_X0Y105_AO6;
  assign CLBLM_R_X5Y100_SLICE_X7Y100_B1 = 1'b1;
  assign CLBLM_R_X5Y100_SLICE_X7Y100_B2 = 1'b1;
  assign CLBLM_R_X5Y100_SLICE_X7Y100_B3 = 1'b1;
  assign CLBLM_R_X5Y100_SLICE_X7Y100_B5 = 1'b1;
  assign LIOI3_SING_X0Y100_ILOGIC_X0Y100_D = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign LIOB33_X0Y143_IOB_X0Y143_O = CLBLL_L_X2Y106_SLICE_X0Y106_BO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_C4 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_C5 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_C6 = CLBLL_L_X4Y108_SLICE_X4Y108_BO6;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_D1 = CLBLL_L_X2Y108_SLICE_X0Y108_CO6;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_T1 = 1'b1;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_A1 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_A2 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_A3 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_A4 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_A5 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_A6 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_B1 = 1'b1;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_B2 = 1'b1;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_B3 = 1'b1;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_B4 = 1'b1;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_B5 = 1'b1;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_B6 = 1'b1;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_C1 = 1'b1;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_C2 = 1'b1;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_C3 = 1'b1;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_C4 = 1'b1;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_C5 = 1'b1;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_C6 = 1'b1;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_D1 = 1'b1;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_D2 = 1'b1;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_D3 = 1'b1;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_D4 = 1'b1;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_D5 = 1'b1;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_D6 = 1'b1;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_A1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_A2 = 1'b1;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_A3 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_A4 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_A5 = 1'b1;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_A6 = 1'b1;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_B1 = CLBLM_L_X8Y102_SLICE_X10Y102_DO6;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_B2 = CLBLM_L_X8Y101_SLICE_X10Y101_AO6;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_B3 = CLBLM_L_X10Y102_SLICE_X13Y102_AO6;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_B4 = CLBLM_R_X5Y102_SLICE_X6Y102_BO6;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_B5 = CLBLM_L_X10Y102_SLICE_X12Y102_AO6;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_B6 = CLBLL_L_X4Y101_SLICE_X5Y101_AO6;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_C1 = CLBLM_L_X10Y103_SLICE_X13Y103_CO6;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_C2 = CLBLM_L_X10Y103_SLICE_X12Y103_AO5;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_C3 = CLBLM_L_X8Y100_SLICE_X10Y100_DO6;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_C4 = CLBLM_L_X10Y102_SLICE_X12Y102_AO5;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_C5 = CLBLM_L_X10Y102_SLICE_X12Y102_DO6;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_C6 = CLBLM_L_X10Y102_SLICE_X12Y102_BO6;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_D1 = CLBLM_L_X10Y102_SLICE_X12Y102_AO6;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_D2 = CLBLM_L_X10Y102_SLICE_X13Y102_AO6;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_D3 = CLBLM_L_X8Y101_SLICE_X10Y101_AO6;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_D4 = CLBLM_R_X5Y102_SLICE_X6Y102_BO6;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_D5 = CLBLM_L_X8Y102_SLICE_X10Y102_DO6;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_D6 = CLBLL_L_X4Y101_SLICE_X5Y101_AO6;
  assign LIOB33_X0Y145_IOB_X0Y146_O = CLBLM_R_X3Y104_SLICE_X3Y104_BO6;
  assign LIOB33_X0Y145_IOB_X0Y145_O = CLBLM_R_X3Y104_SLICE_X3Y104_DO6;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_A1 = CLBLM_L_X10Y103_SLICE_X13Y103_BO6;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_A2 = CLBLM_L_X10Y102_SLICE_X13Y102_AO6;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_A3 = CLBLM_L_X10Y104_SLICE_X13Y104_AO6;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_A4 = CLBLM_R_X5Y102_SLICE_X6Y102_BO6;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_A5 = CLBLM_R_X5Y102_SLICE_X6Y102_AO6;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_A6 = CLBLM_L_X10Y103_SLICE_X12Y103_AO6;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_B2 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_B3 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_B4 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_B5 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_B6 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_C1 = CLBLM_R_X5Y102_SLICE_X6Y102_BO6;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_C2 = CLBLM_L_X10Y102_SLICE_X13Y102_AO6;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_C3 = CLBLM_R_X5Y102_SLICE_X6Y102_AO6;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_C4 = CLBLM_L_X10Y104_SLICE_X13Y104_AO6;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_C5 = CLBLM_L_X10Y103_SLICE_X12Y103_AO6;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_C6 = CLBLM_L_X10Y103_SLICE_X13Y103_BO6;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_D1 = CLBLM_L_X10Y104_SLICE_X13Y104_AO6;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_D2 = CLBLM_L_X10Y102_SLICE_X13Y102_AO6;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_D3 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_D4 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_D5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_D6 = CLBLM_L_X10Y103_SLICE_X13Y103_BO6;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_A1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_A2 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_A3 = 1'b1;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_A4 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_A5 = 1'b1;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_A6 = 1'b1;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_B1 = CLBLM_L_X10Y104_SLICE_X13Y104_CO6;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_B2 = CLBLM_L_X8Y103_SLICE_X10Y103_AO5;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_B3 = CLBLM_L_X10Y102_SLICE_X12Y102_CO6;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_B4 = CLBLM_L_X8Y104_SLICE_X10Y104_AO6;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_B5 = CLBLM_L_X8Y102_SLICE_X11Y102_AO6;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_B6 = CLBLM_L_X10Y104_SLICE_X12Y104_AO5;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_C1 = CLBLM_L_X8Y102_SLICE_X11Y102_AO6;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_C2 = CLBLM_L_X10Y102_SLICE_X12Y102_CO6;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_C3 = CLBLM_L_X8Y103_SLICE_X10Y103_AO5;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_C4 = CLBLM_L_X10Y104_SLICE_X12Y104_AO5;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_C5 = CLBLM_L_X10Y104_SLICE_X13Y104_CO6;
endmodule
