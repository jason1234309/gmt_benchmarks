module top(
  input LIOB33_SING_X0Y50_IOB_X0Y50_IPAD,
  input LIOB33_X0Y51_IOB_X0Y51_IPAD,
  input LIOB33_X0Y51_IOB_X0Y52_IPAD,
  input LIOB33_X0Y53_IOB_X0Y53_IPAD,
  input LIOB33_X0Y53_IOB_X0Y54_IPAD,
  input LIOB33_X0Y55_IOB_X0Y55_IPAD,
  input LIOB33_X0Y55_IOB_X0Y56_IPAD,
  input LIOB33_X0Y57_IOB_X0Y57_IPAD,
  input LIOB33_X0Y57_IOB_X0Y58_IPAD,
  input LIOB33_X0Y59_IOB_X0Y59_IPAD,
  input LIOB33_X0Y59_IOB_X0Y60_IPAD,
  input LIOB33_X0Y61_IOB_X0Y61_IPAD,
  input LIOB33_X0Y61_IOB_X0Y62_IPAD,
  input LIOB33_X0Y63_IOB_X0Y63_IPAD,
  input LIOB33_X0Y63_IOB_X0Y64_IPAD,
  input LIOB33_X0Y65_IOB_X0Y65_IPAD,
  input LIOB33_X0Y65_IOB_X0Y66_IPAD,
  input LIOB33_X0Y67_IOB_X0Y67_IPAD,
  input LIOB33_X0Y67_IOB_X0Y68_IPAD,
  input LIOB33_X0Y69_IOB_X0Y69_IPAD,
  input LIOB33_X0Y69_IOB_X0Y70_IPAD,
  input LIOB33_X0Y71_IOB_X0Y71_IPAD,
  input LIOB33_X0Y71_IOB_X0Y72_IPAD,
  input LIOB33_X0Y73_IOB_X0Y73_IPAD,
  input LIOB33_X0Y73_IOB_X0Y74_IPAD,
  input LIOB33_X0Y75_IOB_X0Y75_IPAD,
  input LIOB33_X0Y75_IOB_X0Y76_IPAD,
  input LIOB33_X0Y77_IOB_X0Y77_IPAD,
  input LIOB33_X0Y77_IOB_X0Y78_IPAD,
  input LIOB33_X0Y79_IOB_X0Y79_IPAD,
  input RIOB33_SING_X105Y100_IOB_X1Y100_IPAD,
  input RIOB33_SING_X105Y149_IOB_X1Y149_IPAD,
  input RIOB33_X105Y101_IOB_X1Y101_IPAD,
  input RIOB33_X105Y101_IOB_X1Y102_IPAD,
  input RIOB33_X105Y103_IOB_X1Y103_IPAD,
  input RIOB33_X105Y103_IOB_X1Y104_IPAD,
  input RIOB33_X105Y105_IOB_X1Y105_IPAD,
  input RIOB33_X105Y105_IOB_X1Y106_IPAD,
  input RIOB33_X105Y107_IOB_X1Y107_IPAD,
  input RIOB33_X105Y107_IOB_X1Y108_IPAD,
  input RIOB33_X105Y109_IOB_X1Y109_IPAD,
  input RIOB33_X105Y109_IOB_X1Y110_IPAD,
  input RIOB33_X105Y111_IOB_X1Y111_IPAD,
  input RIOB33_X105Y111_IOB_X1Y112_IPAD,
  input RIOB33_X105Y113_IOB_X1Y113_IPAD,
  input RIOB33_X105Y113_IOB_X1Y114_IPAD,
  input RIOB33_X105Y115_IOB_X1Y115_IPAD,
  input RIOB33_X105Y115_IOB_X1Y116_IPAD,
  input RIOB33_X105Y117_IOB_X1Y117_IPAD,
  input RIOB33_X105Y117_IOB_X1Y118_IPAD,
  input RIOB33_X105Y119_IOB_X1Y119_IPAD,
  input RIOB33_X105Y119_IOB_X1Y120_IPAD,
  input RIOB33_X105Y121_IOB_X1Y121_IPAD,
  input RIOB33_X105Y121_IOB_X1Y122_IPAD,
  input RIOB33_X105Y123_IOB_X1Y123_IPAD,
  input RIOB33_X105Y123_IOB_X1Y124_IPAD,
  input RIOB33_X105Y125_IOB_X1Y125_IPAD,
  input RIOB33_X105Y125_IOB_X1Y126_IPAD,
  input RIOB33_X105Y127_IOB_X1Y127_IPAD,
  input RIOB33_X105Y127_IOB_X1Y128_IPAD,
  input RIOB33_X105Y129_IOB_X1Y129_IPAD,
  input RIOB33_X105Y129_IOB_X1Y130_IPAD,
  input RIOB33_X105Y131_IOB_X1Y131_IPAD,
  input RIOB33_X105Y131_IOB_X1Y132_IPAD,
  input RIOB33_X105Y133_IOB_X1Y133_IPAD,
  input RIOB33_X105Y133_IOB_X1Y134_IPAD,
  input RIOB33_X105Y135_IOB_X1Y135_IPAD,
  input RIOB33_X105Y135_IOB_X1Y136_IPAD,
  input RIOB33_X105Y137_IOB_X1Y137_IPAD,
  input RIOB33_X105Y137_IOB_X1Y138_IPAD,
  input RIOB33_X105Y139_IOB_X1Y139_IPAD,
  input RIOB33_X105Y139_IOB_X1Y140_IPAD,
  input RIOB33_X105Y141_IOB_X1Y141_IPAD,
  input RIOB33_X105Y141_IOB_X1Y142_IPAD,
  input RIOB33_X105Y143_IOB_X1Y143_IPAD,
  input RIOB33_X105Y143_IOB_X1Y144_IPAD,
  input RIOB33_X105Y145_IOB_X1Y145_IPAD,
  input RIOB33_X105Y145_IOB_X1Y146_IPAD,
  input RIOB33_X105Y147_IOB_X1Y147_IPAD,
  input RIOB33_X105Y147_IOB_X1Y148_IPAD,
  output LIOB33_SING_X0Y100_IOB_X0Y100_OPAD,
  output LIOB33_SING_X0Y149_IOB_X0Y149_OPAD,
  output LIOB33_SING_X0Y150_IOB_X0Y150_OPAD,
  output LIOB33_SING_X0Y199_IOB_X0Y199_OPAD,
  output LIOB33_X0Y101_IOB_X0Y101_OPAD,
  output LIOB33_X0Y101_IOB_X0Y102_OPAD,
  output LIOB33_X0Y103_IOB_X0Y103_OPAD,
  output LIOB33_X0Y103_IOB_X0Y104_OPAD,
  output LIOB33_X0Y105_IOB_X0Y105_OPAD,
  output LIOB33_X0Y105_IOB_X0Y106_OPAD,
  output LIOB33_X0Y107_IOB_X0Y107_OPAD,
  output LIOB33_X0Y107_IOB_X0Y108_OPAD,
  output LIOB33_X0Y109_IOB_X0Y109_OPAD,
  output LIOB33_X0Y109_IOB_X0Y110_OPAD,
  output LIOB33_X0Y111_IOB_X0Y111_OPAD,
  output LIOB33_X0Y111_IOB_X0Y112_OPAD,
  output LIOB33_X0Y113_IOB_X0Y113_OPAD,
  output LIOB33_X0Y113_IOB_X0Y114_OPAD,
  output LIOB33_X0Y115_IOB_X0Y115_OPAD,
  output LIOB33_X0Y115_IOB_X0Y116_OPAD,
  output LIOB33_X0Y117_IOB_X0Y117_OPAD,
  output LIOB33_X0Y117_IOB_X0Y118_OPAD,
  output LIOB33_X0Y119_IOB_X0Y119_OPAD,
  output LIOB33_X0Y119_IOB_X0Y120_OPAD,
  output LIOB33_X0Y121_IOB_X0Y121_OPAD,
  output LIOB33_X0Y121_IOB_X0Y122_OPAD,
  output LIOB33_X0Y123_IOB_X0Y123_OPAD,
  output LIOB33_X0Y123_IOB_X0Y124_OPAD,
  output LIOB33_X0Y125_IOB_X0Y125_OPAD,
  output LIOB33_X0Y125_IOB_X0Y126_OPAD,
  output LIOB33_X0Y127_IOB_X0Y127_OPAD,
  output LIOB33_X0Y127_IOB_X0Y128_OPAD,
  output LIOB33_X0Y129_IOB_X0Y129_OPAD,
  output LIOB33_X0Y129_IOB_X0Y130_OPAD,
  output LIOB33_X0Y131_IOB_X0Y131_OPAD,
  output LIOB33_X0Y131_IOB_X0Y132_OPAD,
  output LIOB33_X0Y133_IOB_X0Y133_OPAD,
  output LIOB33_X0Y133_IOB_X0Y134_OPAD,
  output LIOB33_X0Y135_IOB_X0Y135_OPAD,
  output LIOB33_X0Y135_IOB_X0Y136_OPAD,
  output LIOB33_X0Y137_IOB_X0Y137_OPAD,
  output LIOB33_X0Y137_IOB_X0Y138_OPAD,
  output LIOB33_X0Y139_IOB_X0Y139_OPAD,
  output LIOB33_X0Y139_IOB_X0Y140_OPAD,
  output LIOB33_X0Y141_IOB_X0Y141_OPAD,
  output LIOB33_X0Y141_IOB_X0Y142_OPAD,
  output LIOB33_X0Y143_IOB_X0Y143_OPAD,
  output LIOB33_X0Y145_IOB_X0Y145_OPAD,
  output LIOB33_X0Y145_IOB_X0Y146_OPAD,
  output LIOB33_X0Y147_IOB_X0Y147_OPAD,
  output LIOB33_X0Y147_IOB_X0Y148_OPAD,
  output LIOB33_X0Y151_IOB_X0Y151_OPAD,
  output LIOB33_X0Y151_IOB_X0Y152_OPAD,
  output LIOB33_X0Y153_IOB_X0Y153_OPAD,
  output LIOB33_X0Y153_IOB_X0Y154_OPAD,
  output LIOB33_X0Y155_IOB_X0Y155_OPAD,
  output LIOB33_X0Y155_IOB_X0Y156_OPAD,
  output LIOB33_X0Y157_IOB_X0Y157_OPAD,
  output LIOB33_X0Y157_IOB_X0Y158_OPAD,
  output LIOB33_X0Y159_IOB_X0Y159_OPAD,
  output LIOB33_X0Y159_IOB_X0Y160_OPAD,
  output LIOB33_X0Y161_IOB_X0Y161_OPAD,
  output LIOB33_X0Y161_IOB_X0Y162_OPAD,
  output LIOB33_X0Y163_IOB_X0Y163_OPAD,
  output LIOB33_X0Y163_IOB_X0Y164_OPAD,
  output LIOB33_X0Y165_IOB_X0Y165_OPAD,
  output LIOB33_X0Y165_IOB_X0Y166_OPAD,
  output LIOB33_X0Y167_IOB_X0Y167_OPAD,
  output LIOB33_X0Y167_IOB_X0Y168_OPAD,
  output LIOB33_X0Y169_IOB_X0Y169_OPAD,
  output LIOB33_X0Y169_IOB_X0Y170_OPAD,
  output LIOB33_X0Y171_IOB_X0Y171_OPAD,
  output LIOB33_X0Y171_IOB_X0Y172_OPAD,
  output LIOB33_X0Y173_IOB_X0Y173_OPAD,
  output LIOB33_X0Y173_IOB_X0Y174_OPAD,
  output LIOB33_X0Y175_IOB_X0Y175_OPAD,
  output LIOB33_X0Y175_IOB_X0Y176_OPAD,
  output LIOB33_X0Y177_IOB_X0Y177_OPAD,
  output LIOB33_X0Y177_IOB_X0Y178_OPAD,
  output LIOB33_X0Y179_IOB_X0Y179_OPAD,
  output LIOB33_X0Y179_IOB_X0Y180_OPAD,
  output LIOB33_X0Y181_IOB_X0Y181_OPAD,
  output LIOB33_X0Y181_IOB_X0Y182_OPAD,
  output LIOB33_X0Y183_IOB_X0Y183_OPAD,
  output LIOB33_X0Y183_IOB_X0Y184_OPAD,
  output LIOB33_X0Y185_IOB_X0Y185_OPAD,
  output LIOB33_X0Y185_IOB_X0Y186_OPAD,
  output LIOB33_X0Y187_IOB_X0Y187_OPAD,
  output LIOB33_X0Y187_IOB_X0Y188_OPAD,
  output LIOB33_X0Y189_IOB_X0Y189_OPAD,
  output LIOB33_X0Y189_IOB_X0Y190_OPAD,
  output LIOB33_X0Y191_IOB_X0Y191_OPAD,
  output LIOB33_X0Y191_IOB_X0Y192_OPAD,
  output LIOB33_X0Y193_IOB_X0Y193_OPAD,
  output LIOB33_X0Y193_IOB_X0Y194_OPAD,
  output LIOB33_X0Y195_IOB_X0Y195_OPAD,
  output LIOB33_X0Y195_IOB_X0Y196_OPAD,
  output LIOB33_X0Y197_IOB_X0Y197_OPAD,
  output LIOB33_X0Y197_IOB_X0Y198_OPAD,
  output LIOB33_X0Y79_IOB_X0Y80_OPAD,
  output RIOB33_SING_X105Y150_IOB_X1Y150_OPAD,
  output RIOB33_SING_X105Y199_IOB_X1Y199_OPAD,
  output RIOB33_X105Y151_IOB_X1Y151_OPAD,
  output RIOB33_X105Y151_IOB_X1Y152_OPAD,
  output RIOB33_X105Y153_IOB_X1Y153_OPAD,
  output RIOB33_X105Y153_IOB_X1Y154_OPAD,
  output RIOB33_X105Y155_IOB_X1Y155_OPAD,
  output RIOB33_X105Y155_IOB_X1Y156_OPAD,
  output RIOB33_X105Y157_IOB_X1Y157_OPAD,
  output RIOB33_X105Y157_IOB_X1Y158_OPAD,
  output RIOB33_X105Y159_IOB_X1Y159_OPAD,
  output RIOB33_X105Y159_IOB_X1Y160_OPAD,
  output RIOB33_X105Y161_IOB_X1Y161_OPAD,
  output RIOB33_X105Y161_IOB_X1Y162_OPAD,
  output RIOB33_X105Y163_IOB_X1Y163_OPAD,
  output RIOB33_X105Y163_IOB_X1Y164_OPAD,
  output RIOB33_X105Y165_IOB_X1Y165_OPAD,
  output RIOB33_X105Y165_IOB_X1Y166_OPAD,
  output RIOB33_X105Y167_IOB_X1Y167_OPAD,
  output RIOB33_X105Y167_IOB_X1Y168_OPAD,
  output RIOB33_X105Y169_IOB_X1Y169_OPAD,
  output RIOB33_X105Y169_IOB_X1Y170_OPAD,
  output RIOB33_X105Y171_IOB_X1Y171_OPAD,
  output RIOB33_X105Y171_IOB_X1Y172_OPAD,
  output RIOB33_X105Y173_IOB_X1Y173_OPAD,
  output RIOB33_X105Y173_IOB_X1Y174_OPAD,
  output RIOB33_X105Y175_IOB_X1Y175_OPAD,
  output RIOB33_X105Y175_IOB_X1Y176_OPAD,
  output RIOB33_X105Y177_IOB_X1Y177_OPAD,
  output RIOB33_X105Y177_IOB_X1Y178_OPAD,
  output RIOB33_X105Y179_IOB_X1Y179_OPAD,
  output RIOB33_X105Y179_IOB_X1Y180_OPAD,
  output RIOB33_X105Y181_IOB_X1Y181_OPAD,
  output RIOB33_X105Y181_IOB_X1Y182_OPAD,
  output RIOB33_X105Y183_IOB_X1Y183_OPAD,
  output RIOB33_X105Y183_IOB_X1Y184_OPAD,
  output RIOB33_X105Y185_IOB_X1Y185_OPAD,
  output RIOB33_X105Y185_IOB_X1Y186_OPAD,
  output RIOB33_X105Y187_IOB_X1Y187_OPAD,
  output RIOB33_X105Y187_IOB_X1Y188_OPAD,
  output RIOB33_X105Y189_IOB_X1Y189_OPAD,
  output RIOB33_X105Y189_IOB_X1Y190_OPAD,
  output RIOB33_X105Y191_IOB_X1Y191_OPAD,
  output RIOB33_X105Y191_IOB_X1Y192_OPAD,
  output RIOB33_X105Y193_IOB_X1Y193_OPAD,
  output RIOB33_X105Y193_IOB_X1Y194_OPAD,
  output RIOB33_X105Y195_IOB_X1Y195_OPAD,
  output RIOB33_X105Y195_IOB_X1Y196_OPAD,
  output RIOB33_X105Y197_IOB_X1Y197_OPAD,
  output RIOB33_X105Y197_IOB_X1Y198_OPAD
  );
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_AO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_AO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_BO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_BO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_CO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_CO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_DO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_DO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_AO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_AO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_BO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_BO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_CO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_CO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_DO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_DO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D_XOR;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_A;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_A1;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_A2;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_A3;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_A4;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_A5;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_A6;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_AMUX;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_AO5;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_AO6;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_A_CY;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_A_XOR;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_B;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_B1;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_B2;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_B3;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_B4;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_B5;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_B6;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_BO5;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_BO6;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_B_CY;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_B_XOR;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_C;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_C1;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_C2;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_C3;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_C4;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_C5;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_C6;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_CO5;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_CO6;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_C_CY;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_C_XOR;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_D;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_D1;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_D2;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_D3;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_D4;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_D5;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_D6;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_DO5;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_DO6;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_D_CY;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_D_XOR;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_A;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_A1;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_A2;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_A3;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_A4;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_A5;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_A6;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_AO5;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_AO6;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_A_CY;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_A_XOR;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_B;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_B1;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_B2;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_B3;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_B4;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_B5;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_B6;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_BO5;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_BO6;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_B_CY;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_B_XOR;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_C;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_C1;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_C2;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_C3;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_C4;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_C5;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_C6;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_CO5;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_CO6;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_C_CY;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_C_XOR;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_D;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_D1;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_D2;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_D3;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_D4;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_D5;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_D6;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_DO5;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_DO6;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_D_CY;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_D_XOR;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_A;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_A1;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_A2;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_A3;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_A4;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_A5;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_A6;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_AMUX;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_AO5;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_AO6;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_A_CY;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_A_XOR;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_B;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_B1;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_B2;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_B3;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_B4;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_B5;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_B6;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_BMUX;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_BO5;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_BO6;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_B_CY;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_B_XOR;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_C;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_C1;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_C2;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_C3;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_C4;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_C5;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_C6;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_CMUX;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_CO5;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_CO6;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_C_CY;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_C_XOR;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_D;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_D1;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_D2;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_D3;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_D4;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_D5;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_D6;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_DO5;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_DO6;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_D_CY;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_D_XOR;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_A;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_A1;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_A2;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_A3;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_A4;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_A5;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_A6;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_AO5;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_AO6;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_A_CY;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_A_XOR;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_B;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_B1;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_B2;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_B3;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_B4;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_B5;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_B6;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_BO5;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_BO6;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_B_CY;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_B_XOR;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_C;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_C1;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_C2;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_C3;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_C4;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_C5;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_C6;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_CO5;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_CO6;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_C_CY;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_C_XOR;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_D;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_D1;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_D2;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_D3;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_D4;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_D5;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_D6;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_DO5;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_DO6;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_D_CY;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_D_XOR;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_A;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_A1;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_A2;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_A3;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_A4;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_A5;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_A6;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_AMUX;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_AO5;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_AO6;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_A_CY;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_A_XOR;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_B;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_B1;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_B2;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_B3;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_B4;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_B5;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_B6;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_BO5;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_BO6;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_B_CY;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_B_XOR;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_C;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_C1;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_C2;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_C3;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_C4;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_C5;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_C6;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_CO5;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_CO6;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_C_CY;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_C_XOR;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_D;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_D1;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_D2;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_D3;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_D4;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_D5;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_D6;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_DO5;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_DO6;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_D_CY;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X0Y141_D_XOR;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_A;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_A1;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_A2;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_A3;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_A4;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_A5;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_A6;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_AO5;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_AO6;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_A_CY;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_A_XOR;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_B;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_B1;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_B2;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_B3;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_B4;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_B5;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_B6;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_BO5;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_BO6;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_B_CY;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_B_XOR;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_C;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_C1;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_C2;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_C3;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_C4;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_C5;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_C6;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_CO5;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_CO6;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_C_CY;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_C_XOR;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_D;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_D1;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_D2;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_D3;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_D4;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_D5;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_D6;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_DO5;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_DO6;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_D_CY;
  wire [0:0] CLBLL_L_X2Y141_SLICE_X1Y141_D_XOR;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_A;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_A1;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_A2;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_A3;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_A4;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_A5;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_A6;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_AO5;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_AO6;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_A_CY;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_A_XOR;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_B;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_B1;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_B2;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_B3;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_B4;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_B5;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_B6;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_BO5;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_BO6;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_B_CY;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_B_XOR;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_C;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_C1;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_C2;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_C3;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_C4;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_C5;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_C6;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_CO5;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_CO6;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_C_CY;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_C_XOR;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_D;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_D1;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_D2;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_D3;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_D4;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_D5;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_D6;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_DO5;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_DO6;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_D_CY;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X0Y142_D_XOR;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_A;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_A1;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_A2;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_A3;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_A4;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_A5;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_A6;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_AO5;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_AO6;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_A_CY;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_A_XOR;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_B;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_B1;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_B2;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_B3;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_B4;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_B5;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_B6;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_BO5;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_BO6;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_B_CY;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_B_XOR;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_C;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_C1;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_C2;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_C3;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_C4;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_C5;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_C6;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_CO5;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_CO6;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_C_CY;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_C_XOR;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_D;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_D1;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_D2;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_D3;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_D4;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_D5;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_D6;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_DO5;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_DO6;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_D_CY;
  wire [0:0] CLBLL_L_X2Y142_SLICE_X1Y142_D_XOR;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_A;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_A1;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_A2;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_A3;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_A4;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_A5;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_A6;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_AO5;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_AO6;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_A_CY;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_A_XOR;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_B;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_B1;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_B2;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_B3;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_B4;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_B5;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_B6;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_BO5;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_BO6;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_B_CY;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_B_XOR;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_C;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_C1;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_C2;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_C3;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_C4;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_C5;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_C6;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_CO5;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_CO6;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_C_CY;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_C_XOR;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_D;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_D1;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_D2;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_D3;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_D4;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_D5;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_D6;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_DO5;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_DO6;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_D_CY;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_D_XOR;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_A;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_A1;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_A2;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_A3;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_A4;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_A5;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_A6;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_AO5;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_AO6;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_AQ;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_A_CY;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_A_XOR;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_B;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_B1;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_B2;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_B3;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_B4;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_B5;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_B6;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_BO5;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_BO6;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_BQ;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_B_CY;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_B_XOR;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_C;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_C1;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_C2;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_C3;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_C4;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_C5;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_C6;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_CLK;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_CO5;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_CO6;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_C_CY;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_C_XOR;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_D;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_D1;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_D2;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_D3;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_D4;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_D5;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_D6;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_DO5;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_DO6;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_D_CY;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_D_XOR;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_A;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_A1;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_A2;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_A3;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_A4;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_A5;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_A6;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_AO5;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_AO6;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_A_CY;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_A_XOR;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_B;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_B1;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_B2;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_B3;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_B4;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_B5;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_B6;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_BO5;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_BO6;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_B_CY;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_B_XOR;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_C;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_C1;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_C2;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_C3;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_C4;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_C5;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_C6;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_CO5;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_CO6;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_C_CY;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_C_XOR;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_D;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_D1;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_D2;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_D3;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_D4;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_D5;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_D6;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_DO5;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_DO6;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_D_CY;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_D_XOR;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_A;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_A1;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_A2;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_A3;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_A4;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_A5;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_A6;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_AO5;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_AO6;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_AQ;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_A_CY;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_A_XOR;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_B;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_B1;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_B2;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_B3;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_B4;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_B5;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_B6;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_BO5;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_BO6;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_BQ;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_B_CY;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_B_XOR;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_C;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_C1;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_C2;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_C3;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_C4;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_C5;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_C6;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_CLK;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_CO5;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_CO6;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_CQ;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_C_CY;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_C_XOR;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_D;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_D1;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_D2;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_D3;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_D4;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_D5;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_D6;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_DO5;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_DO6;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_D_CY;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_D_XOR;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_A;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_A1;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_A2;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_A3;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_A4;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_A5;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_A6;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_AO5;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_AO6;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_A_CY;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_A_XOR;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_B;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_B1;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_B2;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_B3;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_B4;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_B5;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_B6;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_BO5;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_BO6;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_B_CY;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_B_XOR;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_C;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_C1;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_C2;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_C3;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_C4;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_C5;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_C6;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_CO5;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_CO6;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_C_CY;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_C_XOR;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_D;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_D1;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_D2;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_D3;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_D4;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_D5;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_D6;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_DO5;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_DO6;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_D_CY;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_D_XOR;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_A;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_A1;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_A2;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_A3;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_A4;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_A5;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_A6;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_AMUX;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_AO5;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_AO6;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_AQ;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_AX;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_A_CY;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_A_XOR;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_B;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_B1;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_B2;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_B3;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_B4;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_B5;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_B6;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_BMUX;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_BO5;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_BO6;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_B_CY;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_B_XOR;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_C;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_C1;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_C2;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_C3;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_C4;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_C5;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_C6;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_CLK;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_CMUX;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_CO5;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_CO6;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_C_CY;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_C_XOR;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_D;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_D1;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_D2;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_D3;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_D4;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_D5;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_D6;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_DO5;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_DO6;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_D_CY;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_D_XOR;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_A;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_A1;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_A2;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_A3;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_A4;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_A5;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_A6;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_AO5;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_AO6;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_A_CY;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_A_XOR;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_B;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_B1;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_B2;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_B3;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_B4;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_B5;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_B6;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_BO5;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_BO6;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_B_CY;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_B_XOR;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_C;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_C1;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_C2;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_C3;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_C4;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_C5;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_C6;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_CO5;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_CO6;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_C_CY;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_C_XOR;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_D;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_D1;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_D2;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_D3;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_D4;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_D5;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_D6;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_DO5;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_DO6;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_D_CY;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_D_XOR;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_A;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_A1;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_A2;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_A3;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_A4;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_A5;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_A6;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_AO5;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_AO6;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_AQ;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_A_CY;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_A_XOR;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_B;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_B1;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_B2;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_B3;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_B4;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_B5;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_B6;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_BO5;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_BO6;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_B_CY;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_B_XOR;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_C;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_C1;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_C2;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_C3;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_C4;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_C5;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_C6;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_CLK;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_CO5;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_CO6;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_C_CY;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_C_XOR;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_D;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_D1;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_D2;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_D3;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_D4;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_D5;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_D6;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_DO5;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_DO6;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_D_CY;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_D_XOR;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_A;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_A1;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_A2;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_A3;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_A4;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_A5;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_A6;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_AO5;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_AO6;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_A_CY;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_A_XOR;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_B;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_B1;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_B2;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_B3;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_B4;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_B5;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_B6;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_BO5;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_BO6;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_B_CY;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_B_XOR;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_C;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_C1;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_C2;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_C3;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_C4;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_C5;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_C6;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_CO5;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_CO6;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_C_CY;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_C_XOR;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_D;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_D1;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_D2;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_D3;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_D4;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_D5;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_D6;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_DO5;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_DO6;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_D_CY;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_D_XOR;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_A;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_A1;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_A2;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_A3;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_A4;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_A5;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_A6;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_AO5;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_AO6;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_A_CY;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_A_XOR;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_B;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_B1;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_B2;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_B3;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_B4;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_B5;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_B6;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_BO5;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_BO6;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_B_CY;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_B_XOR;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_C;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_C1;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_C2;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_C3;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_C4;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_C5;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_C6;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_CO5;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_CO6;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_C_CY;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_C_XOR;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_D;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_D1;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_D2;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_D3;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_D4;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_D5;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_D6;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_DO5;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_DO6;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_D_CY;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_D_XOR;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_A;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_A1;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_A2;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_A3;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_A4;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_A5;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_A6;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_AMUX;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_AO5;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_AO6;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_A_CY;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_A_XOR;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_B;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_B1;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_B2;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_B3;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_B4;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_B5;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_B6;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_BO5;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_BO6;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_B_CY;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_B_XOR;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_C;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_C1;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_C2;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_C3;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_C4;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_C5;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_C6;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_CO5;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_CO6;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_C_CY;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_C_XOR;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_D;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_D1;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_D2;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_D3;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_D4;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_D5;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_D6;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_DO5;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_DO6;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_D_CY;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_D_XOR;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_A;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_A1;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_A2;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_A3;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_A4;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_A5;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_A6;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_AO5;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_AO6;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_A_CY;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_A_XOR;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_B;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_B1;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_B2;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_B3;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_B4;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_B5;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_B6;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_BO5;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_BO6;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_B_CY;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_B_XOR;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_C;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_C1;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_C2;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_C3;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_C4;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_C5;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_C6;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_CO5;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_CO6;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_C_CY;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_C_XOR;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_D;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_D1;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_D2;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_D3;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_D4;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_D5;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_D6;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_DO5;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_DO6;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_D_CY;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_D_XOR;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_A;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_A1;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_A2;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_A3;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_A4;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_A5;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_A6;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_AMUX;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_AO5;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_AO6;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_A_CY;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_A_XOR;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_B;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_B1;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_B2;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_B3;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_B4;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_B5;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_B6;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_BMUX;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_BO5;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_BO6;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_B_CY;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_B_XOR;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_C;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_C1;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_C2;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_C3;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_C4;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_C5;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_C6;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_CMUX;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_CO5;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_CO6;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_C_CY;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_C_XOR;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_D;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_D1;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_D2;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_D3;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_D4;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_D5;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_D6;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_DMUX;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_DO5;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_DO6;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_D_CY;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_D_XOR;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_A;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_A1;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_A2;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_A3;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_A4;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_A5;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_A6;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_AMUX;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_AO5;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_AO6;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_A_CY;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_A_XOR;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_B;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_B1;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_B2;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_B3;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_B4;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_B5;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_B6;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_BO5;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_BO6;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_B_CY;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_B_XOR;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_C;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_C1;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_C2;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_C3;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_C4;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_C5;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_C6;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_CO5;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_CO6;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_C_CY;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_C_XOR;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_D;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_D1;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_D2;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_D3;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_D4;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_D5;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_D6;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_DO5;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_DO6;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_D_CY;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_D_XOR;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_A;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_A1;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_A2;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_A3;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_A4;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_A5;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_A6;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_AO5;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_AO6;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_A_CY;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_A_XOR;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_B;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_B1;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_B2;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_B3;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_B4;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_B5;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_B6;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_BO5;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_BO6;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_B_CY;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_B_XOR;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_C;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_C1;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_C2;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_C3;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_C4;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_C5;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_C6;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_CO5;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_CO6;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_C_CY;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_C_XOR;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_D;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_D1;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_D2;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_D3;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_D4;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_D5;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_D6;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_DO5;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_DO6;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_D_CY;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_D_XOR;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_A;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_A1;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_A2;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_A3;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_A4;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_A5;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_A6;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_AMUX;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_AO5;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_AO6;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_A_CY;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_A_XOR;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_B;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_B1;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_B2;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_B3;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_B4;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_B5;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_B6;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_BMUX;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_BO5;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_BO6;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_B_CY;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_B_XOR;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_C;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_C1;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_C2;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_C3;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_C4;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_C5;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_C6;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_CO5;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_CO6;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_C_CY;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_C_XOR;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_D;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_D1;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_D2;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_D3;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_D4;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_D5;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_D6;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_DO5;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_DO6;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_D_CY;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_D_XOR;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_A;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_A1;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_A2;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_A3;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_A4;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_A5;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_A6;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_AO5;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_AO6;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_A_CY;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_A_XOR;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_B;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_B1;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_B2;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_B3;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_B4;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_B5;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_B6;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_BO5;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_BO6;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_B_CY;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_B_XOR;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_C;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_C1;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_C2;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_C3;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_C4;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_C5;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_C6;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_CO5;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_CO6;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_C_CY;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_C_XOR;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_D;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_D1;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_D2;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_D3;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_D4;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_D5;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_D6;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_DO5;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_DO6;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_D_CY;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_D_XOR;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_A;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_A1;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_A2;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_A3;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_A4;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_A5;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_A6;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_AMUX;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_AO5;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_AO6;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_A_CY;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_A_XOR;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_B;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_B1;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_B2;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_B3;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_B4;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_B5;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_B6;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_BO5;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_BO6;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_B_CY;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_B_XOR;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_C;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_C1;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_C2;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_C3;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_C4;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_C5;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_C6;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_CMUX;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_CO5;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_CO6;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_C_CY;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_C_XOR;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_D;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_D1;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_D2;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_D3;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_D4;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_D5;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_D6;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_DO5;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_DO6;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_D_CY;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_D_XOR;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_A;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_A1;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_A2;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_A3;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_A4;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_A5;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_A6;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_AO5;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_AO6;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_A_CY;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_A_XOR;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_B;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_B1;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_B2;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_B3;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_B4;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_B5;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_B6;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_BO5;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_BO6;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_B_CY;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_B_XOR;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_C;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_C1;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_C2;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_C3;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_C4;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_C5;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_C6;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_CO5;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_CO6;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_C_CY;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_C_XOR;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_D;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_D1;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_D2;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_D3;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_D4;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_D5;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_D6;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_DO5;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_DO6;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_D_CY;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_D_XOR;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_A;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_A1;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_A2;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_A3;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_A4;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_A5;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_A6;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_AMUX;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_AO5;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_AO6;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_A_CY;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_A_XOR;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_B;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_B1;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_B2;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_B3;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_B4;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_B5;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_B6;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_BMUX;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_BO5;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_BO6;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_B_CY;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_B_XOR;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_C;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_C1;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_C2;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_C3;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_C4;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_C5;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_C6;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_CMUX;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_CO5;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_CO6;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_C_CY;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_C_XOR;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_D;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_D1;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_D2;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_D3;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_D4;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_D5;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_D6;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_DO5;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_DO6;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_D_CY;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_D_XOR;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_A;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_A1;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_A2;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_A3;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_A4;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_A5;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_A6;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_AO5;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_AO6;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_A_CY;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_A_XOR;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_B;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_B1;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_B2;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_B3;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_B4;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_B5;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_B6;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_BO5;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_BO6;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_B_CY;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_B_XOR;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_C;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_C1;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_C2;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_C3;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_C4;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_C5;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_C6;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_CO5;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_CO6;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_C_CY;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_C_XOR;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_D;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_D1;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_D2;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_D3;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_D4;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_D5;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_D6;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_DO5;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_DO6;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_D_CY;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_D_XOR;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_A;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_A1;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_A2;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_A3;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_A4;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_A5;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_A6;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_AO5;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_AO6;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_A_CY;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_A_XOR;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_B;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_B1;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_B2;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_B3;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_B4;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_B5;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_B6;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_BO5;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_BO6;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_B_CY;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_B_XOR;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_C;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_C1;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_C2;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_C3;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_C4;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_C5;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_C6;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_CO5;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_CO6;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_C_CY;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_C_XOR;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_D;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_D1;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_D2;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_D3;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_D4;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_D5;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_D6;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_DO5;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_DO6;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_D_CY;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_D_XOR;
  wire [0:0] CLBLL_L_X36Y146_SLICE_X54Y146_A;
  wire [0:0] CLBLL_L_X36Y146_SLICE_X54Y146_A1;
  wire [0:0] CLBLL_L_X36Y146_SLICE_X54Y146_A2;
  wire [0:0] CLBLL_L_X36Y146_SLICE_X54Y146_A3;
  wire [0:0] CLBLL_L_X36Y146_SLICE_X54Y146_A4;
  wire [0:0] CLBLL_L_X36Y146_SLICE_X54Y146_A5;
  wire [0:0] CLBLL_L_X36Y146_SLICE_X54Y146_A6;
  wire [0:0] CLBLL_L_X36Y146_SLICE_X54Y146_AO5;
  wire [0:0] CLBLL_L_X36Y146_SLICE_X54Y146_AO6;
  wire [0:0] CLBLL_L_X36Y146_SLICE_X54Y146_A_CY;
  wire [0:0] CLBLL_L_X36Y146_SLICE_X54Y146_A_XOR;
  wire [0:0] CLBLL_L_X36Y146_SLICE_X54Y146_B;
  wire [0:0] CLBLL_L_X36Y146_SLICE_X54Y146_B1;
  wire [0:0] CLBLL_L_X36Y146_SLICE_X54Y146_B2;
  wire [0:0] CLBLL_L_X36Y146_SLICE_X54Y146_B3;
  wire [0:0] CLBLL_L_X36Y146_SLICE_X54Y146_B4;
  wire [0:0] CLBLL_L_X36Y146_SLICE_X54Y146_B5;
  wire [0:0] CLBLL_L_X36Y146_SLICE_X54Y146_B6;
  wire [0:0] CLBLL_L_X36Y146_SLICE_X54Y146_BO5;
  wire [0:0] CLBLL_L_X36Y146_SLICE_X54Y146_BO6;
  wire [0:0] CLBLL_L_X36Y146_SLICE_X54Y146_B_CY;
  wire [0:0] CLBLL_L_X36Y146_SLICE_X54Y146_B_XOR;
  wire [0:0] CLBLL_L_X36Y146_SLICE_X54Y146_C;
  wire [0:0] CLBLL_L_X36Y146_SLICE_X54Y146_C1;
  wire [0:0] CLBLL_L_X36Y146_SLICE_X54Y146_C2;
  wire [0:0] CLBLL_L_X36Y146_SLICE_X54Y146_C3;
  wire [0:0] CLBLL_L_X36Y146_SLICE_X54Y146_C4;
  wire [0:0] CLBLL_L_X36Y146_SLICE_X54Y146_C5;
  wire [0:0] CLBLL_L_X36Y146_SLICE_X54Y146_C6;
  wire [0:0] CLBLL_L_X36Y146_SLICE_X54Y146_CO5;
  wire [0:0] CLBLL_L_X36Y146_SLICE_X54Y146_CO6;
  wire [0:0] CLBLL_L_X36Y146_SLICE_X54Y146_C_CY;
  wire [0:0] CLBLL_L_X36Y146_SLICE_X54Y146_C_XOR;
  wire [0:0] CLBLL_L_X36Y146_SLICE_X54Y146_D;
  wire [0:0] CLBLL_L_X36Y146_SLICE_X54Y146_D1;
  wire [0:0] CLBLL_L_X36Y146_SLICE_X54Y146_D2;
  wire [0:0] CLBLL_L_X36Y146_SLICE_X54Y146_D3;
  wire [0:0] CLBLL_L_X36Y146_SLICE_X54Y146_D4;
  wire [0:0] CLBLL_L_X36Y146_SLICE_X54Y146_D5;
  wire [0:0] CLBLL_L_X36Y146_SLICE_X54Y146_D6;
  wire [0:0] CLBLL_L_X36Y146_SLICE_X54Y146_DO5;
  wire [0:0] CLBLL_L_X36Y146_SLICE_X54Y146_DO6;
  wire [0:0] CLBLL_L_X36Y146_SLICE_X54Y146_D_CY;
  wire [0:0] CLBLL_L_X36Y146_SLICE_X54Y146_D_XOR;
  wire [0:0] CLBLL_L_X36Y146_SLICE_X55Y146_A;
  wire [0:0] CLBLL_L_X36Y146_SLICE_X55Y146_A1;
  wire [0:0] CLBLL_L_X36Y146_SLICE_X55Y146_A2;
  wire [0:0] CLBLL_L_X36Y146_SLICE_X55Y146_A3;
  wire [0:0] CLBLL_L_X36Y146_SLICE_X55Y146_A4;
  wire [0:0] CLBLL_L_X36Y146_SLICE_X55Y146_A5;
  wire [0:0] CLBLL_L_X36Y146_SLICE_X55Y146_A6;
  wire [0:0] CLBLL_L_X36Y146_SLICE_X55Y146_AO5;
  wire [0:0] CLBLL_L_X36Y146_SLICE_X55Y146_AO6;
  wire [0:0] CLBLL_L_X36Y146_SLICE_X55Y146_A_CY;
  wire [0:0] CLBLL_L_X36Y146_SLICE_X55Y146_A_XOR;
  wire [0:0] CLBLL_L_X36Y146_SLICE_X55Y146_B;
  wire [0:0] CLBLL_L_X36Y146_SLICE_X55Y146_B1;
  wire [0:0] CLBLL_L_X36Y146_SLICE_X55Y146_B2;
  wire [0:0] CLBLL_L_X36Y146_SLICE_X55Y146_B3;
  wire [0:0] CLBLL_L_X36Y146_SLICE_X55Y146_B4;
  wire [0:0] CLBLL_L_X36Y146_SLICE_X55Y146_B5;
  wire [0:0] CLBLL_L_X36Y146_SLICE_X55Y146_B6;
  wire [0:0] CLBLL_L_X36Y146_SLICE_X55Y146_BO5;
  wire [0:0] CLBLL_L_X36Y146_SLICE_X55Y146_BO6;
  wire [0:0] CLBLL_L_X36Y146_SLICE_X55Y146_B_CY;
  wire [0:0] CLBLL_L_X36Y146_SLICE_X55Y146_B_XOR;
  wire [0:0] CLBLL_L_X36Y146_SLICE_X55Y146_C;
  wire [0:0] CLBLL_L_X36Y146_SLICE_X55Y146_C1;
  wire [0:0] CLBLL_L_X36Y146_SLICE_X55Y146_C2;
  wire [0:0] CLBLL_L_X36Y146_SLICE_X55Y146_C3;
  wire [0:0] CLBLL_L_X36Y146_SLICE_X55Y146_C4;
  wire [0:0] CLBLL_L_X36Y146_SLICE_X55Y146_C5;
  wire [0:0] CLBLL_L_X36Y146_SLICE_X55Y146_C6;
  wire [0:0] CLBLL_L_X36Y146_SLICE_X55Y146_CO5;
  wire [0:0] CLBLL_L_X36Y146_SLICE_X55Y146_CO6;
  wire [0:0] CLBLL_L_X36Y146_SLICE_X55Y146_C_CY;
  wire [0:0] CLBLL_L_X36Y146_SLICE_X55Y146_C_XOR;
  wire [0:0] CLBLL_L_X36Y146_SLICE_X55Y146_D;
  wire [0:0] CLBLL_L_X36Y146_SLICE_X55Y146_D1;
  wire [0:0] CLBLL_L_X36Y146_SLICE_X55Y146_D2;
  wire [0:0] CLBLL_L_X36Y146_SLICE_X55Y146_D3;
  wire [0:0] CLBLL_L_X36Y146_SLICE_X55Y146_D4;
  wire [0:0] CLBLL_L_X36Y146_SLICE_X55Y146_D5;
  wire [0:0] CLBLL_L_X36Y146_SLICE_X55Y146_D6;
  wire [0:0] CLBLL_L_X36Y146_SLICE_X55Y146_DO5;
  wire [0:0] CLBLL_L_X36Y146_SLICE_X55Y146_DO6;
  wire [0:0] CLBLL_L_X36Y146_SLICE_X55Y146_D_CY;
  wire [0:0] CLBLL_L_X36Y146_SLICE_X55Y146_D_XOR;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_A;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_A1;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_A2;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_A3;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_A4;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_A5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_A6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_AO5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_AO6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_A_CY;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_A_XOR;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_B;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_B1;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_B2;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_B3;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_B4;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_B5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_B6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_BO5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_BO6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_B_CY;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_B_XOR;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_C;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_C1;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_C2;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_C3;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_C4;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_C5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_C6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_CO5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_CO6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_C_CY;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_C_XOR;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_D;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_D1;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_D2;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_D3;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_D4;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_D5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_D6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_DO5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_DO6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_D_CY;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_D_XOR;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_A;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_A1;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_A2;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_A3;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_A4;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_A5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_A6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_AMUX;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_AO5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_AO6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_AQ;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_A_CY;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_A_XOR;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_B;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_B1;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_B2;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_B3;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_B4;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_B5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_B6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_BO5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_BO6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_B_CY;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_B_XOR;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_C;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_C1;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_C2;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_C3;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_C4;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_C5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_C6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_CLK;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_CO5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_CO6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_C_CY;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_C_XOR;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_D;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_D1;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_D2;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_D3;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_D4;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_D5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_D6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_DO5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_DO6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_D_CY;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_D_XOR;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_A;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_A1;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_A2;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_A3;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_A4;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_A5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_A6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_AO5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_AO6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_AQ;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_A_CY;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_A_XOR;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_B;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_B1;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_B2;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_B3;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_B4;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_B5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_B6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_BO5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_BO6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_BQ;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_B_CY;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_B_XOR;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_C;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_C1;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_C2;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_C3;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_C4;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_C5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_C6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_CLK;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_CMUX;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_CO5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_CO6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_C_CY;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_C_XOR;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_D;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_D1;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_D2;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_D3;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_D4;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_D5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_D6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_DO5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_DO6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_D_CY;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_D_XOR;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_A;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_A1;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_A2;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_A3;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_A4;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_A5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_A6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_AO5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_AO6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_A_CY;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_A_XOR;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_B;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_B1;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_B2;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_B3;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_B4;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_B5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_B6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_BO5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_BO6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_B_CY;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_B_XOR;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_C;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_C1;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_C2;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_C3;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_C4;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_C5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_C6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_CO5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_CO6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_C_CY;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_C_XOR;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_D;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_D1;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_D2;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_D3;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_D4;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_D5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_D6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_DO5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_DO6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_D_CY;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_D_XOR;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_A;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_A1;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_A2;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_A3;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_A4;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_A5;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_A6;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_AO5;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_AO6;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_AQ;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_A_CY;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_A_XOR;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_B;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_B1;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_B2;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_B3;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_B4;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_B5;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_B6;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_BO5;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_BO6;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_BQ;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_B_CY;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_B_XOR;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_C;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_C1;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_C2;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_C3;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_C4;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_C5;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_C6;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_CLK;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_CMUX;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_CO5;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_CO6;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_C_CY;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_C_XOR;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_D;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_D1;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_D2;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_D3;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_D4;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_D5;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_D6;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_DO5;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_DO6;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_D_CY;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_D_XOR;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_A;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_A1;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_A2;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_A3;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_A4;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_A5;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_A5Q;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_A6;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_AMUX;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_AO5;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_AO6;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_AQ;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_AX;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_A_CY;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_A_XOR;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_B;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_B1;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_B2;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_B3;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_B4;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_B5;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_B6;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_BO5;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_BO6;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_BQ;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_B_CY;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_B_XOR;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_C;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_C1;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_C2;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_C3;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_C4;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_C5;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_C6;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_CLK;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_CMUX;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_CO5;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_CO6;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_C_CY;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_C_XOR;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_D;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_D1;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_D2;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_D3;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_D4;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_D5;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_D6;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_DO5;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_DO6;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_D_CY;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_D_XOR;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_A;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_A1;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_A2;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_A3;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_A4;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_A5;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_A5Q;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_A6;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_AMUX;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_AO5;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_AO6;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_AQ;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_AX;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_A_CY;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_A_XOR;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_B;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_B1;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_B2;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_B3;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_B4;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_B5;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_B6;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_BMUX;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_BO5;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_BO6;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_BQ;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_B_CY;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_B_XOR;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_C;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_C1;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_C2;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_C3;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_C4;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_C5;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_C6;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_CLK;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_CO5;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_CO6;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_CQ;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_C_CY;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_C_XOR;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_D;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_D1;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_D2;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_D3;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_D4;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_D5;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_D6;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_DO5;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_DO6;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_D_CY;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_D_XOR;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_A;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_A1;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_A2;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_A3;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_A4;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_A5;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_A6;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_AO5;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_AO6;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_AQ;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_A_CY;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_A_XOR;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_B;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_B1;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_B2;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_B3;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_B4;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_B5;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_B6;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_BMUX;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_BO5;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_BO6;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_B_CY;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_B_XOR;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_C;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_C1;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_C2;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_C3;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_C4;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_C5;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_C6;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_CLK;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_CO5;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_CO6;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_C_CY;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_C_XOR;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_D;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_D1;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_D2;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_D3;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_D4;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_D5;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_D6;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_DO5;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_DO6;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_D_CY;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_D_XOR;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_A;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_A1;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_A2;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_A3;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_A4;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_A5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_A5Q;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_A6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_AMUX;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_AO5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_AO6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_AQ;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_AX;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_A_CY;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_A_XOR;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_B;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_B1;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_B2;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_B3;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_B4;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_B5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_B6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_BO5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_BO6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_BQ;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_B_CY;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_B_XOR;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_C;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_C1;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_C2;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_C3;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_C4;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_C5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_C6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_CLK;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_CMUX;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_CO5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_CO6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_C_CY;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_C_XOR;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_D;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_D1;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_D2;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_D3;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_D4;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_D5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_D6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_DO5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_DO6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_D_CY;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_D_XOR;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_A;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_A1;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_A2;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_A3;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_A4;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_A5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_A5Q;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_A6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_AMUX;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_AO5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_AO6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_AQ;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_AX;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_A_CY;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_A_XOR;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_B;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_B1;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_B2;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_B3;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_B4;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_B5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_B6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_BMUX;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_BO5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_BO6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_B_CY;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_B_XOR;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_C;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_C1;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_C2;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_C3;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_C4;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_C5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_C6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_CLK;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_CO5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_CO6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_CQ;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_C_CY;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_C_XOR;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_D;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_D1;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_D2;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_D3;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_D4;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_D5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_D6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_DO5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_DO6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_D_CY;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_D_XOR;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_A;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_A1;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_A2;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_A3;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_A4;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_A5;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_A6;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_AO5;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_AO6;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_AQ;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_A_CY;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_A_XOR;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_B;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_B1;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_B2;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_B3;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_B4;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_B5;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_B6;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_BO5;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_BO6;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_BQ;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_B_CY;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_B_XOR;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_C;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_C1;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_C2;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_C3;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_C4;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_C5;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_C6;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_CLK;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_CO5;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_CO6;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_CQ;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_C_CY;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_C_XOR;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_D;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_D1;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_D2;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_D3;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_D4;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_D5;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_D6;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_DO5;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_DO6;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_D_CY;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_D_XOR;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_A;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_A1;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_A2;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_A3;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_A4;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_A5;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_A6;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_AO5;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_AO6;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_AQ;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_A_CY;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_A_XOR;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_B;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_B1;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_B2;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_B3;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_B4;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_B5;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_B5Q;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_B6;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_BMUX;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_BO5;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_BO6;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_BQ;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_B_CY;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_B_XOR;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_C;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_C1;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_C2;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_C3;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_C4;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_C5;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_C6;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_CLK;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_CO5;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_CO6;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_CQ;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_C_CY;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_C_XOR;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_D;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_D1;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_D2;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_D3;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_D4;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_D5;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_D6;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_DO5;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_DO6;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_D_CY;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_D_XOR;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_A;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_A1;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_A2;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_A3;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_A4;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_A5;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_A6;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_AO5;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_AO6;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_AQ;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_A_CY;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_A_XOR;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_B;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_B1;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_B2;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_B3;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_B4;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_B5;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_B6;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_BO5;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_BO6;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_BQ;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_B_CY;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_B_XOR;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_C;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_C1;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_C2;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_C3;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_C4;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_C5;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_C5Q;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_C6;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_CLK;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_CMUX;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_CO5;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_CO6;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_CQ;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_C_CY;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_C_XOR;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_D;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_D1;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_D2;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_D3;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_D4;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_D5;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_D6;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_DO5;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_DO6;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_DQ;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_D_CY;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_D_XOR;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_A;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_A1;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_A2;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_A3;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_A4;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_A5;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_A6;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_AO5;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_AO6;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_AQ;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_A_CY;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_A_XOR;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_B;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_B1;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_B2;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_B3;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_B4;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_B5;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_B6;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_BO5;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_BO6;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_BQ;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_B_CY;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_B_XOR;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_C;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_C1;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_C2;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_C3;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_C4;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_C5;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_C6;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_CLK;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_CO5;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_CO6;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_CQ;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_C_CY;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_C_XOR;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_D;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_D1;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_D2;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_D3;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_D4;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_D5;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_D6;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_DO5;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_DO6;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_D_CY;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_D_XOR;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_A;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_A1;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_A2;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_A3;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_A4;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_A5;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_A6;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_AO5;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_AO6;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_AQ;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_A_CY;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_A_XOR;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_B;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_B1;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_B2;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_B3;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_B4;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_B5;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_B6;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_BO5;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_BO6;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_BQ;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_B_CY;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_B_XOR;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_C;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_C1;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_C2;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_C3;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_C4;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_C5;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_C6;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_CLK;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_CO5;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_CO6;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_CQ;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_C_CY;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_C_XOR;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_D;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_D1;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_D2;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_D3;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_D4;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_D5;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_D6;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_DO5;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_DO6;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_DQ;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_D_CY;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_D_XOR;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_A;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_A1;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_A2;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_A3;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_A4;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_A5;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_A5Q;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_A6;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_AMUX;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_AO5;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_AO6;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_AQ;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_AX;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_A_CY;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_A_XOR;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_B;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_B1;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_B2;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_B3;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_B4;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_B5;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_B6;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_BMUX;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_BO5;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_BO6;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_B_CY;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_B_XOR;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_C;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_C1;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_C2;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_C3;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_C4;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_C5;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_C6;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_CLK;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_CO5;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_CO6;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_CQ;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_C_CY;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_C_XOR;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_D;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_D1;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_D2;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_D3;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_D4;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_D5;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_D6;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_DO5;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_DO6;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_DQ;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_D_CY;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_D_XOR;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_A;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_A1;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_A2;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_A3;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_A4;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_A5;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_A6;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_AO5;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_AO6;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_AQ;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_A_CY;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_A_XOR;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_B;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_B1;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_B2;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_B3;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_B4;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_B5;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_B5Q;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_B6;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_BMUX;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_BO5;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_BO6;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_BQ;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_B_CY;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_B_XOR;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_C;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_C1;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_C2;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_C3;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_C4;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_C5;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_C6;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_CLK;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_CO5;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_CO6;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_C_CY;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_C_XOR;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_D;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_D1;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_D2;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_D3;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_D4;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_D5;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_D6;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_DO5;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_DO6;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_D_CY;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_D_XOR;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_A;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_A1;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_A2;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_A3;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_A4;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_A5;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_A6;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_AO5;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_AO6;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_AQ;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_A_CY;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_A_XOR;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_B;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_B1;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_B2;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_B3;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_B4;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_B5;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_B6;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_BO5;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_BO6;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_BQ;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_B_CY;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_B_XOR;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_C;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_C1;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_C2;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_C3;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_C4;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_C5;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_C6;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_CLK;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_CO5;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_CO6;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_C_CY;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_C_XOR;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_D;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_D1;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_D2;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_D3;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_D4;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_D5;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_D6;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_DO5;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_DO6;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_D_CY;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_D_XOR;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_A;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_A1;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_A2;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_A3;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_A4;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_A5;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_A5Q;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_A6;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_AMUX;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_AO5;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_AO6;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_AQ;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_AX;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_A_CY;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_A_XOR;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_B;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_B1;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_B2;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_B3;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_B4;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_B5;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_B6;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_BO5;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_BO6;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_B_CY;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_B_XOR;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_C;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_C1;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_C2;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_C3;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_C4;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_C5;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_C6;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_CLK;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_CO5;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_CO6;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_C_CY;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_C_XOR;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_D;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_D1;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_D2;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_D3;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_D4;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_D5;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_D6;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_DO5;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_DO6;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_D_CY;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_D_XOR;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_A;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_A1;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_A2;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_A3;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_A4;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_A5;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_A6;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_AO5;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_AO6;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_AQ;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_A_CY;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_A_XOR;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_B;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_B1;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_B2;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_B3;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_B4;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_B5;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_B5Q;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_B6;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_BMUX;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_BO5;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_BO6;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_BQ;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_B_CY;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_B_XOR;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_C;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_C1;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_C2;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_C3;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_C4;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_C5;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_C6;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_CLK;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_CO5;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_CO6;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_C_CY;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_C_XOR;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_D;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_D1;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_D2;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_D3;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_D4;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_D5;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_D6;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_DMUX;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_DO5;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_DO6;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_D_CY;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_D_XOR;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_A;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_A1;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_A2;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_A3;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_A4;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_A5;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_A6;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_AMUX;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_AO5;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_AO6;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_A_CY;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_A_XOR;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_B;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_B1;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_B2;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_B3;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_B4;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_B5;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_B6;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_BO5;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_BO6;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_B_CY;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_B_XOR;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_C;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_C1;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_C2;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_C3;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_C4;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_C5;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_C6;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_CMUX;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_CO5;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_CO6;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_C_CY;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_C_XOR;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_D;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_D1;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_D2;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_D3;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_D4;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_D5;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_D6;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_DO5;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_DO6;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_D_CY;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_D_XOR;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_A;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_A1;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_A2;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_A3;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_A4;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_A5;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_A6;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_AMUX;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_AO5;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_AO6;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_A_CY;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_A_XOR;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_B;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_B1;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_B2;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_B3;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_B4;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_B5;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_B6;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_BO5;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_BO6;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_B_CY;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_B_XOR;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_C;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_C1;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_C2;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_C3;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_C4;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_C5;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_C6;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_CO5;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_CO6;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_C_CY;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_C_XOR;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_D;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_D1;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_D2;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_D3;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_D4;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_D5;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_D6;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_DO5;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_DO6;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_D_CY;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_D_XOR;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_A;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_A1;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_A2;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_A3;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_A4;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_A5;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_A6;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_AO5;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_AO6;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_A_CY;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_A_XOR;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_B;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_B1;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_B2;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_B3;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_B4;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_B5;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_B6;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_BO5;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_BO6;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_B_CY;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_B_XOR;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_C;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_C1;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_C2;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_C3;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_C4;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_C5;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_C6;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_CO5;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_CO6;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_C_CY;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_C_XOR;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_D;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_D1;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_D2;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_D3;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_D4;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_D5;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_D6;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_DO5;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_DO6;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_D_CY;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_D_XOR;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_A;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_A1;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_A2;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_A3;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_A4;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_A5;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_A6;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_AO5;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_AO6;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_AQ;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_A_CY;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_A_XOR;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_B;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_B1;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_B2;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_B3;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_B4;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_B5;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_B6;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_BO5;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_BO6;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_B_CY;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_B_XOR;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_C;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_C1;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_C2;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_C3;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_C4;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_C5;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_C6;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_CLK;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_CO5;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_CO6;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_C_CY;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_C_XOR;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_D;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_D1;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_D2;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_D3;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_D4;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_D5;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_D6;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_DO5;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_DO6;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_D_CY;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_D_XOR;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_A;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_A1;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_A2;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_A3;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_A4;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_A5;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_A6;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_AMUX;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_AO5;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_AO6;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_A_CY;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_A_XOR;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_B;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_B1;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_B2;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_B3;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_B4;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_B5;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_B6;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_BO5;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_BO6;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_B_CY;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_B_XOR;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_C;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_C1;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_C2;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_C3;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_C4;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_C5;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_C6;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_CO5;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_CO6;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_C_CY;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_C_XOR;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_D;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_D1;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_D2;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_D3;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_D4;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_D5;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_D6;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_DO5;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_DO6;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_D_CY;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_D_XOR;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_A;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_A1;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_A2;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_A3;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_A4;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_A5;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_A6;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_AO5;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_AO6;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_AQ;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_A_CY;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_A_XOR;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_B;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_B1;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_B2;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_B3;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_B4;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_B5;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_B6;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_BO5;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_BO6;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_BQ;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_B_CY;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_B_XOR;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_C;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_C1;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_C2;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_C3;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_C4;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_C5;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_C6;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_CLK;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_CMUX;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_CO5;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_CO6;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_C_CY;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_C_XOR;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_D;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_D1;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_D2;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_D3;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_D4;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_D5;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_D6;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_DO5;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_DO6;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_D_CY;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_D_XOR;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_A;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_A1;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_A2;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_A3;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_A4;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_A5;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_A6;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_AMUX;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_AO5;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_AO6;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_A_CY;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_A_XOR;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_B;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_B1;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_B2;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_B3;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_B4;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_B5;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_B6;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_BMUX;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_BO5;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_BO6;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_B_CY;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_B_XOR;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_C;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_C1;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_C2;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_C3;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_C4;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_C5;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_C6;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_CO5;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_CO6;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_C_CY;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_C_XOR;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_D;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_D1;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_D2;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_D3;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_D4;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_D5;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_D6;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_DO5;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_DO6;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_D_CY;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_D_XOR;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_A;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_A1;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_A2;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_A3;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_A4;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_A5;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_A6;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_AMUX;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_AO5;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_AO6;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_A_CY;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_A_XOR;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_B;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_B1;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_B2;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_B3;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_B4;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_B5;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_B6;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_BO5;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_BO6;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_B_CY;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_B_XOR;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_C;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_C1;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_C2;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_C3;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_C4;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_C5;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_C6;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_CO5;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_CO6;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_C_CY;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_C_XOR;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_D;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_D1;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_D2;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_D3;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_D4;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_D5;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_D6;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_DO5;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_DO6;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_D_CY;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_D_XOR;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A1;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A2;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A3;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A4;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_AO5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_AO6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A_CY;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A_XOR;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B1;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B2;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B3;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B4;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_BO5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_BO6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B_CY;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B_XOR;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C1;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C2;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C3;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C4;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_CO5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_CO6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C_CY;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C_XOR;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D1;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D2;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D3;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D4;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_DO5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_DO6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D_CY;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D_XOR;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A1;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A2;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A3;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A4;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_AO5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_AO6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A_CY;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A_XOR;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B1;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B2;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B3;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B4;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_BO5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_BO6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B_CY;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B_XOR;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C1;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C2;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C3;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C4;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_CO5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_CO6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C_CY;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C_XOR;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D1;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D2;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D3;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D4;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_DO5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_DO6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D_CY;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D_XOR;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_A;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_A1;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_A2;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_A3;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_A4;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_A5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_A6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_AMUX;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_AO5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_AO6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_A_CY;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_A_XOR;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_B;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_B1;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_B2;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_B3;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_B4;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_B5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_B6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_BMUX;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_BO5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_BO6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_B_CY;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_B_XOR;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_C;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_C1;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_C2;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_C3;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_C4;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_C5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_C6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_CO5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_CO6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_C_CY;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_C_XOR;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_D;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_D1;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_D2;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_D3;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_D4;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_D5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_D6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_DO5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_DO6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_D_CY;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_D_XOR;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_A;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_A1;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_A2;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_A3;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_A4;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_A5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_A6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_AO5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_AO6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_A_CY;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_A_XOR;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_B;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_B1;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_B2;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_B3;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_B4;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_B5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_B6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_BO5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_BO6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_B_CY;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_B_XOR;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_C;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_C1;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_C2;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_C3;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_C4;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_C5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_C6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_CO5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_CO6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_C_CY;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_C_XOR;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_D;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_D1;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_D2;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_D3;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_D4;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_D5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_D6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_DO5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_DO6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_D_CY;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_D_XOR;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_A;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_A1;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_A2;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_A3;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_A4;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_A5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_A6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_AO5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_AO6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_A_CY;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_A_XOR;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_B;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_B1;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_B2;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_B3;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_B4;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_B5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_B6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_BO5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_BO6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_B_CY;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_B_XOR;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_C;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_C1;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_C2;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_C3;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_C4;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_C5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_C6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_CO5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_CO6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_C_CY;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_C_XOR;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_D;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_D1;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_D2;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_D3;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_D4;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_D5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_D6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_DO5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_DO6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_D_CY;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_D_XOR;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_A;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_A1;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_A2;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_A3;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_A4;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_A5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_A6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_AO5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_AO6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_AQ;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_A_CY;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_A_XOR;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_B;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_B1;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_B2;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_B3;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_B4;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_B5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_B6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_BMUX;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_BO5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_BO6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_B_CY;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_B_XOR;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_C;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_C1;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_C2;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_C3;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_C4;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_C5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_C6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_CLK;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_CMUX;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_CO5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_CO6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_C_CY;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_C_XOR;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_D;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_D1;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_D2;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_D3;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_D4;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_D5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_D6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_DMUX;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_DO5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_DO6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_D_CY;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_D_XOR;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_A;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_A1;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_A2;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_A3;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_A4;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_A5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_A6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_AO5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_AO6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_A_CY;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_A_XOR;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_B;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_B1;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_B2;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_B3;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_B4;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_B5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_B6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_BO5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_BO6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_B_CY;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_B_XOR;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_C;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_C1;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_C2;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_C3;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_C4;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_C5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_C6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_CO5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_CO6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_C_CY;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_C_XOR;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_D;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_D1;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_D2;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_D3;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_D4;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_D5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_D6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_DO5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_DO6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_D_CY;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_D_XOR;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_A;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_A1;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_A2;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_A3;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_A4;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_A5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_A6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_AO5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_AO6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_AQ;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_A_CY;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_A_XOR;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_B;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_B1;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_B2;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_B3;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_B4;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_B5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_B6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_BO5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_BO6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_BQ;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_B_CY;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_B_XOR;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_C;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_C1;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_C2;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_C3;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_C4;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_C5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_C6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_CLK;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_CMUX;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_CO5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_CO6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_C_CY;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_C_XOR;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_D;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_D1;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_D2;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_D3;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_D4;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_D5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_D6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_DMUX;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_DO5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_DO6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_D_CY;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_D_XOR;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_A;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_A1;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_A2;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_A3;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_A4;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_A5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_A6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_AO5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_AO6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_AQ;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_A_CY;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_A_XOR;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_B;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_B1;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_B2;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_B3;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_B4;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_B5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_B6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_BO5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_BO6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_BQ;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_B_CY;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_B_XOR;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_C;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_C1;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_C2;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_C3;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_C4;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_C5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_C6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_CLK;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_CO5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_CO6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_CQ;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_C_CY;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_C_XOR;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_D;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_D1;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_D2;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_D3;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_D4;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_D5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_D6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_DO5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_DO6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_D_CY;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_D_XOR;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_A;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_A1;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_A2;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_A3;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_A4;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_A5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_A6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_AO5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_AO6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_AQ;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_A_CY;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_A_XOR;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_B;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_B1;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_B2;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_B3;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_B4;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_B5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_B6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_BO5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_BO6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_BQ;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_B_CY;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_B_XOR;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_C;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_C1;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_C2;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_C3;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_C4;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_C5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_C6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_CLK;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_CO5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_CO6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_CQ;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_C_CY;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_C_XOR;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_D;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_D1;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_D2;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_D3;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_D4;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_D5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_D6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_DO5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_DO6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_D_CY;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_D_XOR;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_A;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_A1;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_A2;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_A3;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_A4;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_A5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_A6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_AO5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_AO6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_AQ;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_A_CY;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_A_XOR;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_B;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_B1;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_B2;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_B3;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_B4;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_B5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_B6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_BO5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_BO6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_BQ;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_B_CY;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_B_XOR;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_C;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_C1;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_C2;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_C3;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_C4;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_C5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_C5Q;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_C6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_CLK;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_CMUX;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_CO5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_CO6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_CQ;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_C_CY;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_C_XOR;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_D;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_D1;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_D2;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_D3;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_D4;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_D5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_D6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_DO5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_DO6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_DQ;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_D_CY;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_D_XOR;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_A;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_A1;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_A2;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_A3;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_A4;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_A5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_A5Q;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_A6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_AMUX;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_AO5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_AO6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_AQ;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_A_CY;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_A_XOR;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_B;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_B1;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_B2;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_B3;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_B4;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_B5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_B6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_BO5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_BO6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_BQ;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_B_CY;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_B_XOR;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_C;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_C1;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_C2;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_C3;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_C4;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_C5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_C6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_CLK;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_CO5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_CO6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_CQ;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_C_CY;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_C_XOR;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_D;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_D1;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_D2;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_D3;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_D4;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_D5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_D6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_DO5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_DO6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_D_CY;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_D_XOR;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_A;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_A1;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_A2;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_A3;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_A4;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_A5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_A5Q;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_A6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_AMUX;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_AO5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_AO6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_AQ;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_AX;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_A_CY;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_A_XOR;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_B;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_B1;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_B2;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_B3;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_B4;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_B5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_B5Q;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_B6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_BMUX;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_BO5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_BO6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_BQ;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_BX;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_B_CY;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_B_XOR;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_C;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_C1;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_C2;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_C3;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_C4;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_C5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_C5Q;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_C6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_CLK;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_CMUX;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_CO5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_CO6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_CQ;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_C_CY;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_C_XOR;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_D;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_D1;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_D2;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_D3;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_D4;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_D5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_D5Q;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_D6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_DMUX;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_DO5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_DO6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_DQ;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_D_CY;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_D_XOR;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_A;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_A1;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_A2;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_A3;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_A4;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_A5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_A5Q;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_A6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_AMUX;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_AO5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_AO6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_AQ;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_A_CY;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_A_XOR;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_B;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_B1;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_B2;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_B3;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_B4;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_B5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_B5Q;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_B6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_BMUX;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_BO5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_BO6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_BQ;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_B_CY;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_B_XOR;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_C;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_C1;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_C2;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_C3;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_C4;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_C5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_C6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_CLK;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_CO5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_CO6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_CQ;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_C_CY;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_C_XOR;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_D;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_D1;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_D2;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_D3;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_D4;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_D5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_D6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_DO5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_DO6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_D_CY;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_D_XOR;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_A;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_A1;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_A2;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_A3;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_A4;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_A5;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_A5Q;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_A6;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_AMUX;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_AO5;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_AO6;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_AQ;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_AX;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_A_CY;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_A_XOR;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_B;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_B1;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_B2;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_B3;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_B4;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_B5;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_B6;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_BMUX;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_BO5;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_BO6;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_B_CY;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_B_XOR;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_C;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_C1;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_C2;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_C3;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_C4;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_C5;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_C6;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_CLK;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_CO5;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_CO6;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_CQ;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_C_CY;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_C_XOR;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_D;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_D1;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_D2;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_D3;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_D4;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_D5;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_D6;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_DMUX;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_DO5;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_DO6;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_D_CY;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_D_XOR;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_A;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_A1;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_A2;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_A3;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_A4;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_A5;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_A6;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_AO5;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_AO6;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_AQ;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_A_CY;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_A_XOR;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_B;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_B1;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_B2;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_B3;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_B4;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_B5;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_B6;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_BO5;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_BO6;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_BQ;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_B_CY;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_B_XOR;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_C;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_C1;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_C2;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_C3;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_C4;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_C5;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_C6;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_CLK;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_CO5;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_CO6;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_C_CY;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_C_XOR;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_D;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_D1;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_D2;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_D3;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_D4;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_D5;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_D6;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_DO5;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_DO6;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_D_CY;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_D_XOR;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_A;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_A1;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_A2;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_A3;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_A4;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_A5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_A6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_AMUX;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_AO5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_AO6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_A_CY;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_A_XOR;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_B;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_B1;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_B2;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_B3;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_B4;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_B5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_B6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_BO5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_BO6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_BQ;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_B_CY;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_B_XOR;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_C;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_C1;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_C2;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_C3;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_C4;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_C5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_C6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_CLK;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_CO5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_CO6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_CQ;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_C_CY;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_C_XOR;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_D;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_D1;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_D2;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_D3;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_D4;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_D5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_D6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_DO5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_DO6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_D_CY;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_D_XOR;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_A;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_A1;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_A2;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_A3;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_A4;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_A5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_A6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_AO5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_AO6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_AQ;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_A_CY;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_A_XOR;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_B;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_B1;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_B2;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_B3;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_B4;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_B5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_B6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_BO5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_BO6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_BQ;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_B_CY;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_B_XOR;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_C;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_C1;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_C2;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_C3;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_C4;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_C5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_C6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_CLK;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_CMUX;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_CO5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_CO6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_C_CY;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_C_XOR;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_D;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_D1;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_D2;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_D3;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_D4;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_D5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_D6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_DO5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_DO6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_D_CY;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_D_XOR;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_A;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_A1;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_A2;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_A3;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_A4;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_A5;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_A6;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_AMUX;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_AO5;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_AO6;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_AQ;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_AX;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_A_CY;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_A_XOR;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_B;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_B1;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_B2;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_B3;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_B4;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_B5;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_B6;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_BMUX;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_BO5;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_BO6;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_B_CY;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_B_XOR;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_C;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_C1;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_C2;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_C3;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_C4;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_C5;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_C6;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_CE;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_CLK;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_CO5;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_CO6;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_C_CY;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_C_XOR;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_D;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_D1;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_D2;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_D3;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_D4;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_D5;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_D6;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_DO5;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_DO6;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_D_CY;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_D_XOR;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_SR;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_A;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_A1;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_A2;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_A3;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_A4;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_A5;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_A5Q;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_A6;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_AMUX;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_AO5;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_AO6;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_AQ;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_AX;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_A_CY;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_A_XOR;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_B;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_B1;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_B2;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_B3;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_B4;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_B5;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_B6;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_BO5;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_BO6;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_BQ;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_B_CY;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_B_XOR;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_C;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_C1;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_C2;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_C3;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_C4;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_C5;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_C6;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_CLK;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_CMUX;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_CO5;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_CO6;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_C_CY;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_C_XOR;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_D;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_D1;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_D2;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_D3;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_D4;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_D5;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_D6;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_DO5;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_DO6;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_DQ;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_D_CY;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_D_XOR;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_A;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_A1;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_A2;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_A3;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_A4;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_A5;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_A5Q;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_A6;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_AMUX;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_AO5;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_AO6;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_AQ;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_AX;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_A_CY;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_A_XOR;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_B;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_B1;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_B2;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_B3;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_B4;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_B5;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_B5Q;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_B6;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_BMUX;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_BO5;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_BO6;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_BQ;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_BX;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_B_CY;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_B_XOR;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_C;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_C1;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_C2;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_C3;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_C4;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_C5;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_C5Q;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_C6;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_CLK;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_CMUX;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_CO5;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_CO6;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_CQ;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_CX;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_C_CY;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_C_XOR;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_D;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_D1;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_D2;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_D3;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_D4;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_D5;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_D6;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_DO5;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_DO6;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_DQ;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_D_CY;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_D_XOR;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_A;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_A1;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_A2;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_A3;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_A4;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_A5;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_A5Q;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_A6;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_AMUX;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_AO5;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_AO6;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_AQ;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_AX;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_A_CY;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_A_XOR;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_B;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_B1;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_B2;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_B3;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_B4;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_B5;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_B6;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_BO5;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_BO6;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_BQ;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_B_CY;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_B_XOR;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_C;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_C1;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_C2;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_C3;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_C4;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_C5;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_C6;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_CLK;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_CO5;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_CO6;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_CQ;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_C_CY;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_C_XOR;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_D;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_D1;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_D2;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_D3;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_D4;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_D5;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_D6;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_DMUX;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_DO5;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_DO6;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_D_CY;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_D_XOR;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_A;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_A1;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_A2;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_A3;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_A4;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_A5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_A6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_AO5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_AO6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_AQ;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_A_CY;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_A_XOR;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_B;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_B1;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_B2;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_B3;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_B4;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_B5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_B6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_BO5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_BO6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_BQ;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_B_CY;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_B_XOR;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_C;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_C1;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_C2;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_C3;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_C4;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_C5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_C6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_CLK;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_CO5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_CO6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_CQ;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_C_CY;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_C_XOR;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_D;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_D1;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_D2;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_D3;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_D4;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_D5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_D6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_DO5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_DO6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_DQ;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_D_CY;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_D_XOR;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_A;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_A1;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_A2;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_A3;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_A4;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_A5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_A6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_AO5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_AO6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_AQ;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_A_CY;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_A_XOR;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_B;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_B1;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_B2;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_B3;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_B4;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_B5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_B6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_BO5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_BO6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_BQ;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_B_CY;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_B_XOR;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_C;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_C1;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_C2;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_C3;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_C4;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_C5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_C6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_CLK;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_CO5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_CO6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_CQ;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_C_CY;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_C_XOR;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_D;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_D1;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_D2;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_D3;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_D4;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_D5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_D6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_DO5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_DO6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_DQ;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_D_CY;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_D_XOR;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_A;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_A1;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_A2;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_A3;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_A4;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_A5;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_A6;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_AO5;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_AO6;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_AQ;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_A_CY;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_A_XOR;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_B;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_B1;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_B2;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_B3;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_B4;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_B5;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_B6;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_BO5;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_BO6;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_BQ;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_B_CY;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_B_XOR;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_C;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_C1;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_C2;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_C3;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_C4;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_C5;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_C6;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_CLK;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_CMUX;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_CO5;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_CO6;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_C_CY;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_C_XOR;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_D;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_D1;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_D2;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_D3;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_D4;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_D5;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_D5Q;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_D6;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_DMUX;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_DO5;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_DO6;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_DQ;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_D_CY;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_D_XOR;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_A;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_A1;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_A2;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_A3;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_A4;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_A5;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_A6;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_AO5;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_AO6;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_AQ;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_A_CY;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_A_XOR;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_B;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_B1;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_B2;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_B3;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_B4;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_B5;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_B6;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_BO5;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_BO6;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_BQ;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_B_CY;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_B_XOR;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_C;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_C1;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_C2;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_C3;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_C4;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_C5;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_C6;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_CLK;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_CMUX;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_CO5;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_CO6;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_C_CY;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_C_XOR;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_D;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_D1;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_D2;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_D3;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_D4;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_D5;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_D6;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_DO5;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_DO6;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_D_CY;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_D_XOR;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_A;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_A1;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_A2;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_A3;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_A4;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_A5;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_A6;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_AO5;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_AO6;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_AQ;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_A_CY;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_A_XOR;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_B;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_B1;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_B2;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_B3;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_B4;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_B5;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_B6;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_BO5;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_BO6;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_BQ;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_B_CY;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_B_XOR;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_C;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_C1;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_C2;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_C3;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_C4;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_C5;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_C6;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_CLK;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_CO5;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_CO6;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_CQ;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_C_CY;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_C_XOR;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_D;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_D1;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_D2;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_D3;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_D4;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_D5;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_D6;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_DO5;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_DO6;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_DQ;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_D_CY;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_D_XOR;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_A;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_A1;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_A2;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_A3;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_A4;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_A5;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_A6;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_AO5;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_AO6;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_AQ;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_A_CY;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_A_XOR;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_B;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_B1;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_B2;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_B3;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_B4;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_B5;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_B6;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_BO5;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_BO6;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_BQ;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_B_CY;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_B_XOR;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_C;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_C1;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_C2;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_C3;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_C4;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_C5;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_C6;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_CLK;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_CO5;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_CO6;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_CQ;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_C_CY;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_C_XOR;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_D;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_D1;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_D2;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_D3;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_D4;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_D5;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_D6;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_DO5;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_DO6;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_DQ;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_D_CY;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_D_XOR;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_A;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_A1;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_A2;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_A3;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_A4;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_A5;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_A6;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_AO5;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_AO6;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_AQ;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_A_CY;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_A_XOR;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_B;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_B1;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_B2;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_B3;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_B4;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_B5;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_B6;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_BO5;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_BO6;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_BQ;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_B_CY;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_B_XOR;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_C;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_C1;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_C2;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_C3;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_C4;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_C5;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_C6;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_CLK;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_CO5;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_CO6;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_CQ;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_C_CY;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_C_XOR;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_D;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_D1;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_D2;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_D3;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_D4;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_D5;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_D6;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_DO5;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_DO6;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_DQ;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_D_CY;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_D_XOR;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_A;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_A1;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_A2;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_A3;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_A4;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_A5;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_A6;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_AO5;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_AO6;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_AQ;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_A_CY;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_A_XOR;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_B;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_B1;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_B2;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_B3;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_B4;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_B5;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_B6;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_BO5;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_BO6;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_BQ;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_B_CY;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_B_XOR;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_C;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_C1;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_C2;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_C3;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_C4;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_C5;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_C6;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_CLK;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_CMUX;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_CO5;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_CO6;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_C_CY;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_C_XOR;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_D;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_D1;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_D2;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_D3;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_D4;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_D5;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_D6;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_DO5;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_DO6;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_D_CY;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_D_XOR;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_A;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_A1;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_A2;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_A3;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_A4;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_A5;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_A6;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_AO5;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_AO6;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_AQ;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_A_CY;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_A_XOR;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_B;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_B1;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_B2;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_B3;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_B4;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_B5;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_B6;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_BO5;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_BO6;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_B_CY;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_B_XOR;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_C;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_C1;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_C2;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_C3;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_C4;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_C5;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_C6;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_CLK;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_CO5;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_CO6;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_C_CY;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_C_XOR;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_D;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_D1;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_D2;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_D3;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_D4;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_D5;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_D6;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_DO5;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_DO6;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_D_CY;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_D_XOR;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_A;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_A1;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_A2;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_A3;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_A4;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_A5;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_A6;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_AO5;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_AO6;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_AQ;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_A_CY;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_A_XOR;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_B;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_B1;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_B2;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_B3;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_B4;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_B5;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_B6;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_BO5;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_BO6;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_BQ;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_B_CY;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_B_XOR;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_C;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_C1;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_C2;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_C3;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_C4;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_C5;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_C6;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_CLK;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_CO5;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_CO6;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_CQ;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_C_CY;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_C_XOR;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_D;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_D1;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_D2;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_D3;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_D4;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_D5;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_D6;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_DO5;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_DO6;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_D_CY;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_D_XOR;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X12Y156_A;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X12Y156_A1;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X12Y156_A2;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X12Y156_A3;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X12Y156_A4;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X12Y156_A5;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X12Y156_A6;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X12Y156_AMUX;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X12Y156_AO5;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X12Y156_AO6;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X12Y156_A_CY;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X12Y156_A_XOR;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X12Y156_B;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X12Y156_B1;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X12Y156_B2;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X12Y156_B3;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X12Y156_B4;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X12Y156_B5;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X12Y156_B6;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X12Y156_BO5;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X12Y156_BO6;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X12Y156_B_CY;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X12Y156_B_XOR;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X12Y156_C;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X12Y156_C1;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X12Y156_C2;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X12Y156_C3;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X12Y156_C4;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X12Y156_C5;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X12Y156_C6;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X12Y156_CO5;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X12Y156_CO6;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X12Y156_C_CY;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X12Y156_C_XOR;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X12Y156_D;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X12Y156_D1;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X12Y156_D2;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X12Y156_D3;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X12Y156_D4;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X12Y156_D5;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X12Y156_D6;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X12Y156_DO5;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X12Y156_DO6;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X12Y156_D_CY;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X12Y156_D_XOR;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X13Y156_A;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X13Y156_A1;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X13Y156_A2;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X13Y156_A3;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X13Y156_A4;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X13Y156_A5;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X13Y156_A6;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X13Y156_AO5;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X13Y156_AO6;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X13Y156_A_CY;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X13Y156_A_XOR;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X13Y156_B;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X13Y156_B1;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X13Y156_B2;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X13Y156_B3;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X13Y156_B4;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X13Y156_B5;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X13Y156_B6;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X13Y156_BO5;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X13Y156_BO6;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X13Y156_B_CY;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X13Y156_B_XOR;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X13Y156_C;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X13Y156_C1;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X13Y156_C2;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X13Y156_C3;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X13Y156_C4;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X13Y156_C5;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X13Y156_C6;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X13Y156_CO5;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X13Y156_CO6;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X13Y156_C_CY;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X13Y156_C_XOR;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X13Y156_D;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X13Y156_D1;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X13Y156_D2;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X13Y156_D3;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X13Y156_D4;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X13Y156_D5;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X13Y156_D6;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X13Y156_DO5;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X13Y156_DO6;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X13Y156_D_CY;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X13Y156_D_XOR;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_A;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_A1;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_A2;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_A3;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_A4;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_A5;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_A6;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_AMUX;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_AO5;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_AO6;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_AQ;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_A_CY;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_A_XOR;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_B;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_B1;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_B2;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_B3;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_B4;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_B5;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_B6;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_BO5;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_BO6;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_BQ;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_B_CY;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_B_XOR;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_C;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_C1;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_C2;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_C3;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_C4;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_C5;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_C6;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_CLK;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_CO5;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_CO6;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_CQ;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_C_CY;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_C_XOR;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_D;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_D1;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_D2;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_D3;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_D4;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_D5;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_D6;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_DMUX;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_DO5;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_DO6;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_D_CY;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_D_XOR;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_A;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_A1;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_A2;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_A3;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_A4;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_A5;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_A6;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_AO5;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_AO6;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_A_CY;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_A_XOR;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_B;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_B1;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_B2;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_B3;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_B4;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_B5;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_B6;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_BO5;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_BO6;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_B_CY;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_B_XOR;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_C;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_C1;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_C2;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_C3;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_C4;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_C5;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_C6;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_CO5;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_CO6;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_C_CY;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_C_XOR;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_D;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_D1;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_D2;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_D3;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_D4;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_D5;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_D6;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_DO5;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_DO6;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_D_CY;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_D_XOR;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_A;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_A1;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_A2;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_A3;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_A4;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_A5;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_A6;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_AO5;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_AO6;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_AQ;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_A_CY;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_A_XOR;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_B;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_B1;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_B2;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_B3;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_B4;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_B5;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_B6;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_BO5;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_BO6;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_BQ;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_B_CY;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_B_XOR;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_C;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_C1;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_C2;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_C3;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_C4;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_C5;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_C6;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_CLK;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_CMUX;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_CO5;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_CO6;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_C_CY;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_C_XOR;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_D;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_D1;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_D2;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_D3;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_D4;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_D5;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_D6;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_DO5;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_DO6;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_D_CY;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_D_XOR;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_A;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_A1;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_A2;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_A3;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_A4;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_A5;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_A6;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_AO5;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_A_CY;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_A_XOR;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_B;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_B1;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_B2;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_B3;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_B4;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_B5;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_B6;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_BO5;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_BO6;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_B_CY;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_B_XOR;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_C;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_C1;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_C2;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_C3;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_C4;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_C5;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_C6;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_CO5;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_CO6;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_C_CY;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_C_XOR;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_D;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_D1;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_D2;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_D3;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_D4;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_D5;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_D6;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_DO5;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_DO6;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_D_CY;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_D_XOR;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_A;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_A1;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_A2;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_A3;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_A4;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_A5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_A6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_AO5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_AO6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_AQ;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_A_CY;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_A_XOR;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_B;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_B1;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_B2;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_B3;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_B4;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_B5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_B6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_BO5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_BO6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_B_CY;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_B_XOR;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_C;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_C1;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_C2;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_C3;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_C4;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_C5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_C6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_CLK;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_CO5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_CO6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_C_CY;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_C_XOR;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_D;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_D1;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_D2;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_D3;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_D4;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_D5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_D6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_DO5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_DO6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_D_CY;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_D_XOR;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_A;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_A1;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_A2;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_A3;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_A4;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_A5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_A6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_AO5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_AO6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_A_CY;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_A_XOR;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_B;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_B1;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_B2;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_B3;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_B4;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_B5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_B6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_BO5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_BO6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_B_CY;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_B_XOR;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_C;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_C1;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_C2;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_C3;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_C4;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_C5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_C6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_CO5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_CO6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_C_CY;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_C_XOR;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_D;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_D1;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_D2;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_D3;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_D4;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_D5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_D6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_DO5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_DO6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_D_CY;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_D_XOR;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_A;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_A1;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_A2;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_A3;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_A4;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_A5;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_A6;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_AO5;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_AO6;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_AQ;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_A_CY;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_A_XOR;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_B;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_B1;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_B2;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_B3;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_B4;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_B5;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_B6;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_BO5;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_BO6;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_B_CY;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_B_XOR;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_C;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_C1;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_C2;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_C3;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_C4;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_C5;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_C6;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_CLK;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_CO5;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_CO6;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_C_CY;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_C_XOR;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_D;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_D1;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_D2;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_D3;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_D4;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_D5;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_D6;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_DO5;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_DO6;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_D_CY;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_D_XOR;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_A;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_A1;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_A2;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_A3;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_A4;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_A5;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_A6;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_AO5;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_AO6;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_A_CY;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_A_XOR;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_B;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_B1;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_B2;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_B3;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_B4;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_B5;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_B6;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_BO5;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_BO6;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_B_CY;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_B_XOR;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_C;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_C1;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_C2;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_C3;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_C4;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_C5;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_C6;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_CO5;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_CO6;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_C_CY;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_C_XOR;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_D;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_D1;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_D2;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_D3;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_D4;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_D5;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_D6;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_DO5;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_DO6;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_D_CY;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_D_XOR;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_A;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_A1;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_A2;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_A3;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_A4;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_A5;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_A6;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_AO5;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_AO6;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_AQ;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_A_CY;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_A_XOR;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_B;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_B1;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_B2;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_B3;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_B4;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_B5;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_B6;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_BO5;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_BO6;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_BQ;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_B_CY;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_B_XOR;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_C;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_C1;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_C2;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_C3;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_C4;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_C5;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_C6;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_CLK;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_CO5;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_CO6;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_C_CY;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_C_XOR;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_D;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_D1;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_D2;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_D3;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_D4;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_D5;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_D6;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_DO5;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_DO6;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_D_CY;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_D_XOR;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_A;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_A1;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_A2;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_A3;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_A4;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_A5;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_A6;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_AO5;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_AO6;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_A_CY;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_A_XOR;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_B;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_B1;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_B2;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_B3;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_B4;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_B5;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_B6;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_BO5;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_BO6;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_B_CY;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_B_XOR;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_C;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_C1;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_C2;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_C3;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_C4;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_C5;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_C6;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_CO5;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_CO6;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_C_CY;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_C_XOR;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_D;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_D1;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_D2;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_D3;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_D4;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_D5;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_D6;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_DO5;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_DO6;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_D_CY;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_D_XOR;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_A;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_A1;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_A2;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_A3;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_A4;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_A5;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_A6;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_AO5;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_AO6;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_AQ;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_A_CY;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_A_XOR;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_B;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_B1;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_B2;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_B3;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_B4;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_B5;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_B6;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_BO5;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_BO6;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_B_CY;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_B_XOR;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_C;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_C1;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_C2;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_C3;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_C4;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_C5;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_C6;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_CLK;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_CO5;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_CO6;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_C_CY;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_C_XOR;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_D;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_D1;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_D2;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_D3;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_D4;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_D5;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_D6;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_DO5;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_DO6;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_D_CY;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_D_XOR;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_A;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_A1;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_A2;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_A3;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_A4;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_A5;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_A6;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_AO5;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_AO6;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_AQ;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_A_CY;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_A_XOR;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_B;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_B1;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_B2;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_B3;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_B4;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_B5;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_B6;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_BO5;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_BO6;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_BQ;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_B_CY;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_B_XOR;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_C;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_C1;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_C2;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_C3;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_C4;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_C5;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_C6;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_CLK;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_CO5;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_CO6;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_CQ;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_C_CY;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_C_XOR;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_D;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_D1;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_D2;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_D3;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_D4;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_D5;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_D6;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_DO5;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_DO6;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_D_CY;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_D_XOR;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_A;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_A1;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_A2;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_A3;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_A4;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_A5;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_A6;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_AO5;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_AO6;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_AQ;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_A_CY;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_A_XOR;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_B;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_B1;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_B2;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_B3;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_B4;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_B5;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_B6;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_BO5;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_BO6;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_BQ;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_B_CY;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_B_XOR;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_C;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_C1;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_C2;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_C3;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_C4;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_C5;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_C6;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_CLK;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_CO5;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_CO6;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_CQ;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_C_CY;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_C_XOR;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_D;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_D1;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_D2;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_D3;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_D4;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_D5;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_D6;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_DMUX;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_DO5;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_DO6;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_D_CY;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_D_XOR;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_A;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_A1;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_A2;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_A3;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_A4;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_A5;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_A6;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_AO5;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_AO6;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_A_CY;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_A_XOR;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_B;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_B1;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_B2;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_B3;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_B4;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_B5;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_B6;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_BO5;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_BO6;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_B_CY;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_B_XOR;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_C;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_C1;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_C2;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_C3;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_C4;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_C5;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_C6;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_CO5;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_CO6;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_C_CY;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_C_XOR;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_D;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_D1;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_D2;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_D3;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_D4;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_D5;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_D6;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_DO5;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_DO6;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_D_CY;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_D_XOR;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_A;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_A1;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_A2;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_A3;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_A4;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_A5;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_A6;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_AO5;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_AO6;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_AQ;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_A_CY;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_A_XOR;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_B;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_B1;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_B2;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_B3;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_B4;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_B5;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_B6;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_BO5;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_BO6;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_BQ;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_B_CY;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_B_XOR;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_C;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_C1;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_C2;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_C3;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_C4;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_C5;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_C6;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_CLK;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_CO5;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_CO6;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_CQ;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_C_CY;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_C_XOR;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_D;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_D1;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_D2;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_D3;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_D4;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_D5;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_D6;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_DMUX;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_DO5;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_DO6;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_D_CY;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_D_XOR;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_A;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_A1;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_A2;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_A3;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_A4;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_A5;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_A6;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_AO5;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_AO6;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_A_CY;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_A_XOR;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_B;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_B1;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_B2;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_B3;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_B4;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_B5;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_B6;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_BO5;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_BO6;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_B_CY;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_B_XOR;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_C;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_C1;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_C2;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_C3;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_C4;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_C5;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_C6;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_CO5;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_CO6;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_C_CY;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_C_XOR;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_D;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_D1;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_D2;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_D3;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_D4;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_D5;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_D6;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_DO5;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_DO6;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_D_CY;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_D_XOR;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_A;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_A1;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_A2;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_A3;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_A4;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_A5;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_A6;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_AO5;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_AO6;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_AQ;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_A_CY;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_A_XOR;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_B;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_B1;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_B2;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_B3;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_B4;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_B5;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_B6;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_BO5;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_BO6;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_BQ;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_B_CY;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_B_XOR;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_C;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_C1;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_C2;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_C3;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_C4;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_C5;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_C6;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_CLK;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_CO5;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_CO6;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_C_CY;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_C_XOR;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_D;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_D1;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_D2;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_D3;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_D4;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_D5;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_D6;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_DO5;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_DO6;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_D_CY;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_D_XOR;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_A;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_A1;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_A2;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_A3;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_A4;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_A5;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_A6;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_AO5;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_AO6;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_AQ;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_A_CY;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_A_XOR;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_B;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_B1;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_B2;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_B3;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_B4;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_B5;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_B6;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_BO5;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_BO6;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_BQ;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_B_CY;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_B_XOR;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_C;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_C1;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_C2;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_C3;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_C4;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_C5;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_C6;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_CLK;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_CO5;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_CO6;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_CQ;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_C_CY;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_C_XOR;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_D;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_D1;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_D2;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_D3;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_D4;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_D5;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_D6;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_DO5;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_DO6;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_D_CY;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_D_XOR;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_A;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_A1;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_A2;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_A3;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_A4;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_A5;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_A6;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_AO5;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_AO6;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_AQ;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_A_CY;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_A_XOR;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_B;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_B1;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_B2;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_B3;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_B4;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_B5;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_B6;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_BO5;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_BO6;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_B_CY;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_B_XOR;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_C;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_C1;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_C2;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_C3;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_C4;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_C5;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_C6;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_CLK;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_CO5;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_CO6;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_C_CY;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_C_XOR;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_D;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_D1;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_D2;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_D3;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_D4;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_D5;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_D6;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_DO5;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_DO6;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_D_CY;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_D_XOR;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_A;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_A1;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_A2;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_A3;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_A4;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_A5;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_A6;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_AO5;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_AO6;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_AQ;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_A_CY;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_A_XOR;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_B;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_B1;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_B2;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_B3;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_B4;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_B5;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_B6;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_BO5;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_BO6;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_B_CY;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_B_XOR;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_C;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_C1;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_C2;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_C3;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_C4;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_C5;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_C6;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_CLK;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_CO5;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_CO6;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_C_CY;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_C_XOR;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_D;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_D1;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_D2;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_D3;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_D4;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_D5;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_D6;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_DO5;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_DO6;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_D_CY;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_D_XOR;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_A;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_A1;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_A2;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_A3;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_A4;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_A5;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_A6;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_AO5;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_AO6;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_AQ;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_A_CY;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_A_XOR;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_B;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_B1;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_B2;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_B3;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_B4;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_B5;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_B6;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_BMUX;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_BO5;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_BO6;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_B_CY;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_B_XOR;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_C;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_C1;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_C2;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_C3;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_C4;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_C5;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_C6;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_CLK;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_CO5;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_CO6;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_C_CY;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_C_XOR;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_D;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_D1;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_D2;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_D3;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_D4;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_D5;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_D6;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_DO5;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_DO6;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_D_CY;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_D_XOR;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_A;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_A1;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_A2;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_A3;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_A4;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_A5;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_A6;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_AO5;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_AO6;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_A_CY;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_A_XOR;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_B;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_B1;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_B2;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_B3;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_B4;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_B5;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_B6;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_BO5;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_BO6;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_B_CY;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_B_XOR;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_C;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_C1;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_C2;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_C3;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_C4;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_C5;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_C6;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_CO5;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_CO6;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_C_CY;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_C_XOR;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_D;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_D1;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_D2;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_D3;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_D4;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_D5;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_D6;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_DO5;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_DO6;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_D_CY;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_D_XOR;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X16Y155_A;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X16Y155_A1;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X16Y155_A2;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X16Y155_A3;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X16Y155_A4;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X16Y155_A5;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X16Y155_A6;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X16Y155_AO5;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X16Y155_AO6;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X16Y155_A_CY;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X16Y155_A_XOR;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X16Y155_B;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X16Y155_B1;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X16Y155_B2;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X16Y155_B3;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X16Y155_B4;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X16Y155_B5;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X16Y155_B6;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X16Y155_BO5;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X16Y155_BO6;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X16Y155_B_CY;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X16Y155_B_XOR;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X16Y155_C;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X16Y155_C1;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X16Y155_C2;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X16Y155_C3;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X16Y155_C4;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X16Y155_C5;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X16Y155_C6;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X16Y155_CO5;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X16Y155_CO6;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X16Y155_C_CY;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X16Y155_C_XOR;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X16Y155_D;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X16Y155_D1;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X16Y155_D2;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X16Y155_D3;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X16Y155_D4;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X16Y155_D5;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X16Y155_D6;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X16Y155_DO5;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X16Y155_DO6;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X16Y155_D_CY;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X16Y155_D_XOR;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X17Y155_A;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X17Y155_A1;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X17Y155_A2;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X17Y155_A3;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X17Y155_A4;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X17Y155_A5;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X17Y155_A6;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X17Y155_AO5;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X17Y155_AO6;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X17Y155_AQ;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X17Y155_A_CY;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X17Y155_A_XOR;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X17Y155_B;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X17Y155_B1;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X17Y155_B2;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X17Y155_B3;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X17Y155_B4;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X17Y155_B5;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X17Y155_B6;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X17Y155_BO5;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X17Y155_BO6;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X17Y155_B_CY;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X17Y155_B_XOR;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X17Y155_C;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X17Y155_C1;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X17Y155_C2;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X17Y155_C3;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X17Y155_C4;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X17Y155_C5;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X17Y155_C6;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X17Y155_CLK;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X17Y155_CO5;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X17Y155_CO6;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X17Y155_C_CY;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X17Y155_C_XOR;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X17Y155_D;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X17Y155_D1;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X17Y155_D2;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X17Y155_D3;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X17Y155_D4;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X17Y155_D5;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X17Y155_D6;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X17Y155_DO5;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X17Y155_DO6;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X17Y155_D_CY;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X17Y155_D_XOR;
  wire [0:0] CLBLM_L_X16Y158_SLICE_X22Y158_A;
  wire [0:0] CLBLM_L_X16Y158_SLICE_X22Y158_A1;
  wire [0:0] CLBLM_L_X16Y158_SLICE_X22Y158_A2;
  wire [0:0] CLBLM_L_X16Y158_SLICE_X22Y158_A3;
  wire [0:0] CLBLM_L_X16Y158_SLICE_X22Y158_A4;
  wire [0:0] CLBLM_L_X16Y158_SLICE_X22Y158_A5;
  wire [0:0] CLBLM_L_X16Y158_SLICE_X22Y158_A6;
  wire [0:0] CLBLM_L_X16Y158_SLICE_X22Y158_AMUX;
  wire [0:0] CLBLM_L_X16Y158_SLICE_X22Y158_AO5;
  wire [0:0] CLBLM_L_X16Y158_SLICE_X22Y158_AO6;
  wire [0:0] CLBLM_L_X16Y158_SLICE_X22Y158_A_CY;
  wire [0:0] CLBLM_L_X16Y158_SLICE_X22Y158_A_XOR;
  wire [0:0] CLBLM_L_X16Y158_SLICE_X22Y158_B;
  wire [0:0] CLBLM_L_X16Y158_SLICE_X22Y158_B1;
  wire [0:0] CLBLM_L_X16Y158_SLICE_X22Y158_B2;
  wire [0:0] CLBLM_L_X16Y158_SLICE_X22Y158_B3;
  wire [0:0] CLBLM_L_X16Y158_SLICE_X22Y158_B4;
  wire [0:0] CLBLM_L_X16Y158_SLICE_X22Y158_B5;
  wire [0:0] CLBLM_L_X16Y158_SLICE_X22Y158_B6;
  wire [0:0] CLBLM_L_X16Y158_SLICE_X22Y158_BO5;
  wire [0:0] CLBLM_L_X16Y158_SLICE_X22Y158_BO6;
  wire [0:0] CLBLM_L_X16Y158_SLICE_X22Y158_B_CY;
  wire [0:0] CLBLM_L_X16Y158_SLICE_X22Y158_B_XOR;
  wire [0:0] CLBLM_L_X16Y158_SLICE_X22Y158_C;
  wire [0:0] CLBLM_L_X16Y158_SLICE_X22Y158_C1;
  wire [0:0] CLBLM_L_X16Y158_SLICE_X22Y158_C2;
  wire [0:0] CLBLM_L_X16Y158_SLICE_X22Y158_C3;
  wire [0:0] CLBLM_L_X16Y158_SLICE_X22Y158_C4;
  wire [0:0] CLBLM_L_X16Y158_SLICE_X22Y158_C5;
  wire [0:0] CLBLM_L_X16Y158_SLICE_X22Y158_C6;
  wire [0:0] CLBLM_L_X16Y158_SLICE_X22Y158_CO5;
  wire [0:0] CLBLM_L_X16Y158_SLICE_X22Y158_CO6;
  wire [0:0] CLBLM_L_X16Y158_SLICE_X22Y158_C_CY;
  wire [0:0] CLBLM_L_X16Y158_SLICE_X22Y158_C_XOR;
  wire [0:0] CLBLM_L_X16Y158_SLICE_X22Y158_D;
  wire [0:0] CLBLM_L_X16Y158_SLICE_X22Y158_D1;
  wire [0:0] CLBLM_L_X16Y158_SLICE_X22Y158_D2;
  wire [0:0] CLBLM_L_X16Y158_SLICE_X22Y158_D3;
  wire [0:0] CLBLM_L_X16Y158_SLICE_X22Y158_D4;
  wire [0:0] CLBLM_L_X16Y158_SLICE_X22Y158_D5;
  wire [0:0] CLBLM_L_X16Y158_SLICE_X22Y158_D6;
  wire [0:0] CLBLM_L_X16Y158_SLICE_X22Y158_DO5;
  wire [0:0] CLBLM_L_X16Y158_SLICE_X22Y158_DO6;
  wire [0:0] CLBLM_L_X16Y158_SLICE_X22Y158_D_CY;
  wire [0:0] CLBLM_L_X16Y158_SLICE_X22Y158_D_XOR;
  wire [0:0] CLBLM_L_X16Y158_SLICE_X23Y158_A;
  wire [0:0] CLBLM_L_X16Y158_SLICE_X23Y158_A1;
  wire [0:0] CLBLM_L_X16Y158_SLICE_X23Y158_A2;
  wire [0:0] CLBLM_L_X16Y158_SLICE_X23Y158_A3;
  wire [0:0] CLBLM_L_X16Y158_SLICE_X23Y158_A4;
  wire [0:0] CLBLM_L_X16Y158_SLICE_X23Y158_A5;
  wire [0:0] CLBLM_L_X16Y158_SLICE_X23Y158_A6;
  wire [0:0] CLBLM_L_X16Y158_SLICE_X23Y158_AO5;
  wire [0:0] CLBLM_L_X16Y158_SLICE_X23Y158_AO6;
  wire [0:0] CLBLM_L_X16Y158_SLICE_X23Y158_A_CY;
  wire [0:0] CLBLM_L_X16Y158_SLICE_X23Y158_A_XOR;
  wire [0:0] CLBLM_L_X16Y158_SLICE_X23Y158_B;
  wire [0:0] CLBLM_L_X16Y158_SLICE_X23Y158_B1;
  wire [0:0] CLBLM_L_X16Y158_SLICE_X23Y158_B2;
  wire [0:0] CLBLM_L_X16Y158_SLICE_X23Y158_B3;
  wire [0:0] CLBLM_L_X16Y158_SLICE_X23Y158_B4;
  wire [0:0] CLBLM_L_X16Y158_SLICE_X23Y158_B5;
  wire [0:0] CLBLM_L_X16Y158_SLICE_X23Y158_B6;
  wire [0:0] CLBLM_L_X16Y158_SLICE_X23Y158_BO5;
  wire [0:0] CLBLM_L_X16Y158_SLICE_X23Y158_BO6;
  wire [0:0] CLBLM_L_X16Y158_SLICE_X23Y158_B_CY;
  wire [0:0] CLBLM_L_X16Y158_SLICE_X23Y158_B_XOR;
  wire [0:0] CLBLM_L_X16Y158_SLICE_X23Y158_C;
  wire [0:0] CLBLM_L_X16Y158_SLICE_X23Y158_C1;
  wire [0:0] CLBLM_L_X16Y158_SLICE_X23Y158_C2;
  wire [0:0] CLBLM_L_X16Y158_SLICE_X23Y158_C3;
  wire [0:0] CLBLM_L_X16Y158_SLICE_X23Y158_C4;
  wire [0:0] CLBLM_L_X16Y158_SLICE_X23Y158_C5;
  wire [0:0] CLBLM_L_X16Y158_SLICE_X23Y158_C6;
  wire [0:0] CLBLM_L_X16Y158_SLICE_X23Y158_CO5;
  wire [0:0] CLBLM_L_X16Y158_SLICE_X23Y158_CO6;
  wire [0:0] CLBLM_L_X16Y158_SLICE_X23Y158_C_CY;
  wire [0:0] CLBLM_L_X16Y158_SLICE_X23Y158_C_XOR;
  wire [0:0] CLBLM_L_X16Y158_SLICE_X23Y158_D;
  wire [0:0] CLBLM_L_X16Y158_SLICE_X23Y158_D1;
  wire [0:0] CLBLM_L_X16Y158_SLICE_X23Y158_D2;
  wire [0:0] CLBLM_L_X16Y158_SLICE_X23Y158_D3;
  wire [0:0] CLBLM_L_X16Y158_SLICE_X23Y158_D4;
  wire [0:0] CLBLM_L_X16Y158_SLICE_X23Y158_D5;
  wire [0:0] CLBLM_L_X16Y158_SLICE_X23Y158_D6;
  wire [0:0] CLBLM_L_X16Y158_SLICE_X23Y158_DO5;
  wire [0:0] CLBLM_L_X16Y158_SLICE_X23Y158_DO6;
  wire [0:0] CLBLM_L_X16Y158_SLICE_X23Y158_D_CY;
  wire [0:0] CLBLM_L_X16Y158_SLICE_X23Y158_D_XOR;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_A;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_A1;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_A2;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_A3;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_A4;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_A5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_A5Q;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_A6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_AMUX;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_AO5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_AO6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_AQ;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_A_CY;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_A_XOR;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_B;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_B1;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_B2;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_B3;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_B4;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_B5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_B6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_BO5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_BO6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_B_CY;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_B_XOR;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_C;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_C1;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_C2;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_C3;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_C4;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_C5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_C6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_CLK;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_CO5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_CO6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_C_CY;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_C_XOR;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_D;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_D1;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_D2;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_D3;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_D4;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_D5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_D6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_DO5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_DO6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_D_CY;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_D_XOR;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_A;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_A1;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_A2;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_A3;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_A4;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_A5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_A6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_AO5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_AO6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_A_CY;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_A_XOR;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_B;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_B1;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_B2;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_B3;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_B4;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_B5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_B6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_BO5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_BO6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_B_CY;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_B_XOR;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_C;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_C1;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_C2;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_C3;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_C4;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_C5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_C6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_CO5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_CO6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_C_CY;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_C_XOR;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_D;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_D1;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_D2;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_D3;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_D4;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_D5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_D6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_DO5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_DO6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_D_CY;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_D_XOR;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_A;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_A1;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_A2;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_A3;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_A4;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_A5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_A6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_AO5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_AO6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_A_CY;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_A_XOR;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_B;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_B1;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_B2;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_B3;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_B4;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_B5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_B6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_BO5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_BO6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_BQ;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_B_CY;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_B_XOR;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_C;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_C1;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_C2;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_C3;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_C4;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_C5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_C6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_CLK;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_CO5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_CO6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_C_CY;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_C_XOR;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_D;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_D1;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_D2;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_D3;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_D4;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_D5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_D6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_DO5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_DO6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_D_CY;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_D_XOR;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_A;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_A1;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_A2;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_A3;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_A4;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_A5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_A6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_AO5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_AO6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_AQ;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_A_CY;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_A_XOR;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_B;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_B1;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_B2;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_B3;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_B4;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_B5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_B6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_BMUX;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_BO5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_BO6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_B_CY;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_B_XOR;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_C;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_C1;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_C2;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_C3;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_C4;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_C5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_C6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_CLK;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_CO5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_CO6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_C_CY;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_C_XOR;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_D;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_D1;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_D2;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_D3;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_D4;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_D5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_D6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_DO5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_DO6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_D_CY;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_D_XOR;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_A;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_A1;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_A2;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_A3;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_A4;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_A5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_A6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_AO5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_AO6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_AQ;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_A_CY;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_A_XOR;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_B;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_B1;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_B2;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_B3;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_B4;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_B5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_B6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_BO5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_BO6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_BQ;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_B_CY;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_B_XOR;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_C;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_C1;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_C2;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_C3;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_C4;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_C5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_C6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_CLK;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_CO5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_CO6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_CQ;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_C_CY;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_C_XOR;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_D;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_D1;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_D2;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_D3;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_D4;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_D5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_D6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_DO5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_DO6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_D_CY;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_D_XOR;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_A;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_A1;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_A2;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_A3;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_A4;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_A5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_A6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_AO5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_AO6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_AQ;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_A_CY;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_A_XOR;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_B;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_B1;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_B2;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_B3;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_B4;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_B5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_B6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_BO5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_BO6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_B_CY;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_B_XOR;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_C;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_C1;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_C2;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_C3;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_C4;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_C5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_C6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_CLK;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_CO5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_CO6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_C_CY;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_C_XOR;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_D;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_D1;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_D2;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_D3;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_D4;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_D5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_D6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_DO5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_DO6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_D_CY;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_D_XOR;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_A;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_A1;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_A2;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_A3;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_A4;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_A5;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_A5Q;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_A6;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_AMUX;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_AO5;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_AO6;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_AQ;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_AX;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_A_CY;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_A_XOR;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_B;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_B1;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_B2;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_B3;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_B4;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_B5;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_B6;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_BO5;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_BO6;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_BQ;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_B_CY;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_B_XOR;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_C;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_C1;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_C2;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_C3;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_C4;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_C5;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_C6;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_CLK;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_CMUX;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_CO5;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_CO6;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_C_CY;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_C_XOR;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_D;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_D1;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_D2;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_D3;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_D4;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_D5;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_D6;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_DO5;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_DO6;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_D_CY;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_D_XOR;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_A;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_A1;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_A2;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_A3;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_A4;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_A5;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_A5Q;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_A6;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_AMUX;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_AO5;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_AO6;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_AQ;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_A_CY;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_A_XOR;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_B;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_B1;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_B2;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_B3;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_B4;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_B5;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_B5Q;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_B6;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_BMUX;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_BO5;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_BO6;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_BQ;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_B_CY;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_B_XOR;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_C;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_C1;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_C2;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_C3;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_C4;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_C5;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_C6;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_CLK;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_CO5;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_CO6;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_CQ;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_C_CY;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_C_XOR;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_D;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_D1;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_D2;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_D3;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_D4;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_D5;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_D6;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_DO5;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_DO6;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_DQ;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_D_CY;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_D_XOR;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_A;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_A1;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_A2;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_A3;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_A4;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_A5;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_A6;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_AO5;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_AO6;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_AQ;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_A_CY;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_A_XOR;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_B;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_B1;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_B2;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_B3;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_B4;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_B5;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_B5Q;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_B6;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_BMUX;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_BO5;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_BO6;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_BQ;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_B_CY;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_B_XOR;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_C;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_C1;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_C2;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_C3;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_C4;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_C5;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_C6;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_CLK;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_CO5;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_CO6;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_CQ;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_C_CY;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_C_XOR;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_D;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_D1;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_D2;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_D3;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_D4;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_D5;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_D6;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_DO5;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_DO6;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_D_CY;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_D_XOR;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_A;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_A1;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_A2;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_A3;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_A4;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_A5;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_A6;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_AO5;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_AO6;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_AQ;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_A_CY;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_A_XOR;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_B;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_B1;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_B2;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_B3;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_B4;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_B5;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_B6;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_BO5;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_BO6;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_BQ;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_B_CY;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_B_XOR;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_C;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_C1;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_C2;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_C3;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_C4;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_C5;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_C6;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_CLK;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_CO5;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_CO6;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_C_CY;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_C_XOR;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_D;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_D1;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_D2;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_D3;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_D4;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_D5;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_D6;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_DO5;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_DO6;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_D_CY;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_D_XOR;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_A;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_A1;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_A2;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_A3;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_A4;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_A5;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_A6;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_AO5;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_AO6;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_AQ;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_A_CY;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_A_XOR;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_B;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_B1;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_B2;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_B3;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_B4;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_B5;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_B6;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_BO5;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_BO6;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_BQ;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_B_CY;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_B_XOR;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_C;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_C1;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_C2;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_C3;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_C4;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_C5;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_C6;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_CLK;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_CO5;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_CO6;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_CQ;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_C_CY;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_C_XOR;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_D;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_D1;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_D2;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_D3;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_D4;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_D5;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_D6;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_DO5;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_DO6;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_DQ;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_D_CY;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_D_XOR;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_A;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_A1;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_A2;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_A3;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_A4;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_A5;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_A6;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_AMUX;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_AO5;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_AO6;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_A_CY;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_A_XOR;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_B;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_B1;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_B2;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_B3;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_B4;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_B5;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_B6;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_BMUX;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_BO5;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_BO6;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_B_CY;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_B_XOR;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_C;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_C1;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_C2;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_C3;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_C4;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_C5;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_C6;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_CMUX;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_CO5;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_CO6;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_C_CY;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_C_XOR;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_D;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_D1;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_D2;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_D3;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_D4;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_D5;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_D6;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_DO5;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_DO6;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_D_CY;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_D_XOR;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_A;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_A1;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_A2;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_A3;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_A4;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_A5;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_A5Q;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_A6;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_AMUX;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_AO5;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_AO6;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_AQ;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_A_CY;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_A_XOR;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_B;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_B1;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_B2;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_B3;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_B4;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_B5;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_B6;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_BMUX;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_BO5;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_BO6;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_BQ;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_BX;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_B_CY;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_B_XOR;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_C;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_C1;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_C2;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_C3;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_C4;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_C5;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_C6;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_CLK;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_CMUX;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_CO5;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_CO6;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_C_CY;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_C_XOR;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_D;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_D1;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_D2;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_D3;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_D4;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_D5;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_D6;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_DMUX;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_DO5;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_DO6;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_D_CY;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_D_XOR;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_A;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_A1;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_A2;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_A3;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_A4;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_A5;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_A6;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_AO5;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_AO6;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_AQ;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_A_CY;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_A_XOR;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_B;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_B1;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_B2;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_B3;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_B4;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_B5;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_B6;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_BO5;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_BO6;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_B_CY;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_B_XOR;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_C;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_C1;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_C2;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_C3;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_C4;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_C5;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_C6;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_CLK;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_CMUX;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_CO5;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_CO6;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_C_CY;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_C_XOR;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_D;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_D1;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_D2;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_D3;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_D4;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_D5;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_D6;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_DO5;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_DO6;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_D_CY;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_D_XOR;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_A;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_A1;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_A2;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_A3;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_A4;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_A5;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_A6;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_AMUX;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_AO5;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_AO6;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_A_CY;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_A_XOR;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_B;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_B1;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_B2;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_B3;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_B4;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_B5;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_B6;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_BO5;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_BO6;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_B_CY;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_B_XOR;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_C;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_C1;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_C2;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_C3;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_C4;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_C5;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_C6;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_CO5;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_CO6;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_C_CY;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_C_XOR;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_D;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_D1;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_D2;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_D3;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_D4;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_D5;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_D6;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_DO5;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_DO6;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_D_CY;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_D_XOR;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_A;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_A1;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_A2;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_A3;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_A4;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_A5;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_A6;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_AO5;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_AO6;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_AQ;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_A_CY;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_A_XOR;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_B;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_B1;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_B2;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_B3;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_B4;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_B5;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_B5Q;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_B6;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_BMUX;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_BO5;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_BO6;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_BQ;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_B_CY;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_B_XOR;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_C;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_C1;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_C2;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_C3;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_C4;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_C5;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_C6;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_CLK;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_CO5;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_CO6;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_CQ;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_C_CY;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_C_XOR;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_D;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_D1;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_D2;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_D3;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_D4;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_D5;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_D6;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_DO5;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_DO6;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_D_CY;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_D_XOR;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_A;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_A1;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_A2;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_A3;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_A4;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_A5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_A6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_AO5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_AO6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_AQ;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_A_CY;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_A_XOR;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_B;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_B1;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_B2;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_B3;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_B4;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_B5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_B6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_BO5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_BO6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_BQ;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_B_CY;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_B_XOR;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_C;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_C1;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_C2;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_C3;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_C4;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_C5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_C6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_CLK;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_CO5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_CO6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_CQ;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_C_CY;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_C_XOR;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_D;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_D1;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_D2;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_D3;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_D4;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_D5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_D6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_DO5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_DO6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_D_CY;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_D_XOR;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_A;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_A1;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_A2;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_A3;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_A4;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_A5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_A6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_AO5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_AO6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_AQ;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_A_CY;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_A_XOR;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_B;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_B1;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_B2;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_B3;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_B4;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_B5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_B6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_BO5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_BO6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_BQ;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_B_CY;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_B_XOR;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_C;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_C1;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_C2;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_C3;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_C4;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_C5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_C6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_CLK;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_CO5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_CO6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_C_CY;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_C_XOR;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_D;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_D1;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_D2;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_D3;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_D4;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_D5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_D6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_DO5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_DO6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_D_CY;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_D_XOR;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_A;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_A1;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_A2;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_A3;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_A4;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_A5;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_A6;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_AO5;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_AO6;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_AQ;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_A_CY;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_A_XOR;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_B;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_B1;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_B2;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_B3;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_B4;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_B5;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_B5Q;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_B6;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_BMUX;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_BO5;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_BO6;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_BQ;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_B_CY;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_B_XOR;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_C;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_C1;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_C2;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_C3;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_C4;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_C5;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_C6;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_CLK;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_CO5;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_CO6;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_CQ;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_C_CY;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_C_XOR;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_D;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_D1;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_D2;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_D3;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_D4;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_D5;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_D6;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_DO5;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_DO6;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_DQ;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_D_CY;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_D_XOR;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_A;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_A1;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_A2;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_A3;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_A4;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_A5;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_A6;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_AO5;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_AO6;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_AQ;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_A_CY;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_A_XOR;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_B;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_B1;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_B2;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_B3;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_B4;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_B5;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_B6;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_BO5;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_BO6;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_BQ;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_B_CY;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_B_XOR;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_C;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_C1;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_C2;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_C3;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_C4;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_C5;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_C6;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_CLK;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_CO5;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_CO6;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_CQ;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_C_CY;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_C_XOR;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_D;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_D1;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_D2;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_D3;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_D4;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_D5;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_D6;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_DO5;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_DO6;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_DQ;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_D_CY;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_D_XOR;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_A;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_A1;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_A2;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_A3;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_A4;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_A5;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_A6;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_AO5;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_AO6;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_AQ;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_A_CY;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_A_XOR;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_B;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_B1;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_B2;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_B3;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_B4;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_B5;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_B6;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_BO5;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_BO6;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_BQ;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_B_CY;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_B_XOR;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_C;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_C1;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_C2;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_C3;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_C4;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_C5;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_C6;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_CLK;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_CO5;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_CO6;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_CQ;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_C_CY;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_C_XOR;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_D;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_D1;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_D2;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_D3;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_D4;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_D5;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_D6;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_DO5;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_DO6;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_DQ;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_D_CY;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_D_XOR;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_A;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_A1;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_A2;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_A3;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_A4;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_A5;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_A6;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_AO5;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_AO6;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_AQ;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_A_CY;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_A_XOR;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_B;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_B1;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_B2;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_B3;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_B4;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_B5;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_B6;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_BMUX;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_BO5;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_BO6;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_B_CY;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_B_XOR;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_C;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_C1;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_C2;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_C3;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_C4;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_C5;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_C6;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_CLK;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_CO5;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_CO6;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_C_CY;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_C_XOR;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_D;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_D1;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_D2;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_D3;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_D4;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_D5;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_D6;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_DO5;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_DO6;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_D_CY;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_D_XOR;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_A;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_A1;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_A2;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_A3;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_A4;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_A5;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_A6;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_AO5;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_AO6;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_AQ;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_A_CY;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_A_XOR;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_B;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_B1;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_B2;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_B3;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_B4;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_B5;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_B6;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_BO5;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_BO6;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_BQ;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_B_CY;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_B_XOR;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_C;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_C1;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_C2;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_C3;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_C4;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_C5;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_C6;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_CLK;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_CMUX;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_CO5;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_CO6;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_C_CY;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_C_XOR;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_D;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_D1;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_D2;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_D3;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_D4;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_D5;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_D6;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_DMUX;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_DO5;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_DO6;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_D_CY;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_D_XOR;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_A;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_A1;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_A2;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_A3;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_A4;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_A5;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_A6;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_AO5;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_AO6;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_AQ;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_A_CY;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_A_XOR;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_B;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_B1;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_B2;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_B3;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_B4;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_B5;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_B6;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_BO5;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_BO6;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_BQ;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_B_CY;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_B_XOR;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_C;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_C1;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_C2;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_C3;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_C4;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_C5;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_C6;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_CLK;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_CO5;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_CO6;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_CQ;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_C_CY;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_C_XOR;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_D;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_D1;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_D2;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_D3;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_D4;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_D5;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_D6;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_DO5;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_DO6;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_DQ;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_D_CY;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_D_XOR;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_A;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_A1;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_A2;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_A3;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_A4;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_A5;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_A6;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_AO5;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_AO6;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_AQ;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_A_CY;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_A_XOR;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_B;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_B1;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_B2;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_B3;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_B4;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_B5;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_B6;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_BMUX;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_BO5;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_BO6;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_B_CY;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_B_XOR;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_C;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_C1;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_C2;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_C3;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_C4;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_C5;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_C6;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_CLK;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_CO5;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_CO6;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_C_CY;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_C_XOR;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_D;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_D1;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_D2;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_D3;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_D4;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_D5;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_D6;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_DMUX;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_DO5;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_DO6;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_D_CY;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_D_XOR;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_A;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_A1;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_A2;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_A3;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_A4;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_A5;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_A6;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_AMUX;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_AO5;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_AO6;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_A_CY;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_A_XOR;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_B;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_B1;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_B2;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_B3;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_B4;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_B5;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_B6;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_BO5;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_BO6;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_B_CY;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_B_XOR;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_C;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_C1;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_C2;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_C3;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_C4;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_C5;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_C6;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_CO5;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_CO6;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_C_CY;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_C_XOR;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_D;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_D1;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_D2;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_D3;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_D4;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_D5;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_D6;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_DO5;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_DO6;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_D_CY;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_D_XOR;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_A;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_A1;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_A2;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_A3;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_A4;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_A5;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_A6;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_AO5;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_AO6;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_AQ;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_A_CY;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_A_XOR;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_B;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_B1;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_B2;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_B3;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_B4;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_B5;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_B6;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_BO5;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_BO6;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_BQ;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_B_CY;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_B_XOR;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_C;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_C1;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_C2;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_C3;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_C4;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_C5;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_C6;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_CLK;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_CMUX;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_CO5;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_CO6;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_C_CY;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_C_XOR;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_D;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_D1;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_D2;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_D3;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_D4;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_D5;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_D6;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_DO5;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_DO6;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_D_CY;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_D_XOR;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X11Y155_A;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X11Y155_A1;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X11Y155_A2;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X11Y155_A3;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X11Y155_A4;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X11Y155_A5;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X11Y155_A6;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X11Y155_AO5;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X11Y155_AO6;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X11Y155_A_CY;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X11Y155_A_XOR;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X11Y155_B;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X11Y155_B1;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X11Y155_B2;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X11Y155_B3;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X11Y155_B4;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X11Y155_B5;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X11Y155_B6;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X11Y155_BO5;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X11Y155_BO6;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X11Y155_B_CY;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X11Y155_B_XOR;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X11Y155_C;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X11Y155_C1;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X11Y155_C2;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X11Y155_C3;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X11Y155_C4;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X11Y155_C5;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X11Y155_C6;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X11Y155_CO5;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X11Y155_CO6;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X11Y155_C_CY;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X11Y155_C_XOR;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X11Y155_D;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X11Y155_D1;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X11Y155_D2;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X11Y155_D3;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X11Y155_D4;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X11Y155_D5;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X11Y155_D6;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X11Y155_DO5;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X11Y155_DO6;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X11Y155_D_CY;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X11Y155_D_XOR;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X10Y159_A;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X10Y159_A1;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X10Y159_A2;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X10Y159_A3;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X10Y159_A4;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X10Y159_A5;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X10Y159_A6;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X10Y159_AO5;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X10Y159_AO6;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X10Y159_A_CY;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X10Y159_A_XOR;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X10Y159_B;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X10Y159_B1;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X10Y159_B2;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X10Y159_B3;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X10Y159_B4;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X10Y159_B5;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X10Y159_B6;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X10Y159_BO5;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X10Y159_BO6;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X10Y159_B_CY;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X10Y159_B_XOR;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X10Y159_C;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X10Y159_C1;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X10Y159_C2;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X10Y159_C3;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X10Y159_C4;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X10Y159_C5;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X10Y159_C6;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X10Y159_CO5;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X10Y159_CO6;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X10Y159_C_CY;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X10Y159_C_XOR;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X10Y159_D;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X10Y159_D1;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X10Y159_D2;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X10Y159_D3;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X10Y159_D4;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X10Y159_D5;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X10Y159_D6;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X10Y159_DO5;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X10Y159_DO6;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X10Y159_D_CY;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X10Y159_D_XOR;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X11Y159_A;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X11Y159_A1;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X11Y159_A2;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X11Y159_A3;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X11Y159_A4;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X11Y159_A5;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X11Y159_A6;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X11Y159_AO5;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X11Y159_AO6;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X11Y159_A_CY;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X11Y159_A_XOR;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X11Y159_B;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X11Y159_B1;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X11Y159_B2;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X11Y159_B3;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X11Y159_B4;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X11Y159_B5;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X11Y159_B6;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X11Y159_BO5;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X11Y159_BO6;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X11Y159_B_CY;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X11Y159_B_XOR;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X11Y159_C;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X11Y159_C1;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X11Y159_C2;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X11Y159_C3;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X11Y159_C4;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X11Y159_C5;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X11Y159_C6;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X11Y159_CO5;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X11Y159_CO6;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X11Y159_C_CY;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X11Y159_C_XOR;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X11Y159_D;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X11Y159_D1;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X11Y159_D2;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X11Y159_D3;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X11Y159_D4;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X11Y159_D5;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X11Y159_D6;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X11Y159_DO5;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X11Y159_DO6;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X11Y159_D_CY;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X11Y159_D_XOR;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_A;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_A1;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_A2;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_A3;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_A4;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_A5;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_A6;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_AO5;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_AO6;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_A_CY;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_A_XOR;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_B;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_B1;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_B2;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_B3;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_B4;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_B5;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_B6;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_BO5;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_BO6;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_B_CY;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_B_XOR;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_C;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_C1;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_C2;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_C3;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_C4;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_C5;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_C6;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_CO5;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_CO6;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_C_CY;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_C_XOR;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_D;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_D1;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_D2;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_D3;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_D4;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_D5;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_D6;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_DO5;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_DO6;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_D_CY;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_D_XOR;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_A;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_A1;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_A2;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_A3;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_A4;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_A5;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_A6;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_AMUX;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_AO5;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_AO6;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_A_CY;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_A_XOR;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_B;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_B1;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_B2;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_B3;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_B4;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_B5;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_B6;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_BO5;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_BO6;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_B_CY;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_B_XOR;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_C;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_C1;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_C2;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_C3;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_C4;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_C5;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_C6;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_CO5;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_CO6;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_C_CY;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_C_XOR;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_D;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_D1;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_D2;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_D3;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_D4;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_D5;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_D6;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_DO5;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_DO6;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_D_CY;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_D_XOR;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A1;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A2;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A3;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A4;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_AO5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_AO6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A_CY;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A_XOR;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B1;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B2;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B3;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B4;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_BO5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_BO6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B_CY;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B_XOR;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C1;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C2;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C3;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C4;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_CO5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_CO6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C_CY;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C_XOR;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D1;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D2;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D3;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D4;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_DO5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_DO6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D_CY;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D_XOR;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A1;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A2;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A3;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A4;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_AO5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_AO6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A_CY;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A_XOR;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B1;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B2;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B3;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B4;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_BO5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_BO6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B_CY;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B_XOR;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C1;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C2;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C3;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C4;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_CO5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_CO6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C_CY;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C_XOR;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D1;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D2;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D3;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D4;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_DO5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_DO6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D_CY;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D_XOR;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_A;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_A1;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_A2;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_A3;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_A4;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_A5;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_A6;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_AO5;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_AO6;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_A_CY;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_A_XOR;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_B;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_B1;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_B2;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_B3;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_B4;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_B5;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_B6;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_BO5;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_BO6;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_B_CY;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_B_XOR;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_C;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_C1;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_C2;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_C3;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_C4;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_C5;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_C6;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_CO5;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_CO6;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_C_CY;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_C_XOR;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_D;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_D1;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_D2;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_D3;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_D4;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_D5;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_D6;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_DO5;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_DO6;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_D_CY;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_D_XOR;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_A;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_A1;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_A2;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_A3;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_A4;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_A5;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_A6;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_AMUX;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_AO5;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_AO6;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_A_CY;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_A_XOR;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_B;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_B1;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_B2;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_B3;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_B4;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_B5;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_B6;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_BO5;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_BO6;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_B_CY;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_B_XOR;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_C;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_C1;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_C2;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_C3;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_C4;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_C5;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_C6;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_CO5;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_CO6;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_C_CY;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_C_XOR;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_D;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_D1;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_D2;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_D3;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_D4;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_D5;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_D6;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_DO5;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_DO6;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_D_CY;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_D_XOR;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_A;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_A1;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_A2;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_A3;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_A4;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_A5;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_A6;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_AO5;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_AO6;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_A_CY;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_A_XOR;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_B;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_B1;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_B2;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_B3;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_B4;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_B5;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_B6;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_BO5;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_BO6;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_B_CY;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_B_XOR;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_C;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_C1;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_C2;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_C3;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_C4;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_C5;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_C6;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_CO5;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_CO6;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_C_CY;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_C_XOR;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_D;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_D1;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_D2;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_D3;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_D4;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_D5;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_D6;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_DO5;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_DO6;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_D_CY;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_D_XOR;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_A;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_A1;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_A2;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_A3;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_A4;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_A5;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_A6;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_AMUX;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_AO5;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_AO6;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_A_CY;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_A_XOR;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_B;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_B1;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_B2;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_B3;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_B4;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_B5;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_B6;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_BO5;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_BO6;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_B_CY;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_B_XOR;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_C;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_C1;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_C2;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_C3;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_C4;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_C5;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_C6;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_CO5;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_CO6;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_C_CY;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_C_XOR;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_D;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_D1;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_D2;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_D3;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_D4;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_D5;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_D6;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_DO5;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_DO6;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_D_CY;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_D_XOR;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_A;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_A1;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_A2;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_A3;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_A4;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_A5;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_A6;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_AO5;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_AO6;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_A_CY;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_A_XOR;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_B;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_B1;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_B2;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_B3;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_B4;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_B5;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_B6;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_BO5;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_BO6;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_B_CY;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_B_XOR;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_C;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_C1;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_C2;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_C3;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_C4;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_C5;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_C6;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_CO5;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_CO6;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_C_CY;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_C_XOR;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_D;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_D1;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_D2;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_D3;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_D4;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_D5;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_D6;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_DO5;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_DO6;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_D_CY;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X162Y176_D_XOR;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_A;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_A1;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_A2;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_A3;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_A4;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_A5;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_A6;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_AMUX;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_AO5;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_AO6;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_A_CY;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_A_XOR;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_B;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_B1;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_B2;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_B3;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_B4;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_B5;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_B6;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_BO5;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_BO6;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_B_CY;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_B_XOR;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_C;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_C1;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_C2;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_C3;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_C4;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_C5;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_C6;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_CO5;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_CO6;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_C_CY;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_C_XOR;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_D;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_D1;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_D2;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_D3;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_D4;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_D5;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_D6;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_DO5;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_DO6;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_D_CY;
  wire [0:0] CLBLM_R_X103Y176_SLICE_X163Y176_D_XOR;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_A;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_A1;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_A2;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_A3;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_A4;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_A5;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_A6;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_AO5;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_AO6;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_A_CY;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_A_XOR;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_B;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_B1;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_B2;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_B3;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_B4;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_B5;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_B6;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_BO5;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_BO6;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_B_CY;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_B_XOR;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_C;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_C1;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_C2;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_C3;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_C4;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_C5;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_C6;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_CO5;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_CO6;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_C_CY;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_C_XOR;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_D;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_D1;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_D2;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_D3;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_D4;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_D5;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_D6;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_DO5;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_DO6;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_D_CY;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_D_XOR;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_A;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_A1;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_A2;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_A3;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_A4;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_A5;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_A6;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_AMUX;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_AO5;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_AO6;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_A_CY;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_A_XOR;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_B;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_B1;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_B2;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_B3;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_B4;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_B5;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_B6;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_BO5;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_BO6;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_B_CY;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_B_XOR;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_C;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_C1;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_C2;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_C3;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_C4;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_C5;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_C6;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_CO5;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_CO6;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_C_CY;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_C_XOR;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_D;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_D1;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_D2;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_D3;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_D4;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_D5;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_D6;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_DO5;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_DO6;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_D_CY;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_D_XOR;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_A;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_A1;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_A2;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_A3;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_A4;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_A5;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_A6;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_AO5;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_AO6;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_AQ;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_A_CY;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_A_XOR;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_B;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_B1;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_B2;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_B3;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_B4;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_B5;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_B6;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_BO5;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_BO6;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_BQ;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_B_CY;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_B_XOR;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_C;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_C1;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_C2;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_C3;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_C4;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_C5;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_C6;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_CLK;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_CMUX;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_CO5;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_CO6;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_C_CY;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_C_XOR;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_D;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_D1;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_D2;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_D3;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_D4;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_D5;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_D6;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_DO5;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_DO6;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_D_CY;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_D_XOR;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_A;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_A1;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_A2;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_A3;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_A4;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_A5;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_A6;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_AO5;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_AO6;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_A_CY;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_A_XOR;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_B;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_B1;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_B2;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_B3;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_B4;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_B5;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_B6;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_BO5;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_BO6;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_B_CY;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_B_XOR;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_C;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_C1;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_C2;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_C3;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_C4;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_C5;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_C6;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_CO5;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_CO6;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_C_CY;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_C_XOR;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_D;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_D1;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_D2;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_D3;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_D4;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_D5;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_D6;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_DO5;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_DO6;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_D_CY;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_D_XOR;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_A;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_A1;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_A2;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_A3;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_A4;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_A5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_A6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_AO5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_AO6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_AQ;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_A_CY;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_A_XOR;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_B;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_B1;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_B2;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_B3;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_B4;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_B5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_B6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_BO5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_BO6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_BQ;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_B_CY;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_B_XOR;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_C;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_C1;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_C2;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_C3;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_C4;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_C5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_C6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_CLK;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_CO5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_CO6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_C_CY;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_C_XOR;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_D;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_D1;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_D2;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_D3;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_D4;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_D5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_D6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_DO5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_DO6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_D_CY;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_D_XOR;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_A;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_A1;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_A2;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_A3;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_A4;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_A5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_A6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_AMUX;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_AO5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_AO6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_A_CY;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_A_XOR;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_B;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_B1;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_B2;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_B3;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_B4;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_B5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_B6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_BO5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_BO6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_B_CY;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_B_XOR;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_C;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_C1;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_C2;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_C3;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_C4;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_C5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_C6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_CO5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_CO6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_C_CY;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_C_XOR;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_D;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_D1;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_D2;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_D3;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_D4;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_D5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_D6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_DO5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_DO6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_D_CY;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_D_XOR;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_A;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_A1;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_A2;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_A3;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_A4;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_A5;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_A6;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_AO5;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_AO6;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_AQ;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_A_CY;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_A_XOR;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_B;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_B1;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_B2;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_B3;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_B4;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_B5;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_B6;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_BO5;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_BO6;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_BQ;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_B_CY;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_B_XOR;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_C;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_C1;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_C2;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_C3;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_C4;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_C5;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_C6;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_CLK;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_CO5;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_CO6;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_C_CY;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_C_XOR;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_D;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_D1;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_D2;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_D3;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_D4;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_D5;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_D6;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_DO5;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_DO6;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_D_CY;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_D_XOR;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_A;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_A1;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_A2;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_A3;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_A4;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_A5;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_A6;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_AO5;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_AO6;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_AQ;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_A_CY;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_A_XOR;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_B;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_B1;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_B2;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_B3;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_B4;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_B5;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_B6;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_BO5;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_BO6;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_BQ;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_B_CY;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_B_XOR;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_C;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_C1;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_C2;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_C3;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_C4;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_C5;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_C6;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_CLK;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_CO5;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_CO6;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_C_CY;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_C_XOR;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_D;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_D1;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_D2;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_D3;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_D4;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_D5;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_D6;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_DO5;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_DO6;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_D_CY;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_D_XOR;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_A;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_A1;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_A2;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_A3;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_A4;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_A5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_A6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_AO5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_AO6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_AQ;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_A_CY;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_A_XOR;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_B;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_B1;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_B2;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_B3;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_B4;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_B5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_B6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_BO5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_BO6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_BQ;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_B_CY;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_B_XOR;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_C;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_C1;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_C2;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_C3;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_C4;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_C5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_C6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_CLK;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_CO5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_CO6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_CQ;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_C_CY;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_C_XOR;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_D;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_D1;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_D2;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_D3;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_D4;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_D5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_D6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_DO5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_DO6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_DQ;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_D_CY;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_D_XOR;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_A;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_A1;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_A2;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_A3;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_A4;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_A5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_A6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_AO5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_AO6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_AQ;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_A_CY;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_A_XOR;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_B;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_B1;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_B2;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_B3;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_B4;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_B5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_B6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_BO5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_BO6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_BQ;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_B_CY;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_B_XOR;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_C;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_C1;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_C2;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_C3;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_C4;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_C5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_C6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_CLK;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_CO5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_CO6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_CQ;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_C_CY;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_C_XOR;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_D;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_D1;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_D2;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_D3;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_D4;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_D5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_D6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_DO5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_DO6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_DQ;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_D_CY;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_D_XOR;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_A;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_A1;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_A2;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_A3;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_A4;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_A5;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_A6;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_AO5;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_AO6;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_AQ;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_A_CY;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_A_XOR;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_B;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_B1;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_B2;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_B3;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_B4;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_B5;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_B6;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_BO5;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_BO6;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_BQ;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_B_CY;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_B_XOR;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_C;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_C1;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_C2;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_C3;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_C4;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_C5;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_C6;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_CLK;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_CO5;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_CO6;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_C_CY;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_C_XOR;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_D;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_D1;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_D2;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_D3;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_D4;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_D5;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_D6;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_DO5;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_DO6;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_D_CY;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_D_XOR;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_A;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_A1;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_A2;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_A3;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_A4;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_A5;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_A6;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_AO5;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_AO6;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_AQ;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_A_CY;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_A_XOR;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_B;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_B1;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_B2;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_B3;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_B4;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_B5;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_B6;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_BO5;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_BO6;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_BQ;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_B_CY;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_B_XOR;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_C;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_C1;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_C2;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_C3;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_C4;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_C5;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_C6;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_CLK;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_CO5;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_CO6;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_CQ;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_C_CY;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_C_XOR;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_D;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_D1;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_D2;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_D3;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_D4;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_D5;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_D6;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_DO5;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_DO6;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_DQ;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_D_CY;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_D_XOR;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_A;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_A1;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_A2;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_A3;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_A4;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_A5;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_A6;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_AO5;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_AO6;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_AQ;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_A_CY;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_A_XOR;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_B;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_B1;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_B2;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_B3;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_B4;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_B5;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_B6;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_BO5;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_BO6;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_BQ;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_B_CY;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_B_XOR;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_C;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_C1;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_C2;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_C3;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_C4;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_C5;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_C6;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_CLK;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_CO5;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_CO6;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_CQ;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_C_CY;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_C_XOR;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_D;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_D1;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_D2;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_D3;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_D4;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_D5;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_D6;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_DO5;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_DO6;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_DQ;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_D_CY;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_D_XOR;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_A;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_A1;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_A2;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_A3;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_A4;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_A5;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_A5Q;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_A6;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_AMUX;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_AO5;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_AO6;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_AQ;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_AX;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_A_CY;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_A_XOR;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_B;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_B1;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_B2;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_B3;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_B4;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_B5;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_B5Q;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_B6;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_BMUX;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_BO5;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_BO6;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_BQ;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_B_CY;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_B_XOR;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_C;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_C1;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_C2;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_C3;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_C4;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_C5;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_C6;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_CLK;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_CO5;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_CO6;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_CQ;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_C_CY;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_C_XOR;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_D;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_D1;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_D2;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_D3;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_D4;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_D5;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_D6;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_DO5;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_DO6;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_D_CY;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_D_XOR;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_A;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_A1;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_A2;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_A3;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_A4;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_A5;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_A6;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_AO5;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_AO6;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_AQ;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_A_CY;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_A_XOR;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_B;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_B1;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_B2;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_B3;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_B4;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_B5;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_B6;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_BO5;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_BO6;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_BQ;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_B_CY;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_B_XOR;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_C;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_C1;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_C2;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_C3;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_C4;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_C5;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_C6;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_CLK;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_CO5;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_CO6;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_CQ;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_C_CY;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_C_XOR;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_D;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_D1;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_D2;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_D3;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_D4;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_D5;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_D6;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_DMUX;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_DO5;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_DO6;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_D_CY;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_D_XOR;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_A;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_A1;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_A2;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_A3;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_A4;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_A5;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_A6;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_AO5;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_AO6;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_A_CY;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_A_XOR;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_B;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_B1;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_B2;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_B3;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_B4;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_B5;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_B6;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_BO5;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_BO6;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_B_CY;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_B_XOR;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_C;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_C1;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_C2;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_C3;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_C4;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_C5;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_C6;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_CO5;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_CO6;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_C_CY;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_C_XOR;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_D;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_D1;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_D2;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_D3;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_D4;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_D5;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_D6;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_DO5;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_DO6;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_D_CY;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_D_XOR;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_A;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_A1;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_A2;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_A3;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_A4;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_A5;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_A6;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_AO5;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_AO6;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_A_CY;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_A_XOR;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_B;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_B1;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_B2;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_B3;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_B4;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_B5;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_B6;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_BO5;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_BO6;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_B_CY;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_B_XOR;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_C;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_C1;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_C2;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_C3;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_C4;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_C5;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_C6;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_CO5;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_CO6;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_C_CY;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_C_XOR;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_D;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_D1;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_D2;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_D3;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_D4;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_D5;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_D6;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_DO5;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_DO6;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_D_CY;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_D_XOR;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_A;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_A1;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_A2;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_A3;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_A4;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_A5;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_A6;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_AO5;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_AO6;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_AQ;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_A_CY;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_A_XOR;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_B;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_B1;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_B2;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_B3;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_B4;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_B5;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_B6;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_BO5;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_BO6;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_BQ;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_B_CY;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_B_XOR;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_C;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_C1;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_C2;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_C3;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_C4;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_C5;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_C6;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_CLK;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_CO5;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_CO6;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_CQ;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_C_CY;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_C_XOR;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_D;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_D1;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_D2;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_D3;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_D4;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_D5;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_D6;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_DMUX;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_DO5;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_DO6;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_D_CY;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_D_XOR;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_A;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_A1;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_A2;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_A3;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_A4;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_A5;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_A6;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_AMUX;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_AO5;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_AO6;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_AQ;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_AX;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_A_CY;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_A_XOR;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_B;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_B1;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_B2;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_B3;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_B4;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_B5;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_B6;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_BMUX;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_BO5;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_BO6;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_BQ;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_BX;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_B_CY;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_B_XOR;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_C;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_C1;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_C2;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_C3;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_C4;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_C5;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_C6;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_CE;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_CLK;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_CMUX;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_CO5;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_CO6;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_C_CY;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_C_XOR;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_D;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_D1;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_D2;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_D3;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_D4;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_D5;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_D6;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_DMUX;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_DO5;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_DO6;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_D_CY;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_D_XOR;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_SR;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_A;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_A1;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_A2;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_A3;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_A4;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_A5;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_A5Q;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_A6;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_AMUX;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_AO5;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_AO6;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_AQ;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_AX;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_A_CY;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_A_XOR;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_B;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_B1;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_B2;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_B3;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_B4;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_B5;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_B6;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_BO5;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_BO6;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_BQ;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_B_CY;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_B_XOR;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_C;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_C1;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_C2;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_C3;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_C4;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_C5;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_C6;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_CLK;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_CMUX;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_CO5;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_CO6;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_C_CY;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_C_XOR;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_D;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_D1;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_D2;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_D3;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_D4;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_D5;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_D6;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_DO5;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_DO6;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_D_CY;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_D_XOR;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_A;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_A1;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_A2;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_A3;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_A4;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_A5;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_A6;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_AO5;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_AO6;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_AQ;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_A_CY;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_A_XOR;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_B;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_B1;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_B2;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_B3;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_B4;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_B5;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_B6;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_BO5;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_BO6;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_BQ;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_B_CY;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_B_XOR;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_C;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_C1;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_C2;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_C3;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_C4;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_C5;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_C6;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_CLK;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_CO5;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_CO6;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_CQ;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_C_CY;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_C_XOR;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_D;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_D1;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_D2;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_D3;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_D4;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_D5;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_D6;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_DO5;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_DO6;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_DQ;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_D_CY;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_D_XOR;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_A;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_A1;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_A2;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_A3;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_A4;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_A5;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_A6;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_AO5;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_AO6;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_AQ;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_A_CY;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_A_XOR;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_B;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_B1;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_B2;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_B3;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_B4;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_B5;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_B6;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_BO5;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_BO6;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_BQ;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_B_CY;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_B_XOR;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_C;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_C1;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_C2;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_C3;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_C4;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_C5;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_C6;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_CLK;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_CO5;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_CO6;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_C_CY;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_C_XOR;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_D;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_D1;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_D2;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_D3;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_D4;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_D5;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_D6;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_DO5;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_DO6;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_D_CY;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_D_XOR;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_A;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_A1;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_A2;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_A3;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_A4;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_A5;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_A6;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_AMUX;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_AO5;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_AO6;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_AQ;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_AX;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_A_CY;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_A_XOR;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_B;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_B1;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_B2;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_B3;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_B4;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_B5;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_B6;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_BMUX;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_BO5;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_BO6;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_BQ;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_BX;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_B_CY;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_B_XOR;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_C;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_C1;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_C2;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_C3;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_C4;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_C5;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_C6;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_CE;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_CLK;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_CMUX;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_CO5;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_CO6;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_CQ;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_CX;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_C_CY;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_C_XOR;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_D;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_D1;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_D2;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_D3;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_D4;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_D5;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_D6;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_DMUX;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_DO5;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_DO6;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_D_CY;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_D_XOR;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_SR;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_A;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_A1;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_A2;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_A3;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_A4;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_A5;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_A6;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_AO5;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_AO6;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_AQ;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_A_CY;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_A_XOR;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_B;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_B1;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_B2;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_B3;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_B4;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_B5;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_B6;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_BO5;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_BO6;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_BQ;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_B_CY;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_B_XOR;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_C;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_C1;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_C2;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_C3;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_C4;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_C5;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_C6;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_CLK;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_CMUX;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_CO5;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_CO6;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_C_CY;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_C_XOR;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_D;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_D1;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_D2;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_D3;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_D4;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_D5;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_D6;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_DO5;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_DO6;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_D_CY;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_D_XOR;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_A;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_A1;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_A2;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_A3;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_A4;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_A5;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_A6;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_AO5;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_AO6;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_AQ;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_A_CY;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_A_XOR;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_B;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_B1;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_B2;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_B3;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_B4;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_B5;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_B6;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_BMUX;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_BO5;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_BO6;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_B_CY;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_B_XOR;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_C;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_C1;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_C2;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_C3;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_C4;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_C5;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_C6;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_CLK;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_CMUX;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_CO5;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_CO6;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_C_CY;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_C_XOR;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_D;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_D1;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_D2;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_D3;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_D4;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_D5;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_D6;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_DO5;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_DO6;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_D_CY;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_D_XOR;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X15Y154_A;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X15Y154_A1;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X15Y154_A2;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X15Y154_A3;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X15Y154_A4;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X15Y154_A5;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X15Y154_A6;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X15Y154_AO5;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X15Y154_AO6;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X15Y154_AQ;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X15Y154_A_CY;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X15Y154_A_XOR;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X15Y154_B;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X15Y154_B1;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X15Y154_B2;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X15Y154_B3;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X15Y154_B4;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X15Y154_B5;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X15Y154_B6;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X15Y154_BO5;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X15Y154_BO6;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X15Y154_BQ;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X15Y154_B_CY;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X15Y154_B_XOR;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X15Y154_C;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X15Y154_C1;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X15Y154_C2;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X15Y154_C3;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X15Y154_C4;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X15Y154_C5;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X15Y154_C6;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X15Y154_CLK;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X15Y154_CMUX;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X15Y154_CO5;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X15Y154_CO6;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X15Y154_C_CY;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X15Y154_C_XOR;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X15Y154_D;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X15Y154_D1;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X15Y154_D2;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X15Y154_D3;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X15Y154_D4;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X15Y154_D5;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X15Y154_D6;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X15Y154_DO5;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X15Y154_DO6;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X15Y154_D_CY;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X15Y154_D_XOR;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X14Y157_A;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X14Y157_A1;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X14Y157_A2;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X14Y157_A3;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X14Y157_A4;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X14Y157_A5;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X14Y157_A6;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X14Y157_AMUX;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X14Y157_AO5;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X14Y157_AO6;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X14Y157_A_CY;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X14Y157_A_XOR;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X14Y157_B;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X14Y157_B1;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X14Y157_B2;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X14Y157_B3;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X14Y157_B4;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X14Y157_B5;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X14Y157_B6;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X14Y157_BO5;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X14Y157_BO6;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X14Y157_B_CY;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X14Y157_B_XOR;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X14Y157_C;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X14Y157_C1;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X14Y157_C2;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X14Y157_C3;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X14Y157_C4;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X14Y157_C5;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X14Y157_C6;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X14Y157_CO5;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X14Y157_CO6;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X14Y157_C_CY;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X14Y157_C_XOR;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X14Y157_D;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X14Y157_D1;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X14Y157_D2;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X14Y157_D3;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X14Y157_D4;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X14Y157_D5;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X14Y157_D6;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X14Y157_DO5;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X14Y157_DO6;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X14Y157_D_CY;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X14Y157_D_XOR;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X15Y157_A;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X15Y157_A1;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X15Y157_A2;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X15Y157_A3;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X15Y157_A4;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X15Y157_A5;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X15Y157_A6;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X15Y157_AO5;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X15Y157_AO6;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X15Y157_A_CY;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X15Y157_A_XOR;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X15Y157_B;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X15Y157_B1;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X15Y157_B2;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X15Y157_B3;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X15Y157_B4;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X15Y157_B5;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X15Y157_B6;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X15Y157_BO5;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X15Y157_BO6;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X15Y157_B_CY;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X15Y157_B_XOR;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X15Y157_C;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X15Y157_C1;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X15Y157_C2;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X15Y157_C3;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X15Y157_C4;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X15Y157_C5;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X15Y157_C6;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X15Y157_CO5;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X15Y157_CO6;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X15Y157_C_CY;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X15Y157_C_XOR;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X15Y157_D;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X15Y157_D1;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X15Y157_D2;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X15Y157_D3;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X15Y157_D4;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X15Y157_D5;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X15Y157_D6;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X15Y157_DO5;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X15Y157_DO6;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X15Y157_D_CY;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X15Y157_D_XOR;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_A;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_A1;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_A2;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_A3;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_A4;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_A5;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_A6;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_AO5;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_AO6;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_A_CY;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_A_XOR;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_B;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_B1;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_B2;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_B3;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_B4;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_B5;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_B6;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_BO5;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_BO6;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_B_CY;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_B_XOR;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_C;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_C1;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_C2;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_C3;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_C4;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_C5;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_C6;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_CO5;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_CO6;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_C_CY;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_C_XOR;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_D;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_D1;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_D2;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_D3;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_D4;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_D5;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_D6;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_DO5;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_DO6;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_D_CY;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_D_XOR;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_A;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_A1;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_A2;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_A3;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_A4;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_A5;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_A6;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_AO5;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_AO6;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_A_CY;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_A_XOR;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_B;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_B1;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_B2;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_B3;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_B4;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_B5;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_B6;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_BO5;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_BO6;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_B_CY;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_B_XOR;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_C;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_C1;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_C2;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_C3;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_C4;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_C5;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_C6;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_CO5;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_CO6;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_C_CY;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_C_XOR;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_D;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_D1;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_D2;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_D3;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_D4;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_D5;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_D6;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_DO5;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_DO6;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_D_CY;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_D_XOR;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_A;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_A1;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_A2;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_A3;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_A4;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_A5;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_A6;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_AO5;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_AO6;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_A_CY;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_A_XOR;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_B;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_B1;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_B2;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_B3;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_B4;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_B5;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_B6;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_BO5;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_BO6;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_B_CY;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_B_XOR;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_C;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_C1;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_C2;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_C3;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_C4;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_C5;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_C6;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_CO5;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_CO6;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_C_CY;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_C_XOR;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_D;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_D1;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_D2;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_D3;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_D4;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_D5;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_D6;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_DO5;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_DO6;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_D_CY;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_D_XOR;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_A;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_A1;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_A2;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_A3;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_A4;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_A5;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_A6;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_AO5;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_AO6;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_A_CY;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_A_XOR;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_B;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_B1;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_B2;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_B3;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_B4;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_B5;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_B6;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_BO5;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_BO6;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_B_CY;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_B_XOR;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_C;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_C1;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_C2;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_C3;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_C4;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_C5;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_C6;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_CO5;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_CO6;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_C_CY;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_C_XOR;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_D;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_D1;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_D2;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_D3;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_D4;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_D5;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_D6;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_DO5;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_DO6;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_D_CY;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_D_XOR;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_A;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_A1;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_A2;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_A3;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_A4;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_A5;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_A6;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_AO5;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_AO6;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_AQ;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_AX;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_A_CY;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_A_XOR;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_B;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_B1;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_B2;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_B3;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_B4;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_B5;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_B6;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_BO5;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_BO6;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_B_CY;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_B_XOR;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_C;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_C1;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_C2;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_C3;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_C4;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_C5;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_C6;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_CLK;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_CO5;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_CO6;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_C_CY;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_C_XOR;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_D;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_D1;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_D2;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_D3;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_D4;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_D5;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_D6;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_DO5;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_DO6;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_D_CY;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X20Y151_D_XOR;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_A;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_A1;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_A2;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_A3;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_A4;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_A5;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_A6;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_AO5;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_AO6;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_A_CY;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_A_XOR;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_B;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_B1;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_B2;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_B3;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_B4;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_B5;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_B6;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_BO5;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_BO6;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_B_CY;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_B_XOR;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_C;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_C1;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_C2;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_C3;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_C4;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_C5;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_C6;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_CO5;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_CO6;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_C_CY;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_C_XOR;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_D;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_D1;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_D2;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_D3;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_D4;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_D5;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_D6;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_DO5;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_DO6;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_D_CY;
  wire [0:0] CLBLM_R_X15Y151_SLICE_X21Y151_D_XOR;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X20Y153_A;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X20Y153_A1;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X20Y153_A2;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X20Y153_A3;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X20Y153_A4;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X20Y153_A5;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X20Y153_A6;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X20Y153_AMUX;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X20Y153_AO5;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X20Y153_AO6;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X20Y153_A_CY;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X20Y153_A_XOR;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X20Y153_B;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X20Y153_B1;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X20Y153_B2;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X20Y153_B3;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X20Y153_B4;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X20Y153_B5;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X20Y153_B6;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X20Y153_BO5;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X20Y153_BO6;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X20Y153_B_CY;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X20Y153_B_XOR;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X20Y153_C;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X20Y153_C1;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X20Y153_C2;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X20Y153_C3;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X20Y153_C4;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X20Y153_C5;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X20Y153_C6;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X20Y153_CO5;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X20Y153_CO6;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X20Y153_C_CY;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X20Y153_C_XOR;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X20Y153_D;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X20Y153_D1;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X20Y153_D2;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X20Y153_D3;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X20Y153_D4;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X20Y153_D5;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X20Y153_D6;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X20Y153_DO5;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X20Y153_DO6;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X20Y153_D_CY;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X20Y153_D_XOR;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X21Y153_A;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X21Y153_A1;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X21Y153_A2;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X21Y153_A3;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X21Y153_A4;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X21Y153_A5;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X21Y153_A6;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X21Y153_AO5;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X21Y153_AO6;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X21Y153_A_CY;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X21Y153_A_XOR;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X21Y153_B;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X21Y153_B1;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X21Y153_B2;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X21Y153_B3;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X21Y153_B4;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X21Y153_B5;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X21Y153_B6;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X21Y153_BO5;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X21Y153_BO6;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X21Y153_B_CY;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X21Y153_B_XOR;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X21Y153_C;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X21Y153_C1;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X21Y153_C2;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X21Y153_C3;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X21Y153_C4;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X21Y153_C5;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X21Y153_C6;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X21Y153_CO5;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X21Y153_CO6;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X21Y153_C_CY;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X21Y153_C_XOR;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X21Y153_D;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X21Y153_D1;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X21Y153_D2;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X21Y153_D3;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X21Y153_D4;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X21Y153_D5;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X21Y153_D6;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X21Y153_DO5;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X21Y153_DO6;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X21Y153_D_CY;
  wire [0:0] CLBLM_R_X15Y153_SLICE_X21Y153_D_XOR;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_A;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_A1;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_A2;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_A3;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_A4;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_A5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_A6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_AO5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_AO6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_A_CY;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_A_XOR;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_B;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_B1;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_B2;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_B3;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_B4;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_B5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_B6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_BO5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_BO6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_B_CY;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_B_XOR;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_C;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_C1;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_C2;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_C3;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_C4;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_C5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_C6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_CO5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_CO6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_C_CY;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_C_XOR;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_D;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_D1;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_D2;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_D3;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_D4;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_D5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_D6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_DO5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_DO6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_D_CY;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_D_XOR;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_A;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_A1;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_A2;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_A3;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_A4;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_A5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_A6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_AO5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_AO6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_A_CY;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_A_XOR;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_B;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_B1;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_B2;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_B3;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_B4;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_B5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_B6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_BO5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_BO6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_B_CY;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_B_XOR;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_C;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_C1;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_C2;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_C3;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_C4;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_C5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_C6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_CO5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_CO6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_C_CY;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_C_XOR;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_D;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_D1;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_D2;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_D3;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_D4;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_D5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_D6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_DO5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_DO6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_D_CY;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_D_XOR;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_A;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_A1;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_A2;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_A3;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_A4;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_A5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_A6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_AO5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_AO6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_AQ;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_A_CY;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_A_XOR;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_B;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_B1;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_B2;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_B3;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_B4;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_B5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_B6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_BO5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_BO6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_BQ;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_B_CY;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_B_XOR;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_C;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_C1;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_C2;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_C3;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_C4;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_C5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_C6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_CLK;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_CO5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_CO6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_CQ;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_C_CY;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_C_XOR;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_D;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_D1;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_D2;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_D3;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_D4;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_D5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_D6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_DMUX;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_DO5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_DO6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_D_CY;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_D_XOR;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_A;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_A1;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_A2;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_A3;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_A4;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_A5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_A6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_AO5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_AO6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_A_CY;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_A_XOR;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_B;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_B1;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_B2;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_B3;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_B4;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_B5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_B6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_BO5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_BO6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_B_CY;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_B_XOR;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_C;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_C1;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_C2;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_C3;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_C4;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_C5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_C6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_CO5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_CO6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_C_CY;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_C_XOR;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_D;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_D1;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_D2;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_D3;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_D4;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_D5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_D6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_DO5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_DO6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_D_CY;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_D_XOR;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_A;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_A1;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_A2;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_A3;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_A4;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_A5;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_A6;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_AO5;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_AO6;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_AQ;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_A_CY;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_A_XOR;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_B;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_B1;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_B2;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_B3;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_B4;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_B5;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_B6;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_BO5;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_BO6;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_BQ;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_B_CY;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_B_XOR;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_C;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_C1;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_C2;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_C3;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_C4;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_C5;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_C6;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_CLK;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_CO5;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_CO6;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_CQ;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_C_CY;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_C_XOR;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_D;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_D1;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_D2;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_D3;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_D4;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_D5;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_D6;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_DO5;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_DO6;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_DQ;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_D_CY;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_D_XOR;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_A;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_A1;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_A2;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_A3;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_A4;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_A5;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_A5Q;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_A6;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_AMUX;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_AO5;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_AO6;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_AQ;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_AX;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_A_CY;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_A_XOR;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_B;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_B1;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_B2;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_B3;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_B4;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_B5;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_B5Q;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_B6;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_BMUX;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_BO5;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_BO6;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_BQ;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_BX;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_B_CY;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_B_XOR;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_C;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_C1;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_C2;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_C3;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_C4;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_C5;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_C6;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_CLK;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_CMUX;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_CO5;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_CO6;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_C_CY;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_C_XOR;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_D;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_D1;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_D2;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_D3;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_D4;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_D5;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_D6;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_DMUX;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_DO5;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_DO6;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_D_CY;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_D_XOR;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_A;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_A1;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_A2;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_A3;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_A4;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_A5;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_A5Q;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_A6;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_AMUX;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_AO5;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_AO6;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_AQ;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_A_CY;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_A_XOR;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_B;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_B1;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_B2;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_B3;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_B4;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_B5;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_B5Q;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_B6;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_BMUX;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_BO5;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_BO6;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_BQ;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_B_CY;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_B_XOR;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_C;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_C1;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_C2;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_C3;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_C4;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_C5;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_C6;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_CLK;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_CO5;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_CO6;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_C_CY;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_C_XOR;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_D;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_D1;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_D2;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_D3;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_D4;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_D5;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_D6;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_DO5;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_DO6;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_D_CY;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_D_XOR;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_A;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_A1;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_A2;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_A3;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_A4;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_A5;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_A6;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_AO5;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_AO6;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_AQ;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_A_CY;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_A_XOR;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_B;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_B1;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_B2;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_B3;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_B4;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_B5;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_B6;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_BMUX;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_BO5;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_BO6;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_B_CY;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_B_XOR;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_C;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_C1;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_C2;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_C3;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_C4;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_C5;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_C6;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_CLK;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_CO5;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_CO6;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_C_CY;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_C_XOR;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_D;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_D1;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_D2;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_D3;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_D4;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_D5;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_D6;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_DO5;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_DO6;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_D_CY;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_D_XOR;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_A;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_A1;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_A2;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_A3;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_A4;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_A5;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_A5Q;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_A6;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_AMUX;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_AO5;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_AO6;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_AQ;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_AX;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_A_CY;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_A_XOR;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_B;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_B1;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_B2;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_B3;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_B4;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_B5;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_B6;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_BO5;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_BO6;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_BQ;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_B_CY;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_B_XOR;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_C;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_C1;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_C2;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_C3;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_C4;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_C5;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_C6;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_CLK;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_CMUX;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_CO5;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_CO6;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_C_CY;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_C_XOR;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_D;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_D1;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_D2;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_D3;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_D4;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_D5;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_D6;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_DO5;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_DO6;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_D_CY;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_D_XOR;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_A;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_A1;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_A2;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_A3;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_A4;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_A5;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_A5Q;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_A6;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_AMUX;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_AO5;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_AO6;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_AQ;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_A_CY;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_A_XOR;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_B;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_B1;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_B2;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_B3;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_B4;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_B5;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_B6;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_BO5;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_BO6;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_BQ;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_B_CY;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_B_XOR;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_C;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_C1;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_C2;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_C3;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_C4;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_C5;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_C6;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_CLK;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_CO5;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_CO6;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_CQ;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_C_CY;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_C_XOR;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_D;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_D1;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_D2;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_D3;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_D4;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_D5;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_D5Q;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_D6;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_DMUX;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_DO5;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_DO6;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_DQ;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_D_CY;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_D_XOR;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_A;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_A1;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_A2;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_A3;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_A4;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_A5;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_A6;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_AO5;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_AO6;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_AQ;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_A_CY;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_A_XOR;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_B;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_B1;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_B2;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_B3;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_B4;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_B5;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_B6;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_BO5;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_BO6;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_BQ;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_B_CY;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_B_XOR;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_C;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_C1;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_C2;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_C3;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_C4;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_C5;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_C6;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_CLK;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_CO5;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_CO6;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_C_CY;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_C_XOR;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_D;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_D1;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_D2;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_D3;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_D4;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_D5;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_D6;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_DO5;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_DO6;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_D_CY;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_D_XOR;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_A;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_A1;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_A2;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_A3;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_A4;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_A5;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_A6;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_AO5;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_AO6;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_AQ;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_A_CY;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_A_XOR;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_B;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_B1;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_B2;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_B3;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_B4;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_B5;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_B6;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_BO5;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_BO6;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_BQ;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_B_CY;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_B_XOR;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_C;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_C1;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_C2;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_C3;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_C4;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_C5;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_C6;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_CLK;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_CO5;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_CO6;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_CQ;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_C_CY;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_C_XOR;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_D;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_D1;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_D2;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_D3;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_D4;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_D5;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_D6;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_DMUX;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_DO5;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_DO6;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_D_CY;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_D_XOR;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_A;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_A1;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_A2;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_A3;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_A4;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_A5;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_A5Q;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_A6;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_AMUX;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_AO5;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_AO6;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_AQ;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_AX;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_A_CY;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_A_XOR;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_B;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_B1;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_B2;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_B3;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_B4;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_B5;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_B6;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_BMUX;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_BO5;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_BO6;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_B_CY;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_B_XOR;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_C;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_C1;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_C2;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_C3;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_C4;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_C5;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_C6;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_CLK;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_CO5;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_CO6;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_CQ;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_C_CY;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_C_XOR;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_D;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_D1;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_D2;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_D3;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_D4;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_D5;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_D6;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_DO5;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_DO6;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_DQ;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_D_CY;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_D_XOR;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_A;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_A1;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_A2;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_A3;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_A4;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_A5;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_A6;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_AO5;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_AO6;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_AQ;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_A_CY;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_A_XOR;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_B;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_B1;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_B2;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_B3;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_B4;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_B5;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_B6;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_BO5;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_BO6;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_BQ;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_B_CY;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_B_XOR;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_C;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_C1;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_C2;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_C3;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_C4;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_C5;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_C5Q;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_C6;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_CLK;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_CMUX;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_CO5;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_CO6;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_CQ;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_C_CY;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_C_XOR;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_D;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_D1;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_D2;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_D3;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_D4;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_D5;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_D6;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_DO5;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_DO6;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_DQ;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_D_CY;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_D_XOR;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_A;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_A1;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_A2;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_A3;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_A4;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_A5;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_A6;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_AMUX;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_AO5;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_AO6;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_AQ;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_A_CY;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_A_XOR;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_B;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_B1;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_B2;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_B3;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_B4;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_B5;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_B6;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_BO5;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_BO6;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_BQ;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_B_CY;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_B_XOR;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_C;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_C1;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_C2;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_C3;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_C4;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_C5;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_C6;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_CLK;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_CO5;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_CO6;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_CQ;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_C_CY;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_C_XOR;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_D;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_D1;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_D2;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_D3;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_D4;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_D5;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_D6;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_DO5;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_DO6;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_DQ;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_D_CY;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_D_XOR;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_A;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_A1;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_A2;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_A3;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_A4;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_A5;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_A6;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_AO5;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_AO6;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_AQ;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_A_CY;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_A_XOR;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_B;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_B1;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_B2;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_B3;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_B4;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_B5;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_B5Q;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_B6;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_BMUX;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_BO5;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_BO6;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_BQ;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_B_CY;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_B_XOR;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_C;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_C1;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_C2;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_C3;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_C4;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_C5;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_C6;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_CLK;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_CO5;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_CO6;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_CQ;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_C_CY;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_C_XOR;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_D;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_D1;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_D2;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_D3;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_D4;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_D5;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_D6;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_DMUX;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_DO5;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_DO6;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_D_CY;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_D_XOR;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_A;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_A1;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_A2;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_A3;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_A4;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_A5;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_A6;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_AO5;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_AO6;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_AQ;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_A_CY;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_A_XOR;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_B;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_B1;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_B2;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_B3;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_B4;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_B5;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_B6;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_BO5;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_BO6;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_BQ;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_B_CY;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_B_XOR;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_C;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_C1;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_C2;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_C3;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_C4;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_C5;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_C6;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_CLK;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_CO5;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_CO6;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_CQ;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_C_CY;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_C_XOR;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_D;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_D1;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_D2;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_D3;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_D4;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_D5;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_D6;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_DO5;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_DO6;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_D_CY;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_D_XOR;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_A;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_A1;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_A2;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_A3;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_A4;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_A5;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_A6;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_AO5;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_AO6;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_AQ;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_A_CY;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_A_XOR;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_B;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_B1;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_B2;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_B3;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_B4;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_B5;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_B5Q;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_B6;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_BMUX;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_BO5;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_BO6;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_BQ;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_B_CY;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_B_XOR;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_C;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_C1;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_C2;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_C3;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_C4;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_C5;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_C6;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_CLK;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_CO5;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_CO6;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_CQ;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_C_CY;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_C_XOR;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_D;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_D1;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_D2;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_D3;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_D4;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_D5;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_D6;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_DO5;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_DO6;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_DQ;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_D_CY;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_D_XOR;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_A;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_A1;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_A2;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_A3;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_A4;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_A5;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_A6;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_AO5;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_AO6;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_A_CY;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_A_XOR;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_B;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_B1;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_B2;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_B3;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_B4;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_B5;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_B6;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_BO5;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_BO6;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_B_CY;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_B_XOR;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_C;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_C1;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_C2;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_C3;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_C4;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_C5;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_C6;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_CO5;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_CO6;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_C_CY;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_C_XOR;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_D;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_D1;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_D2;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_D3;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_D4;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_D5;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_D6;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_DO5;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_DO6;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_D_CY;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_D_XOR;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_A;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_A1;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_A2;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_A3;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_A4;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_A5;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_A5Q;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_A6;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_AMUX;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_AO5;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_AQ;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_A_CY;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_A_XOR;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_B;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_B1;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_B2;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_B3;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_B4;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_B5;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_B6;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_BO5;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_BO6;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_BQ;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_B_CY;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_B_XOR;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_C;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_C1;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_C2;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_C3;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_C4;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_C5;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_C6;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_CLK;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_CO5;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_CO6;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_C_CY;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_C_XOR;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_D;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_D1;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_D2;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_D3;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_D4;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_D5;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_D6;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_DO5;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_DO6;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_D_CY;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_D_XOR;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_A;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_A1;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_A2;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_A3;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_A4;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_A5;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_A6;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_AO5;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_AO6;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_A_CY;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_A_XOR;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_B;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_B1;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_B2;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_B3;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_B4;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_B5;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_B6;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_BO5;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_BO6;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_B_CY;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_B_XOR;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_C;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_C1;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_C2;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_C3;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_C4;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_C5;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_C6;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_CMUX;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_CO5;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_CO6;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_C_CY;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_C_XOR;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_D;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_D1;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_D2;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_D3;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_D4;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_D5;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_D6;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_DO5;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_DO6;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_D_CY;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_D_XOR;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_A;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_A1;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_A2;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_A3;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_A4;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_A5;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_A6;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_AO5;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_AO6;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_A_CY;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_A_XOR;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_B;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_B1;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_B2;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_B3;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_B4;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_B5;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_B6;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_BO5;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_BO6;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_B_CY;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_B_XOR;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_C;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_C1;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_C2;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_C3;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_C4;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_C5;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_C6;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_CO5;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_CO6;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_C_CY;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_C_XOR;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_D;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_D1;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_D2;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_D3;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_D4;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_D5;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_D6;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_DO5;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_DO6;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_D_CY;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_D_XOR;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_A;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_A1;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_A2;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_A3;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_A4;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_A5;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_A6;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_AMUX;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_AO5;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_AO6;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_A_CY;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_A_XOR;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_B;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_B1;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_B2;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_B3;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_B4;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_B5;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_B6;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_BMUX;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_BO5;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_BO6;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_B_CY;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_B_XOR;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_C;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_C1;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_C2;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_C3;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_C4;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_C5;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_C6;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_CO5;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_CO6;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_C_CY;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_C_XOR;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_D;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_D1;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_D2;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_D3;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_D4;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_D5;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_D6;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_DO5;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_DO6;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_D_CY;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_D_XOR;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_A;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_A1;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_A2;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_A3;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_A4;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_A5;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_A6;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_AO5;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_AO6;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_A_CY;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_A_XOR;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_B;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_B1;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_B2;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_B3;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_B4;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_B5;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_B6;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_BO5;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_BO6;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_B_CY;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_B_XOR;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_C;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_C1;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_C2;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_C3;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_C4;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_C5;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_C6;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_CMUX;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_CO5;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_CO6;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_C_CY;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_C_XOR;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_D;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_D1;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_D2;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_D3;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_D4;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_D5;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_D6;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_DO5;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_DO6;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_D_CY;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_D_XOR;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_A;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_A1;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_A2;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_A3;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_A4;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_A5;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_A6;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_AO5;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_AO6;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_A_CY;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_A_XOR;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_B;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_B1;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_B2;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_B3;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_B4;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_B5;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_B6;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_BO5;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_BO6;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_B_CY;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_B_XOR;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_C;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_C1;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_C2;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_C3;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_C4;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_C5;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_C6;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_CO5;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_CO6;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_C_CY;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_C_XOR;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_D;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_D1;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_D2;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_D3;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_D4;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_D5;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_D6;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_DO5;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_DO6;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_D_CY;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_D_XOR;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_A;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_A1;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_A2;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_A3;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_A4;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_A5;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_A6;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_AO5;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_AO6;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_A_CY;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_A_XOR;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_B;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_B1;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_B2;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_B3;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_B4;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_B5;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_B6;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_BO5;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_BO6;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_B_CY;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_B_XOR;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_C;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_C1;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_C2;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_C3;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_C4;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_C5;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_C6;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_CMUX;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_CO5;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_CO6;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_C_CY;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_C_XOR;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_D;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_D1;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_D2;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_D3;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_D4;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_D5;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_D6;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_DO5;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_DO6;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_D_CY;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_D_XOR;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_A;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_A1;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_A2;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_A3;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_A4;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_A5;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_A6;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_AO5;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_AO6;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_A_CY;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_A_XOR;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_B;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_B1;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_B2;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_B3;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_B4;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_B5;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_B6;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_BO5;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_BO6;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_B_CY;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_B_XOR;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_C;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_C1;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_C2;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_C3;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_C4;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_C5;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_C6;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_CO5;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_CO6;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_C_CY;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_C_XOR;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_D;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_D1;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_D2;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_D3;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_D4;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_D5;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_D6;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_DO5;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_DO6;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_D_CY;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_D_XOR;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_A;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_A1;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_A2;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_A3;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_A4;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_A5;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_A6;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_AO5;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_AO6;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_A_CY;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_A_XOR;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_B;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_B1;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_B2;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_B3;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_B4;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_B5;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_B6;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_BO5;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_BO6;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_B_CY;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_B_XOR;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_C;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_C1;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_C2;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_C3;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_C4;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_C5;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_C6;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_CMUX;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_CO5;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_CO6;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_C_CY;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_C_XOR;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_D;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_D1;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_D2;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_D3;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_D4;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_D5;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_D6;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_DO5;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_DO6;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_D_CY;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_D_XOR;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_A;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_A1;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_A2;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_A3;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_A4;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_A5;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_A6;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_AO5;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_AO6;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_A_CY;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_A_XOR;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_B;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_B1;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_B2;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_B3;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_B4;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_B5;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_B6;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_BO5;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_BO6;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_B_CY;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_B_XOR;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_C;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_C1;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_C2;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_C3;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_C4;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_C5;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_C6;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_CO5;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_CO6;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_C_CY;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_C_XOR;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_D;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_D1;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_D2;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_D3;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_D4;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_D5;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_D6;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_DMUX;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_DO5;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_DO6;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_D_CY;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_D_XOR;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_A;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_A1;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_A2;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_A3;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_A4;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_A5;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_A6;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_AMUX;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_AO5;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_AO6;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_A_CY;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_A_XOR;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_B;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_B1;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_B2;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_B3;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_B4;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_B5;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_B6;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_BO5;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_BO6;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_B_CY;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_B_XOR;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_C;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_C1;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_C2;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_C3;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_C4;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_C5;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_C6;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_CMUX;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_CO5;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_CO6;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_C_CY;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_C_XOR;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_D;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_D1;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_D2;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_D3;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_D4;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_D5;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_D6;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_DO5;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_DO6;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_D_CY;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_D_XOR;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_A;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_A1;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_A2;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_A3;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_A4;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_A5;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_A6;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_AMUX;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_AO5;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_AO6;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_A_CY;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_A_XOR;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_B;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_B1;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_B2;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_B3;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_B4;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_B5;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_B6;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_BO5;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_BO6;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_B_CY;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_B_XOR;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_C;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_C1;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_C2;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_C3;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_C4;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_C5;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_C6;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_CO5;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_CO6;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_C_CY;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_C_XOR;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_D;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_D1;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_D2;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_D3;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_D4;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_D5;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_D6;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_DO5;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_DO6;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_D_CY;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_D_XOR;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_A;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_A1;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_A2;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_A3;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_A4;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_A5;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_A6;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_AO5;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_AO6;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_A_CY;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_A_XOR;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_B;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_B1;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_B2;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_B3;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_B4;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_B5;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_B6;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_BO5;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_BO6;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_B_CY;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_B_XOR;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_C;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_C1;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_C2;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_C3;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_C4;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_C5;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_C6;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_CO5;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_CO6;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_C_CY;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_C_XOR;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_D;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_D1;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_D2;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_D3;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_D4;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_D5;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_D6;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_DO5;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_DO6;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_D_CY;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_D_XOR;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_A;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_A1;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_A2;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_A3;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_A4;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_A5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_A6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_AO5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_AO6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_A_CY;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_A_XOR;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_B;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_B1;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_B2;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_B3;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_B4;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_B5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_B6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_BO5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_BO6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_B_CY;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_B_XOR;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_C;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_C1;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_C2;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_C3;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_C4;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_C5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_C6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_CO5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_CO6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_C_CY;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_C_XOR;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_D;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_D1;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_D2;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_D3;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_D4;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_D5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_D6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_DO5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_DO6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_D_CY;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_D_XOR;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_A;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_A1;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_A2;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_A3;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_A4;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_A5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_A6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_AO5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_AO6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_AQ;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_AX;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_A_CY;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_A_XOR;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_B;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_B1;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_B2;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_B3;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_B4;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_B5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_B6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_BO5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_BO6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_B_CY;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_B_XOR;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_C;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_C1;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_C2;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_C3;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_C4;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_C5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_C6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_CLK;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_CO5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_CO6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_C_CY;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_C_XOR;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_D;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_D1;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_D2;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_D3;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_D4;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_D5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_D6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_DO5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_DO6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_D_CY;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_D_XOR;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_A;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_A1;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_A2;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_A3;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_A4;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_A5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_A6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_AO5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_AO6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_AQ;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_A_CY;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_A_XOR;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_B;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_B1;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_B2;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_B3;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_B4;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_B5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_B6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_BO5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_BO6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_B_CY;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_B_XOR;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_C;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_C1;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_C2;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_C3;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_C4;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_C5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_C6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_CLK;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_CO5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_CO6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_C_CY;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_C_XOR;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_D;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_D1;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_D2;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_D3;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_D4;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_D5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_D6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_DO5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_DO6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_D_CY;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_D_XOR;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_A;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_A1;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_A2;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_A3;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_A4;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_A5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_A6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_AO5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_AO6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_AQ;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_A_CY;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_A_XOR;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_B;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_B1;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_B2;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_B3;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_B4;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_B5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_B6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_BMUX;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_BO5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_BO6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_B_CY;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_B_XOR;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_C;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_C1;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_C2;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_C3;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_C4;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_C5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_C6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_CLK;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_CO5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_CO6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_C_CY;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_C_XOR;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_D;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_D1;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_D2;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_D3;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_D4;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_D5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_D6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_DO5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_DO6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_D_CY;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_D_XOR;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_A;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_A1;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_A2;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_A3;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_A4;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_A5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_A6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_AO5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_AO6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_AQ;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_A_CY;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_A_XOR;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_B;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_B1;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_B2;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_B3;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_B4;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_B5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_B6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_BMUX;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_BO5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_BO6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_B_CY;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_B_XOR;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_C;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_C1;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_C2;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_C3;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_C4;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_C5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_C6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_CLK;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_CO5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_CO6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_C_CY;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_C_XOR;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_D;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_D1;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_D2;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_D3;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_D4;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_D5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_D6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_DO5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_DO6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_D_CY;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_D_XOR;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_A;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_A1;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_A2;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_A3;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_A4;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_A5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_A6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_AO5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_AO6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_AQ;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_A_CY;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_A_XOR;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_B;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_B1;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_B2;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_B3;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_B4;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_B5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_B5Q;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_B6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_BMUX;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_BO5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_BO6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_BQ;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_B_CY;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_B_XOR;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_C;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_C1;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_C2;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_C3;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_C4;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_C5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_C6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_CLK;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_CO5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_CO6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_CQ;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_C_CY;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_C_XOR;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_D;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_D1;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_D2;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_D3;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_D4;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_D5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_D6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_DO5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_DO6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_D_CY;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_D_XOR;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_A;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_A1;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_A2;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_A3;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_A4;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_A5;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_A5Q;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_A6;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_AMUX;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_AO5;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_AO6;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_AQ;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_AX;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_A_CY;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_A_XOR;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_B;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_B1;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_B2;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_B3;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_B4;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_B5;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_B6;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_BMUX;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_BO5;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_BO6;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_B_CY;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_B_XOR;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_C;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_C1;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_C2;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_C3;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_C4;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_C5;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_C6;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_CLK;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_CO5;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_CO6;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_CQ;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_C_CY;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_C_XOR;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_D;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_D1;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_D2;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_D3;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_D4;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_D5;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_D6;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_DMUX;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_DO5;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_DO6;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_D_CY;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_D_XOR;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_A;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_A1;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_A2;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_A3;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_A4;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_A5;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_A6;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_AO5;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_AO6;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_AQ;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_A_CY;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_A_XOR;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_B;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_B1;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_B2;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_B3;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_B4;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_B5;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_B6;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_BO5;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_BO6;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_BQ;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_B_CY;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_B_XOR;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_C;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_C1;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_C2;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_C3;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_C4;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_C5;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_C6;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_CLK;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_CO5;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_CO6;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_CQ;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_C_CY;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_C_XOR;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_D;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_D1;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_D2;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_D3;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_D4;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_D5;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_D6;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_DMUX;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_DO5;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_DO6;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_D_CY;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_D_XOR;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_A;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_A1;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_A2;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_A3;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_A4;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_A5;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_A5Q;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_A6;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_AMUX;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_AO5;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_AO6;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_AQ;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_AX;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_A_CY;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_A_XOR;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_B;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_B1;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_B2;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_B3;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_B4;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_B5;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_B6;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_BMUX;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_BO5;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_BO6;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_B_CY;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_B_XOR;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_C;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_C1;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_C2;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_C3;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_C4;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_C5;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_C6;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_CLK;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_CO5;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_CO6;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_CQ;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_C_CY;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_C_XOR;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_D;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_D1;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_D2;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_D3;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_D4;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_D5;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_D6;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_DO5;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_DO6;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_DQ;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_D_CY;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_D_XOR;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_A;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_A1;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_A2;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_A3;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_A4;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_A5;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_A6;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_AMUX;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_AO5;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_AO6;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_A_CY;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_A_XOR;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_B;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_B1;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_B2;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_B3;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_B4;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_B5;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_B6;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_BO5;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_BO6;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_B_CY;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_B_XOR;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_C;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_C1;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_C2;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_C3;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_C4;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_C5;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_C6;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_CMUX;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_CO5;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_CO6;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_C_CY;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_C_XOR;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_D;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_D1;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_D2;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_D3;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_D4;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_D5;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_D6;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_DMUX;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_DO5;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_DO6;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_D_CY;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_D_XOR;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_A;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_A1;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_A2;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_A3;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_A4;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_A5;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_A6;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_AO5;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_AO6;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_AQ;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_A_CY;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_A_XOR;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_B;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_B1;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_B2;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_B3;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_B4;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_B5;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_B6;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_BO5;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_BO6;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_BQ;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_B_CY;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_B_XOR;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_C;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_C1;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_C2;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_C3;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_C4;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_C5;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_C6;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_CLK;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_CO5;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_CO6;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_CQ;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_C_CY;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_C_XOR;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_D;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_D1;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_D2;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_D3;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_D4;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_D5;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_D6;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_DO5;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_DO6;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_D_CY;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_D_XOR;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_A;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_A1;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_A2;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_A3;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_A4;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_A5;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_A6;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_AO5;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_AO6;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_AQ;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_A_CY;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_A_XOR;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_B;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_B1;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_B2;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_B3;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_B4;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_B5;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_B6;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_BO5;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_BO6;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_BQ;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_B_CY;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_B_XOR;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_C;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_C1;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_C2;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_C3;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_C4;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_C5;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_C6;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_CLK;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_CO5;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_CO6;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_CQ;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_C_CY;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_C_XOR;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_D;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_D1;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_D2;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_D3;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_D4;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_D5;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_D5Q;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_D6;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_DMUX;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_DO5;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_DO6;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_DQ;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_D_CY;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_D_XOR;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_A;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_A1;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_A2;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_A3;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_A4;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_A5;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_A6;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_AO5;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_AO6;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_AQ;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_A_CY;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_A_XOR;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_B;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_B1;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_B2;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_B3;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_B4;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_B5;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_B6;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_BO5;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_BO6;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_BQ;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_B_CY;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_B_XOR;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_C;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_C1;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_C2;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_C3;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_C4;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_C5;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_C6;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_CLK;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_CO5;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_CO6;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_C_CY;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_C_XOR;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_D;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_D1;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_D2;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_D3;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_D4;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_D5;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_D6;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_DO5;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_DO6;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_D_CY;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_D_XOR;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_A;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_A1;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_A2;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_A3;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_A4;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_A5;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_A6;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_AO5;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_AO6;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_AQ;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_A_CY;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_A_XOR;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_B;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_B1;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_B2;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_B3;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_B4;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_B5;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_B6;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_BO5;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_BO6;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_BQ;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_B_CY;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_B_XOR;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_C;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_C1;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_C2;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_C3;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_C4;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_C5;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_C5Q;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_C6;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_CLK;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_CMUX;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_CO5;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_CO6;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_CQ;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_C_CY;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_C_XOR;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_D;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_D1;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_D2;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_D3;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_D4;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_D5;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_D6;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_DO5;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_DO6;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_D_CY;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_D_XOR;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_A;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_A1;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_A2;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_A3;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_A4;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_A5;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_A6;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_AO5;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_AO6;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_AQ;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_A_CY;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_A_XOR;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_B;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_B1;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_B2;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_B3;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_B4;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_B5;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_B6;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_BO5;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_BO6;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_BQ;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_B_CY;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_B_XOR;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_C;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_C1;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_C2;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_C3;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_C4;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_C5;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_C6;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_CLK;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_CMUX;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_CO5;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_CO6;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_C_CY;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_C_XOR;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_D;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_D1;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_D2;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_D3;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_D4;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_D5;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_D6;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_DO5;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_DO6;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_D_CY;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_D_XOR;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_A;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_A1;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_A2;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_A3;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_A4;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_A5;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_A6;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_AO5;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_AO6;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_AQ;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_A_CY;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_A_XOR;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_B;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_B1;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_B2;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_B3;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_B4;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_B5;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_B6;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_BO5;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_BO6;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_BQ;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_B_CY;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_B_XOR;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_C;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_C1;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_C2;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_C3;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_C4;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_C5;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_C6;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_CLK;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_CO5;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_CO6;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_CQ;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_C_CY;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_C_XOR;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_D;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_D1;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_D2;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_D3;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_D4;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_D5;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_D6;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_DO5;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_DO6;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_D_CY;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_D_XOR;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_A;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_A1;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_A2;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_A3;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_A4;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_A5;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_A5Q;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_A6;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_AMUX;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_AO5;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_AO6;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_AQ;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_A_CY;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_A_XOR;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_B;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_B1;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_B2;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_B3;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_B4;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_B5;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_B6;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_BO5;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_BO6;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_BQ;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_B_CY;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_B_XOR;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_C;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_C1;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_C2;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_C3;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_C4;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_C5;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_C6;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_CLK;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_CO5;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_CO6;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_CQ;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_C_CY;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_C_XOR;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_D;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_D1;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_D2;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_D3;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_D4;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_D5;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_D6;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_DO5;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_DO6;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_DQ;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_D_CY;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_D_XOR;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_A;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_A1;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_A2;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_A3;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_A4;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_A5;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_A6;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_AO5;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_AO6;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_AQ;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_A_CY;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_A_XOR;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_B;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_B1;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_B2;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_B3;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_B4;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_B5;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_B6;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_BO5;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_BO6;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_BQ;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_B_CY;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_B_XOR;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_C;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_C1;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_C2;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_C3;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_C4;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_C5;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_C6;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_CLK;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_CO5;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_CO6;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_C_CY;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_C_XOR;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_D;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_D1;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_D2;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_D3;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_D4;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_D5;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_D6;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_DMUX;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_DO5;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_DO6;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_D_CY;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_D_XOR;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_A;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_A1;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_A2;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_A3;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_A4;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_A5;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_A6;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_AO5;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_AO6;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_AQ;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_A_CY;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_A_XOR;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_B;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_B1;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_B2;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_B3;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_B4;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_B5;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_B6;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_BO5;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_BO6;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_BQ;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_B_CY;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_B_XOR;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_C;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_C1;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_C2;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_C3;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_C4;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_C5;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_C6;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_CLK;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_CO5;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_CO6;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_CQ;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_C_CY;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_C_XOR;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_D;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_D1;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_D2;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_D3;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_D4;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_D5;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_D6;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_DO5;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_DO6;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_DQ;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_D_CY;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_D_XOR;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_A;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_A1;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_A2;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_A3;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_A4;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_A5;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_A6;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_AO5;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_AO6;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_AQ;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_A_CY;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_A_XOR;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_B;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_B1;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_B2;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_B3;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_B4;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_B5;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_B6;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_BO5;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_BO6;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_BQ;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_B_CY;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_B_XOR;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_C;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_C1;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_C2;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_C3;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_C4;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_C5;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_C6;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_CLK;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_CO5;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_CO6;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_CQ;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_C_CY;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_C_XOR;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_D;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_D1;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_D2;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_D3;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_D4;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_D5;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_D6;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_DMUX;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_DO5;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_DO6;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_D_CY;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_D_XOR;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_A;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_A1;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_A2;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_A3;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_A4;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_A5;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_A5Q;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_A6;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_AMUX;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_AO5;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_AO6;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_AQ;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_AX;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_A_CY;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_A_XOR;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_B;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_B1;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_B2;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_B3;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_B4;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_B5;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_B6;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_BO5;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_BO6;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_BQ;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_B_CY;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_B_XOR;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_C;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_C1;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_C2;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_C3;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_C4;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_C5;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_C6;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_CLK;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_CO5;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_CO6;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_CQ;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_C_CY;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_C_XOR;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_D;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_D1;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_D2;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_D3;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_D4;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_D5;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_D6;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_DO5;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_DO6;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_D_CY;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_D_XOR;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_A;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_A1;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_A2;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_A3;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_A4;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_A5;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_A6;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_AO5;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_AO6;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_AQ;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_A_CY;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_A_XOR;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_B;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_B1;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_B2;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_B3;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_B4;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_B5;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_B5Q;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_B6;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_BMUX;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_BO5;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_BO6;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_BQ;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_B_CY;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_B_XOR;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_C;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_C1;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_C2;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_C3;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_C4;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_C5;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_C6;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_CLK;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_CO5;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_CO6;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_CQ;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_C_CY;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_C_XOR;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_D;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_D1;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_D2;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_D3;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_D4;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_D5;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_D6;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_DMUX;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_DO5;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_DO6;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_D_CY;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_D_XOR;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_A;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_A1;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_A2;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_A3;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_A4;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_A5;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_A5Q;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_A6;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_AMUX;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_AO5;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_AO6;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_AQ;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_AX;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_A_CY;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_A_XOR;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_B;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_B1;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_B2;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_B3;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_B4;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_B5;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_B6;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_BO5;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_BO6;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_BQ;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_B_CY;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_B_XOR;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_C;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_C1;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_C2;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_C3;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_C4;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_C5;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_C6;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_CLK;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_CMUX;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_CO5;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_CO6;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_C_CY;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_C_XOR;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_D;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_D1;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_D2;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_D3;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_D4;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_D5;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_D6;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_DO5;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_DO6;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_D_CY;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_D_XOR;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_A;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_A1;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_A2;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_A3;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_A4;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_A5;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_A6;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_AO5;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_AO6;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_AQ;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_A_CY;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_A_XOR;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_B;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_B1;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_B2;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_B3;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_B4;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_B5;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_B6;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_BO5;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_BO6;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_BQ;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_B_CY;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_B_XOR;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_C;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_C1;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_C2;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_C3;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_C4;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_C5;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_C6;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_CLK;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_CO5;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_CO6;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_C_CY;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_C_XOR;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_D;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_D1;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_D2;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_D3;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_D4;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_D5;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_D6;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_DO5;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_DO6;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_D_CY;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_D_XOR;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_A;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_A1;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_A2;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_A3;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_A4;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_A5;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_A6;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_AO5;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_AO6;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_AQ;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_A_CY;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_A_XOR;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_B;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_B1;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_B2;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_B3;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_B4;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_B5;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_B6;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_BO5;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_BO6;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_B_CY;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_B_XOR;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_C;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_C1;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_C2;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_C3;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_C4;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_C5;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_C6;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_CLK;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_CO5;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_CO6;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_C_CY;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_C_XOR;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_D;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_D1;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_D2;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_D3;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_D4;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_D5;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_D6;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_DO5;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_DO6;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_D_CY;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_D_XOR;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_A;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_A1;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_A2;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_A3;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_A4;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_A5;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_A6;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_AMUX;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_AO5;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_AO6;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_A_CY;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_A_XOR;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_B;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_B1;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_B2;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_B3;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_B4;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_B5;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_B6;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_BO5;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_BO6;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_B_CY;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_B_XOR;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_C;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_C1;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_C2;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_C3;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_C4;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_C5;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_C6;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_CO5;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_CO6;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_C_CY;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_C_XOR;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_D;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_D1;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_D2;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_D3;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_D4;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_D5;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_D6;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_DO5;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_DO6;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_D_CY;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_D_XOR;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X6Y155_A;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X6Y155_A1;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X6Y155_A2;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X6Y155_A3;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X6Y155_A4;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X6Y155_A5;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X6Y155_A6;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X6Y155_AO5;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X6Y155_AO6;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X6Y155_AQ;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X6Y155_A_CY;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X6Y155_A_XOR;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X6Y155_B;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X6Y155_B1;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X6Y155_B2;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X6Y155_B3;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X6Y155_B4;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X6Y155_B5;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X6Y155_B6;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X6Y155_BO5;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X6Y155_BO6;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X6Y155_BQ;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X6Y155_B_CY;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X6Y155_B_XOR;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X6Y155_C;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X6Y155_C1;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X6Y155_C2;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X6Y155_C3;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X6Y155_C4;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X6Y155_C5;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X6Y155_C6;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X6Y155_CLK;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X6Y155_CO5;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X6Y155_CO6;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X6Y155_C_CY;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X6Y155_C_XOR;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X6Y155_D;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X6Y155_D1;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X6Y155_D2;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X6Y155_D3;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X6Y155_D4;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X6Y155_D5;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X6Y155_D6;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X6Y155_DO5;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X6Y155_DO6;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X6Y155_D_CY;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X6Y155_D_XOR;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X7Y155_A;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X7Y155_A1;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X7Y155_A2;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X7Y155_A3;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X7Y155_A4;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X7Y155_A5;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X7Y155_A6;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X7Y155_AO5;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X7Y155_AO6;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X7Y155_AQ;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X7Y155_A_CY;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X7Y155_A_XOR;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X7Y155_B;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X7Y155_B1;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X7Y155_B2;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X7Y155_B3;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X7Y155_B4;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X7Y155_B5;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X7Y155_B6;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X7Y155_BMUX;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X7Y155_BO5;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X7Y155_BO6;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X7Y155_B_CY;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X7Y155_B_XOR;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X7Y155_C;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X7Y155_C1;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X7Y155_C2;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X7Y155_C3;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X7Y155_C4;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X7Y155_C5;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X7Y155_C6;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X7Y155_CLK;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X7Y155_CO5;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X7Y155_CO6;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X7Y155_C_CY;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X7Y155_C_XOR;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X7Y155_D;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X7Y155_D1;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X7Y155_D2;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X7Y155_D3;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X7Y155_D4;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X7Y155_D5;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X7Y155_D6;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X7Y155_DO5;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X7Y155_DO6;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X7Y155_D_CY;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X7Y155_D_XOR;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_A;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_A1;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_A2;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_A3;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_A4;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_A5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_A6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_AMUX;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_AO5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_AO6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_A_CY;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_A_XOR;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_B;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_B1;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_B2;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_B3;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_B4;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_B5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_B6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_BO5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_BO6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_BQ;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_B_CY;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_B_XOR;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_C;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_C1;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_C2;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_C3;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_C4;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_C5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_C6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_CLK;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_CO5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_CO6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_CQ;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_C_CY;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_C_XOR;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_D;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_D1;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_D2;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_D3;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_D4;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_D5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_D6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_DMUX;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_DO5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_DO6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_D_CY;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_D_XOR;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_A;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_A1;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_A2;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_A3;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_A4;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_A5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_A6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_AO5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_AO6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_A_CY;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_A_XOR;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_B;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_B1;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_B2;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_B3;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_B4;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_B5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_B6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_BO5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_BO6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_B_CY;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_B_XOR;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_C;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_C1;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_C2;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_C3;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_C4;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_C5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_C6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_CO5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_CO6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_C_CY;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_C_XOR;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_D;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_D1;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_D2;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_D3;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_D4;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_D5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_D6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_DO5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_DO6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_D_CY;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_D_XOR;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_A;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_A1;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_A2;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_A3;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_A4;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_A5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_A6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_AO5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_AO6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_AQ;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_A_CY;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_A_XOR;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_B;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_B1;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_B2;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_B3;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_B4;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_B5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_B5Q;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_B6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_BMUX;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_BO5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_BO6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_BQ;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_B_CY;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_B_XOR;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_C;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_C1;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_C2;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_C3;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_C4;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_C5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_C6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_CLK;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_CO5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_CO6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_CQ;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_C_CY;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_C_XOR;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_D;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_D1;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_D2;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_D3;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_D4;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_D5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_D6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_DO5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_DO6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_D_CY;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_D_XOR;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_A;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_A1;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_A2;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_A3;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_A4;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_A5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_A6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_AO5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_AO6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_AQ;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_A_CY;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_A_XOR;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_B;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_B1;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_B2;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_B3;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_B4;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_B5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_B6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_BO5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_BO6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_BQ;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_B_CY;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_B_XOR;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_C;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_C1;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_C2;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_C3;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_C4;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_C5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_C6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_CLK;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_CO5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_CO6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_CQ;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_C_CY;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_C_XOR;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_D;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_D1;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_D2;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_D3;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_D4;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_D5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_D6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_DO5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_DO6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_D_CY;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_D_XOR;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_A;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_A1;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_A2;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_A3;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_A4;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_A5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_A6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_AO5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_AO6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_AQ;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_A_CY;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_A_XOR;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_B;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_B1;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_B2;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_B3;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_B4;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_B5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_B6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_BO5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_BO6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_BQ;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_B_CY;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_B_XOR;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_C;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_C1;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_C2;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_C3;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_C4;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_C5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_C6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_CLK;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_CO5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_CO6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_CQ;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_C_CY;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_C_XOR;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_D;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_D1;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_D2;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_D3;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_D4;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_D5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_D6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_DO5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_DO6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_DQ;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_D_CY;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_D_XOR;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_A;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_A1;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_A2;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_A3;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_A4;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_A5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_A5Q;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_A6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_AMUX;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_AO5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_AO6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_AQ;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_AX;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_A_CY;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_A_XOR;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_B;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_B1;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_B2;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_B3;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_B4;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_B5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_B6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_BO5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_BO6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_BQ;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_B_CY;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_B_XOR;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_C;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_C1;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_C2;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_C3;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_C4;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_C5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_C6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_CLK;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_CO5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_CO6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_CQ;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_C_CY;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_C_XOR;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_D;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_D1;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_D2;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_D3;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_D4;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_D5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_D6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_DMUX;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_DO5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_DO6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_D_CY;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_D_XOR;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_A;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_A1;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_A2;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_A3;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_A4;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_A5;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_A6;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_AO5;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_AO6;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_AQ;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_A_CY;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_A_XOR;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_B;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_B1;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_B2;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_B3;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_B4;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_B5;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_B6;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_BO5;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_BO6;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_BQ;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_B_CY;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_B_XOR;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_C;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_C1;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_C2;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_C3;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_C4;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_C5;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_C5Q;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_C6;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_CLK;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_CMUX;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_CO5;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_CO6;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_CQ;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_C_CY;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_C_XOR;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_D;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_D1;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_D2;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_D3;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_D4;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_D5;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_D6;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_DMUX;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_DO5;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_DO6;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_D_CY;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_D_XOR;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_A;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_A1;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_A2;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_A3;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_A4;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_A5;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_A6;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_AO5;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_AO6;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_AQ;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_A_CY;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_A_XOR;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_B;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_B1;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_B2;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_B3;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_B4;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_B5;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_B6;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_BO5;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_BO6;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_BQ;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_B_CY;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_B_XOR;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_C;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_C1;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_C2;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_C3;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_C4;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_C5;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_C5Q;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_C6;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_CLK;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_CMUX;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_CO5;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_CO6;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_CQ;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_C_CY;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_C_XOR;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_D;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_D1;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_D2;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_D3;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_D4;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_D5;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_D6;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_DO5;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_DO6;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_D_CY;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_D_XOR;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_A;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_A1;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_A2;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_A3;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_A4;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_A5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_A6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_AO5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_AO6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_A_CY;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_A_XOR;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_B;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_B1;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_B2;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_B3;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_B4;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_B5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_B6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_BMUX;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_BO5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_BO6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_B_CY;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_B_XOR;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_C;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_C1;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_C2;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_C3;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_C4;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_C5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_C5Q;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_C6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_CLK;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_CMUX;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_CO5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_CO6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_CQ;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_C_CY;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_C_XOR;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_D;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_D1;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_D2;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_D3;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_D4;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_D5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_D6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_DO5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_DO6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_DQ;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_D_CY;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_D_XOR;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_A;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_A1;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_A2;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_A3;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_A4;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_A5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_A6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_AO5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_AO6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_AQ;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_A_CY;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_A_XOR;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_B;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_B1;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_B2;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_B3;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_B4;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_B5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_B6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_BO5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_BO6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_BQ;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_B_CY;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_B_XOR;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_C;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_C1;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_C2;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_C3;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_C4;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_C5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_C6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_CLK;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_CO5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_CO6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_CQ;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_C_CY;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_C_XOR;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_D;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_D1;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_D2;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_D3;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_D4;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_D5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_D6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_DO5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_DO6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_D_CY;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_D_XOR;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_A;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_A1;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_A2;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_A3;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_A4;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_A5;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_A6;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_AO5;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_AO6;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_AQ;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_A_CY;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_A_XOR;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_B;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_B1;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_B2;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_B3;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_B4;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_B5;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_B5Q;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_B6;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_BMUX;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_BO5;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_BO6;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_BQ;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_B_CY;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_B_XOR;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_C;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_C1;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_C2;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_C3;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_C4;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_C5;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_C5Q;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_C6;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_CLK;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_CMUX;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_CO5;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_CO6;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_CQ;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_C_CY;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_C_XOR;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_D;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_D1;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_D2;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_D3;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_D4;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_D5;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_D6;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_DO5;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_DO6;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_DQ;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_D_CY;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_D_XOR;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_A;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_A1;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_A2;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_A3;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_A4;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_A5;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_A6;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_AO5;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_AO6;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_AQ;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_A_CY;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_A_XOR;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_B;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_B1;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_B2;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_B3;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_B4;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_B5;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_B6;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_BO5;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_BO6;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_BQ;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_B_CY;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_B_XOR;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_C;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_C1;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_C2;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_C3;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_C4;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_C5;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_C6;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_CLK;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_CMUX;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_CO5;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_CO6;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_C_CY;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_C_XOR;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_D;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_D1;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_D2;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_D3;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_D4;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_D5;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_D6;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_DO5;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_DO6;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_D_CY;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_D_XOR;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_A;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_A1;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_A2;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_A3;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_A4;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_A5;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_A6;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_AO5;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_AO6;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_AQ;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_A_CY;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_A_XOR;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_B;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_B1;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_B2;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_B3;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_B4;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_B5;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_B6;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_BMUX;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_BO5;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_BO6;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_B_CY;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_B_XOR;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_C;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_C1;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_C2;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_C3;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_C4;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_C5;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_C6;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_CLK;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_CO5;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_CO6;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_CQ;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_C_CY;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_C_XOR;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_D;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_D1;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_D2;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_D3;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_D4;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_D5;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_D5Q;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_D6;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_DMUX;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_DO5;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_DO6;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_DQ;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_D_CY;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_D_XOR;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_A;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_A1;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_A2;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_A3;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_A4;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_A5;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_A6;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_AO5;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_AO6;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_AQ;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_A_CY;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_A_XOR;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_B;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_B1;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_B2;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_B3;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_B4;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_B5;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_B6;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_BO5;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_BO6;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_BQ;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_B_CY;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_B_XOR;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_C;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_C1;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_C2;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_C3;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_C4;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_C5;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_C6;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_CLK;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_CO5;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_CO6;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_CQ;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_C_CY;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_C_XOR;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_D;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_D1;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_D2;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_D3;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_D4;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_D5;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_D6;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_DO5;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_DO6;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_DQ;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_D_CY;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_D_XOR;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_A;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_A1;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_A2;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_A3;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_A4;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_A5;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_A6;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_AO5;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_AO6;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_AQ;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_A_CY;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_A_XOR;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_B;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_B1;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_B2;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_B3;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_B4;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_B5;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_B6;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_BO5;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_BO6;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_BQ;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_B_CY;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_B_XOR;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_C;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_C1;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_C2;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_C3;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_C4;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_C5;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_C6;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_CLK;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_CO5;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_CO6;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_CQ;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_C_CY;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_C_XOR;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_D;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_D1;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_D2;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_D3;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_D4;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_D5;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_D6;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_DO5;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_DO6;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_DQ;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_D_CY;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_D_XOR;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_A;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_A1;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_A2;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_A3;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_A4;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_A5;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_A6;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_AO5;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_AO6;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_A_CY;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_A_XOR;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_B;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_B1;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_B2;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_B3;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_B4;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_B5;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_B6;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_BO5;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_BO6;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_B_CY;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_B_XOR;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_C;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_C1;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_C2;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_C3;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_C4;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_C5;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_C6;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_CLK;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_CO5;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_CO6;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_C_CY;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_C_XOR;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_D;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_D1;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_D2;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_D3;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_D4;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_D5;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_D6;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_DO5;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_DO6;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_D_CY;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_D_XOR;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_A;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_A1;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_A2;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_A3;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_A4;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_A5;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_A6;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_AO5;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_AO6;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_AQ;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_A_CY;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_A_XOR;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_B;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_B1;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_B2;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_B3;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_B4;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_B5;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_B6;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_BO5;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_BO6;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_BQ;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_B_CY;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_B_XOR;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_C;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_C1;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_C2;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_C3;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_C4;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_C5;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_C6;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_CLK;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_CO5;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_CO6;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_CQ;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_C_CY;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_C_XOR;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_D;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_D1;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_D2;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_D3;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_D4;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_D5;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_D6;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_DO5;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_DO6;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_D_CY;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_D_XOR;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_A;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_A1;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_A2;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_A3;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_A4;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_A5;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_A5Q;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_A6;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_AMUX;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_AO5;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_AO6;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_AQ;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_AX;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_A_CY;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_A_XOR;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_B;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_B1;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_B2;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_B3;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_B4;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_B5;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_B6;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_BMUX;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_BO5;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_BO6;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_B_CY;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_B_XOR;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_C;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_C1;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_C2;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_C3;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_C4;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_C5;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_C6;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_CLK;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_CMUX;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_CO5;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_CO6;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_C_CY;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_C_XOR;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_D;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_D1;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_D2;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_D3;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_D4;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_D5;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_D6;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_DO5;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_DO6;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_D_CY;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_D_XOR;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_A;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_A1;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_A2;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_A3;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_A4;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_A5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_A5Q;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_A6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_AMUX;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_AO5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_AO6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_AQ;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_AX;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_A_CY;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_A_XOR;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_B;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_B1;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_B2;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_B3;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_B4;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_B5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_B6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_BO5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_BO6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_BQ;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_B_CY;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_B_XOR;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_C;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_C1;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_C2;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_C3;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_C4;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_C5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_C6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_CLK;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_CMUX;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_CO5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_CO6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_C_CY;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_C_XOR;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_D;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_D1;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_D2;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_D3;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_D4;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_D5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_D6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_DMUX;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_DO5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_DO6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_D_CY;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_D_XOR;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_A;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_A1;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_A2;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_A3;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_A4;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_A5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_A6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_AO5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_AO6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_AQ;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_A_CY;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_A_XOR;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_B;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_B1;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_B2;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_B3;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_B4;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_B5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_B6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_BO5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_BO6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_BQ;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_B_CY;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_B_XOR;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_C;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_C1;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_C2;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_C3;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_C4;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_C5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_C6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_CLK;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_CO5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_CO6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_CQ;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_C_CY;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_C_XOR;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_D;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_D1;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_D2;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_D3;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_D4;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_D5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_D6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_DMUX;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_DO5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_DO6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_D_CY;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_D_XOR;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_A;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_A1;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_A2;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_A3;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_A4;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_A5;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_A6;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_AO5;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_AO6;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_AQ;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_A_CY;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_A_XOR;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_B;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_B1;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_B2;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_B3;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_B4;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_B5;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_B6;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_BO5;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_BO6;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_BQ;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_B_CY;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_B_XOR;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_C;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_C1;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_C2;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_C3;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_C4;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_C5;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_C6;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_CLK;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_CO5;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_CO6;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_CQ;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_C_CY;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_C_XOR;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_D;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_D1;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_D2;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_D3;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_D4;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_D5;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_D6;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_DO5;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_DO6;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_DQ;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_D_CY;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_D_XOR;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_A;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_A1;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_A2;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_A3;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_A4;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_A5;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_A6;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_AO5;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_AO6;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_AQ;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_A_CY;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_A_XOR;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_B;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_B1;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_B2;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_B3;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_B4;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_B5;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_B6;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_BO5;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_BO6;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_BQ;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_B_CY;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_B_XOR;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_C;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_C1;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_C2;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_C3;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_C4;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_C5;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_C6;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_CLK;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_CO5;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_CO6;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_CQ;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_C_CY;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_C_XOR;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_D;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_D1;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_D2;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_D3;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_D4;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_D5;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_D6;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_DO5;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_DO6;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_D_CY;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_D_XOR;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_A;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_A1;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_A2;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_A3;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_A4;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_A5;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_A6;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_AO5;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_AO6;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_AQ;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_A_CY;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_A_XOR;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_B;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_B1;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_B2;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_B3;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_B4;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_B5;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_B6;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_BO5;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_BO6;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_BQ;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_B_CY;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_B_XOR;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_C;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_C1;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_C2;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_C3;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_C4;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_C5;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_C6;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_CLK;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_CO5;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_CO6;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_CQ;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_C_CY;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_C_XOR;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_D;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_D1;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_D2;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_D3;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_D4;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_D5;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_D6;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_DO5;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_DO6;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_DQ;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_D_CY;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_D_XOR;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_A;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_A1;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_A2;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_A3;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_A4;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_A5;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_A5Q;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_A6;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_AMUX;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_AO5;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_AO6;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_AQ;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_AX;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_A_CY;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_A_XOR;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_B;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_B1;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_B2;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_B3;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_B4;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_B5;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_B6;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_BO5;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_BO6;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_BQ;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_B_CY;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_B_XOR;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_C;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_C1;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_C2;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_C3;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_C4;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_C5;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_C6;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_CLK;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_CMUX;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_CO5;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_CO6;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_C_CY;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_C_XOR;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_D;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_D1;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_D2;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_D3;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_D4;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_D5;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_D6;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_DO5;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_DO6;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_DQ;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_D_CY;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_D_XOR;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_A;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_A1;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_A2;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_A3;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_A4;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_A5;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_A6;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_AO5;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_AO6;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_AQ;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_A_CY;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_A_XOR;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_B;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_B1;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_B2;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_B3;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_B4;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_B5;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_B6;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_BO5;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_BO6;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_BQ;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_B_CY;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_B_XOR;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_C;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_C1;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_C2;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_C3;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_C4;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_C5;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_C6;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_CLK;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_CO5;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_CO6;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_CQ;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_C_CY;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_C_XOR;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_D;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_D1;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_D2;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_D3;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_D4;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_D5;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_D6;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_DO5;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_DO6;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_D_CY;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_D_XOR;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_A;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_A1;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_A2;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_A3;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_A4;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_A5;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_A6;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_AO5;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_AO6;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_AQ;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_A_CY;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_A_XOR;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_B;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_B1;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_B2;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_B3;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_B4;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_B5;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_B6;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_BO5;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_BO6;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_BQ;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_B_CY;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_B_XOR;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_C;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_C1;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_C2;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_C3;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_C4;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_C5;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_C6;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_CLK;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_CO5;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_CO6;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_C_CY;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_C_XOR;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_D;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_D1;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_D2;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_D3;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_D4;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_D5;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_D6;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_DO5;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_DO6;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_D_CY;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_D_XOR;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_A;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_A1;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_A2;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_A3;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_A4;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_A5;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_A5Q;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_A6;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_AMUX;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_AO5;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_AO6;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_AQ;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_A_CY;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_A_XOR;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_B;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_B1;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_B2;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_B3;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_B4;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_B5;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_B6;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_BMUX;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_BO5;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_BO6;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_B_CY;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_B_XOR;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_C;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_C1;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_C2;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_C3;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_C4;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_C5;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_C6;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_CLK;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_CMUX;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_CO5;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_CO6;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_C_CY;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_C_XOR;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_D;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_D1;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_D2;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_D3;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_D4;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_D5;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_D6;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_DO5;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_DO6;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_D_CY;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_D_XOR;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_A;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_A1;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_A2;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_A3;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_A4;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_A5;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_A6;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_AO5;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_AO6;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_AQ;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_A_CY;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_A_XOR;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_B;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_B1;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_B2;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_B3;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_B4;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_B5;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_B6;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_BO5;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_BO6;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_B_CY;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_B_XOR;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_C;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_C1;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_C2;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_C3;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_C4;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_C5;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_C6;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_CLK;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_CO5;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_CO6;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_C_CY;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_C_XOR;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_D;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_D1;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_D2;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_D3;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_D4;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_D5;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_D6;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_DO5;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_DO6;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_D_CY;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_D_XOR;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X8Y157_A;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X8Y157_A1;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X8Y157_A2;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X8Y157_A3;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X8Y157_A4;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X8Y157_A5;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X8Y157_A6;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X8Y157_AO5;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X8Y157_AO6;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X8Y157_AQ;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X8Y157_AX;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X8Y157_A_CY;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X8Y157_A_XOR;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X8Y157_B;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X8Y157_B1;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X8Y157_B2;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X8Y157_B3;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X8Y157_B4;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X8Y157_B5;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X8Y157_B6;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X8Y157_BO5;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X8Y157_BO6;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X8Y157_B_CY;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X8Y157_B_XOR;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X8Y157_C;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X8Y157_C1;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X8Y157_C2;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X8Y157_C3;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X8Y157_C4;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X8Y157_C5;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X8Y157_C6;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X8Y157_CLK;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X8Y157_CO5;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X8Y157_CO6;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X8Y157_C_CY;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X8Y157_C_XOR;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X8Y157_D;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X8Y157_D1;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X8Y157_D2;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X8Y157_D3;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X8Y157_D4;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X8Y157_D5;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X8Y157_D6;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X8Y157_DO5;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X8Y157_DO6;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X8Y157_D_CY;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X8Y157_D_XOR;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X9Y157_A;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X9Y157_A1;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X9Y157_A2;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X9Y157_A3;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X9Y157_A4;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X9Y157_A5;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X9Y157_A6;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X9Y157_AO5;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X9Y157_AO6;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X9Y157_A_CY;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X9Y157_A_XOR;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X9Y157_B;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X9Y157_B1;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X9Y157_B2;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X9Y157_B3;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X9Y157_B4;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X9Y157_B5;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X9Y157_B6;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X9Y157_BO5;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X9Y157_BO6;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X9Y157_B_CY;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X9Y157_B_XOR;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X9Y157_C;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X9Y157_C1;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X9Y157_C2;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X9Y157_C3;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X9Y157_C4;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X9Y157_C5;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X9Y157_C6;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X9Y157_CO5;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X9Y157_CO6;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X9Y157_C_CY;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X9Y157_C_XOR;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X9Y157_D;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X9Y157_D1;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X9Y157_D2;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X9Y157_D3;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X9Y157_D4;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X9Y157_D5;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X9Y157_D6;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X9Y157_DO5;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X9Y157_DO6;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X9Y157_D_CY;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X9Y157_D_XOR;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE1;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I1;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE1;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S1;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_CE;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_I;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  wire [0:0] CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_CE;
  wire [0:0] CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_I;
  wire [0:0] CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  wire [0:0] LIOB33_SING_X0Y100_IOB_X0Y100_O;
  wire [0:0] LIOB33_SING_X0Y149_IOB_X0Y149_O;
  wire [0:0] LIOB33_SING_X0Y150_IOB_X0Y150_O;
  wire [0:0] LIOB33_SING_X0Y199_IOB_X0Y199_O;
  wire [0:0] LIOB33_SING_X0Y50_IOB_X0Y50_I;
  wire [0:0] LIOB33_X0Y101_IOB_X0Y101_O;
  wire [0:0] LIOB33_X0Y101_IOB_X0Y102_O;
  wire [0:0] LIOB33_X0Y103_IOB_X0Y103_O;
  wire [0:0] LIOB33_X0Y103_IOB_X0Y104_O;
  wire [0:0] LIOB33_X0Y105_IOB_X0Y105_O;
  wire [0:0] LIOB33_X0Y105_IOB_X0Y106_O;
  wire [0:0] LIOB33_X0Y107_IOB_X0Y107_O;
  wire [0:0] LIOB33_X0Y107_IOB_X0Y108_O;
  wire [0:0] LIOB33_X0Y109_IOB_X0Y109_O;
  wire [0:0] LIOB33_X0Y109_IOB_X0Y110_O;
  wire [0:0] LIOB33_X0Y111_IOB_X0Y111_O;
  wire [0:0] LIOB33_X0Y111_IOB_X0Y112_O;
  wire [0:0] LIOB33_X0Y113_IOB_X0Y113_O;
  wire [0:0] LIOB33_X0Y113_IOB_X0Y114_O;
  wire [0:0] LIOB33_X0Y115_IOB_X0Y115_O;
  wire [0:0] LIOB33_X0Y115_IOB_X0Y116_O;
  wire [0:0] LIOB33_X0Y117_IOB_X0Y117_O;
  wire [0:0] LIOB33_X0Y117_IOB_X0Y118_O;
  wire [0:0] LIOB33_X0Y119_IOB_X0Y119_O;
  wire [0:0] LIOB33_X0Y119_IOB_X0Y120_O;
  wire [0:0] LIOB33_X0Y121_IOB_X0Y121_O;
  wire [0:0] LIOB33_X0Y121_IOB_X0Y122_O;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y123_O;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y124_O;
  wire [0:0] LIOB33_X0Y125_IOB_X0Y125_O;
  wire [0:0] LIOB33_X0Y125_IOB_X0Y126_O;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y127_O;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y128_O;
  wire [0:0] LIOB33_X0Y129_IOB_X0Y129_O;
  wire [0:0] LIOB33_X0Y129_IOB_X0Y130_O;
  wire [0:0] LIOB33_X0Y131_IOB_X0Y131_O;
  wire [0:0] LIOB33_X0Y131_IOB_X0Y132_O;
  wire [0:0] LIOB33_X0Y133_IOB_X0Y133_O;
  wire [0:0] LIOB33_X0Y133_IOB_X0Y134_O;
  wire [0:0] LIOB33_X0Y135_IOB_X0Y135_O;
  wire [0:0] LIOB33_X0Y135_IOB_X0Y136_O;
  wire [0:0] LIOB33_X0Y137_IOB_X0Y137_O;
  wire [0:0] LIOB33_X0Y137_IOB_X0Y138_O;
  wire [0:0] LIOB33_X0Y139_IOB_X0Y139_O;
  wire [0:0] LIOB33_X0Y139_IOB_X0Y140_O;
  wire [0:0] LIOB33_X0Y141_IOB_X0Y141_O;
  wire [0:0] LIOB33_X0Y141_IOB_X0Y142_O;
  wire [0:0] LIOB33_X0Y143_IOB_X0Y143_O;
  wire [0:0] LIOB33_X0Y145_IOB_X0Y145_O;
  wire [0:0] LIOB33_X0Y145_IOB_X0Y146_O;
  wire [0:0] LIOB33_X0Y147_IOB_X0Y147_O;
  wire [0:0] LIOB33_X0Y147_IOB_X0Y148_O;
  wire [0:0] LIOB33_X0Y151_IOB_X0Y151_O;
  wire [0:0] LIOB33_X0Y151_IOB_X0Y152_O;
  wire [0:0] LIOB33_X0Y153_IOB_X0Y153_O;
  wire [0:0] LIOB33_X0Y153_IOB_X0Y154_O;
  wire [0:0] LIOB33_X0Y155_IOB_X0Y155_O;
  wire [0:0] LIOB33_X0Y155_IOB_X0Y156_O;
  wire [0:0] LIOB33_X0Y157_IOB_X0Y157_O;
  wire [0:0] LIOB33_X0Y157_IOB_X0Y158_O;
  wire [0:0] LIOB33_X0Y159_IOB_X0Y159_O;
  wire [0:0] LIOB33_X0Y159_IOB_X0Y160_O;
  wire [0:0] LIOB33_X0Y161_IOB_X0Y161_O;
  wire [0:0] LIOB33_X0Y161_IOB_X0Y162_O;
  wire [0:0] LIOB33_X0Y163_IOB_X0Y163_O;
  wire [0:0] LIOB33_X0Y163_IOB_X0Y164_O;
  wire [0:0] LIOB33_X0Y165_IOB_X0Y165_O;
  wire [0:0] LIOB33_X0Y165_IOB_X0Y166_O;
  wire [0:0] LIOB33_X0Y167_IOB_X0Y167_O;
  wire [0:0] LIOB33_X0Y167_IOB_X0Y168_O;
  wire [0:0] LIOB33_X0Y169_IOB_X0Y169_O;
  wire [0:0] LIOB33_X0Y169_IOB_X0Y170_O;
  wire [0:0] LIOB33_X0Y171_IOB_X0Y171_O;
  wire [0:0] LIOB33_X0Y171_IOB_X0Y172_O;
  wire [0:0] LIOB33_X0Y173_IOB_X0Y173_O;
  wire [0:0] LIOB33_X0Y173_IOB_X0Y174_O;
  wire [0:0] LIOB33_X0Y175_IOB_X0Y175_O;
  wire [0:0] LIOB33_X0Y175_IOB_X0Y176_O;
  wire [0:0] LIOB33_X0Y177_IOB_X0Y177_O;
  wire [0:0] LIOB33_X0Y177_IOB_X0Y178_O;
  wire [0:0] LIOB33_X0Y179_IOB_X0Y179_O;
  wire [0:0] LIOB33_X0Y179_IOB_X0Y180_O;
  wire [0:0] LIOB33_X0Y181_IOB_X0Y181_O;
  wire [0:0] LIOB33_X0Y181_IOB_X0Y182_O;
  wire [0:0] LIOB33_X0Y183_IOB_X0Y183_O;
  wire [0:0] LIOB33_X0Y183_IOB_X0Y184_O;
  wire [0:0] LIOB33_X0Y185_IOB_X0Y185_O;
  wire [0:0] LIOB33_X0Y185_IOB_X0Y186_O;
  wire [0:0] LIOB33_X0Y187_IOB_X0Y187_O;
  wire [0:0] LIOB33_X0Y187_IOB_X0Y188_O;
  wire [0:0] LIOB33_X0Y189_IOB_X0Y189_O;
  wire [0:0] LIOB33_X0Y189_IOB_X0Y190_O;
  wire [0:0] LIOB33_X0Y191_IOB_X0Y191_O;
  wire [0:0] LIOB33_X0Y191_IOB_X0Y192_O;
  wire [0:0] LIOB33_X0Y193_IOB_X0Y193_O;
  wire [0:0] LIOB33_X0Y193_IOB_X0Y194_O;
  wire [0:0] LIOB33_X0Y195_IOB_X0Y195_O;
  wire [0:0] LIOB33_X0Y195_IOB_X0Y196_O;
  wire [0:0] LIOB33_X0Y197_IOB_X0Y197_O;
  wire [0:0] LIOB33_X0Y197_IOB_X0Y198_O;
  wire [0:0] LIOB33_X0Y51_IOB_X0Y51_I;
  wire [0:0] LIOB33_X0Y51_IOB_X0Y52_I;
  wire [0:0] LIOB33_X0Y53_IOB_X0Y53_I;
  wire [0:0] LIOB33_X0Y53_IOB_X0Y54_I;
  wire [0:0] LIOB33_X0Y55_IOB_X0Y55_I;
  wire [0:0] LIOB33_X0Y55_IOB_X0Y56_I;
  wire [0:0] LIOB33_X0Y57_IOB_X0Y57_I;
  wire [0:0] LIOB33_X0Y57_IOB_X0Y58_I;
  wire [0:0] LIOB33_X0Y59_IOB_X0Y59_I;
  wire [0:0] LIOB33_X0Y59_IOB_X0Y60_I;
  wire [0:0] LIOB33_X0Y61_IOB_X0Y61_I;
  wire [0:0] LIOB33_X0Y61_IOB_X0Y62_I;
  wire [0:0] LIOB33_X0Y63_IOB_X0Y63_I;
  wire [0:0] LIOB33_X0Y63_IOB_X0Y64_I;
  wire [0:0] LIOB33_X0Y65_IOB_X0Y65_I;
  wire [0:0] LIOB33_X0Y65_IOB_X0Y66_I;
  wire [0:0] LIOB33_X0Y67_IOB_X0Y67_I;
  wire [0:0] LIOB33_X0Y67_IOB_X0Y68_I;
  wire [0:0] LIOB33_X0Y69_IOB_X0Y69_I;
  wire [0:0] LIOB33_X0Y69_IOB_X0Y70_I;
  wire [0:0] LIOB33_X0Y71_IOB_X0Y71_I;
  wire [0:0] LIOB33_X0Y71_IOB_X0Y72_I;
  wire [0:0] LIOB33_X0Y73_IOB_X0Y73_I;
  wire [0:0] LIOB33_X0Y73_IOB_X0Y74_I;
  wire [0:0] LIOB33_X0Y75_IOB_X0Y75_I;
  wire [0:0] LIOB33_X0Y75_IOB_X0Y76_I;
  wire [0:0] LIOB33_X0Y77_IOB_X0Y77_I;
  wire [0:0] LIOB33_X0Y77_IOB_X0Y78_I;
  wire [0:0] LIOB33_X0Y79_IOB_X0Y79_I;
  wire [0:0] LIOB33_X0Y79_IOB_X0Y80_O;
  wire [0:0] LIOI3_SING_X0Y100_OLOGIC_X0Y100_D1;
  wire [0:0] LIOI3_SING_X0Y100_OLOGIC_X0Y100_OQ;
  wire [0:0] LIOI3_SING_X0Y100_OLOGIC_X0Y100_T1;
  wire [0:0] LIOI3_SING_X0Y100_OLOGIC_X0Y100_TQ;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_D1;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_OQ;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_T1;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_TQ;
  wire [0:0] LIOI3_SING_X0Y150_OLOGIC_X0Y150_D1;
  wire [0:0] LIOI3_SING_X0Y150_OLOGIC_X0Y150_OQ;
  wire [0:0] LIOI3_SING_X0Y150_OLOGIC_X0Y150_T1;
  wire [0:0] LIOI3_SING_X0Y150_OLOGIC_X0Y150_TQ;
  wire [0:0] LIOI3_SING_X0Y199_OLOGIC_X0Y199_D1;
  wire [0:0] LIOI3_SING_X0Y199_OLOGIC_X0Y199_OQ;
  wire [0:0] LIOI3_SING_X0Y199_OLOGIC_X0Y199_T1;
  wire [0:0] LIOI3_SING_X0Y199_OLOGIC_X0Y199_TQ;
  wire [0:0] LIOI3_SING_X0Y50_ILOGIC_X0Y50_D;
  wire [0:0] LIOI3_SING_X0Y50_ILOGIC_X0Y50_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y57_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y57_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y58_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y58_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y69_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y69_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y70_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y70_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y63_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y63_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y64_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y64_O;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y101_D1;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y101_OQ;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y101_T1;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y101_TQ;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y102_D1;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y102_OQ;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y102_T1;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y102_TQ;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y103_D1;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y103_OQ;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y103_T1;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y103_TQ;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y104_D1;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y104_OQ;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y104_T1;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y104_TQ;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y105_D1;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y105_OQ;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y105_T1;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y105_TQ;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y106_D1;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y106_OQ;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y106_T1;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y106_TQ;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y109_D1;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y109_OQ;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y109_T1;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y109_TQ;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y110_D1;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y110_OQ;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y110_T1;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y110_TQ;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_D1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_OQ;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_T1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_TQ;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y112_D1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y112_OQ;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y112_T1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y112_TQ;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y115_D1;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y115_OQ;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y115_T1;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y115_TQ;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y116_D1;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y116_OQ;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y116_T1;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y116_TQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y117_D1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y117_OQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y117_T1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y117_TQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_D1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_OQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_T1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_TQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_D1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_OQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_T1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_TQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_D1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_OQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_T1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_TQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_D1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_OQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_T1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_TQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_D1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_OQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_T1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_TQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_D1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_OQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_T1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_TQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_D1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_OQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_T1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_TQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_D1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_OQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_T1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_TQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_D1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_OQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_T1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_TQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_D1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_OQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_T1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_TQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_D1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_OQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_T1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_TQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_D1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_OQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_T1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_TQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_D1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_OQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_T1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_TQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_D1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_OQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_T1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_TQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_D1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_OQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_T1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_TQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_D1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_OQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_T1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_TQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_D1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_OQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_T1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_TQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_D1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_OQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_T1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_TQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_D1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_OQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_T1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_TQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_D1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_OQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_T1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_TQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_D1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_OQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_T1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_TQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_D1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_OQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_T1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_TQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_D1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_OQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_T1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_TQ;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y151_D1;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y151_OQ;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y151_T1;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y151_TQ;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y152_D1;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y152_OQ;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y152_T1;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y152_TQ;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y153_D1;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y153_OQ;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y153_T1;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y153_TQ;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y154_D1;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y154_OQ;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y154_T1;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y154_TQ;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y155_D1;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y155_OQ;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y155_T1;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y155_TQ;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y156_D1;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y156_OQ;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y156_T1;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y156_TQ;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y159_D1;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y159_OQ;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y159_T1;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y159_TQ;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y160_D1;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y160_OQ;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y160_T1;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y160_TQ;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y161_D1;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y161_OQ;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y161_T1;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y161_TQ;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y162_D1;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y162_OQ;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y162_T1;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y162_TQ;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y165_D1;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y165_OQ;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y165_T1;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y165_TQ;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y166_D1;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y166_OQ;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y166_T1;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y166_TQ;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y167_D1;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y167_OQ;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y167_T1;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y167_TQ;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y168_D1;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y168_OQ;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y168_T1;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y168_TQ;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y171_D1;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y171_OQ;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y171_T1;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y171_TQ;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y172_D1;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y172_OQ;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y172_T1;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y172_TQ;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y173_D1;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y173_OQ;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y173_T1;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y173_TQ;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y174_D1;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y174_OQ;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y174_T1;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y174_TQ;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y175_D1;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y175_OQ;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y175_T1;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y175_TQ;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y176_D1;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y176_OQ;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y176_T1;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y176_TQ;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y177_D1;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y177_OQ;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y177_T1;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y177_TQ;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y178_D1;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y178_OQ;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y178_T1;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y178_TQ;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y179_D1;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y179_OQ;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y179_T1;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y179_TQ;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y180_D1;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y180_OQ;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y180_T1;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y180_TQ;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y183_D1;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y183_OQ;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y183_T1;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y183_TQ;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y184_D1;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y184_OQ;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y184_T1;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y184_TQ;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y185_D1;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y185_OQ;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y185_T1;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y185_TQ;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y186_D1;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y186_OQ;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y186_T1;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y186_TQ;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y189_D1;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y189_OQ;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y189_T1;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y189_TQ;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y190_D1;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y190_OQ;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y190_T1;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y190_TQ;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y191_D1;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y191_OQ;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y191_T1;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y191_TQ;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y192_D1;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y192_OQ;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y192_T1;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y192_TQ;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y195_D1;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y195_OQ;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y195_T1;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y195_TQ;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y196_D1;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y196_OQ;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y196_T1;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y196_TQ;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y197_D1;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y197_OQ;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y197_T1;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y197_TQ;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y198_D1;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y198_OQ;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y198_T1;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y198_TQ;
  wire [0:0] LIOI3_X0Y51_ILOGIC_X0Y51_D;
  wire [0:0] LIOI3_X0Y51_ILOGIC_X0Y51_O;
  wire [0:0] LIOI3_X0Y51_ILOGIC_X0Y52_D;
  wire [0:0] LIOI3_X0Y51_ILOGIC_X0Y52_O;
  wire [0:0] LIOI3_X0Y53_ILOGIC_X0Y53_D;
  wire [0:0] LIOI3_X0Y53_ILOGIC_X0Y53_O;
  wire [0:0] LIOI3_X0Y53_ILOGIC_X0Y54_D;
  wire [0:0] LIOI3_X0Y53_ILOGIC_X0Y54_O;
  wire [0:0] LIOI3_X0Y55_ILOGIC_X0Y55_D;
  wire [0:0] LIOI3_X0Y55_ILOGIC_X0Y55_O;
  wire [0:0] LIOI3_X0Y55_ILOGIC_X0Y56_D;
  wire [0:0] LIOI3_X0Y55_ILOGIC_X0Y56_O;
  wire [0:0] LIOI3_X0Y59_ILOGIC_X0Y59_D;
  wire [0:0] LIOI3_X0Y59_ILOGIC_X0Y59_O;
  wire [0:0] LIOI3_X0Y59_ILOGIC_X0Y60_D;
  wire [0:0] LIOI3_X0Y59_ILOGIC_X0Y60_O;
  wire [0:0] LIOI3_X0Y61_ILOGIC_X0Y61_D;
  wire [0:0] LIOI3_X0Y61_ILOGIC_X0Y61_O;
  wire [0:0] LIOI3_X0Y61_ILOGIC_X0Y62_D;
  wire [0:0] LIOI3_X0Y61_ILOGIC_X0Y62_O;
  wire [0:0] LIOI3_X0Y65_ILOGIC_X0Y65_D;
  wire [0:0] LIOI3_X0Y65_ILOGIC_X0Y65_O;
  wire [0:0] LIOI3_X0Y65_ILOGIC_X0Y66_D;
  wire [0:0] LIOI3_X0Y65_ILOGIC_X0Y66_O;
  wire [0:0] LIOI3_X0Y67_ILOGIC_X0Y67_D;
  wire [0:0] LIOI3_X0Y67_ILOGIC_X0Y67_O;
  wire [0:0] LIOI3_X0Y67_ILOGIC_X0Y68_D;
  wire [0:0] LIOI3_X0Y67_ILOGIC_X0Y68_O;
  wire [0:0] LIOI3_X0Y71_ILOGIC_X0Y71_D;
  wire [0:0] LIOI3_X0Y71_ILOGIC_X0Y71_O;
  wire [0:0] LIOI3_X0Y71_ILOGIC_X0Y72_D;
  wire [0:0] LIOI3_X0Y71_ILOGIC_X0Y72_O;
  wire [0:0] LIOI3_X0Y73_ILOGIC_X0Y73_D;
  wire [0:0] LIOI3_X0Y73_ILOGIC_X0Y73_O;
  wire [0:0] LIOI3_X0Y73_ILOGIC_X0Y74_D;
  wire [0:0] LIOI3_X0Y73_ILOGIC_X0Y74_O;
  wire [0:0] LIOI3_X0Y75_ILOGIC_X0Y75_D;
  wire [0:0] LIOI3_X0Y75_ILOGIC_X0Y75_O;
  wire [0:0] LIOI3_X0Y75_ILOGIC_X0Y76_D;
  wire [0:0] LIOI3_X0Y75_ILOGIC_X0Y76_O;
  wire [0:0] LIOI3_X0Y77_ILOGIC_X0Y77_D;
  wire [0:0] LIOI3_X0Y77_ILOGIC_X0Y77_O;
  wire [0:0] LIOI3_X0Y77_ILOGIC_X0Y78_D;
  wire [0:0] LIOI3_X0Y77_ILOGIC_X0Y78_O;
  wire [0:0] LIOI3_X0Y79_ILOGIC_X0Y79_D;
  wire [0:0] LIOI3_X0Y79_ILOGIC_X0Y79_O;
  wire [0:0] LIOI3_X0Y79_OLOGIC_X0Y80_D1;
  wire [0:0] LIOI3_X0Y79_OLOGIC_X0Y80_OQ;
  wire [0:0] LIOI3_X0Y79_OLOGIC_X0Y80_T1;
  wire [0:0] LIOI3_X0Y79_OLOGIC_X0Y80_TQ;
  wire [0:0] RIOB33_SING_X105Y100_IOB_X1Y100_I;
  wire [0:0] RIOB33_SING_X105Y149_IOB_X1Y149_I;
  wire [0:0] RIOB33_SING_X105Y150_IOB_X1Y150_O;
  wire [0:0] RIOB33_SING_X105Y199_IOB_X1Y199_O;
  wire [0:0] RIOB33_X105Y101_IOB_X1Y101_I;
  wire [0:0] RIOB33_X105Y101_IOB_X1Y102_I;
  wire [0:0] RIOB33_X105Y103_IOB_X1Y103_I;
  wire [0:0] RIOB33_X105Y103_IOB_X1Y104_I;
  wire [0:0] RIOB33_X105Y105_IOB_X1Y105_I;
  wire [0:0] RIOB33_X105Y105_IOB_X1Y106_I;
  wire [0:0] RIOB33_X105Y107_IOB_X1Y107_I;
  wire [0:0] RIOB33_X105Y107_IOB_X1Y108_I;
  wire [0:0] RIOB33_X105Y109_IOB_X1Y109_I;
  wire [0:0] RIOB33_X105Y109_IOB_X1Y110_I;
  wire [0:0] RIOB33_X105Y111_IOB_X1Y111_I;
  wire [0:0] RIOB33_X105Y111_IOB_X1Y112_I;
  wire [0:0] RIOB33_X105Y113_IOB_X1Y113_I;
  wire [0:0] RIOB33_X105Y113_IOB_X1Y114_I;
  wire [0:0] RIOB33_X105Y115_IOB_X1Y115_I;
  wire [0:0] RIOB33_X105Y115_IOB_X1Y116_I;
  wire [0:0] RIOB33_X105Y117_IOB_X1Y117_I;
  wire [0:0] RIOB33_X105Y117_IOB_X1Y118_I;
  wire [0:0] RIOB33_X105Y119_IOB_X1Y119_I;
  wire [0:0] RIOB33_X105Y119_IOB_X1Y120_I;
  wire [0:0] RIOB33_X105Y121_IOB_X1Y121_I;
  wire [0:0] RIOB33_X105Y121_IOB_X1Y122_I;
  wire [0:0] RIOB33_X105Y123_IOB_X1Y123_I;
  wire [0:0] RIOB33_X105Y123_IOB_X1Y124_I;
  wire [0:0] RIOB33_X105Y125_IOB_X1Y125_I;
  wire [0:0] RIOB33_X105Y125_IOB_X1Y126_I;
  wire [0:0] RIOB33_X105Y127_IOB_X1Y127_I;
  wire [0:0] RIOB33_X105Y127_IOB_X1Y128_I;
  wire [0:0] RIOB33_X105Y129_IOB_X1Y129_I;
  wire [0:0] RIOB33_X105Y129_IOB_X1Y130_I;
  wire [0:0] RIOB33_X105Y131_IOB_X1Y131_I;
  wire [0:0] RIOB33_X105Y131_IOB_X1Y132_I;
  wire [0:0] RIOB33_X105Y133_IOB_X1Y133_I;
  wire [0:0] RIOB33_X105Y133_IOB_X1Y134_I;
  wire [0:0] RIOB33_X105Y135_IOB_X1Y135_I;
  wire [0:0] RIOB33_X105Y135_IOB_X1Y136_I;
  wire [0:0] RIOB33_X105Y137_IOB_X1Y137_I;
  wire [0:0] RIOB33_X105Y137_IOB_X1Y138_I;
  wire [0:0] RIOB33_X105Y139_IOB_X1Y139_I;
  wire [0:0] RIOB33_X105Y139_IOB_X1Y140_I;
  wire [0:0] RIOB33_X105Y141_IOB_X1Y141_I;
  wire [0:0] RIOB33_X105Y141_IOB_X1Y142_I;
  wire [0:0] RIOB33_X105Y143_IOB_X1Y143_I;
  wire [0:0] RIOB33_X105Y143_IOB_X1Y144_I;
  wire [0:0] RIOB33_X105Y145_IOB_X1Y145_I;
  wire [0:0] RIOB33_X105Y145_IOB_X1Y146_I;
  wire [0:0] RIOB33_X105Y147_IOB_X1Y147_I;
  wire [0:0] RIOB33_X105Y147_IOB_X1Y148_I;
  wire [0:0] RIOB33_X105Y151_IOB_X1Y151_O;
  wire [0:0] RIOB33_X105Y151_IOB_X1Y152_O;
  wire [0:0] RIOB33_X105Y153_IOB_X1Y153_O;
  wire [0:0] RIOB33_X105Y153_IOB_X1Y154_O;
  wire [0:0] RIOB33_X105Y155_IOB_X1Y155_O;
  wire [0:0] RIOB33_X105Y155_IOB_X1Y156_O;
  wire [0:0] RIOB33_X105Y157_IOB_X1Y157_O;
  wire [0:0] RIOB33_X105Y157_IOB_X1Y158_O;
  wire [0:0] RIOB33_X105Y159_IOB_X1Y159_O;
  wire [0:0] RIOB33_X105Y159_IOB_X1Y160_O;
  wire [0:0] RIOB33_X105Y161_IOB_X1Y161_O;
  wire [0:0] RIOB33_X105Y161_IOB_X1Y162_O;
  wire [0:0] RIOB33_X105Y163_IOB_X1Y163_O;
  wire [0:0] RIOB33_X105Y163_IOB_X1Y164_O;
  wire [0:0] RIOB33_X105Y165_IOB_X1Y165_O;
  wire [0:0] RIOB33_X105Y165_IOB_X1Y166_O;
  wire [0:0] RIOB33_X105Y167_IOB_X1Y167_O;
  wire [0:0] RIOB33_X105Y167_IOB_X1Y168_O;
  wire [0:0] RIOB33_X105Y169_IOB_X1Y169_O;
  wire [0:0] RIOB33_X105Y169_IOB_X1Y170_O;
  wire [0:0] RIOB33_X105Y171_IOB_X1Y171_O;
  wire [0:0] RIOB33_X105Y171_IOB_X1Y172_O;
  wire [0:0] RIOB33_X105Y173_IOB_X1Y173_O;
  wire [0:0] RIOB33_X105Y173_IOB_X1Y174_O;
  wire [0:0] RIOB33_X105Y175_IOB_X1Y175_O;
  wire [0:0] RIOB33_X105Y175_IOB_X1Y176_O;
  wire [0:0] RIOB33_X105Y177_IOB_X1Y177_O;
  wire [0:0] RIOB33_X105Y177_IOB_X1Y178_O;
  wire [0:0] RIOB33_X105Y179_IOB_X1Y179_O;
  wire [0:0] RIOB33_X105Y179_IOB_X1Y180_O;
  wire [0:0] RIOB33_X105Y181_IOB_X1Y181_O;
  wire [0:0] RIOB33_X105Y181_IOB_X1Y182_O;
  wire [0:0] RIOB33_X105Y183_IOB_X1Y183_O;
  wire [0:0] RIOB33_X105Y183_IOB_X1Y184_O;
  wire [0:0] RIOB33_X105Y185_IOB_X1Y185_O;
  wire [0:0] RIOB33_X105Y185_IOB_X1Y186_O;
  wire [0:0] RIOB33_X105Y187_IOB_X1Y187_O;
  wire [0:0] RIOB33_X105Y187_IOB_X1Y188_O;
  wire [0:0] RIOB33_X105Y189_IOB_X1Y189_O;
  wire [0:0] RIOB33_X105Y189_IOB_X1Y190_O;
  wire [0:0] RIOB33_X105Y191_IOB_X1Y191_O;
  wire [0:0] RIOB33_X105Y191_IOB_X1Y192_O;
  wire [0:0] RIOB33_X105Y193_IOB_X1Y193_O;
  wire [0:0] RIOB33_X105Y193_IOB_X1Y194_O;
  wire [0:0] RIOB33_X105Y195_IOB_X1Y195_O;
  wire [0:0] RIOB33_X105Y195_IOB_X1Y196_O;
  wire [0:0] RIOB33_X105Y197_IOB_X1Y197_O;
  wire [0:0] RIOB33_X105Y197_IOB_X1Y198_O;
  wire [0:0] RIOI3_SING_X105Y100_ILOGIC_X1Y100_D;
  wire [0:0] RIOI3_SING_X105Y100_ILOGIC_X1Y100_O;
  wire [0:0] RIOI3_SING_X105Y149_ILOGIC_X1Y149_D;
  wire [0:0] RIOI3_SING_X105Y149_ILOGIC_X1Y149_O;
  wire [0:0] RIOI3_SING_X105Y150_OLOGIC_X1Y150_D1;
  wire [0:0] RIOI3_SING_X105Y150_OLOGIC_X1Y150_OQ;
  wire [0:0] RIOI3_SING_X105Y150_OLOGIC_X1Y150_T1;
  wire [0:0] RIOI3_SING_X105Y150_OLOGIC_X1Y150_TQ;
  wire [0:0] RIOI3_SING_X105Y199_OLOGIC_X1Y199_D1;
  wire [0:0] RIOI3_SING_X105Y199_OLOGIC_X1Y199_OQ;
  wire [0:0] RIOI3_SING_X105Y199_OLOGIC_X1Y199_T1;
  wire [0:0] RIOI3_SING_X105Y199_OLOGIC_X1Y199_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y131_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y131_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y132_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y132_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y143_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y143_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y144_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y144_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y114_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y114_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y137_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y137_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y138_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y138_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_TQ;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y101_D;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y101_O;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y102_D;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y102_O;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y103_D;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y103_O;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y104_D;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y104_O;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y105_D;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y105_O;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y106_D;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y106_O;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y109_D;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y109_O;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y110_D;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y110_O;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y111_D;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y111_O;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y112_D;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y112_O;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y115_D;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y115_O;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y116_D;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y116_O;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y117_D;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y117_O;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y118_D;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y118_O;
  wire [0:0] RIOI3_X105Y121_ILOGIC_X1Y121_D;
  wire [0:0] RIOI3_X105Y121_ILOGIC_X1Y121_O;
  wire [0:0] RIOI3_X105Y121_ILOGIC_X1Y122_D;
  wire [0:0] RIOI3_X105Y121_ILOGIC_X1Y122_O;
  wire [0:0] RIOI3_X105Y123_ILOGIC_X1Y123_D;
  wire [0:0] RIOI3_X105Y123_ILOGIC_X1Y123_O;
  wire [0:0] RIOI3_X105Y123_ILOGIC_X1Y124_D;
  wire [0:0] RIOI3_X105Y123_ILOGIC_X1Y124_O;
  wire [0:0] RIOI3_X105Y125_ILOGIC_X1Y125_D;
  wire [0:0] RIOI3_X105Y125_ILOGIC_X1Y125_O;
  wire [0:0] RIOI3_X105Y125_ILOGIC_X1Y126_D;
  wire [0:0] RIOI3_X105Y125_ILOGIC_X1Y126_O;
  wire [0:0] RIOI3_X105Y127_ILOGIC_X1Y127_D;
  wire [0:0] RIOI3_X105Y127_ILOGIC_X1Y127_O;
  wire [0:0] RIOI3_X105Y127_ILOGIC_X1Y128_D;
  wire [0:0] RIOI3_X105Y127_ILOGIC_X1Y128_O;
  wire [0:0] RIOI3_X105Y129_ILOGIC_X1Y129_D;
  wire [0:0] RIOI3_X105Y129_ILOGIC_X1Y129_O;
  wire [0:0] RIOI3_X105Y129_ILOGIC_X1Y130_D;
  wire [0:0] RIOI3_X105Y129_ILOGIC_X1Y130_O;
  wire [0:0] RIOI3_X105Y133_ILOGIC_X1Y133_D;
  wire [0:0] RIOI3_X105Y133_ILOGIC_X1Y133_O;
  wire [0:0] RIOI3_X105Y133_ILOGIC_X1Y134_D;
  wire [0:0] RIOI3_X105Y133_ILOGIC_X1Y134_O;
  wire [0:0] RIOI3_X105Y135_ILOGIC_X1Y135_D;
  wire [0:0] RIOI3_X105Y135_ILOGIC_X1Y135_O;
  wire [0:0] RIOI3_X105Y135_ILOGIC_X1Y136_D;
  wire [0:0] RIOI3_X105Y135_ILOGIC_X1Y136_O;
  wire [0:0] RIOI3_X105Y139_ILOGIC_X1Y139_D;
  wire [0:0] RIOI3_X105Y139_ILOGIC_X1Y139_O;
  wire [0:0] RIOI3_X105Y139_ILOGIC_X1Y140_D;
  wire [0:0] RIOI3_X105Y139_ILOGIC_X1Y140_O;
  wire [0:0] RIOI3_X105Y141_ILOGIC_X1Y141_D;
  wire [0:0] RIOI3_X105Y141_ILOGIC_X1Y141_O;
  wire [0:0] RIOI3_X105Y141_ILOGIC_X1Y142_D;
  wire [0:0] RIOI3_X105Y141_ILOGIC_X1Y142_O;
  wire [0:0] RIOI3_X105Y145_ILOGIC_X1Y145_D;
  wire [0:0] RIOI3_X105Y145_ILOGIC_X1Y145_O;
  wire [0:0] RIOI3_X105Y145_ILOGIC_X1Y146_D;
  wire [0:0] RIOI3_X105Y145_ILOGIC_X1Y146_O;
  wire [0:0] RIOI3_X105Y147_ILOGIC_X1Y147_D;
  wire [0:0] RIOI3_X105Y147_ILOGIC_X1Y147_O;
  wire [0:0] RIOI3_X105Y147_ILOGIC_X1Y148_D;
  wire [0:0] RIOI3_X105Y147_ILOGIC_X1Y148_O;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y151_D1;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y151_OQ;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y151_T1;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y151_TQ;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y152_D1;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y152_OQ;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y152_T1;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y152_TQ;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y153_D1;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y153_OQ;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y153_T1;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y153_TQ;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y154_D1;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y154_OQ;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y154_T1;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y154_TQ;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y155_D1;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y155_OQ;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y155_T1;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y155_TQ;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y156_D1;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y156_OQ;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y156_T1;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y156_TQ;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y159_D1;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y159_OQ;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y159_T1;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y159_TQ;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y160_D1;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y160_OQ;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y160_T1;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y160_TQ;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y161_D1;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y161_OQ;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y161_T1;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y161_TQ;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y162_D1;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y162_OQ;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y162_T1;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y162_TQ;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y165_D1;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y165_OQ;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y165_T1;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y165_TQ;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y166_D1;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y166_OQ;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y166_T1;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y166_TQ;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y167_D1;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y167_OQ;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y167_T1;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y167_TQ;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y168_D1;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y168_OQ;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y168_T1;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y168_TQ;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y171_D1;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y171_OQ;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y171_T1;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y171_TQ;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y172_D1;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y172_OQ;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y172_T1;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y172_TQ;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y173_D1;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y173_OQ;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y173_T1;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y173_TQ;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y174_D1;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y174_OQ;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y174_T1;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y174_TQ;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y175_D1;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y175_OQ;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y175_T1;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y175_TQ;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y176_D1;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y176_OQ;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y176_T1;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y176_TQ;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y177_D1;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y177_OQ;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y177_T1;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y177_TQ;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y178_D1;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y178_OQ;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y178_T1;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y178_TQ;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y179_D1;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y179_OQ;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y179_T1;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y179_TQ;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y180_D1;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y180_OQ;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y180_T1;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y180_TQ;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y183_D1;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y183_OQ;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y183_T1;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y183_TQ;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y184_D1;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y184_OQ;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y184_T1;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y184_TQ;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y185_D1;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y185_OQ;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y185_T1;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y185_TQ;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y186_D1;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y186_OQ;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y186_T1;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y186_TQ;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y189_D1;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y189_OQ;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y189_T1;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y189_TQ;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y190_D1;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y190_OQ;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y190_T1;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y190_TQ;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y191_D1;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y191_OQ;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y191_T1;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y191_TQ;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y192_D1;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y192_OQ;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y192_T1;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y192_TQ;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y195_D1;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y195_OQ;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y195_T1;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y195_TQ;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y196_D1;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y196_OQ;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y196_T1;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y196_TQ;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y197_D1;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y197_OQ;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y197_T1;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y197_TQ;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y198_D1;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y198_OQ;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y198_T1;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y198_TQ;


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y120_SLICE_X0Y120_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y120_SLICE_X0Y120_DO5),
.O6(CLBLL_L_X2Y120_SLICE_X0Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y120_SLICE_X0Y120_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y120_SLICE_X0Y120_CO5),
.O6(CLBLL_L_X2Y120_SLICE_X0Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y120_SLICE_X0Y120_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y120_SLICE_X0Y120_BO5),
.O6(CLBLL_L_X2Y120_SLICE_X0Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00ff00ff00ff)
  ) CLBLL_L_X2Y120_SLICE_X0Y120_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLL_L_X2Y141_SLICE_X0Y141_BO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y120_SLICE_X0Y120_AO5),
.O6(CLBLL_L_X2Y120_SLICE_X0Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y120_SLICE_X1Y120_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y120_SLICE_X1Y120_DO5),
.O6(CLBLL_L_X2Y120_SLICE_X1Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y120_SLICE_X1Y120_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y120_SLICE_X1Y120_CO5),
.O6(CLBLL_L_X2Y120_SLICE_X1Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y120_SLICE_X1Y120_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y120_SLICE_X1Y120_BO5),
.O6(CLBLL_L_X2Y120_SLICE_X1Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y120_SLICE_X1Y120_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y120_SLICE_X1Y120_AO5),
.O6(CLBLL_L_X2Y120_SLICE_X1Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y134_SLICE_X0Y134_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y134_SLICE_X0Y134_DO5),
.O6(CLBLL_L_X2Y134_SLICE_X0Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y134_SLICE_X0Y134_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y134_SLICE_X0Y134_CO5),
.O6(CLBLL_L_X2Y134_SLICE_X0Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y134_SLICE_X0Y134_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y134_SLICE_X0Y134_BO5),
.O6(CLBLL_L_X2Y134_SLICE_X0Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0ff00ff030303030)
  ) CLBLL_L_X2Y134_SLICE_X0Y134_ALUT (
.I0(1'b1),
.I1(CLBLL_L_X2Y141_SLICE_X0Y141_BO6),
.I2(CLBLL_L_X2Y147_SLICE_X0Y147_AO6),
.I3(CLBLM_R_X5Y145_SLICE_X6Y145_DO5),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y134_SLICE_X0Y134_AO5),
.O6(CLBLL_L_X2Y134_SLICE_X0Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y134_SLICE_X1Y134_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y134_SLICE_X1Y134_DO5),
.O6(CLBLL_L_X2Y134_SLICE_X1Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y134_SLICE_X1Y134_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y134_SLICE_X1Y134_CO5),
.O6(CLBLL_L_X2Y134_SLICE_X1Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y134_SLICE_X1Y134_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y134_SLICE_X1Y134_BO5),
.O6(CLBLL_L_X2Y134_SLICE_X1Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y134_SLICE_X1Y134_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y134_SLICE_X1Y134_AO5),
.O6(CLBLL_L_X2Y134_SLICE_X1Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y138_SLICE_X0Y138_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y138_SLICE_X0Y138_DO5),
.O6(CLBLL_L_X2Y138_SLICE_X0Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffbfffbfffffbfb)
  ) CLBLL_L_X2Y138_SLICE_X0Y138_CLUT (
.I0(RIOB33_X105Y127_IOB_X1Y128_I),
.I1(RIOB33_X105Y137_IOB_X1Y137_I),
.I2(RIOB33_X105Y129_IOB_X1Y129_I),
.I3(CLBLM_R_X3Y152_SLICE_X3Y152_CO6),
.I4(CLBLM_R_X3Y153_SLICE_X2Y153_DO6),
.I5(1'b1),
.O5(CLBLL_L_X2Y138_SLICE_X0Y138_CO5),
.O6(CLBLL_L_X2Y138_SLICE_X0Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffdfffdfffffdfd)
  ) CLBLL_L_X2Y138_SLICE_X0Y138_BLUT (
.I0(RIOB33_X105Y137_IOB_X1Y137_I),
.I1(RIOB33_X105Y129_IOB_X1Y129_I),
.I2(RIOB33_X105Y127_IOB_X1Y128_I),
.I3(CLBLL_L_X2Y151_SLICE_X1Y151_BO6),
.I4(CLBLM_R_X3Y151_SLICE_X3Y151_AO6),
.I5(1'b1),
.O5(CLBLL_L_X2Y138_SLICE_X0Y138_BO5),
.O6(CLBLL_L_X2Y138_SLICE_X0Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffafffefffeff)
  ) CLBLL_L_X2Y138_SLICE_X0Y138_ALUT (
.I0(RIOB33_X105Y129_IOB_X1Y129_I),
.I1(CLBLM_R_X3Y154_SLICE_X2Y154_BO6),
.I2(RIOB33_X105Y127_IOB_X1Y128_I),
.I3(RIOB33_X105Y137_IOB_X1Y137_I),
.I4(CLBLL_L_X2Y153_SLICE_X1Y153_DO6),
.I5(1'b1),
.O5(CLBLL_L_X2Y138_SLICE_X0Y138_AO5),
.O6(CLBLL_L_X2Y138_SLICE_X0Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y138_SLICE_X1Y138_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y138_SLICE_X1Y138_DO5),
.O6(CLBLL_L_X2Y138_SLICE_X1Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y138_SLICE_X1Y138_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y138_SLICE_X1Y138_CO5),
.O6(CLBLL_L_X2Y138_SLICE_X1Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y138_SLICE_X1Y138_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y138_SLICE_X1Y138_BO5),
.O6(CLBLL_L_X2Y138_SLICE_X1Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y138_SLICE_X1Y138_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y138_SLICE_X1Y138_AO5),
.O6(CLBLL_L_X2Y138_SLICE_X1Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y141_SLICE_X0Y141_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y141_SLICE_X0Y141_DO5),
.O6(CLBLL_L_X2Y141_SLICE_X0Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y141_SLICE_X0Y141_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y141_SLICE_X0Y141_CO5),
.O6(CLBLL_L_X2Y141_SLICE_X0Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000eac00000)
  ) CLBLL_L_X2Y141_SLICE_X0Y141_BLUT (
.I0(CLBLL_L_X4Y154_SLICE_X4Y154_CO6),
.I1(CLBLL_L_X2Y151_SLICE_X1Y151_BO6),
.I2(LIOB33_X0Y51_IOB_X0Y51_I),
.I3(CLBLM_R_X3Y148_SLICE_X3Y148_BQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X3Y141_SLICE_X2Y141_BO6),
.O5(CLBLL_L_X2Y141_SLICE_X0Y141_BO5),
.O6(CLBLL_L_X2Y141_SLICE_X0Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffff3fffffbfb)
  ) CLBLL_L_X2Y141_SLICE_X0Y141_ALUT (
.I0(CLBLL_L_X4Y154_SLICE_X4Y154_CO6),
.I1(RIOB33_X105Y137_IOB_X1Y137_I),
.I2(RIOB33_X105Y127_IOB_X1Y128_I),
.I3(CLBLM_R_X3Y150_SLICE_X2Y150_BO6),
.I4(RIOB33_X105Y129_IOB_X1Y129_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y141_SLICE_X0Y141_AO5),
.O6(CLBLL_L_X2Y141_SLICE_X0Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y141_SLICE_X1Y141_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y141_SLICE_X1Y141_DO5),
.O6(CLBLL_L_X2Y141_SLICE_X1Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y141_SLICE_X1Y141_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y141_SLICE_X1Y141_CO5),
.O6(CLBLL_L_X2Y141_SLICE_X1Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y141_SLICE_X1Y141_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y141_SLICE_X1Y141_BO5),
.O6(CLBLL_L_X2Y141_SLICE_X1Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y141_SLICE_X1Y141_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y141_SLICE_X1Y141_AO5),
.O6(CLBLL_L_X2Y141_SLICE_X1Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y142_SLICE_X0Y142_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y142_SLICE_X0Y142_DO5),
.O6(CLBLL_L_X2Y142_SLICE_X0Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y142_SLICE_X0Y142_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y142_SLICE_X0Y142_CO5),
.O6(CLBLL_L_X2Y142_SLICE_X0Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y142_SLICE_X0Y142_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y142_SLICE_X0Y142_BO5),
.O6(CLBLL_L_X2Y142_SLICE_X0Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y142_SLICE_X0Y142_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y142_SLICE_X0Y142_AO5),
.O6(CLBLL_L_X2Y142_SLICE_X0Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y142_SLICE_X1Y142_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y142_SLICE_X1Y142_DO5),
.O6(CLBLL_L_X2Y142_SLICE_X1Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y142_SLICE_X1Y142_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y142_SLICE_X1Y142_CO5),
.O6(CLBLL_L_X2Y142_SLICE_X1Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y142_SLICE_X1Y142_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y142_SLICE_X1Y142_BO5),
.O6(CLBLL_L_X2Y142_SLICE_X1Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8888888800000000)
  ) CLBLL_L_X2Y142_SLICE_X1Y142_ALUT (
.I0(CLBLM_R_X3Y143_SLICE_X3Y143_A5Q),
.I1(CLBLM_R_X3Y143_SLICE_X2Y143_CQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X3Y142_SLICE_X2Y142_BQ),
.O5(CLBLL_L_X2Y142_SLICE_X1Y142_AO5),
.O6(CLBLL_L_X2Y142_SLICE_X1Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y145_SLICE_X0Y145_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y145_SLICE_X0Y145_DO5),
.O6(CLBLL_L_X2Y145_SLICE_X0Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y145_SLICE_X0Y145_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y145_SLICE_X0Y145_CO5),
.O6(CLBLL_L_X2Y145_SLICE_X0Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y145_SLICE_X0Y145_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y145_SLICE_X0Y145_BO5),
.O6(CLBLL_L_X2Y145_SLICE_X0Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y145_SLICE_X0Y145_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y145_SLICE_X0Y145_AO5),
.O6(CLBLL_L_X2Y145_SLICE_X0Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y145_SLICE_X1Y145_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y145_SLICE_X1Y145_AO6),
.Q(CLBLL_L_X2Y145_SLICE_X1Y145_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y145_SLICE_X1Y145_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y145_SLICE_X1Y145_BO6),
.Q(CLBLL_L_X2Y145_SLICE_X1Y145_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y145_SLICE_X1Y145_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y145_SLICE_X1Y145_DO5),
.O6(CLBLL_L_X2Y145_SLICE_X1Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y145_SLICE_X1Y145_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y145_SLICE_X1Y145_CO5),
.O6(CLBLL_L_X2Y145_SLICE_X1Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haf05af05ae04ae04)
  ) CLBLL_L_X2Y145_SLICE_X1Y145_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLL_L_X2Y145_SLICE_X1Y145_BQ),
.I2(CLBLM_R_X3Y144_SLICE_X2Y144_CO6),
.I3(CLBLM_R_X5Y146_SLICE_X6Y146_CQ),
.I4(1'b1),
.I5(CLBLL_L_X4Y145_SLICE_X4Y145_A5Q),
.O5(CLBLL_L_X2Y145_SLICE_X1Y145_BO5),
.O6(CLBLL_L_X2Y145_SLICE_X1Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h888d88d888888888)
  ) CLBLL_L_X2Y145_SLICE_X1Y145_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y152_SLICE_X6Y152_BQ),
.I2(CLBLL_L_X2Y145_SLICE_X1Y145_AQ),
.I3(CLBLM_R_X3Y145_SLICE_X3Y145_D5Q),
.I4(CLBLL_L_X2Y142_SLICE_X1Y142_AO6),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLL_L_X2Y145_SLICE_X1Y145_AO5),
.O6(CLBLL_L_X2Y145_SLICE_X1Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y146_SLICE_X0Y146_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y146_SLICE_X0Y146_DO5),
.O6(CLBLL_L_X2Y146_SLICE_X0Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y146_SLICE_X0Y146_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y146_SLICE_X0Y146_CO5),
.O6(CLBLL_L_X2Y146_SLICE_X0Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y146_SLICE_X0Y146_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y146_SLICE_X0Y146_BO5),
.O6(CLBLL_L_X2Y146_SLICE_X0Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y146_SLICE_X0Y146_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y146_SLICE_X0Y146_AO5),
.O6(CLBLL_L_X2Y146_SLICE_X0Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y146_SLICE_X1Y146_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y146_SLICE_X1Y146_AO6),
.Q(CLBLL_L_X2Y146_SLICE_X1Y146_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y146_SLICE_X1Y146_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y146_SLICE_X1Y146_BO6),
.Q(CLBLL_L_X2Y146_SLICE_X1Y146_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y146_SLICE_X1Y146_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y146_SLICE_X1Y146_CO6),
.Q(CLBLL_L_X2Y146_SLICE_X1Y146_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y146_SLICE_X1Y146_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y146_SLICE_X1Y146_DO5),
.O6(CLBLL_L_X2Y146_SLICE_X1Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0028288888)
  ) CLBLL_L_X2Y146_SLICE_X1Y146_CLUT (
.I0(CLBLM_R_X3Y144_SLICE_X3Y144_BO6),
.I1(CLBLL_L_X2Y146_SLICE_X1Y146_CQ),
.I2(CLBLL_L_X4Y144_SLICE_X4Y144_DO6),
.I3(CLBLL_L_X4Y146_SLICE_X5Y146_CQ),
.I4(CLBLL_L_X2Y146_SLICE_X1Y146_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLL_L_X2Y146_SLICE_X1Y146_CO5),
.O6(CLBLL_L_X2Y146_SLICE_X1Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaac0cf0000)
  ) CLBLL_L_X2Y146_SLICE_X1Y146_BLUT (
.I0(CLBLL_L_X4Y146_SLICE_X4Y146_BQ),
.I1(CLBLL_L_X2Y146_SLICE_X1Y146_BQ),
.I2(CLBLM_R_X3Y144_SLICE_X2Y144_DO6),
.I3(CLBLL_L_X2Y147_SLICE_X1Y147_BO6),
.I4(CLBLM_R_X3Y144_SLICE_X3Y144_BO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLL_L_X2Y146_SLICE_X1Y146_BO5),
.O6(CLBLL_L_X2Y146_SLICE_X1Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc5a005a00)
  ) CLBLL_L_X2Y146_SLICE_X1Y146_ALUT (
.I0(CLBLL_L_X4Y144_SLICE_X4Y144_DO6),
.I1(CLBLL_L_X2Y146_SLICE_X1Y146_BQ),
.I2(CLBLL_L_X2Y146_SLICE_X1Y146_AQ),
.I3(CLBLM_R_X3Y144_SLICE_X3Y144_BO6),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLL_L_X2Y146_SLICE_X1Y146_AO5),
.O6(CLBLL_L_X2Y146_SLICE_X1Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y147_SLICE_X0Y147_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y147_SLICE_X0Y147_DO5),
.O6(CLBLL_L_X2Y147_SLICE_X0Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y147_SLICE_X0Y147_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y147_SLICE_X0Y147_CO5),
.O6(CLBLL_L_X2Y147_SLICE_X0Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y147_SLICE_X0Y147_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y147_SLICE_X0Y147_BO5),
.O6(CLBLL_L_X2Y147_SLICE_X0Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h000f0f0fbbbbbbbb)
  ) CLBLL_L_X2Y147_SLICE_X0Y147_ALUT (
.I0(CLBLM_R_X3Y147_SLICE_X2Y147_BO5),
.I1(CLBLL_L_X2Y153_SLICE_X1Y153_DO6),
.I2(CLBLL_L_X2Y147_SLICE_X1Y147_CO6),
.I3(CLBLL_L_X4Y154_SLICE_X4Y154_CO6),
.I4(CLBLL_L_X4Y150_SLICE_X4Y150_B5Q),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLL_L_X2Y147_SLICE_X0Y147_AO5),
.O6(CLBLL_L_X2Y147_SLICE_X0Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y147_SLICE_X1Y147_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y147_SLICE_X1Y147_BO5),
.Q(CLBLL_L_X2Y147_SLICE_X1Y147_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y147_SLICE_X1Y147_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y147_SLICE_X1Y147_DO5),
.O6(CLBLL_L_X2Y147_SLICE_X1Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8fff8f8f88ff8888)
  ) CLBLL_L_X2Y147_SLICE_X1Y147_CLUT (
.I0(CLBLM_R_X3Y143_SLICE_X2Y143_BQ),
.I1(CLBLM_R_X3Y154_SLICE_X2Y154_BO6),
.I2(CLBLM_R_X11Y147_SLICE_X15Y147_AQ),
.I3(CLBLL_L_X2Y147_SLICE_X1Y147_AO5),
.I4(CLBLM_R_X3Y152_SLICE_X3Y152_CO6),
.I5(CLBLM_R_X3Y153_SLICE_X2Y153_DO6),
.O5(CLBLL_L_X2Y147_SLICE_X1Y147_CO5),
.O6(CLBLL_L_X2Y147_SLICE_X1Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0000000e0c0c0c0)
  ) CLBLL_L_X2Y147_SLICE_X1Y147_BLUT (
.I0(CLBLL_L_X2Y146_SLICE_X1Y146_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X3Y144_SLICE_X3Y144_AQ),
.I3(CLBLL_L_X2Y146_SLICE_X1Y146_BQ),
.I4(CLBLL_L_X2Y146_SLICE_X1Y146_CQ),
.I5(1'b1),
.O5(CLBLL_L_X2Y147_SLICE_X1Y147_BO5),
.O6(CLBLL_L_X2Y147_SLICE_X1Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha2aaa0aaddddffff)
  ) CLBLL_L_X2Y147_SLICE_X1Y147_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X5Y144_SLICE_X7Y144_BQ),
.I2(CLBLL_L_X4Y150_SLICE_X4Y150_B5Q),
.I3(CLBLM_R_X5Y152_SLICE_X7Y152_BQ),
.I4(CLBLM_R_X3Y148_SLICE_X3Y148_AQ),
.I5(1'b1),
.O5(CLBLL_L_X2Y147_SLICE_X1Y147_AO5),
.O6(CLBLL_L_X2Y147_SLICE_X1Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y148_SLICE_X0Y148_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y148_SLICE_X0Y148_DO5),
.O6(CLBLL_L_X2Y148_SLICE_X0Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y148_SLICE_X0Y148_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y148_SLICE_X0Y148_CO5),
.O6(CLBLL_L_X2Y148_SLICE_X0Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y148_SLICE_X0Y148_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y148_SLICE_X0Y148_BO5),
.O6(CLBLL_L_X2Y148_SLICE_X0Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y148_SLICE_X0Y148_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y148_SLICE_X0Y148_AO5),
.O6(CLBLL_L_X2Y148_SLICE_X0Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y148_SLICE_X1Y148_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y148_SLICE_X1Y148_AO6),
.Q(CLBLL_L_X2Y148_SLICE_X1Y148_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y148_SLICE_X1Y148_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y148_SLICE_X1Y148_DO5),
.O6(CLBLL_L_X2Y148_SLICE_X1Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y148_SLICE_X1Y148_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y148_SLICE_X1Y148_CO5),
.O6(CLBLL_L_X2Y148_SLICE_X1Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaafffffabaffff)
  ) CLBLL_L_X2Y148_SLICE_X1Y148_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X3Y148_SLICE_X3Y148_AQ),
.I2(CLBLM_R_X5Y152_SLICE_X7Y152_BQ),
.I3(CLBLM_R_X5Y144_SLICE_X7Y144_BQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLL_L_X4Y150_SLICE_X4Y150_B5Q),
.O5(CLBLL_L_X2Y148_SLICE_X1Y148_BO5),
.O6(CLBLL_L_X2Y148_SLICE_X1Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hd8ddd8ddd888d888)
  ) CLBLL_L_X2Y148_SLICE_X1Y148_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X12Y153_SLICE_X16Y153_AQ),
.I2(CLBLL_L_X2Y148_SLICE_X1Y148_AQ),
.I3(CLBLM_R_X3Y144_SLICE_X2Y144_CO6),
.I4(1'b1),
.I5(CLBLM_R_X3Y144_SLICE_X2Y144_AQ),
.O5(CLBLL_L_X2Y148_SLICE_X1Y148_AO5),
.O6(CLBLL_L_X2Y148_SLICE_X1Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y149_SLICE_X0Y149_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y149_SLICE_X0Y149_DO5),
.O6(CLBLL_L_X2Y149_SLICE_X0Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0011004000000040)
  ) CLBLL_L_X2Y149_SLICE_X0Y149_CLUT (
.I0(CLBLL_L_X2Y152_SLICE_X1Y152_AO5),
.I1(RIOB33_X105Y133_IOB_X1Y133_I),
.I2(LIOB33_X0Y63_IOB_X0Y63_I),
.I3(CLBLM_R_X5Y149_SLICE_X6Y149_CO5),
.I4(RIOB33_X105Y133_IOB_X1Y134_I),
.I5(LIOB33_X0Y57_IOB_X0Y58_I),
.O5(CLBLL_L_X2Y149_SLICE_X0Y149_CO5),
.O6(CLBLL_L_X2Y149_SLICE_X0Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000050040004)
  ) CLBLL_L_X2Y149_SLICE_X0Y149_BLUT (
.I0(CLBLL_L_X2Y152_SLICE_X1Y152_AO5),
.I1(CLBLM_R_X3Y143_SLICE_X2Y143_DQ),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(LIOB33_X0Y57_IOB_X0Y57_I),
.I5(CLBLL_L_X2Y150_SLICE_X0Y150_AO5),
.O5(CLBLL_L_X2Y149_SLICE_X0Y149_BO5),
.O6(CLBLL_L_X2Y149_SLICE_X0Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0044000000100010)
  ) CLBLL_L_X2Y149_SLICE_X0Y149_ALUT (
.I0(CLBLL_L_X2Y152_SLICE_X1Y152_AO5),
.I1(RIOB33_X105Y131_IOB_X1Y132_I),
.I2(CLBLL_L_X2Y148_SLICE_X1Y148_AQ),
.I3(CLBLL_L_X2Y150_SLICE_X0Y150_AO5),
.I4(LIOB33_X0Y55_IOB_X0Y55_I),
.I5(RIOB33_X105Y131_IOB_X1Y131_I),
.O5(CLBLL_L_X2Y149_SLICE_X0Y149_AO5),
.O6(CLBLL_L_X2Y149_SLICE_X0Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000020000)
  ) CLBLL_L_X2Y149_SLICE_X1Y149_DLUT (
.I0(CLBLL_L_X2Y145_SLICE_X1Y145_BQ),
.I1(RIOB33_X105Y131_IOB_X1Y132_I),
.I2(CLBLL_L_X2Y152_SLICE_X1Y152_AO5),
.I3(RIOB33_X105Y133_IOB_X1Y133_I),
.I4(RIOB33_X105Y133_IOB_X1Y134_I),
.I5(RIOB33_X105Y131_IOB_X1Y131_I),
.O5(CLBLL_L_X2Y149_SLICE_X1Y149_DO5),
.O6(CLBLL_L_X2Y149_SLICE_X1Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000373300000500)
  ) CLBLL_L_X2Y149_SLICE_X1Y149_CLUT (
.I0(RIOB33_X105Y131_IOB_X1Y132_I),
.I1(CLBLL_L_X4Y155_SLICE_X4Y155_BO6),
.I2(CLBLL_L_X2Y151_SLICE_X1Y151_AO5),
.I3(CLBLL_L_X4Y146_SLICE_X5Y146_CQ),
.I4(CLBLL_L_X2Y152_SLICE_X1Y152_AO5),
.I5(CLBLL_L_X2Y146_SLICE_X1Y146_BQ),
.O5(CLBLL_L_X2Y149_SLICE_X1Y149_CO5),
.O6(CLBLL_L_X2Y149_SLICE_X1Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haf00af00af00efcc)
  ) CLBLL_L_X2Y149_SLICE_X1Y149_BLUT (
.I0(RIOB33_X105Y129_IOB_X1Y129_I),
.I1(CLBLM_R_X3Y148_SLICE_X3Y148_CQ),
.I2(RIOB33_X105Y137_IOB_X1Y137_I),
.I3(CLBLM_R_X3Y145_SLICE_X3Y145_AQ),
.I4(CLBLL_L_X2Y151_SLICE_X0Y151_CO5),
.I5(CLBLL_L_X2Y152_SLICE_X1Y152_AO5),
.O5(CLBLL_L_X2Y149_SLICE_X1Y149_BO5),
.O6(CLBLL_L_X2Y149_SLICE_X1Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haf00af00bf33af00)
  ) CLBLL_L_X2Y149_SLICE_X1Y149_ALUT (
.I0(RIOB33_X105Y129_IOB_X1Y129_I),
.I1(CLBLL_L_X4Y155_SLICE_X4Y155_BO6),
.I2(RIOB33_X105Y137_IOB_X1Y137_I),
.I3(CLBLM_R_X5Y150_SLICE_X6Y150_AQ),
.I4(CLBLM_R_X3Y144_SLICE_X3Y144_AQ),
.I5(CLBLL_L_X2Y152_SLICE_X1Y152_AO5),
.O5(CLBLL_L_X2Y149_SLICE_X1Y149_AO5),
.O6(CLBLL_L_X2Y149_SLICE_X1Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y150_SLICE_X0Y150_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y150_SLICE_X0Y150_DO5),
.O6(CLBLL_L_X2Y150_SLICE_X0Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y150_SLICE_X0Y150_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y150_SLICE_X0Y150_CO5),
.O6(CLBLL_L_X2Y150_SLICE_X0Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0404040455045504)
  ) CLBLL_L_X2Y150_SLICE_X0Y150_BLUT (
.I0(CLBLL_L_X2Y152_SLICE_X1Y152_AO5),
.I1(LIOB33_X0Y59_IOB_X0Y59_I),
.I2(CLBLL_L_X2Y154_SLICE_X1Y154_BO5),
.I3(CLBLM_R_X3Y149_SLICE_X2Y149_CQ),
.I4(1'b1),
.I5(CLBLL_L_X2Y151_SLICE_X0Y151_CO5),
.O5(CLBLL_L_X2Y150_SLICE_X0Y150_BO5),
.O6(CLBLL_L_X2Y150_SLICE_X0Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafffaffafafafaf)
  ) CLBLL_L_X2Y150_SLICE_X0Y150_ALUT (
.I0(RIOB33_X105Y133_IOB_X1Y133_I),
.I1(1'b1),
.I2(RIOB33_X105Y133_IOB_X1Y134_I),
.I3(RIOB33_X105Y131_IOB_X1Y132_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y150_SLICE_X0Y150_AO5),
.O6(CLBLL_L_X2Y150_SLICE_X0Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0f0a0f0a0f0ecfc)
  ) CLBLL_L_X2Y150_SLICE_X1Y150_DLUT (
.I0(RIOB33_X105Y129_IOB_X1Y129_I),
.I1(LIOB33_X0Y65_IOB_X0Y65_I),
.I2(CLBLM_R_X5Y150_SLICE_X6Y150_A5Q),
.I3(RIOB33_X105Y137_IOB_X1Y137_I),
.I4(CLBLL_L_X2Y152_SLICE_X1Y152_AO5),
.I5(CLBLL_L_X2Y154_SLICE_X1Y154_BO5),
.O5(CLBLL_L_X2Y150_SLICE_X1Y150_DO5),
.O6(CLBLL_L_X2Y150_SLICE_X1Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffafe)
  ) CLBLL_L_X2Y150_SLICE_X1Y150_CLUT (
.I0(CLBLL_L_X2Y149_SLICE_X1Y149_BO6),
.I1(RIOB33_X105Y109_IOB_X1Y109_I),
.I2(CLBLM_R_X3Y150_SLICE_X2Y150_CO6),
.I3(CLBLL_L_X2Y154_SLICE_X1Y154_BO6),
.I4(CLBLL_L_X2Y149_SLICE_X0Y149_CO6),
.I5(CLBLL_L_X2Y149_SLICE_X1Y149_CO6),
.O5(CLBLL_L_X2Y150_SLICE_X1Y150_CO5),
.O6(CLBLL_L_X2Y150_SLICE_X1Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h000a030b000a000a)
  ) CLBLL_L_X2Y150_SLICE_X1Y150_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(RIOB33_X105Y131_IOB_X1Y132_I),
.I2(CLBLL_L_X2Y152_SLICE_X1Y152_AO5),
.I3(CLBLL_L_X2Y154_SLICE_X1Y154_BO5),
.I4(CLBLL_L_X2Y151_SLICE_X1Y151_AO5),
.I5(CLBLM_R_X5Y153_SLICE_X6Y153_A5Q),
.O5(CLBLL_L_X2Y150_SLICE_X1Y150_BO5),
.O6(CLBLL_L_X2Y150_SLICE_X1Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffdfffc)
  ) CLBLL_L_X2Y150_SLICE_X1Y150_ALUT (
.I0(CLBLL_L_X2Y154_SLICE_X1Y154_BO6),
.I1(CLBLM_R_X3Y150_SLICE_X2Y150_AO6),
.I2(CLBLL_L_X2Y149_SLICE_X1Y149_AO6),
.I3(CLBLL_L_X2Y150_SLICE_X1Y150_BO6),
.I4(RIOB33_X105Y107_IOB_X1Y108_I),
.I5(CLBLL_L_X2Y149_SLICE_X0Y149_BO6),
.O5(CLBLL_L_X2Y150_SLICE_X1Y150_AO5),
.O6(CLBLL_L_X2Y150_SLICE_X1Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0aceffff0ace0ace)
  ) CLBLL_L_X2Y151_SLICE_X0Y151_DLUT (
.I0(LIOB33_X0Y53_IOB_X0Y54_I),
.I1(CLBLL_L_X2Y146_SLICE_X1Y146_AQ),
.I2(CLBLL_L_X2Y151_SLICE_X0Y151_AO5),
.I3(CLBLL_L_X2Y151_SLICE_X0Y151_CO6),
.I4(CLBLL_L_X2Y151_SLICE_X0Y151_BO5),
.I5(CLBLM_R_X5Y146_SLICE_X6Y146_A5Q),
.O5(CLBLL_L_X2Y151_SLICE_X0Y151_DO5),
.O6(CLBLL_L_X2Y151_SLICE_X0Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffff7fffdfffd)
  ) CLBLL_L_X2Y151_SLICE_X0Y151_CLUT (
.I0(RIOB33_X105Y133_IOB_X1Y134_I),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(RIOB33_X105Y133_IOB_X1Y133_I),
.I3(RIOB33_X105Y131_IOB_X1Y132_I),
.I4(CLBLL_L_X2Y152_SLICE_X1Y152_AO5),
.I5(1'b1),
.O5(CLBLL_L_X2Y151_SLICE_X0Y151_CO5),
.O6(CLBLL_L_X2Y151_SLICE_X0Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hefffffffffbfffff)
  ) CLBLL_L_X2Y151_SLICE_X0Y151_BLUT (
.I0(CLBLL_L_X2Y152_SLICE_X1Y152_AO5),
.I1(RIOB33_X105Y133_IOB_X1Y134_I),
.I2(RIOB33_X105Y133_IOB_X1Y133_I),
.I3(RIOB33_X105Y131_IOB_X1Y132_I),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y151_SLICE_X0Y151_BO5),
.O6(CLBLL_L_X2Y151_SLICE_X0Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffbfbffffff)
  ) CLBLL_L_X2Y151_SLICE_X0Y151_ALUT (
.I0(CLBLL_L_X2Y152_SLICE_X1Y152_AO5),
.I1(RIOB33_X105Y133_IOB_X1Y134_I),
.I2(RIOB33_X105Y133_IOB_X1Y133_I),
.I3(RIOB33_X105Y131_IOB_X1Y132_I),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y151_SLICE_X0Y151_AO5),
.O6(CLBLL_L_X2Y151_SLICE_X0Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h040404040f0f0404)
  ) CLBLL_L_X2Y151_SLICE_X1Y151_DLUT (
.I0(CLBLL_L_X2Y151_SLICE_X1Y151_AO6),
.I1(LIOB33_X0Y71_IOB_X0Y71_I),
.I2(CLBLL_L_X2Y152_SLICE_X1Y152_AO5),
.I3(1'b1),
.I4(CLBLL_L_X2Y146_SLICE_X1Y146_CQ),
.I5(CLBLL_L_X4Y155_SLICE_X4Y155_BO6),
.O5(CLBLL_L_X2Y151_SLICE_X1Y151_DO5),
.O6(CLBLL_L_X2Y151_SLICE_X1Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffdcdcdc)
  ) CLBLL_L_X2Y151_SLICE_X1Y151_CLUT (
.I0(CLBLL_L_X2Y154_SLICE_X1Y154_CO5),
.I1(CLBLM_R_X3Y156_SLICE_X2Y156_CO6),
.I2(LIOB33_X0Y69_IOB_X0Y70_I),
.I3(CLBLL_L_X4Y151_SLICE_X4Y151_A5Q),
.I4(CLBLM_L_X16Y158_SLICE_X22Y158_AO5),
.I5(CLBLL_L_X2Y150_SLICE_X0Y150_BO6),
.O5(CLBLL_L_X2Y151_SLICE_X1Y151_CO5),
.O6(CLBLL_L_X2Y151_SLICE_X1Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLL_L_X2Y151_SLICE_X1Y151_BLUT (
.I0(CLBLM_R_X3Y150_SLICE_X2Y150_DO6),
.I1(CLBLL_L_X2Y151_SLICE_X0Y151_DO6),
.I2(CLBLM_R_X5Y153_SLICE_X6Y153_DO6),
.I3(CLBLM_R_X3Y152_SLICE_X3Y152_BO6),
.I4(CLBLM_R_X3Y155_SLICE_X2Y155_DO6),
.I5(CLBLL_L_X2Y151_SLICE_X1Y151_CO6),
.O5(CLBLL_L_X2Y151_SLICE_X1Y151_BO5),
.O6(CLBLL_L_X2Y151_SLICE_X1Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff7fff75fff5fff)
  ) CLBLL_L_X2Y151_SLICE_X1Y151_ALUT (
.I0(RIOB33_X105Y133_IOB_X1Y133_I),
.I1(RIOB33_X105Y131_IOB_X1Y132_I),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(RIOB33_X105Y133_IOB_X1Y134_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y151_SLICE_X1Y151_AO5),
.O6(CLBLL_L_X2Y151_SLICE_X1Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y152_SLICE_X0Y152_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y152_SLICE_X0Y152_DO5),
.O6(CLBLL_L_X2Y152_SLICE_X0Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y152_SLICE_X0Y152_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y152_SLICE_X0Y152_CO5),
.O6(CLBLL_L_X2Y152_SLICE_X0Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y152_SLICE_X0Y152_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y152_SLICE_X0Y152_BO5),
.O6(CLBLL_L_X2Y152_SLICE_X0Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y152_SLICE_X0Y152_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y152_SLICE_X0Y152_AO5),
.O6(CLBLL_L_X2Y152_SLICE_X0Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f33bfbb0f00afaa)
  ) CLBLL_L_X2Y152_SLICE_X1Y152_DLUT (
.I0(CLBLL_L_X4Y151_SLICE_X5Y151_AQ),
.I1(CLBLL_L_X4Y155_SLICE_X5Y155_AO6),
.I2(CLBLL_L_X2Y154_SLICE_X1Y154_BO6),
.I3(RIOB33_X105Y111_IOB_X1Y112_I),
.I4(CLBLL_L_X2Y152_SLICE_X1Y152_BO5),
.I5(CLBLM_R_X3Y145_SLICE_X3Y145_BQ),
.O5(CLBLL_L_X2Y152_SLICE_X1Y152_DO5),
.O6(CLBLL_L_X2Y152_SLICE_X1Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h111f1111000f0000)
  ) CLBLL_L_X2Y152_SLICE_X1Y152_CLUT (
.I0(CLBLL_L_X2Y152_SLICE_X1Y152_AO6),
.I1(CLBLL_L_X4Y155_SLICE_X4Y155_BO6),
.I2(CLBLL_L_X2Y154_SLICE_X1Y154_BO5),
.I3(CLBLL_L_X2Y155_SLICE_X1Y155_DO6),
.I4(CLBLM_R_X3Y145_SLICE_X3Y145_BQ),
.I5(CLBLL_L_X4Y151_SLICE_X5Y151_AQ),
.O5(CLBLL_L_X2Y152_SLICE_X1Y152_CO5),
.O6(CLBLL_L_X2Y152_SLICE_X1Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffbfffffffffdf)
  ) CLBLL_L_X2Y152_SLICE_X1Y152_BLUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(RIOB33_X105Y133_IOB_X1Y133_I),
.I2(RIOB33_X105Y133_IOB_X1Y134_I),
.I3(RIOB33_X105Y131_IOB_X1Y132_I),
.I4(CLBLL_L_X2Y152_SLICE_X1Y152_AO6),
.I5(1'b1),
.O5(CLBLL_L_X2Y152_SLICE_X1Y152_BO5),
.O6(CLBLL_L_X2Y152_SLICE_X1Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffefffffefffff)
  ) CLBLL_L_X2Y152_SLICE_X1Y152_ALUT (
.I0(RIOB33_X105Y129_IOB_X1Y129_I),
.I1(RIOB33_X105Y129_IOB_X1Y130_I),
.I2(RIOB33_X105Y137_IOB_X1Y137_I),
.I3(RIOB33_X105Y135_IOB_X1Y136_I),
.I4(RIOB33_X105Y135_IOB_X1Y135_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y152_SLICE_X1Y152_AO5),
.O6(CLBLL_L_X2Y152_SLICE_X1Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y153_SLICE_X0Y153_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y153_SLICE_X0Y153_DO5),
.O6(CLBLL_L_X2Y153_SLICE_X0Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y153_SLICE_X0Y153_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y153_SLICE_X0Y153_CO5),
.O6(CLBLL_L_X2Y153_SLICE_X0Y153_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y153_SLICE_X0Y153_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y153_SLICE_X0Y153_BO5),
.O6(CLBLL_L_X2Y153_SLICE_X0Y153_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y153_SLICE_X0Y153_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y153_SLICE_X0Y153_AO5),
.O6(CLBLL_L_X2Y153_SLICE_X0Y153_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffdcdc)
  ) CLBLL_L_X2Y153_SLICE_X1Y153_DLUT (
.I0(CLBLL_L_X2Y155_SLICE_X1Y155_AO6),
.I1(CLBLL_L_X4Y151_SLICE_X5Y151_CO6),
.I2(CLBLL_L_X2Y152_SLICE_X1Y152_BO5),
.I3(1'b1),
.I4(CLBLL_L_X2Y152_SLICE_X1Y152_DO6),
.I5(CLBLL_L_X2Y153_SLICE_X1Y153_BO6),
.O5(CLBLL_L_X2Y153_SLICE_X1Y153_DO5),
.O6(CLBLL_L_X2Y153_SLICE_X1Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h050f0505000f0000)
  ) CLBLL_L_X2Y153_SLICE_X1Y153_CLUT (
.I0(CLBLL_L_X2Y151_SLICE_X0Y151_CO5),
.I1(1'b1),
.I2(CLBLL_L_X2Y152_SLICE_X1Y152_AO5),
.I3(CLBLL_L_X2Y154_SLICE_X1Y154_BO5),
.I4(LIOB33_X0Y67_IOB_X0Y67_I),
.I5(CLBLM_R_X3Y150_SLICE_X3Y150_BQ),
.O5(CLBLL_L_X2Y153_SLICE_X1Y153_CO5),
.O6(CLBLL_L_X2Y153_SLICE_X1Y153_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffff2fff22)
  ) CLBLL_L_X2Y153_SLICE_X1Y153_BLUT (
.I0(LIOB33_X0Y67_IOB_X0Y67_I),
.I1(CLBLL_L_X2Y151_SLICE_X0Y151_BO6),
.I2(CLBLL_L_X2Y151_SLICE_X0Y151_AO6),
.I3(CLBLL_L_X4Y152_SLICE_X5Y152_BO6),
.I4(CLBLM_R_X3Y150_SLICE_X3Y150_BQ),
.I5(CLBLL_L_X4Y153_SLICE_X4Y153_CO6),
.O5(CLBLL_L_X2Y153_SLICE_X1Y153_BO5),
.O6(CLBLL_L_X2Y153_SLICE_X1Y153_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffff4)
  ) CLBLL_L_X2Y153_SLICE_X1Y153_ALUT (
.I0(CLBLL_L_X2Y154_SLICE_X1Y154_BO6),
.I1(RIOB33_X105Y111_IOB_X1Y112_I),
.I2(CLBLL_L_X2Y152_SLICE_X1Y152_CO6),
.I3(CLBLL_L_X4Y152_SLICE_X5Y152_BO6),
.I4(CLBLL_L_X2Y153_SLICE_X1Y153_CO6),
.I5(CLBLL_L_X4Y153_SLICE_X4Y153_CO6),
.O5(CLBLL_L_X2Y153_SLICE_X1Y153_AO5),
.O6(CLBLL_L_X2Y153_SLICE_X1Y153_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y154_SLICE_X0Y154_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y154_SLICE_X0Y154_DO5),
.O6(CLBLL_L_X2Y154_SLICE_X0Y154_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y154_SLICE_X0Y154_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y154_SLICE_X0Y154_CO5),
.O6(CLBLL_L_X2Y154_SLICE_X0Y154_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y154_SLICE_X0Y154_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y154_SLICE_X0Y154_BO5),
.O6(CLBLL_L_X2Y154_SLICE_X0Y154_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y154_SLICE_X0Y154_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y154_SLICE_X0Y154_AO5),
.O6(CLBLL_L_X2Y154_SLICE_X0Y154_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y154_SLICE_X1Y154_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y154_SLICE_X1Y154_DO5),
.O6(CLBLL_L_X2Y154_SLICE_X1Y154_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h10312000fffffdff)
  ) CLBLL_L_X2Y154_SLICE_X1Y154_CLUT (
.I0(RIOB33_X105Y131_IOB_X1Y132_I),
.I1(CLBLL_L_X2Y152_SLICE_X1Y152_AO5),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(RIOB33_X105Y133_IOB_X1Y133_I),
.I4(RIOB33_X105Y133_IOB_X1Y134_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y154_SLICE_X1Y154_CO5),
.O6(CLBLL_L_X2Y154_SLICE_X1Y154_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbffffffbbffffff)
  ) CLBLL_L_X2Y154_SLICE_X1Y154_BLUT (
.I0(RIOB33_X105Y133_IOB_X1Y134_I),
.I1(RIOB33_X105Y131_IOB_X1Y132_I),
.I2(CLBLL_L_X2Y152_SLICE_X1Y152_AO6),
.I3(RIOB33_X105Y133_IOB_X1Y133_I),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y154_SLICE_X1Y154_BO5),
.O6(CLBLL_L_X2Y154_SLICE_X1Y154_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3fff7fdf7ffffff)
  ) CLBLL_L_X2Y154_SLICE_X1Y154_ALUT (
.I0(RIOB33_X105Y133_IOB_X1Y134_I),
.I1(RIOB33_X105Y131_IOB_X1Y132_I),
.I2(CLBLL_L_X2Y152_SLICE_X1Y152_AO6),
.I3(RIOB33_X105Y133_IOB_X1Y133_I),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y154_SLICE_X1Y154_AO5),
.O6(CLBLL_L_X2Y154_SLICE_X1Y154_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y155_SLICE_X0Y155_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y155_SLICE_X0Y155_DO5),
.O6(CLBLL_L_X2Y155_SLICE_X0Y155_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y155_SLICE_X0Y155_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y155_SLICE_X0Y155_CO5),
.O6(CLBLL_L_X2Y155_SLICE_X0Y155_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y155_SLICE_X0Y155_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y155_SLICE_X0Y155_BO5),
.O6(CLBLL_L_X2Y155_SLICE_X0Y155_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y155_SLICE_X0Y155_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y155_SLICE_X0Y155_AO5),
.O6(CLBLL_L_X2Y155_SLICE_X0Y155_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffefef)
  ) CLBLL_L_X2Y155_SLICE_X1Y155_DLUT (
.I0(RIOB33_X105Y129_IOB_X1Y129_I),
.I1(RIOB33_X105Y135_IOB_X1Y136_I),
.I2(RIOB33_X105Y137_IOB_X1Y137_I),
.I3(1'b1),
.I4(RIOB33_X105Y135_IOB_X1Y135_I),
.I5(RIOB33_X105Y129_IOB_X1Y130_I),
.O5(CLBLL_L_X2Y155_SLICE_X1Y155_DO5),
.O6(CLBLL_L_X2Y155_SLICE_X1Y155_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000ffffffdf)
  ) CLBLL_L_X2Y155_SLICE_X1Y155_CLUT (
.I0(RIOB33_X105Y133_IOB_X1Y133_I),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(CLBLL_L_X2Y152_SLICE_X1Y152_AO5),
.I4(RIOB33_X105Y133_IOB_X1Y134_I),
.I5(CLBLM_L_X16Y158_SLICE_X22Y158_AO5),
.O5(CLBLL_L_X2Y155_SLICE_X1Y155_CO5),
.O6(CLBLL_L_X2Y155_SLICE_X1Y155_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbffffffffffffff)
  ) CLBLL_L_X2Y155_SLICE_X1Y155_BLUT (
.I0(CLBLL_L_X2Y154_SLICE_X1Y154_CO6),
.I1(CLBLL_L_X2Y154_SLICE_X1Y154_AO6),
.I2(CLBLM_R_X3Y156_SLICE_X2Y156_CO6),
.I3(CLBLM_R_X3Y155_SLICE_X3Y155_AO6),
.I4(CLBLL_L_X4Y154_SLICE_X5Y154_CO6),
.I5(CLBLL_L_X2Y155_SLICE_X1Y155_CO6),
.O5(CLBLL_L_X2Y155_SLICE_X1Y155_BO5),
.O6(CLBLL_L_X2Y155_SLICE_X1Y155_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffbfffffff)
  ) CLBLL_L_X2Y155_SLICE_X1Y155_ALUT (
.I0(CLBLL_L_X2Y154_SLICE_X1Y154_CO6),
.I1(CLBLL_L_X2Y154_SLICE_X1Y154_AO6),
.I2(CLBLL_L_X2Y154_SLICE_X1Y154_CO5),
.I3(CLBLM_R_X3Y155_SLICE_X3Y155_AO6),
.I4(CLBLL_L_X4Y154_SLICE_X5Y154_CO6),
.I5(CLBLM_L_X16Y158_SLICE_X22Y158_AO5),
.O5(CLBLL_L_X2Y155_SLICE_X1Y155_AO5),
.O6(CLBLL_L_X2Y155_SLICE_X1Y155_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y142_SLICE_X4Y142_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y142_SLICE_X4Y142_DO5),
.O6(CLBLL_L_X4Y142_SLICE_X4Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y142_SLICE_X4Y142_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y142_SLICE_X4Y142_CO5),
.O6(CLBLL_L_X4Y142_SLICE_X4Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y142_SLICE_X4Y142_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y142_SLICE_X4Y142_BO5),
.O6(CLBLL_L_X4Y142_SLICE_X4Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y142_SLICE_X4Y142_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y142_SLICE_X4Y142_AO5),
.O6(CLBLL_L_X4Y142_SLICE_X4Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y142_SLICE_X5Y142_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y142_SLICE_X5Y142_AO6),
.Q(CLBLL_L_X4Y142_SLICE_X5Y142_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y142_SLICE_X5Y142_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y142_SLICE_X5Y142_DO5),
.O6(CLBLL_L_X4Y142_SLICE_X5Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y142_SLICE_X5Y142_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y142_SLICE_X5Y142_CO5),
.O6(CLBLL_L_X4Y142_SLICE_X5Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y142_SLICE_X5Y142_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y142_SLICE_X5Y142_BO5),
.O6(CLBLL_L_X4Y142_SLICE_X5Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcc00ccf7f7f7f7)
  ) CLBLL_L_X4Y142_SLICE_X5Y142_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLL_L_X4Y147_SLICE_X5Y147_CQ),
.I2(CLBLL_L_X4Y142_SLICE_X5Y142_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X5Y151_SLICE_X6Y151_DQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y142_SLICE_X5Y142_AO5),
.O6(CLBLL_L_X4Y142_SLICE_X5Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y143_SLICE_X4Y143_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y143_SLICE_X4Y143_AO6),
.Q(CLBLL_L_X4Y143_SLICE_X4Y143_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y143_SLICE_X4Y143_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y143_SLICE_X4Y143_BO6),
.Q(CLBLL_L_X4Y143_SLICE_X4Y143_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y143_SLICE_X4Y143_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y143_SLICE_X4Y143_DO5),
.O6(CLBLL_L_X4Y143_SLICE_X4Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hc00000002a000000)
  ) CLBLL_L_X4Y143_SLICE_X4Y143_CLUT (
.I0(CLBLM_R_X7Y142_SLICE_X8Y142_DO6),
.I1(CLBLL_L_X4Y143_SLICE_X4Y143_AQ),
.I2(CLBLL_L_X4Y144_SLICE_X5Y144_BQ),
.I3(CLBLL_L_X4Y144_SLICE_X5Y144_AQ),
.I4(CLBLL_L_X4Y144_SLICE_X5Y144_A5Q),
.I5(1'b1),
.O5(CLBLL_L_X4Y143_SLICE_X4Y143_CO5),
.O6(CLBLL_L_X4Y143_SLICE_X4Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000ffc000c0)
  ) CLBLL_L_X4Y143_SLICE_X4Y143_BLUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y143_SLICE_X4Y143_BQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X3Y142_SLICE_X2Y142_AQ),
.I5(CLBLM_R_X5Y148_SLICE_X7Y148_CQ),
.O5(CLBLL_L_X4Y143_SLICE_X4Y143_BO5),
.O6(CLBLL_L_X4Y143_SLICE_X4Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff04ff4000040040)
  ) CLBLL_L_X4Y143_SLICE_X4Y143_ALUT (
.I0(CLBLM_L_X8Y145_SLICE_X11Y145_AQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLL_L_X4Y143_SLICE_X4Y143_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLL_L_X4Y143_SLICE_X4Y143_CO5),
.I5(CLBLM_R_X3Y143_SLICE_X2Y143_DQ),
.O5(CLBLL_L_X4Y143_SLICE_X4Y143_AO5),
.O6(CLBLL_L_X4Y143_SLICE_X4Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y143_SLICE_X5Y143_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y143_SLICE_X5Y143_DO5),
.O6(CLBLL_L_X4Y143_SLICE_X5Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y143_SLICE_X5Y143_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y143_SLICE_X5Y143_CO5),
.O6(CLBLL_L_X4Y143_SLICE_X5Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y143_SLICE_X5Y143_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y143_SLICE_X5Y143_BO5),
.O6(CLBLL_L_X4Y143_SLICE_X5Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h004400ccff33ff33)
  ) CLBLL_L_X4Y143_SLICE_X5Y143_ALUT (
.I0(CLBLL_L_X4Y144_SLICE_X5Y144_BQ),
.I1(CLBLL_L_X4Y144_SLICE_X5Y144_AQ),
.I2(1'b1),
.I3(CLBLL_L_X4Y145_SLICE_X5Y145_DO6),
.I4(CLBLL_L_X4Y143_SLICE_X4Y143_AQ),
.I5(CLBLL_L_X4Y144_SLICE_X5Y144_A5Q),
.O5(CLBLL_L_X4Y143_SLICE_X5Y143_AO5),
.O6(CLBLL_L_X4Y143_SLICE_X5Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y144_SLICE_X4Y144_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y144_SLICE_X4Y144_AO6),
.Q(CLBLL_L_X4Y144_SLICE_X4Y144_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y144_SLICE_X4Y144_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y144_SLICE_X4Y144_BO6),
.Q(CLBLL_L_X4Y144_SLICE_X4Y144_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0008000000000000)
  ) CLBLL_L_X4Y144_SLICE_X4Y144_DLUT (
.I0(CLBLL_L_X4Y144_SLICE_X5Y144_AQ),
.I1(CLBLL_L_X4Y144_SLICE_X5Y144_A5Q),
.I2(CLBLM_L_X8Y144_SLICE_X11Y144_BO6),
.I3(CLBLM_R_X7Y142_SLICE_X8Y142_DO6),
.I4(CLBLL_L_X4Y143_SLICE_X4Y143_AQ),
.I5(CLBLL_L_X4Y144_SLICE_X5Y144_BQ),
.O5(CLBLL_L_X4Y144_SLICE_X4Y144_DO5),
.O6(CLBLL_L_X4Y144_SLICE_X4Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff153f80008000)
  ) CLBLL_L_X4Y144_SLICE_X4Y144_CLUT (
.I0(CLBLM_R_X3Y145_SLICE_X2Y145_BQ),
.I1(CLBLM_R_X5Y144_SLICE_X6Y144_AQ),
.I2(CLBLM_R_X3Y145_SLICE_X2Y145_A5Q),
.I3(CLBLM_R_X3Y145_SLICE_X3Y145_CQ),
.I4(CLBLM_R_X3Y144_SLICE_X3Y144_CO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y144_SLICE_X4Y144_CO5),
.O6(CLBLL_L_X4Y144_SLICE_X4Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hba30eac0ba30eac0)
  ) CLBLL_L_X4Y144_SLICE_X4Y144_BLUT (
.I0(CLBLL_L_X4Y154_SLICE_X5Y154_AQ),
.I1(CLBLL_L_X4Y144_SLICE_X4Y144_BQ),
.I2(CLBLM_R_X5Y144_SLICE_X6Y144_BO6),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLL_L_X4Y144_SLICE_X4Y144_CO5),
.I5(1'b1),
.O5(CLBLL_L_X4Y144_SLICE_X4Y144_BO5),
.O6(CLBLL_L_X4Y144_SLICE_X4Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa3caaf0aa00aa00)
  ) CLBLL_L_X4Y144_SLICE_X4Y144_ALUT (
.I0(CLBLM_R_X7Y145_SLICE_X9Y145_CQ),
.I1(CLBLL_L_X4Y144_SLICE_X4Y144_BQ),
.I2(CLBLL_L_X4Y144_SLICE_X4Y144_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLL_L_X4Y144_SLICE_X4Y144_CO5),
.I5(CLBLM_R_X5Y144_SLICE_X6Y144_BO5),
.O5(CLBLL_L_X4Y144_SLICE_X4Y144_AO5),
.O6(CLBLL_L_X4Y144_SLICE_X4Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y144_SLICE_X5Y144_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y144_SLICE_X5Y144_CO6),
.Q(CLBLL_L_X4Y144_SLICE_X5Y144_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y144_SLICE_X5Y144_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y144_SLICE_X5Y144_AO6),
.Q(CLBLL_L_X4Y144_SLICE_X5Y144_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y144_SLICE_X5Y144_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y144_SLICE_X5Y144_BO6),
.Q(CLBLL_L_X4Y144_SLICE_X5Y144_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffeff)
  ) CLBLL_L_X4Y144_SLICE_X5Y144_DLUT (
.I0(CLBLM_R_X3Y144_SLICE_X2Y144_A5Q),
.I1(CLBLM_R_X3Y145_SLICE_X3Y145_A5Q),
.I2(CLBLL_L_X4Y145_SLICE_X5Y145_BO5),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X3Y149_SLICE_X3Y149_B5Q),
.I5(CLBLM_R_X7Y145_SLICE_X8Y145_C5Q),
.O5(CLBLL_L_X4Y144_SLICE_X5Y144_DO5),
.O6(CLBLL_L_X4Y144_SLICE_X5Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc05cc00000f0000)
  ) CLBLL_L_X4Y144_SLICE_X5Y144_CLUT (
.I0(CLBLL_L_X4Y143_SLICE_X5Y143_AO6),
.I1(CLBLM_L_X10Y145_SLICE_X12Y145_AQ),
.I2(CLBLM_L_X8Y145_SLICE_X11Y145_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y144_SLICE_X5Y144_CO5),
.O6(CLBLL_L_X4Y144_SLICE_X5Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffecff00ecec0000)
  ) CLBLL_L_X4Y144_SLICE_X5Y144_BLUT (
.I0(CLBLL_L_X4Y143_SLICE_X4Y143_AQ),
.I1(CLBLL_L_X4Y144_SLICE_X5Y144_BQ),
.I2(CLBLL_L_X4Y143_SLICE_X4Y143_CO5),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLL_L_X4Y144_SLICE_X5Y144_CO5),
.I5(CLBLL_L_X4Y149_SLICE_X5Y149_DQ),
.O5(CLBLL_L_X4Y144_SLICE_X5Y144_BO5),
.O6(CLBLL_L_X4Y144_SLICE_X5Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff888888ff88888)
  ) CLBLL_L_X4Y144_SLICE_X5Y144_ALUT (
.I0(CLBLM_R_X5Y155_SLICE_X6Y155_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLL_L_X4Y144_SLICE_X5Y144_AQ),
.I3(CLBLM_R_X7Y142_SLICE_X8Y142_DO6),
.I4(CLBLL_L_X4Y144_SLICE_X5Y144_CO5),
.I5(CLBLL_L_X4Y143_SLICE_X4Y143_CO6),
.O5(CLBLL_L_X4Y144_SLICE_X5Y144_AO5),
.O6(CLBLL_L_X4Y144_SLICE_X5Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y145_SLICE_X4Y145_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y146_SLICE_X4Y146_CO6),
.Q(CLBLL_L_X4Y145_SLICE_X4Y145_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y145_SLICE_X4Y145_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y145_SLICE_X4Y145_AO6),
.Q(CLBLL_L_X4Y145_SLICE_X4Y145_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y145_SLICE_X4Y145_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y145_SLICE_X4Y145_BO6),
.Q(CLBLL_L_X4Y145_SLICE_X4Y145_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y145_SLICE_X4Y145_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y145_SLICE_X4Y145_CO6),
.Q(CLBLL_L_X4Y145_SLICE_X4Y145_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafafafafafafafa)
  ) CLBLL_L_X4Y145_SLICE_X4Y145_DLUT (
.I0(CLBLM_R_X3Y149_SLICE_X3Y149_B5Q),
.I1(1'b1),
.I2(CLBLM_R_X3Y145_SLICE_X3Y145_A5Q),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y145_SLICE_X4Y145_DO5),
.O6(CLBLL_L_X4Y145_SLICE_X4Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff06ff0c0006000c)
  ) CLBLL_L_X4Y145_SLICE_X4Y145_CLUT (
.I0(CLBLM_R_X7Y147_SLICE_X8Y147_AQ),
.I1(CLBLL_L_X4Y145_SLICE_X4Y145_CQ),
.I2(CLBLM_R_X11Y146_SLICE_X14Y146_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLL_L_X4Y145_SLICE_X4Y145_BO5),
.I5(CLBLM_L_X10Y146_SLICE_X12Y146_C5Q),
.O5(CLBLL_L_X4Y145_SLICE_X4Y145_CO5),
.O6(CLBLL_L_X4Y145_SLICE_X4Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000e0e44444444)
  ) CLBLL_L_X4Y145_SLICE_X4Y145_BLUT (
.I0(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_R_X7Y145_SLICE_X8Y145_DO6),
.I3(CLBLM_R_X3Y143_SLICE_X2Y143_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y145_SLICE_X4Y145_BO5),
.O6(CLBLL_L_X4Y145_SLICE_X4Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffccff00fcccf000)
  ) CLBLL_L_X4Y145_SLICE_X4Y145_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLL_L_X4Y145_SLICE_X4Y145_AQ),
.I3(CLBLM_R_X5Y152_SLICE_X7Y152_DO6),
.I4(CLBLM_L_X10Y145_SLICE_X13Y145_AQ),
.I5(CLBLM_R_X7Y149_SLICE_X8Y149_DQ),
.O5(CLBLL_L_X4Y145_SLICE_X4Y145_AO5),
.O6(CLBLL_L_X4Y145_SLICE_X4Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y145_SLICE_X5Y145_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y145_SLICE_X5Y145_AO6),
.Q(CLBLL_L_X4Y145_SLICE_X5Y145_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffeff)
  ) CLBLL_L_X4Y145_SLICE_X5Y145_DLUT (
.I0(CLBLM_R_X7Y145_SLICE_X8Y145_C5Q),
.I1(CLBLM_R_X3Y151_SLICE_X2Y151_AO6),
.I2(CLBLL_L_X4Y145_SLICE_X4Y145_DO6),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X5Y152_SLICE_X7Y152_B5Q),
.I5(CLBLL_L_X4Y145_SLICE_X5Y145_BO6),
.O5(CLBLL_L_X4Y145_SLICE_X5Y145_DO5),
.O6(CLBLL_L_X4Y145_SLICE_X5Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaabbabffffffff)
  ) CLBLL_L_X4Y145_SLICE_X5Y145_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(LIOB33_X0Y53_IOB_X0Y53_I),
.I2(CLBLL_L_X4Y147_SLICE_X5Y147_CQ),
.I3(CLBLL_L_X4Y142_SLICE_X5Y142_AQ),
.I4(CLBLM_R_X5Y145_SLICE_X6Y145_A5Q),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLL_L_X4Y145_SLICE_X5Y145_CO5),
.O6(CLBLL_L_X4Y145_SLICE_X5Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffefffffffa)
  ) CLBLL_L_X4Y145_SLICE_X5Y145_BLUT (
.I0(CLBLM_R_X3Y143_SLICE_X3Y143_B5Q),
.I1(CLBLM_R_X3Y144_SLICE_X2Y144_A5Q),
.I2(CLBLM_R_X3Y144_SLICE_X2Y144_AQ),
.I3(CLBLL_L_X4Y145_SLICE_X4Y145_A5Q),
.I4(CLBLL_L_X4Y148_SLICE_X4Y148_C5Q),
.I5(1'b1),
.O5(CLBLL_L_X4Y145_SLICE_X5Y145_BO5),
.O6(CLBLL_L_X4Y145_SLICE_X5Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffc400c4fff700f7)
  ) CLBLL_L_X4Y145_SLICE_X5Y145_ALUT (
.I0(CLBLL_L_X4Y147_SLICE_X5Y147_CQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLL_L_X4Y142_SLICE_X5Y142_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X11Y145_SLICE_X14Y145_AQ),
.I5(LIOB33_X0Y53_IOB_X0Y53_I),
.O5(CLBLL_L_X4Y145_SLICE_X5Y145_AO5),
.O6(CLBLL_L_X4Y145_SLICE_X5Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y146_SLICE_X4Y146_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y146_SLICE_X8Y146_BO6),
.Q(CLBLL_L_X4Y146_SLICE_X4Y146_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y146_SLICE_X4Y146_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y146_SLICE_X4Y146_AO6),
.Q(CLBLL_L_X4Y146_SLICE_X4Y146_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y146_SLICE_X4Y146_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y146_SLICE_X4Y146_BO6),
.Q(CLBLL_L_X4Y146_SLICE_X4Y146_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0800000000000000)
  ) CLBLL_L_X4Y146_SLICE_X4Y146_DLUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLL_L_X4Y145_SLICE_X4Y145_CQ),
.I2(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.I3(CLBLM_R_X7Y147_SLICE_X8Y147_AQ),
.I4(CLBLM_R_X5Y145_SLICE_X7Y145_AQ),
.I5(CLBLM_R_X7Y145_SLICE_X8Y145_AQ),
.O5(CLBLL_L_X4Y146_SLICE_X4Y146_DO5),
.O6(CLBLL_L_X4Y146_SLICE_X4Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5a0a0333f333f)
  ) CLBLL_L_X4Y146_SLICE_X4Y146_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y121_IOB_X1Y121_I),
.I2(CLBLM_L_X8Y147_SLICE_X10Y147_CQ),
.I3(CLBLM_L_X10Y146_SLICE_X13Y146_B5Q),
.I4(CLBLM_R_X3Y146_SLICE_X2Y146_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y146_SLICE_X4Y146_CO5),
.O6(CLBLL_L_X4Y146_SLICE_X4Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa0faa0caa00aa00)
  ) CLBLL_L_X4Y146_SLICE_X4Y146_BLUT (
.I0(CLBLL_L_X4Y147_SLICE_X5Y147_CQ),
.I1(CLBLL_L_X4Y146_SLICE_X4Y146_BQ),
.I2(RIOB33_X105Y117_IOB_X1Y118_I),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X11Y146_SLICE_X15Y146_DQ),
.I5(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.O5(CLBLL_L_X4Y146_SLICE_X4Y146_BO5),
.O6(CLBLL_L_X4Y146_SLICE_X4Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffe4ffcc00e400cc)
  ) CLBLL_L_X4Y146_SLICE_X4Y146_ALUT (
.I0(CLBLM_L_X8Y149_SLICE_X11Y149_AQ),
.I1(CLBLM_R_X5Y145_SLICE_X7Y145_AQ),
.I2(CLBLL_L_X4Y146_SLICE_X4Y146_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLL_L_X4Y151_SLICE_X4Y151_AQ),
.I5(CLBLM_R_X3Y146_SLICE_X2Y146_AQ),
.O5(CLBLL_L_X4Y146_SLICE_X4Y146_AO5),
.O6(CLBLL_L_X4Y146_SLICE_X4Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y146_SLICE_X5Y146_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y146_SLICE_X5Y146_BO6),
.Q(CLBLL_L_X4Y146_SLICE_X5Y146_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y146_SLICE_X5Y146_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y146_SLICE_X5Y146_AO6),
.Q(CLBLL_L_X4Y146_SLICE_X5Y146_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y146_SLICE_X5Y146_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y146_SLICE_X5Y146_CO6),
.Q(CLBLL_L_X4Y146_SLICE_X5Y146_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fff7fffffffffff)
  ) CLBLL_L_X4Y146_SLICE_X5Y146_DLUT (
.I0(CLBLM_R_X7Y146_SLICE_X8Y146_C5Q),
.I1(CLBLM_R_X11Y147_SLICE_X14Y147_BQ),
.I2(CLBLM_R_X3Y147_SLICE_X3Y147_BQ),
.I3(CLBLM_L_X8Y146_SLICE_X10Y146_BQ),
.I4(1'b1),
.I5(CLBLL_L_X4Y147_SLICE_X5Y147_BQ),
.O5(CLBLL_L_X4Y146_SLICE_X5Y146_DO5),
.O6(CLBLL_L_X4Y146_SLICE_X5Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0cff0c0c0c0c0c)
  ) CLBLL_L_X4Y146_SLICE_X5Y146_CLUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y146_SLICE_X5Y146_CQ),
.I2(CLBLL_L_X4Y145_SLICE_X5Y145_CO6),
.I3(CLBLM_L_X12Y144_SLICE_X16Y144_CQ),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLL_L_X4Y146_SLICE_X5Y146_CO5),
.O6(CLBLL_L_X4Y146_SLICE_X5Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcac0cac0cccc0000)
  ) CLBLL_L_X4Y146_SLICE_X5Y146_BLUT (
.I0(CLBLM_R_X7Y146_SLICE_X8Y146_DQ),
.I1(CLBLL_L_X4Y147_SLICE_X5Y147_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X3Y146_SLICE_X3Y146_BQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y146_SLICE_X5Y146_BO5),
.O6(CLBLL_L_X4Y146_SLICE_X5Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff005454fcfc)
  ) CLBLL_L_X4Y146_SLICE_X5Y146_ALUT (
.I0(CLBLM_L_X8Y149_SLICE_X11Y149_AQ),
.I1(CLBLL_L_X4Y147_SLICE_X5Y147_BQ),
.I2(CLBLL_L_X4Y146_SLICE_X5Y146_AQ),
.I3(CLBLM_R_X7Y146_SLICE_X8Y146_C5Q),
.I4(CLBLL_L_X4Y151_SLICE_X4Y151_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLL_L_X4Y146_SLICE_X5Y146_AO5),
.O6(CLBLL_L_X4Y146_SLICE_X5Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y147_SLICE_X4Y147_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y147_SLICE_X4Y147_AO6),
.Q(CLBLL_L_X4Y147_SLICE_X4Y147_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y147_SLICE_X4Y147_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y147_SLICE_X4Y147_BO6),
.Q(CLBLL_L_X4Y147_SLICE_X4Y147_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y147_SLICE_X4Y147_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y147_SLICE_X4Y147_CO6),
.Q(CLBLL_L_X4Y147_SLICE_X4Y147_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcacfcac0c5c0c5)
  ) CLBLL_L_X4Y147_SLICE_X4Y147_DLUT (
.I0(CLBLL_L_X4Y143_SLICE_X4Y143_BQ),
.I1(CLBLL_L_X4Y148_SLICE_X4Y148_CQ),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLM_L_X8Y148_SLICE_X10Y148_DO5),
.I4(1'b1),
.I5(CLBLM_R_X7Y144_SLICE_X9Y144_CQ),
.O5(CLBLL_L_X4Y147_SLICE_X4Y147_DO5),
.O6(CLBLL_L_X4Y147_SLICE_X4Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff05ff0a0005000a)
  ) CLBLL_L_X4Y147_SLICE_X4Y147_CLUT (
.I0(CLBLM_R_X7Y149_SLICE_X8Y149_AQ),
.I1(1'b1),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLL_L_X4Y147_SLICE_X4Y147_DO6),
.I5(CLBLM_R_X3Y147_SLICE_X3Y147_C5Q),
.O5(CLBLL_L_X4Y147_SLICE_X4Y147_CO5),
.O6(CLBLL_L_X4Y147_SLICE_X4Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0011114444)
  ) CLBLL_L_X4Y147_SLICE_X4Y147_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X8Y148_SLICE_X11Y148_BO6),
.I2(1'b1),
.I3(CLBLM_R_X3Y145_SLICE_X2Y145_BQ),
.I4(CLBLM_L_X8Y150_SLICE_X10Y150_BQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLL_L_X4Y147_SLICE_X4Y147_BO5),
.O6(CLBLL_L_X4Y147_SLICE_X4Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00fafaff00c8c8)
  ) CLBLL_L_X4Y147_SLICE_X4Y147_ALUT (
.I0(CLBLL_L_X4Y147_SLICE_X4Y147_DO6),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLL_L_X4Y147_SLICE_X4Y147_AQ),
.I3(CLBLM_R_X3Y148_SLICE_X2Y148_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.O5(CLBLL_L_X4Y147_SLICE_X4Y147_AO5),
.O6(CLBLL_L_X4Y147_SLICE_X4Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y147_SLICE_X5Y147_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y147_SLICE_X5Y147_BO5),
.Q(CLBLL_L_X4Y147_SLICE_X5Y147_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y147_SLICE_X5Y147_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y147_SLICE_X5Y147_AO6),
.Q(CLBLL_L_X4Y147_SLICE_X5Y147_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y147_SLICE_X5Y147_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y147_SLICE_X5Y147_BO6),
.Q(CLBLL_L_X4Y147_SLICE_X5Y147_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y147_SLICE_X5Y147_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y147_SLICE_X5Y147_CO6),
.Q(CLBLL_L_X4Y147_SLICE_X5Y147_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00006aaa0000aaaa)
  ) CLBLL_L_X4Y147_SLICE_X5Y147_DLUT (
.I0(CLBLL_L_X4Y147_SLICE_X5Y147_BQ),
.I1(CLBLM_L_X10Y147_SLICE_X12Y147_AQ),
.I2(CLBLL_L_X4Y146_SLICE_X4Y146_DO6),
.I3(CLBLM_R_X3Y146_SLICE_X3Y146_BQ),
.I4(CLBLM_R_X11Y146_SLICE_X14Y146_AQ),
.I5(CLBLM_R_X11Y147_SLICE_X14Y147_BQ),
.O5(CLBLL_L_X4Y147_SLICE_X5Y147_DO5),
.O6(CLBLL_L_X4Y147_SLICE_X5Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'heaaaaaaa40000000)
  ) CLBLL_L_X4Y147_SLICE_X5Y147_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y146_SLICE_X6Y146_A5Q),
.I2(CLBLM_R_X5Y153_SLICE_X6Y153_A5Q),
.I3(CLBLL_L_X4Y146_SLICE_X5Y146_CQ),
.I4(CLBLM_R_X7Y151_SLICE_X8Y151_A5Q),
.I5(CLBLM_L_X12Y146_SLICE_X16Y146_AQ),
.O5(CLBLL_L_X4Y147_SLICE_X5Y147_CO5),
.O6(CLBLL_L_X4Y147_SLICE_X5Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa0afa0affffc0c0)
  ) CLBLL_L_X4Y147_SLICE_X5Y147_BLUT (
.I0(CLBLL_L_X4Y147_SLICE_X5Y147_DO6),
.I1(CLBLM_R_X7Y143_SLICE_X9Y143_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y147_SLICE_X8Y147_AQ),
.I4(CLBLM_R_X7Y154_SLICE_X8Y154_DO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y147_SLICE_X5Y147_BO5),
.O6(CLBLL_L_X4Y147_SLICE_X5Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfe32fe32dc10dc10)
  ) CLBLL_L_X4Y147_SLICE_X5Y147_ALUT (
.I0(CLBLM_R_X5Y152_SLICE_X7Y152_DO5),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLL_L_X4Y147_SLICE_X5Y147_AQ),
.I3(CLBLM_L_X8Y146_SLICE_X10Y146_CQ),
.I4(1'b1),
.I5(CLBLM_R_X7Y146_SLICE_X9Y146_AQ),
.O5(CLBLL_L_X4Y147_SLICE_X5Y147_AO5),
.O6(CLBLL_L_X4Y147_SLICE_X5Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y148_SLICE_X4Y148_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y148_SLICE_X4Y148_CO5),
.Q(CLBLL_L_X4Y148_SLICE_X4Y148_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y148_SLICE_X4Y148_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y148_SLICE_X4Y148_AO6),
.Q(CLBLL_L_X4Y148_SLICE_X4Y148_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y148_SLICE_X4Y148_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y148_SLICE_X4Y148_BO6),
.Q(CLBLL_L_X4Y148_SLICE_X4Y148_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y148_SLICE_X4Y148_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y148_SLICE_X4Y148_CO6),
.Q(CLBLL_L_X4Y148_SLICE_X4Y148_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y148_SLICE_X4Y148_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y148_SLICE_X4Y148_DO6),
.Q(CLBLL_L_X4Y148_SLICE_X4Y148_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaff33aaaaf030)
  ) CLBLL_L_X4Y148_SLICE_X4Y148_DLUT (
.I0(CLBLM_R_X3Y146_SLICE_X3Y146_BQ),
.I1(CLBLM_L_X8Y148_SLICE_X10Y148_A5Q),
.I2(CLBLL_L_X4Y148_SLICE_X4Y148_DQ),
.I3(CLBLM_R_X11Y150_SLICE_X14Y150_BO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X10Y147_SLICE_X12Y147_AQ),
.O5(CLBLL_L_X4Y148_SLICE_X4Y148_DO5),
.O6(CLBLL_L_X4Y148_SLICE_X4Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc5500f0f0cccc)
  ) CLBLL_L_X4Y148_SLICE_X4Y148_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLL_L_X4Y144_SLICE_X4Y144_AQ),
.I2(CLBLM_R_X3Y149_SLICE_X3Y149_DQ),
.I3(CLBLM_R_X5Y148_SLICE_X7Y148_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y148_SLICE_X4Y148_CO5),
.O6(CLBLL_L_X4Y148_SLICE_X4Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccceeee00002222)
  ) CLBLL_L_X4Y148_SLICE_X4Y148_BLUT (
.I0(CLBLM_L_X10Y145_SLICE_X12Y145_CQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(1'b1),
.I3(1'b1),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X5Y149_SLICE_X6Y149_BQ),
.O5(CLBLL_L_X4Y148_SLICE_X4Y148_BO5),
.O6(CLBLL_L_X4Y148_SLICE_X4Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffcc00ccf0ccf0)
  ) CLBLL_L_X4Y148_SLICE_X4Y148_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y148_SLICE_X8Y148_D5Q),
.I2(CLBLL_L_X4Y148_SLICE_X4Y148_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X5Y148_SLICE_X6Y148_AQ),
.I5(CLBLM_R_X5Y152_SLICE_X7Y152_DO5),
.O5(CLBLL_L_X4Y148_SLICE_X4Y148_AO5),
.O6(CLBLL_L_X4Y148_SLICE_X4Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y148_SLICE_X5Y148_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y148_SLICE_X5Y148_AO6),
.Q(CLBLL_L_X4Y148_SLICE_X5Y148_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y148_SLICE_X5Y148_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y148_SLICE_X5Y148_BO6),
.Q(CLBLL_L_X4Y148_SLICE_X5Y148_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y148_SLICE_X5Y148_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y148_SLICE_X5Y148_CO6),
.Q(CLBLL_L_X4Y148_SLICE_X5Y148_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff7fffffffffffff)
  ) CLBLL_L_X4Y148_SLICE_X5Y148_DLUT (
.I0(CLBLM_R_X3Y146_SLICE_X3Y146_BQ),
.I1(CLBLL_L_X4Y145_SLICE_X4Y145_CQ),
.I2(CLBLM_R_X7Y145_SLICE_X8Y145_AQ),
.I3(CLBLM_R_X5Y145_SLICE_X7Y145_AQ),
.I4(CLBLM_R_X7Y147_SLICE_X8Y147_AQ),
.I5(CLBLM_L_X10Y147_SLICE_X12Y147_AQ),
.O5(CLBLL_L_X4Y148_SLICE_X5Y148_DO5),
.O6(CLBLL_L_X4Y148_SLICE_X5Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa00000f0f)
  ) CLBLL_L_X4Y148_SLICE_X5Y148_CLUT (
.I0(CLBLL_L_X2Y148_SLICE_X1Y148_AQ),
.I1(1'b1),
.I2(CLBLL_L_X4Y146_SLICE_X5Y146_DO6),
.I3(1'b1),
.I4(CLBLL_L_X4Y148_SLICE_X5Y148_DO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLL_L_X4Y148_SLICE_X5Y148_CO5),
.O6(CLBLL_L_X4Y148_SLICE_X5Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaafffcaaaa000c)
  ) CLBLL_L_X4Y148_SLICE_X5Y148_BLUT (
.I0(CLBLM_R_X3Y148_SLICE_X3Y148_CQ),
.I1(CLBLL_L_X4Y148_SLICE_X5Y148_BQ),
.I2(RIOB33_X105Y117_IOB_X1Y118_I),
.I3(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y144_SLICE_X8Y144_CQ),
.O5(CLBLL_L_X4Y148_SLICE_X5Y148_BO5),
.O6(CLBLL_L_X4Y148_SLICE_X5Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000e2aae2aa)
  ) CLBLL_L_X4Y148_SLICE_X5Y148_ALUT (
.I0(CLBLM_L_X10Y147_SLICE_X12Y147_AQ),
.I1(CLBLM_L_X8Y149_SLICE_X11Y149_AQ),
.I2(CLBLL_L_X4Y148_SLICE_X5Y148_AQ),
.I3(CLBLL_L_X4Y151_SLICE_X4Y151_AQ),
.I4(CLBLL_L_X4Y147_SLICE_X4Y147_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLL_L_X4Y148_SLICE_X5Y148_AO5),
.O6(CLBLL_L_X4Y148_SLICE_X5Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y149_SLICE_X4Y149_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y149_SLICE_X4Y149_AO6),
.Q(CLBLL_L_X4Y149_SLICE_X4Y149_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y149_SLICE_X4Y149_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y149_SLICE_X4Y149_BO6),
.Q(CLBLL_L_X4Y149_SLICE_X4Y149_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y149_SLICE_X4Y149_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y149_SLICE_X4Y149_CO6),
.Q(CLBLL_L_X4Y149_SLICE_X4Y149_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y149_SLICE_X4Y149_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y149_SLICE_X4Y149_DO6),
.Q(CLBLL_L_X4Y149_SLICE_X4Y149_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hd8d8d8d888d888d8)
  ) CLBLL_L_X4Y149_SLICE_X4Y149_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X3Y148_SLICE_X3Y148_B5Q),
.I2(CLBLL_L_X4Y149_SLICE_X4Y149_DQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(1'b1),
.I5(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.O5(CLBLL_L_X4Y149_SLICE_X4Y149_DO5),
.O6(CLBLL_L_X4Y149_SLICE_X4Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55ff4400550044)
  ) CLBLL_L_X4Y149_SLICE_X4Y149_CLUT (
.I0(CLBLM_R_X5Y152_SLICE_X7Y152_DO5),
.I1(CLBLL_L_X4Y149_SLICE_X4Y149_CQ),
.I2(1'b1),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X5Y151_SLICE_X6Y151_CQ),
.I5(CLBLL_L_X4Y149_SLICE_X5Y149_A5Q),
.O5(CLBLL_L_X4Y149_SLICE_X4Y149_CO5),
.O6(CLBLL_L_X4Y149_SLICE_X4Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hafafacaca0a0a0a0)
  ) CLBLL_L_X4Y149_SLICE_X4Y149_BLUT (
.I0(CLBLM_R_X3Y145_SLICE_X3Y145_AQ),
.I1(CLBLL_L_X4Y149_SLICE_X4Y149_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(CLBLM_R_X7Y150_SLICE_X8Y150_CQ),
.I5(CLBLM_L_X8Y152_SLICE_X11Y152_BO6),
.O5(CLBLL_L_X4Y149_SLICE_X4Y149_BO5),
.O6(CLBLL_L_X4Y149_SLICE_X4Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbff1155bafa1050)
  ) CLBLL_L_X4Y149_SLICE_X4Y149_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y148_SLICE_X10Y148_A5Q),
.I2(CLBLL_L_X4Y149_SLICE_X4Y149_AQ),
.I3(CLBLM_R_X11Y150_SLICE_X14Y150_AO6),
.I4(CLBLM_R_X5Y144_SLICE_X7Y144_BQ),
.I5(CLBLM_R_X3Y146_SLICE_X3Y146_BQ),
.O5(CLBLL_L_X4Y149_SLICE_X4Y149_AO5),
.O6(CLBLL_L_X4Y149_SLICE_X4Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y149_SLICE_X5Y149_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y149_SLICE_X5Y149_BO6),
.Q(CLBLL_L_X4Y149_SLICE_X5Y149_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y149_SLICE_X5Y149_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y149_SLICE_X5Y149_AO6),
.Q(CLBLL_L_X4Y149_SLICE_X5Y149_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y149_SLICE_X5Y149_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y149_SLICE_X5Y149_CO6),
.Q(CLBLL_L_X4Y149_SLICE_X5Y149_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y149_SLICE_X5Y149_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y149_SLICE_X5Y149_DO6),
.Q(CLBLL_L_X4Y149_SLICE_X5Y149_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcc3300fedc3210)
  ) CLBLL_L_X4Y149_SLICE_X5Y149_DLUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLL_L_X4Y149_SLICE_X5Y149_DQ),
.I3(CLBLM_R_X7Y149_SLICE_X9Y149_BO6),
.I4(CLBLM_R_X3Y149_SLICE_X3Y149_CQ),
.I5(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.O5(CLBLL_L_X4Y149_SLICE_X5Y149_DO5),
.O6(CLBLL_L_X4Y149_SLICE_X5Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f000f0f0c000c)
  ) CLBLL_L_X4Y149_SLICE_X5Y149_CLUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y149_SLICE_X5Y149_CQ),
.I2(CLBLM_R_X5Y152_SLICE_X7Y152_DO6),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLL_L_X4Y149_SLICE_X5Y149_AQ),
.I5(CLBLM_L_X8Y150_SLICE_X10Y150_BQ),
.O5(CLBLL_L_X4Y149_SLICE_X5Y149_CO5),
.O6(CLBLL_L_X4Y149_SLICE_X5Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f404cccc0000)
  ) CLBLL_L_X4Y149_SLICE_X5Y149_BLUT (
.I0(CLBLM_R_X5Y149_SLICE_X7Y149_DO6),
.I1(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLL_L_X4Y147_SLICE_X4Y147_CQ),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y149_SLICE_X5Y149_BO5),
.O6(CLBLL_L_X4Y149_SLICE_X5Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff005050ff00d8d8)
  ) CLBLL_L_X4Y149_SLICE_X5Y149_ALUT (
.I0(CLBLL_L_X4Y149_SLICE_X5Y149_BO5),
.I1(CLBLM_R_X3Y150_SLICE_X2Y150_BO6),
.I2(CLBLL_L_X4Y149_SLICE_X5Y149_AQ),
.I3(CLBLL_L_X4Y147_SLICE_X5Y147_B5Q),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLL_L_X4Y149_SLICE_X5Y149_AO5),
.O6(CLBLL_L_X4Y149_SLICE_X5Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y150_SLICE_X4Y150_B5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y150_SLICE_X4Y150_BO5),
.Q(CLBLL_L_X4Y150_SLICE_X4Y150_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y150_SLICE_X4Y150_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y150_SLICE_X4Y150_AO6),
.Q(CLBLL_L_X4Y150_SLICE_X4Y150_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y150_SLICE_X4Y150_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y150_SLICE_X4Y150_BO6),
.Q(CLBLL_L_X4Y150_SLICE_X4Y150_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7350ffff73507350)
  ) CLBLL_L_X4Y150_SLICE_X4Y150_DLUT (
.I0(CLBLL_L_X4Y155_SLICE_X5Y155_AO6),
.I1(CLBLL_L_X4Y152_SLICE_X4Y152_AO5),
.I2(CLBLM_R_X5Y149_SLICE_X6Y149_BQ),
.I3(RIOB33_X105Y115_IOB_X1Y116_I),
.I4(CLBLL_L_X4Y152_SLICE_X4Y152_AO6),
.I5(CLBLM_L_X8Y151_SLICE_X10Y151_CQ),
.O5(CLBLL_L_X4Y150_SLICE_X4Y150_DO5),
.O6(CLBLL_L_X4Y150_SLICE_X4Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h30ff3030baffbaba)
  ) CLBLL_L_X4Y150_SLICE_X4Y150_CLUT (
.I0(CLBLL_L_X4Y146_SLICE_X4Y146_AQ),
.I1(CLBLL_L_X4Y152_SLICE_X5Y152_AO5),
.I2(CLBLM_R_X5Y149_SLICE_X6Y149_AQ),
.I3(CLBLL_L_X4Y152_SLICE_X5Y152_AO6),
.I4(CLBLM_L_X8Y147_SLICE_X10Y147_BQ),
.I5(CLBLL_L_X2Y152_SLICE_X1Y152_BO6),
.O5(CLBLL_L_X4Y150_SLICE_X4Y150_CO5),
.O6(CLBLL_L_X4Y150_SLICE_X4Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcc3300e2e2e2e2)
  ) CLBLL_L_X4Y150_SLICE_X4Y150_BLUT (
.I0(CLBLM_R_X11Y150_SLICE_X14Y150_AO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X11Y149_SLICE_X14Y149_BQ),
.I3(CLBLL_L_X2Y153_SLICE_X1Y153_DO6),
.I4(CLBLM_R_X3Y147_SLICE_X2Y147_A5Q),
.I5(1'b1),
.O5(CLBLL_L_X4Y150_SLICE_X4Y150_BO5),
.O6(CLBLL_L_X4Y150_SLICE_X4Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccf000f0f0)
  ) CLBLL_L_X4Y150_SLICE_X4Y150_ALUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y150_SLICE_X4Y150_BQ),
.I2(CLBLL_L_X4Y150_SLICE_X4Y150_AQ),
.I3(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLL_L_X4Y150_SLICE_X4Y150_AO5),
.O6(CLBLL_L_X4Y150_SLICE_X4Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y150_SLICE_X5Y150_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y150_SLICE_X5Y150_AO6),
.Q(CLBLL_L_X4Y150_SLICE_X5Y150_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y150_SLICE_X5Y150_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y150_SLICE_X5Y150_BO6),
.Q(CLBLL_L_X4Y150_SLICE_X5Y150_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333f3f30000f0f0)
  ) CLBLL_L_X4Y150_SLICE_X5Y150_DLUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y152_SLICE_X5Y152_AO5),
.I2(CLBLL_L_X4Y149_SLICE_X5Y149_AQ),
.I3(1'b1),
.I4(CLBLL_L_X2Y154_SLICE_X1Y154_AO5),
.I5(CLBLM_R_X5Y148_SLICE_X7Y148_AQ),
.O5(CLBLL_L_X4Y150_SLICE_X5Y150_DO5),
.O6(CLBLL_L_X4Y150_SLICE_X5Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8800000088000000)
  ) CLBLL_L_X4Y150_SLICE_X5Y150_CLUT (
.I0(CLBLM_R_X5Y150_SLICE_X7Y150_BQ),
.I1(CLBLL_L_X4Y147_SLICE_X4Y147_BQ),
.I2(1'b1),
.I3(CLBLM_R_X5Y152_SLICE_X6Y152_A5Q),
.I4(CLBLM_R_X7Y149_SLICE_X8Y149_DQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y150_SLICE_X5Y150_CO5),
.O6(CLBLL_L_X4Y150_SLICE_X5Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0ffcc00cc)
  ) CLBLL_L_X4Y150_SLICE_X5Y150_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y145_SLICE_X7Y145_CQ),
.I2(CLBLL_L_X4Y148_SLICE_X4Y148_DQ),
.I3(CLBLM_R_X5Y152_SLICE_X7Y152_DO5),
.I4(CLBLL_L_X4Y150_SLICE_X5Y150_BQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLL_L_X4Y150_SLICE_X5Y150_BO5),
.O6(CLBLL_L_X4Y150_SLICE_X5Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000fc30fc30)
  ) CLBLL_L_X4Y150_SLICE_X5Y150_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y152_SLICE_X7Y152_DO5),
.I2(CLBLL_L_X4Y150_SLICE_X5Y150_AQ),
.I3(CLBLM_R_X5Y147_SLICE_X6Y147_CQ),
.I4(CLBLM_R_X7Y150_SLICE_X8Y150_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLL_L_X4Y150_SLICE_X5Y150_AO5),
.O6(CLBLL_L_X4Y150_SLICE_X5Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y151_SLICE_X4Y151_A5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y151_SLICE_X9Y151_DO6),
.Q(CLBLL_L_X4Y151_SLICE_X4Y151_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y151_SLICE_X4Y151_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y151_SLICE_X4Y151_AO6),
.Q(CLBLL_L_X4Y151_SLICE_X4Y151_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000303033003330)
  ) CLBLL_L_X4Y151_SLICE_X4Y151_DLUT (
.I0(1'b1),
.I1(CLBLL_L_X2Y155_SLICE_X1Y155_DO6),
.I2(CLBLM_R_X5Y151_SLICE_X6Y151_AQ),
.I3(CLBLM_R_X5Y151_SLICE_X7Y151_BQ),
.I4(CLBLL_L_X2Y154_SLICE_X1Y154_BO5),
.I5(CLBLL_L_X4Y155_SLICE_X4Y155_BO6),
.O5(CLBLL_L_X4Y151_SLICE_X4Y151_DO5),
.O6(CLBLL_L_X4Y151_SLICE_X4Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000008)
  ) CLBLL_L_X4Y151_SLICE_X4Y151_CLUT (
.I0(RIOB33_X105Y131_IOB_X1Y132_I),
.I1(CLBLM_R_X5Y152_SLICE_X6Y152_CQ),
.I2(CLBLL_L_X2Y155_SLICE_X1Y155_DO6),
.I3(RIOB33_X105Y133_IOB_X1Y133_I),
.I4(RIOB33_X105Y133_IOB_X1Y134_I),
.I5(RIOB33_X105Y131_IOB_X1Y131_I),
.O5(CLBLL_L_X4Y151_SLICE_X4Y151_CO5),
.O6(CLBLL_L_X4Y151_SLICE_X4Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffefffefe)
  ) CLBLL_L_X4Y151_SLICE_X4Y151_BLUT (
.I0(CLBLL_L_X2Y151_SLICE_X1Y151_DO6),
.I1(CLBLL_L_X4Y151_SLICE_X5Y151_DO6),
.I2(CLBLL_L_X2Y149_SLICE_X0Y149_AO6),
.I3(CLBLL_L_X2Y154_SLICE_X1Y154_AO5),
.I4(CLBLM_R_X5Y146_SLICE_X6Y146_AQ),
.I5(CLBLL_L_X4Y151_SLICE_X4Y151_CO6),
.O5(CLBLL_L_X4Y151_SLICE_X4Y151_BO5),
.O6(CLBLL_L_X4Y151_SLICE_X4Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0c0c0cfcf)
  ) CLBLL_L_X4Y151_SLICE_X4Y151_ALUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y151_SLICE_X5Y151_B5Q),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(CLBLM_L_X8Y149_SLICE_X11Y149_AQ),
.I5(CLBLM_R_X3Y150_SLICE_X3Y150_A5Q),
.O5(CLBLL_L_X4Y151_SLICE_X4Y151_AO5),
.O6(CLBLL_L_X4Y151_SLICE_X4Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y151_SLICE_X5Y151_B5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y151_SLICE_X5Y151_BO5),
.Q(CLBLL_L_X4Y151_SLICE_X5Y151_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y151_SLICE_X5Y151_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y151_SLICE_X5Y151_AO6),
.Q(CLBLL_L_X4Y151_SLICE_X5Y151_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y151_SLICE_X5Y151_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y151_SLICE_X5Y151_BO6),
.Q(CLBLL_L_X4Y151_SLICE_X5Y151_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000400)
  ) CLBLL_L_X4Y151_SLICE_X5Y151_DLUT (
.I0(RIOB33_X105Y131_IOB_X1Y132_I),
.I1(CLBLM_L_X8Y152_SLICE_X10Y152_BQ),
.I2(RIOB33_X105Y133_IOB_X1Y134_I),
.I3(RIOB33_X105Y133_IOB_X1Y133_I),
.I4(CLBLL_L_X2Y155_SLICE_X1Y155_DO6),
.I5(RIOB33_X105Y131_IOB_X1Y131_I),
.O5(CLBLL_L_X4Y151_SLICE_X5Y151_DO5),
.O6(CLBLL_L_X4Y151_SLICE_X5Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h55ddf5fd00ccf0fc)
  ) CLBLL_L_X4Y151_SLICE_X5Y151_CLUT (
.I0(CLBLL_L_X4Y152_SLICE_X5Y152_AO6),
.I1(CLBLM_R_X7Y151_SLICE_X9Y151_BQ),
.I2(CLBLM_R_X5Y151_SLICE_X7Y151_AQ),
.I3(CLBLL_L_X2Y152_SLICE_X1Y152_BO6),
.I4(CLBLL_L_X2Y154_SLICE_X1Y154_AO5),
.I5(CLBLM_R_X7Y150_SLICE_X8Y150_BQ),
.O5(CLBLL_L_X4Y151_SLICE_X5Y151_CO5),
.O6(CLBLL_L_X4Y151_SLICE_X5Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0aaf0aaffcc00cc)
  ) CLBLL_L_X4Y151_SLICE_X5Y151_BLUT (
.I0(CLBLM_R_X3Y153_SLICE_X2Y153_DO6),
.I1(CLBLM_R_X3Y154_SLICE_X2Y154_BO6),
.I2(CLBLM_L_X8Y144_SLICE_X10Y144_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLL_L_X4Y148_SLICE_X5Y148_CQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y151_SLICE_X5Y151_BO5),
.O6(CLBLL_L_X4Y151_SLICE_X5Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffbb00bbffb000b0)
  ) CLBLL_L_X4Y151_SLICE_X5Y151_ALUT (
.I0(CLBLM_R_X11Y150_SLICE_X14Y150_BO6),
.I1(CLBLM_L_X8Y148_SLICE_X10Y148_A5Q),
.I2(CLBLL_L_X4Y151_SLICE_X5Y151_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y150_SLICE_X8Y150_BQ),
.I5(CLBLM_R_X7Y147_SLICE_X8Y147_AQ),
.O5(CLBLL_L_X4Y151_SLICE_X5Y151_AO5),
.O6(CLBLL_L_X4Y151_SLICE_X5Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h30303030ffff3030)
  ) CLBLL_L_X4Y152_SLICE_X4Y152_DLUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y152_SLICE_X5Y152_AO5),
.I2(CLBLM_L_X10Y152_SLICE_X12Y152_D5Q),
.I3(1'b1),
.I4(CLBLM_R_X3Y146_SLICE_X3Y146_AQ),
.I5(CLBLL_L_X2Y152_SLICE_X1Y152_BO6),
.O5(CLBLL_L_X4Y152_SLICE_X4Y152_DO5),
.O6(CLBLL_L_X4Y152_SLICE_X4Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000004444ff44)
  ) CLBLL_L_X4Y152_SLICE_X4Y152_CLUT (
.I0(CLBLL_L_X2Y151_SLICE_X0Y151_CO5),
.I1(CLBLL_L_X4Y149_SLICE_X5Y149_CQ),
.I2(1'b1),
.I3(CLBLL_L_X4Y153_SLICE_X5Y153_AQ),
.I4(CLBLL_L_X2Y154_SLICE_X1Y154_BO5),
.I5(CLBLL_L_X2Y155_SLICE_X1Y155_DO6),
.O5(CLBLL_L_X4Y152_SLICE_X4Y152_CO5),
.O6(CLBLL_L_X4Y152_SLICE_X4Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h000c555d000c000c)
  ) CLBLL_L_X4Y152_SLICE_X4Y152_BLUT (
.I0(CLBLL_L_X2Y151_SLICE_X1Y151_AO6),
.I1(CLBLM_R_X5Y147_SLICE_X7Y147_BQ),
.I2(CLBLL_L_X2Y151_SLICE_X0Y151_CO5),
.I3(CLBLL_L_X2Y155_SLICE_X1Y155_DO6),
.I4(CLBLL_L_X2Y152_SLICE_X1Y152_AO6),
.I5(RIOB33_X105Y117_IOB_X1Y117_I),
.O5(CLBLL_L_X4Y152_SLICE_X4Y152_BO5),
.O6(CLBLL_L_X4Y152_SLICE_X4Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffefffffffffdff)
  ) CLBLL_L_X4Y152_SLICE_X4Y152_ALUT (
.I0(RIOB33_X105Y133_IOB_X1Y133_I),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(CLBLL_L_X2Y152_SLICE_X1Y152_AO6),
.I3(RIOB33_X105Y131_IOB_X1Y132_I),
.I4(RIOB33_X105Y133_IOB_X1Y134_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y152_SLICE_X4Y152_AO5),
.O6(CLBLL_L_X4Y152_SLICE_X4Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000040)
  ) CLBLL_L_X4Y152_SLICE_X5Y152_DLUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(CLBLM_L_X8Y150_SLICE_X11Y150_BQ),
.I2(RIOB33_X105Y133_IOB_X1Y133_I),
.I3(RIOB33_X105Y133_IOB_X1Y134_I),
.I4(RIOB33_X105Y131_IOB_X1Y132_I),
.I5(CLBLL_L_X2Y155_SLICE_X1Y155_DO6),
.O5(CLBLL_L_X4Y152_SLICE_X5Y152_DO5),
.O6(CLBLL_L_X4Y152_SLICE_X5Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000004000000000)
  ) CLBLL_L_X4Y152_SLICE_X5Y152_CLUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(RIOB33_X105Y133_IOB_X1Y133_I),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(RIOB33_X105Y133_IOB_X1Y134_I),
.I4(CLBLL_L_X2Y155_SLICE_X1Y155_DO6),
.I5(CLBLL_L_X4Y147_SLICE_X5Y147_AQ),
.O5(CLBLL_L_X4Y152_SLICE_X5Y152_CO5),
.O6(CLBLL_L_X4Y152_SLICE_X5Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000270500002200)
  ) CLBLL_L_X4Y152_SLICE_X5Y152_BLUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(CLBLL_L_X2Y155_SLICE_X1Y155_DO6),
.I2(CLBLL_L_X2Y152_SLICE_X1Y152_AO6),
.I3(CLBLM_R_X5Y152_SLICE_X7Y152_AQ),
.I4(CLBLL_L_X4Y154_SLICE_X5Y154_CO5),
.I5(CLBLM_R_X5Y150_SLICE_X6Y150_BQ),
.O5(CLBLL_L_X4Y152_SLICE_X5Y152_BO5),
.O6(CLBLL_L_X4Y152_SLICE_X5Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffeffffffffbffff)
  ) CLBLL_L_X4Y152_SLICE_X5Y152_ALUT (
.I0(RIOB33_X105Y133_IOB_X1Y134_I),
.I1(RIOB33_X105Y131_IOB_X1Y132_I),
.I2(RIOB33_X105Y133_IOB_X1Y133_I),
.I3(CLBLL_L_X2Y155_SLICE_X1Y155_DO6),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y152_SLICE_X5Y152_AO5),
.O6(CLBLL_L_X4Y152_SLICE_X5Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h44ff4444f4fff4f4)
  ) CLBLL_L_X4Y153_SLICE_X4Y153_DLUT (
.I0(CLBLL_L_X4Y155_SLICE_X5Y155_AO6),
.I1(CLBLM_R_X5Y153_SLICE_X6Y153_BQ),
.I2(CLBLL_L_X4Y154_SLICE_X5Y154_AQ),
.I3(CLBLL_L_X4Y152_SLICE_X4Y152_AO6),
.I4(CLBLL_L_X4Y148_SLICE_X4Y148_DQ),
.I5(CLBLM_R_X3Y152_SLICE_X2Y152_AO5),
.O5(CLBLL_L_X4Y153_SLICE_X4Y153_DO5),
.O6(CLBLL_L_X4Y153_SLICE_X4Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haabaffff00300030)
  ) CLBLL_L_X4Y153_SLICE_X4Y153_CLUT (
.I0(RIOB33_X105Y129_IOB_X1Y129_I),
.I1(CLBLL_L_X2Y152_SLICE_X1Y152_AO5),
.I2(CLBLM_R_X5Y153_SLICE_X7Y153_BQ),
.I3(CLBLL_L_X4Y155_SLICE_X4Y155_BO6),
.I4(RIOB33_X105Y137_IOB_X1Y137_I),
.I5(CLBLL_L_X4Y150_SLICE_X4Y150_BQ),
.O5(CLBLL_L_X4Y153_SLICE_X4Y153_CO5),
.O6(CLBLL_L_X4Y153_SLICE_X4Y153_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0005000400000004)
  ) CLBLL_L_X4Y153_SLICE_X4Y153_BLUT (
.I0(CLBLM_R_X3Y155_SLICE_X3Y155_DO6),
.I1(CLBLL_L_X4Y149_SLICE_X4Y149_BQ),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(CLBLL_L_X2Y155_SLICE_X1Y155_DO6),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(CLBLM_L_X8Y152_SLICE_X10Y152_AQ),
.O5(CLBLL_L_X4Y153_SLICE_X4Y153_BO5),
.O6(CLBLL_L_X4Y153_SLICE_X4Y153_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h000a000a000accce)
  ) CLBLL_L_X4Y153_SLICE_X4Y153_ALUT (
.I0(CLBLL_L_X4Y148_SLICE_X4Y148_DQ),
.I1(CLBLM_R_X5Y153_SLICE_X6Y153_BQ),
.I2(CLBLL_L_X2Y151_SLICE_X0Y151_CO5),
.I3(CLBLL_L_X2Y152_SLICE_X1Y152_AO6),
.I4(CLBLL_L_X2Y154_SLICE_X1Y154_BO5),
.I5(CLBLL_L_X2Y155_SLICE_X1Y155_DO6),
.O5(CLBLL_L_X4Y153_SLICE_X4Y153_AO5),
.O6(CLBLL_L_X4Y153_SLICE_X4Y153_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y153_SLICE_X5Y153_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y153_SLICE_X5Y153_AO6),
.Q(CLBLL_L_X4Y153_SLICE_X5Y153_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h4444ff44f4f4fff4)
  ) CLBLL_L_X4Y153_SLICE_X5Y153_DLUT (
.I0(CLBLL_L_X4Y152_SLICE_X5Y152_AO6),
.I1(CLBLM_L_X8Y152_SLICE_X10Y152_AQ),
.I2(CLBLL_L_X4Y146_SLICE_X5Y146_AQ),
.I3(CLBLL_L_X4Y149_SLICE_X4Y149_BQ),
.I4(CLBLM_R_X5Y154_SLICE_X7Y154_AO6),
.I5(CLBLL_L_X2Y152_SLICE_X1Y152_BO6),
.O5(CLBLL_L_X4Y153_SLICE_X5Y153_DO5),
.O6(CLBLL_L_X4Y153_SLICE_X5Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffff4f44)
  ) CLBLL_L_X4Y153_SLICE_X5Y153_CLUT (
.I0(CLBLL_L_X4Y152_SLICE_X5Y152_AO6),
.I1(CLBLM_R_X5Y153_SLICE_X6Y153_AQ),
.I2(CLBLL_L_X2Y154_SLICE_X1Y154_AO5),
.I3(CLBLM_R_X7Y151_SLICE_X9Y151_AQ),
.I4(CLBLL_L_X4Y152_SLICE_X5Y152_DO6),
.I5(CLBLL_L_X4Y153_SLICE_X5Y153_BO6),
.O5(CLBLL_L_X4Y153_SLICE_X5Y153_CO5),
.O6(CLBLL_L_X4Y153_SLICE_X5Y153_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000040)
  ) CLBLL_L_X4Y153_SLICE_X5Y153_BLUT (
.I0(RIOB33_X105Y133_IOB_X1Y134_I),
.I1(CLBLM_R_X5Y153_SLICE_X7Y153_AQ),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(CLBLL_L_X2Y155_SLICE_X1Y155_DO6),
.I4(RIOB33_X105Y133_IOB_X1Y133_I),
.I5(RIOB33_X105Y131_IOB_X1Y131_I),
.O5(CLBLL_L_X4Y153_SLICE_X5Y153_BO5),
.O6(CLBLL_L_X4Y153_SLICE_X5Y153_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccf0ccaaccf0ccaa)
  ) CLBLL_L_X4Y153_SLICE_X5Y153_ALUT (
.I0(CLBLL_L_X4Y153_SLICE_X5Y153_AQ),
.I1(CLBLM_R_X5Y153_SLICE_X6Y153_AQ),
.I2(CLBLM_R_X5Y151_SLICE_X6Y151_BQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X5Y152_SLICE_X7Y152_DO5),
.I5(1'b1),
.O5(CLBLL_L_X4Y153_SLICE_X5Y153_AO5),
.O6(CLBLL_L_X4Y153_SLICE_X5Y153_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff2fff2fff22ff22)
  ) CLBLL_L_X4Y154_SLICE_X4Y154_DLUT (
.I0(CLBLL_L_X4Y150_SLICE_X5Y150_AQ),
.I1(CLBLL_L_X4Y155_SLICE_X5Y155_AO5),
.I2(CLBLL_L_X2Y152_SLICE_X1Y152_BO5),
.I3(CLBLL_L_X4Y152_SLICE_X4Y152_BO6),
.I4(1'b1),
.I5(CLBLM_R_X3Y148_SLICE_X3Y148_B5Q),
.O5(CLBLL_L_X4Y154_SLICE_X4Y154_DO5),
.O6(CLBLL_L_X4Y154_SLICE_X4Y154_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffefe)
  ) CLBLL_L_X4Y154_SLICE_X4Y154_CLUT (
.I0(CLBLL_L_X2Y150_SLICE_X1Y150_CO6),
.I1(CLBLM_R_X5Y154_SLICE_X7Y154_DO6),
.I2(CLBLL_L_X4Y153_SLICE_X4Y153_DO6),
.I3(1'b1),
.I4(CLBLL_L_X4Y154_SLICE_X4Y154_DO6),
.I5(CLBLM_R_X3Y155_SLICE_X2Y155_DO6),
.O5(CLBLL_L_X4Y154_SLICE_X4Y154_CO5),
.O6(CLBLL_L_X4Y154_SLICE_X4Y154_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffcfffcfc)
  ) CLBLL_L_X4Y154_SLICE_X4Y154_BLUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y152_SLICE_X4Y152_BO6),
.I2(CLBLL_L_X4Y153_SLICE_X4Y153_AO6),
.I3(CLBLM_R_X3Y152_SLICE_X2Y152_AO5),
.I4(CLBLL_L_X4Y154_SLICE_X5Y154_AQ),
.I5(CLBLL_L_X4Y154_SLICE_X4Y154_AO6),
.O5(CLBLL_L_X4Y154_SLICE_X4Y154_BO5),
.O6(CLBLL_L_X4Y154_SLICE_X4Y154_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0537003305050000)
  ) CLBLL_L_X4Y154_SLICE_X4Y154_ALUT (
.I0(CLBLL_L_X2Y155_SLICE_X1Y155_DO6),
.I1(CLBLL_L_X4Y155_SLICE_X4Y155_BO6),
.I2(CLBLL_L_X2Y151_SLICE_X1Y151_AO6),
.I3(CLBLL_L_X2Y152_SLICE_X1Y152_AO6),
.I4(CLBLL_L_X4Y150_SLICE_X5Y150_AQ),
.I5(CLBLM_R_X3Y148_SLICE_X3Y148_B5Q),
.O5(CLBLL_L_X4Y154_SLICE_X4Y154_AO5),
.O6(CLBLL_L_X4Y154_SLICE_X4Y154_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y154_SLICE_X5Y154_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y154_SLICE_X5Y154_AO6),
.Q(CLBLL_L_X4Y154_SLICE_X5Y154_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y154_SLICE_X5Y154_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y154_SLICE_X5Y154_BO6),
.Q(CLBLL_L_X4Y154_SLICE_X5Y154_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000040000000)
  ) CLBLL_L_X4Y154_SLICE_X5Y154_DLUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(RIOB33_X105Y133_IOB_X1Y133_I),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(RIOB33_X105Y133_IOB_X1Y134_I),
.I4(CLBLL_L_X4Y146_SLICE_X5Y146_AQ),
.I5(CLBLL_L_X2Y152_SLICE_X1Y152_AO6),
.O5(CLBLL_L_X4Y154_SLICE_X5Y154_DO5),
.O6(CLBLL_L_X4Y154_SLICE_X5Y154_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffff3cfffcfffcf)
  ) CLBLL_L_X4Y154_SLICE_X5Y154_CLUT (
.I0(1'b1),
.I1(RIOB33_X105Y131_IOB_X1Y132_I),
.I2(RIOB33_X105Y133_IOB_X1Y134_I),
.I3(RIOB33_X105Y133_IOB_X1Y133_I),
.I4(CLBLL_L_X2Y155_SLICE_X1Y155_DO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y154_SLICE_X5Y154_CO5),
.O6(CLBLL_L_X4Y154_SLICE_X5Y154_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ccccff008888)
  ) CLBLL_L_X4Y154_SLICE_X5Y154_BLUT (
.I0(CLBLL_L_X4Y154_SLICE_X5Y154_BQ),
.I1(CLBLM_R_X3Y144_SLICE_X2Y144_CO6),
.I2(1'b1),
.I3(CLBLL_L_X4Y147_SLICE_X5Y147_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y145_SLICE_X8Y145_C5Q),
.O5(CLBLL_L_X4Y154_SLICE_X5Y154_BO5),
.O6(CLBLL_L_X4Y154_SLICE_X5Y154_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffcc00ccf0ccf0)
  ) CLBLL_L_X4Y154_SLICE_X5Y154_ALUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y153_SLICE_X5Y153_AQ),
.I2(CLBLL_L_X4Y154_SLICE_X5Y154_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X5Y150_SLICE_X7Y150_BQ),
.I5(CLBLM_R_X5Y152_SLICE_X7Y152_DO5),
.O5(CLBLL_L_X4Y154_SLICE_X5Y154_AO5),
.O6(CLBLL_L_X4Y154_SLICE_X5Y154_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f30000f3fb00aa)
  ) CLBLL_L_X4Y155_SLICE_X4Y155_DLUT (
.I0(CLBLL_L_X4Y154_SLICE_X5Y154_BQ),
.I1(RIOB33_X105Y137_IOB_X1Y137_I),
.I2(RIOB33_X105Y129_IOB_X1Y129_I),
.I3(CLBLL_L_X2Y152_SLICE_X1Y152_AO5),
.I4(CLBLL_L_X4Y151_SLICE_X5Y151_B5Q),
.I5(CLBLL_L_X4Y155_SLICE_X4Y155_BO6),
.O5(CLBLL_L_X4Y155_SLICE_X4Y155_DO5),
.O6(CLBLL_L_X4Y155_SLICE_X4Y155_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000cffff00ae)
  ) CLBLL_L_X4Y155_SLICE_X4Y155_CLUT (
.I0(CLBLL_L_X4Y154_SLICE_X5Y154_BQ),
.I1(LIOB33_X0Y67_IOB_X0Y68_I),
.I2(CLBLL_L_X2Y154_SLICE_X1Y154_BO5),
.I3(CLBLL_L_X2Y152_SLICE_X1Y152_AO5),
.I4(CLBLL_L_X4Y155_SLICE_X4Y155_AO6),
.I5(CLBLL_L_X4Y155_SLICE_X4Y155_BO6),
.O5(CLBLL_L_X4Y155_SLICE_X4Y155_CO5),
.O6(CLBLL_L_X4Y155_SLICE_X4Y155_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfaffffff20200000)
  ) CLBLL_L_X4Y155_SLICE_X4Y155_BLUT (
.I0(RIOB33_X105Y131_IOB_X1Y132_I),
.I1(CLBLL_L_X2Y152_SLICE_X1Y152_AO6),
.I2(RIOB33_X105Y133_IOB_X1Y133_I),
.I3(RIOB33_X105Y133_IOB_X1Y134_I),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y155_SLICE_X4Y155_BO5),
.O6(CLBLL_L_X4Y155_SLICE_X4Y155_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0aaa0aafcfffcff)
  ) CLBLL_L_X4Y155_SLICE_X4Y155_ALUT (
.I0(CLBLL_L_X4Y151_SLICE_X5Y151_B5Q),
.I1(RIOB33_X105Y129_IOB_X1Y130_I),
.I2(RIOB33_X105Y129_IOB_X1Y129_I),
.I3(RIOB33_X105Y137_IOB_X1Y137_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y155_SLICE_X4Y155_AO5),
.O6(CLBLL_L_X4Y155_SLICE_X4Y155_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y155_SLICE_X5Y155_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y155_SLICE_X5Y155_DO5),
.O6(CLBLL_L_X4Y155_SLICE_X5Y155_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y155_SLICE_X5Y155_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y155_SLICE_X5Y155_CO5),
.O6(CLBLL_L_X4Y155_SLICE_X5Y155_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y155_SLICE_X5Y155_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y155_SLICE_X5Y155_BO5),
.O6(CLBLL_L_X4Y155_SLICE_X5Y155_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffdffffffffdffff)
  ) CLBLL_L_X4Y155_SLICE_X5Y155_ALUT (
.I0(RIOB33_X105Y131_IOB_X1Y132_I),
.I1(RIOB33_X105Y133_IOB_X1Y134_I),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(CLBLL_L_X2Y155_SLICE_X1Y155_DO6),
.I4(RIOB33_X105Y133_IOB_X1Y133_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y155_SLICE_X5Y155_AO5),
.O6(CLBLL_L_X4Y155_SLICE_X5Y155_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X36Y146_SLICE_X54Y146_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X36Y146_SLICE_X54Y146_DO5),
.O6(CLBLL_L_X36Y146_SLICE_X54Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X36Y146_SLICE_X54Y146_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X36Y146_SLICE_X54Y146_CO5),
.O6(CLBLL_L_X36Y146_SLICE_X54Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X36Y146_SLICE_X54Y146_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X36Y146_SLICE_X54Y146_BO5),
.O6(CLBLL_L_X36Y146_SLICE_X54Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h1111000011110000)
  ) CLBLL_L_X36Y146_SLICE_X54Y146_ALUT (
.I0(CLBLM_R_X7Y146_SLICE_X8Y146_CQ),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(1'b1),
.I3(1'b1),
.I4(RIOB33_X105Y119_IOB_X1Y119_I),
.I5(1'b1),
.O5(CLBLL_L_X36Y146_SLICE_X54Y146_AO5),
.O6(CLBLL_L_X36Y146_SLICE_X54Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X36Y146_SLICE_X55Y146_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X36Y146_SLICE_X55Y146_DO5),
.O6(CLBLL_L_X36Y146_SLICE_X55Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X36Y146_SLICE_X55Y146_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X36Y146_SLICE_X55Y146_CO5),
.O6(CLBLL_L_X36Y146_SLICE_X55Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X36Y146_SLICE_X55Y146_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X36Y146_SLICE_X55Y146_BO5),
.O6(CLBLL_L_X36Y146_SLICE_X55Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X36Y146_SLICE_X55Y146_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X36Y146_SLICE_X55Y146_AO5),
.O6(CLBLL_L_X36Y146_SLICE_X55Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y126_SLICE_X78Y126_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y126_SLICE_X78Y126_DO5),
.O6(CLBLL_L_X52Y126_SLICE_X78Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y126_SLICE_X78Y126_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y126_SLICE_X78Y126_CO5),
.O6(CLBLL_L_X52Y126_SLICE_X78Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y126_SLICE_X78Y126_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y126_SLICE_X78Y126_BO5),
.O6(CLBLL_L_X52Y126_SLICE_X78Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00ff00ff00ff)
  ) CLBLL_L_X52Y126_SLICE_X78Y126_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(RIOB33_X105Y123_IOB_X1Y124_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y126_SLICE_X78Y126_AO5),
.O6(CLBLL_L_X52Y126_SLICE_X78Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y126_SLICE_X79Y126_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y126_SLICE_X79Y126_DO5),
.O6(CLBLL_L_X52Y126_SLICE_X79Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y126_SLICE_X79Y126_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y126_SLICE_X79Y126_CO5),
.O6(CLBLL_L_X52Y126_SLICE_X79Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y126_SLICE_X79Y126_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y126_SLICE_X79Y126_BO5),
.O6(CLBLL_L_X52Y126_SLICE_X79Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y126_SLICE_X79Y126_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y126_SLICE_X79Y126_AO5),
.O6(CLBLL_L_X52Y126_SLICE_X79Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y142_SLICE_X10Y142_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y142_SLICE_X10Y142_AO5),
.Q(CLBLM_L_X8Y142_SLICE_X10Y142_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y142_SLICE_X10Y142_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y142_SLICE_X10Y142_AO6),
.Q(CLBLM_L_X8Y142_SLICE_X10Y142_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y142_SLICE_X10Y142_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y142_SLICE_X10Y142_DO5),
.O6(CLBLM_L_X8Y142_SLICE_X10Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y142_SLICE_X10Y142_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y142_SLICE_X10Y142_CO5),
.O6(CLBLM_L_X8Y142_SLICE_X10Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y142_SLICE_X10Y142_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y142_SLICE_X10Y142_BO5),
.O6(CLBLM_L_X8Y142_SLICE_X10Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5a0f5a0ffaa5500)
  ) CLBLM_L_X8Y142_SLICE_X10Y142_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(1'b1),
.I2(CLBLM_R_X3Y142_SLICE_X2Y142_BQ),
.I3(RIOB33_X105Y125_IOB_X1Y126_I),
.I4(CLBLM_R_X11Y152_SLICE_X15Y152_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y142_SLICE_X10Y142_AO5),
.O6(CLBLM_L_X8Y142_SLICE_X10Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y142_SLICE_X11Y142_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y142_SLICE_X11Y142_DO5),
.O6(CLBLM_L_X8Y142_SLICE_X11Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y142_SLICE_X11Y142_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y142_SLICE_X11Y142_CO5),
.O6(CLBLM_L_X8Y142_SLICE_X11Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y142_SLICE_X11Y142_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y142_SLICE_X11Y142_BO5),
.O6(CLBLM_L_X8Y142_SLICE_X11Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y142_SLICE_X11Y142_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y142_SLICE_X11Y142_AO5),
.O6(CLBLM_L_X8Y142_SLICE_X11Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y143_SLICE_X10Y143_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y143_SLICE_X10Y143_AO6),
.Q(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y143_SLICE_X10Y143_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y143_SLICE_X10Y143_BO6),
.Q(CLBLM_L_X8Y143_SLICE_X10Y143_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y143_SLICE_X10Y143_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y143_SLICE_X10Y143_DO5),
.O6(CLBLM_L_X8Y143_SLICE_X10Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000100010)
  ) CLBLM_L_X8Y143_SLICE_X10Y143_CLUT (
.I0(CLBLM_L_X8Y143_SLICE_X10Y143_BQ),
.I1(CLBLM_R_X7Y143_SLICE_X9Y143_CQ),
.I2(CLBLM_L_X8Y143_SLICE_X11Y143_BO6),
.I3(CLBLM_R_X7Y143_SLICE_X9Y143_DO6),
.I4(1'b1),
.I5(CLBLM_L_X8Y145_SLICE_X10Y145_BQ),
.O5(CLBLM_L_X8Y143_SLICE_X10Y143_CO5),
.O6(CLBLM_L_X8Y143_SLICE_X10Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc55555500)
  ) CLBLM_L_X8Y143_SLICE_X10Y143_BLUT (
.I0(CLBLM_R_X5Y143_SLICE_X7Y143_CO6),
.I1(CLBLM_L_X8Y148_SLICE_X10Y148_BQ),
.I2(1'b1),
.I3(CLBLM_R_X5Y143_SLICE_X6Y143_AQ),
.I4(CLBLM_L_X8Y143_SLICE_X10Y143_BQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y143_SLICE_X10Y143_BO5),
.O6(CLBLM_L_X8Y143_SLICE_X10Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0031313131)
  ) CLBLM_L_X8Y143_SLICE_X10Y143_ALUT (
.I0(RIOB33_X105Y141_IOB_X1Y142_I),
.I1(CLBLM_L_X10Y143_SLICE_X12Y143_AO6),
.I2(CLBLM_R_X5Y142_SLICE_X7Y142_AQ),
.I3(CLBLL_L_X4Y149_SLICE_X4Y149_BQ),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y143_SLICE_X10Y143_AO5),
.O6(CLBLM_L_X8Y143_SLICE_X10Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y143_SLICE_X11Y143_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y143_SLICE_X11Y143_AO6),
.Q(CLBLM_L_X8Y143_SLICE_X11Y143_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7d7d7d7dbebebebe)
  ) CLBLM_L_X8Y143_SLICE_X11Y143_DLUT (
.I0(CLBLM_L_X8Y148_SLICE_X10Y148_BQ),
.I1(CLBLM_R_X11Y143_SLICE_X14Y143_AQ),
.I2(CLBLM_R_X7Y145_SLICE_X9Y145_CQ),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X5Y143_SLICE_X6Y143_AQ),
.O5(CLBLM_L_X8Y143_SLICE_X11Y143_DO5),
.O6(CLBLM_L_X8Y143_SLICE_X11Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000c300000000c3)
  ) CLBLM_L_X8Y143_SLICE_X11Y143_CLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y145_SLICE_X10Y145_BQ),
.I2(CLBLM_R_X3Y145_SLICE_X3Y145_DQ),
.I3(CLBLM_R_X15Y151_SLICE_X20Y151_AQ),
.I4(CLBLM_L_X8Y143_SLICE_X11Y143_DO6),
.I5(CLBLM_L_X8Y143_SLICE_X11Y143_AQ),
.O5(CLBLM_L_X8Y143_SLICE_X11Y143_CO5),
.O6(CLBLM_L_X8Y143_SLICE_X11Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000001)
  ) CLBLM_L_X8Y143_SLICE_X11Y143_BLUT (
.I0(CLBLM_L_X8Y144_SLICE_X10Y144_BQ),
.I1(CLBLM_R_X5Y143_SLICE_X6Y143_AQ),
.I2(CLBLM_L_X8Y144_SLICE_X11Y144_AQ),
.I3(CLBLM_L_X10Y145_SLICE_X12Y145_DQ),
.I4(CLBLM_L_X10Y144_SLICE_X12Y144_BQ),
.I5(CLBLM_R_X11Y143_SLICE_X14Y143_AQ),
.O5(CLBLM_L_X8Y143_SLICE_X11Y143_BO5),
.O6(CLBLM_L_X8Y143_SLICE_X11Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haafeaafe00540054)
  ) CLBLM_L_X8Y143_SLICE_X11Y143_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y145_SLICE_X10Y145_BQ),
.I2(CLBLM_L_X8Y143_SLICE_X11Y143_AQ),
.I3(CLBLM_R_X5Y143_SLICE_X7Y143_CO6),
.I4(1'b1),
.I5(CLBLM_L_X10Y143_SLICE_X13Y143_AQ),
.O5(CLBLM_L_X8Y143_SLICE_X11Y143_AO5),
.O6(CLBLM_L_X8Y143_SLICE_X11Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y144_SLICE_X10Y144_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y144_SLICE_X10Y144_AO6),
.Q(CLBLM_L_X8Y144_SLICE_X10Y144_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y144_SLICE_X10Y144_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y144_SLICE_X10Y144_BO6),
.Q(CLBLM_L_X8Y144_SLICE_X10Y144_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y144_SLICE_X10Y144_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y144_SLICE_X10Y144_CO6),
.Q(CLBLM_L_X8Y144_SLICE_X10Y144_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc00330f0f0f0f)
  ) CLBLM_L_X8Y144_SLICE_X10Y144_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y144_SLICE_X10Y144_CQ),
.I2(CLBLM_L_X10Y146_SLICE_X12Y146_CQ),
.I3(CLBLM_L_X8Y143_SLICE_X10Y143_CO6),
.I4(CLBLM_L_X8Y145_SLICE_X11Y145_CQ),
.I5(CLBLL_L_X4Y143_SLICE_X4Y143_CO6),
.O5(CLBLM_L_X8Y144_SLICE_X10Y144_DO5),
.O6(CLBLM_L_X8Y144_SLICE_X10Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0afacafac)
  ) CLBLM_L_X8Y144_SLICE_X10Y144_CLUT (
.I0(CLBLM_L_X8Y150_SLICE_X11Y150_BQ),
.I1(CLBLM_L_X8Y144_SLICE_X10Y144_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y143_SLICE_X9Y143_CQ),
.I4(1'b1),
.I5(CLBLM_R_X5Y143_SLICE_X7Y143_CO6),
.O5(CLBLM_L_X8Y144_SLICE_X10Y144_CO5),
.O6(CLBLM_L_X8Y144_SLICE_X10Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hafacafaca0a0a0a0)
  ) CLBLM_L_X8Y144_SLICE_X10Y144_BLUT (
.I0(CLBLM_R_X7Y145_SLICE_X9Y145_AQ),
.I1(CLBLM_L_X8Y144_SLICE_X10Y144_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y144_SLICE_X12Y144_BQ),
.I4(1'b1),
.I5(CLBLM_R_X7Y142_SLICE_X8Y142_DO6),
.O5(CLBLM_L_X8Y144_SLICE_X10Y144_BO5),
.O6(CLBLM_L_X8Y144_SLICE_X10Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffccfedc33003210)
  ) CLBLM_L_X8Y144_SLICE_X10Y144_ALUT (
.I0(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X8Y144_SLICE_X10Y144_AQ),
.I3(CLBLM_R_X7Y144_SLICE_X9Y144_AQ),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLM_L_X10Y144_SLICE_X12Y144_BQ),
.O5(CLBLM_L_X8Y144_SLICE_X10Y144_AO5),
.O6(CLBLM_L_X8Y144_SLICE_X10Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y144_SLICE_X11Y144_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y144_SLICE_X11Y144_AO6),
.Q(CLBLM_L_X8Y144_SLICE_X11Y144_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000000f0f0f0f)
  ) CLBLM_L_X8Y144_SLICE_X11Y144_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_L_X10Y144_SLICE_X12Y144_DO6),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X5Y143_SLICE_X7Y143_CO6),
.O5(CLBLM_L_X8Y144_SLICE_X11Y144_DO5),
.O6(CLBLM_L_X8Y144_SLICE_X11Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffeeffffffee)
  ) CLBLM_L_X8Y144_SLICE_X11Y144_CLUT (
.I0(CLBLM_R_X11Y144_SLICE_X14Y144_AQ),
.I1(CLBLM_L_X10Y142_SLICE_X13Y142_AQ),
.I2(1'b1),
.I3(CLBLM_L_X8Y147_SLICE_X10Y147_DQ),
.I4(CLBLM_R_X7Y144_SLICE_X9Y144_CQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y144_SLICE_X11Y144_CO5),
.O6(CLBLM_L_X8Y144_SLICE_X11Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0021000021000000)
  ) CLBLM_L_X8Y144_SLICE_X11Y144_BLUT (
.I0(CLBLM_L_X10Y145_SLICE_X13Y145_A5Q),
.I1(CLBLM_L_X10Y143_SLICE_X12Y143_CO6),
.I2(CLBLM_R_X5Y143_SLICE_X7Y143_AQ),
.I3(CLBLM_L_X8Y144_SLICE_X10Y144_DO6),
.I4(CLBLM_L_X8Y143_SLICE_X11Y143_CO6),
.I5(CLBLM_L_X10Y146_SLICE_X12Y146_CQ),
.O5(CLBLM_L_X8Y144_SLICE_X11Y144_BO5),
.O6(CLBLM_L_X8Y144_SLICE_X11Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaa5500faaa5000)
  ) CLBLM_L_X8Y144_SLICE_X11Y144_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(1'b1),
.I2(CLBLM_L_X10Y145_SLICE_X12Y145_DQ),
.I3(CLBLM_R_X7Y142_SLICE_X8Y142_DO6),
.I4(CLBLM_L_X8Y152_SLICE_X10Y152_DQ),
.I5(CLBLM_L_X8Y144_SLICE_X11Y144_AQ),
.O5(CLBLM_L_X8Y144_SLICE_X11Y144_AO5),
.O6(CLBLM_L_X8Y144_SLICE_X11Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y145_SLICE_X10Y145_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y147_SLICE_X12Y147_BO6),
.Q(CLBLM_L_X8Y145_SLICE_X10Y145_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y145_SLICE_X10Y145_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y145_SLICE_X10Y145_AO6),
.Q(CLBLM_L_X8Y145_SLICE_X10Y145_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y145_SLICE_X10Y145_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y145_SLICE_X10Y145_BO6),
.Q(CLBLM_L_X8Y145_SLICE_X10Y145_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000c000d5)
  ) CLBLM_L_X8Y145_SLICE_X10Y145_DLUT (
.I0(CLBLM_L_X10Y144_SLICE_X13Y144_AQ),
.I1(CLBLM_L_X8Y148_SLICE_X10Y148_CO6),
.I2(CLBLL_L_X4Y154_SLICE_X4Y154_CO6),
.I3(CLBLM_L_X8Y145_SLICE_X10Y145_CO6),
.I4(CLBLM_R_X5Y144_SLICE_X7Y144_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y145_SLICE_X10Y145_DO5),
.O6(CLBLM_L_X8Y145_SLICE_X10Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffff2000f000f)
  ) CLBLM_L_X8Y145_SLICE_X10Y145_CLUT (
.I0(CLBLM_L_X10Y144_SLICE_X13Y144_AQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_R_X5Y144_SLICE_X7Y144_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y145_SLICE_X10Y145_CO5),
.O6(CLBLM_L_X8Y145_SLICE_X10Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf4f5f4f504050405)
  ) CLBLM_L_X8Y145_SLICE_X10Y145_BLUT (
.I0(CLBLL_L_X4Y145_SLICE_X5Y145_DO6),
.I1(CLBLM_L_X8Y145_SLICE_X10Y145_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y144_SLICE_X10Y144_DO6),
.I4(1'b1),
.I5(CLBLM_R_X7Y153_SLICE_X9Y153_BQ),
.O5(CLBLM_L_X8Y145_SLICE_X10Y145_BO5),
.O6(CLBLM_L_X8Y145_SLICE_X10Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f02222f0f02222)
  ) CLBLM_L_X8Y145_SLICE_X10Y145_ALUT (
.I0(CLBLM_L_X10Y147_SLICE_X13Y147_AQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLL_L_X4Y144_SLICE_X5Y144_BQ),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y145_SLICE_X10Y145_AO5),
.O6(CLBLM_L_X8Y145_SLICE_X10Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y145_SLICE_X11Y145_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y145_SLICE_X11Y145_AO5),
.Q(CLBLM_L_X8Y145_SLICE_X11Y145_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y145_SLICE_X11Y145_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y145_SLICE_X11Y145_BO5),
.Q(CLBLM_L_X8Y145_SLICE_X11Y145_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y145_SLICE_X11Y145_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y145_SLICE_X11Y145_AO6),
.Q(CLBLM_L_X8Y145_SLICE_X11Y145_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y145_SLICE_X11Y145_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y145_SLICE_X11Y145_BO6),
.Q(CLBLM_L_X8Y145_SLICE_X11Y145_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y145_SLICE_X11Y145_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y145_SLICE_X11Y145_CO6),
.Q(CLBLM_L_X8Y145_SLICE_X11Y145_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y145_SLICE_X11Y145_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y145_SLICE_X11Y145_DO6),
.Q(CLBLM_L_X8Y145_SLICE_X11Y145_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00f0f0d8d8)
  ) CLBLM_L_X8Y145_SLICE_X11Y145_DLUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_R_X7Y145_SLICE_X9Y145_DO6),
.I2(CLBLM_L_X8Y145_SLICE_X11Y145_DQ),
.I3(CLBLM_L_X10Y145_SLICE_X12Y145_DQ),
.I4(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y145_SLICE_X11Y145_DO5),
.O6(CLBLM_L_X8Y145_SLICE_X11Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0ee00ee00)
  ) CLBLM_L_X8Y145_SLICE_X11Y145_CLUT (
.I0(CLBLM_L_X8Y144_SLICE_X10Y144_CQ),
.I1(CLBLM_L_X8Y145_SLICE_X11Y145_CQ),
.I2(CLBLM_L_X8Y144_SLICE_X11Y144_AQ),
.I3(CLBLM_R_X7Y142_SLICE_X8Y142_DO6),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y145_SLICE_X11Y145_CO5),
.O6(CLBLM_L_X8Y145_SLICE_X11Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaf0aaf0ccffcc00)
  ) CLBLM_L_X8Y145_SLICE_X11Y145_BLUT (
.I0(CLBLM_R_X11Y146_SLICE_X14Y146_AQ),
.I1(CLBLM_R_X7Y144_SLICE_X8Y144_BQ),
.I2(CLBLM_L_X10Y150_SLICE_X12Y150_A5Q),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y103_IOB_X1Y103_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y145_SLICE_X11Y145_BO5),
.O6(CLBLM_L_X8Y145_SLICE_X11Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hacacacacc0cfc0c0)
  ) CLBLM_L_X8Y145_SLICE_X11Y145_ALUT (
.I0(CLBLM_L_X8Y145_SLICE_X11Y145_B5Q),
.I1(CLBLM_L_X10Y146_SLICE_X12Y146_AQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_L_X8Y145_SLICE_X11Y145_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X8Y145_SLICE_X11Y145_AO5),
.O6(CLBLM_L_X8Y145_SLICE_X11Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y146_SLICE_X10Y146_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y146_SLICE_X10Y146_BO5),
.Q(CLBLM_L_X8Y146_SLICE_X10Y146_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y146_SLICE_X10Y146_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y146_SLICE_X10Y146_AO6),
.Q(CLBLM_L_X8Y146_SLICE_X10Y146_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y146_SLICE_X10Y146_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y146_SLICE_X10Y146_BO6),
.Q(CLBLM_L_X8Y146_SLICE_X10Y146_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y146_SLICE_X10Y146_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y146_SLICE_X10Y146_CO6),
.Q(CLBLM_L_X8Y146_SLICE_X10Y146_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h55df55df55005500)
  ) CLBLM_L_X8Y146_SLICE_X10Y146_DLUT (
.I0(CLBLM_L_X8Y148_SLICE_X10Y148_CO5),
.I1(CLBLL_L_X2Y153_SLICE_X1Y153_DO6),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X5Y144_SLICE_X7Y144_AQ),
.I4(1'b1),
.I5(CLBLM_L_X10Y144_SLICE_X13Y144_AQ),
.O5(CLBLM_L_X8Y146_SLICE_X10Y146_DO5),
.O6(CLBLM_L_X8Y146_SLICE_X10Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f4f0f400040004)
  ) CLBLM_L_X8Y146_SLICE_X10Y146_CLUT (
.I0(CLBLM_L_X8Y147_SLICE_X11Y147_CO6),
.I1(CLBLM_L_X10Y147_SLICE_X13Y147_AQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(1'b1),
.I5(CLBLM_L_X8Y142_SLICE_X10Y142_A5Q),
.O5(CLBLM_L_X8Y146_SLICE_X10Y146_CO5),
.O6(CLBLM_L_X8Y146_SLICE_X10Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0afa0cacfcacf)
  ) CLBLM_L_X8Y146_SLICE_X10Y146_BLUT (
.I0(CLBLM_R_X7Y146_SLICE_X8Y146_CQ),
.I1(CLBLM_R_X3Y148_SLICE_X2Y148_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y119_IOB_X1Y119_I),
.I4(CLBLM_L_X8Y146_SLICE_X10Y146_BQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y146_SLICE_X10Y146_BO5),
.O6(CLBLM_L_X8Y146_SLICE_X10Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f6f0f600060006)
  ) CLBLM_L_X8Y146_SLICE_X10Y146_ALUT (
.I0(CLBLM_L_X8Y147_SLICE_X11Y147_AO5),
.I1(CLBLM_L_X8Y152_SLICE_X10Y152_DQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(1'b1),
.I5(CLBLM_R_X7Y146_SLICE_X8Y146_DQ),
.O5(CLBLM_L_X8Y146_SLICE_X10Y146_AO5),
.O6(CLBLM_L_X8Y146_SLICE_X10Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y146_SLICE_X11Y146_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y146_SLICE_X11Y146_AO6),
.Q(CLBLM_L_X8Y146_SLICE_X11Y146_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y146_SLICE_X11Y146_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y146_SLICE_X11Y146_BO6),
.Q(CLBLM_L_X8Y146_SLICE_X11Y146_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000001100000011)
  ) CLBLM_L_X8Y146_SLICE_X11Y146_DLUT (
.I0(CLBLL_L_X4Y150_SLICE_X4Y150_AQ),
.I1(CLBLL_L_X4Y149_SLICE_X4Y149_DQ),
.I2(1'b1),
.I3(CLBLM_L_X8Y146_SLICE_X11Y146_AQ),
.I4(CLBLM_R_X11Y146_SLICE_X14Y146_BQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y146_SLICE_X11Y146_DO5),
.O6(CLBLM_L_X8Y146_SLICE_X11Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa22aaaaaa22aaa0)
  ) CLBLM_L_X8Y146_SLICE_X11Y146_CLUT (
.I0(RIOB33_X105Y121_IOB_X1Y121_I),
.I1(CLBLM_L_X8Y145_SLICE_X11Y145_DQ),
.I2(CLBLM_R_X5Y149_SLICE_X6Y149_CO6),
.I3(CLBLM_L_X10Y147_SLICE_X13Y147_AQ),
.I4(CLBLM_L_X8Y146_SLICE_X11Y146_DO6),
.I5(CLBLM_R_X3Y153_SLICE_X2Y153_DO6),
.O5(CLBLM_L_X8Y146_SLICE_X11Y146_CO5),
.O6(CLBLM_L_X8Y146_SLICE_X11Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f05500f0f04400)
  ) CLBLM_L_X8Y146_SLICE_X11Y146_BLUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_L_X8Y146_SLICE_X11Y146_BQ),
.I2(CLBLM_L_X8Y146_SLICE_X11Y146_AQ),
.I3(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y146_SLICE_X10Y146_DO6),
.O5(CLBLM_L_X8Y146_SLICE_X11Y146_BO5),
.O6(CLBLM_L_X8Y146_SLICE_X11Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcca0cca0ccf0ccf0)
  ) CLBLM_L_X8Y146_SLICE_X11Y146_ALUT (
.I0(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.I1(CLBLM_L_X8Y145_SLICE_X11Y145_DQ),
.I2(CLBLM_L_X8Y146_SLICE_X11Y146_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_L_X8Y146_SLICE_X11Y146_AO5),
.O6(CLBLM_L_X8Y146_SLICE_X11Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y147_SLICE_X10Y147_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y147_SLICE_X10Y147_AO6),
.Q(CLBLM_L_X8Y147_SLICE_X10Y147_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y147_SLICE_X10Y147_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y147_SLICE_X10Y147_BO6),
.Q(CLBLM_L_X8Y147_SLICE_X10Y147_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y147_SLICE_X10Y147_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y147_SLICE_X10Y147_CO6),
.Q(CLBLM_L_X8Y147_SLICE_X10Y147_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y147_SLICE_X10Y147_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y147_SLICE_X10Y147_DO6),
.Q(CLBLM_L_X8Y147_SLICE_X10Y147_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haa30aa30aa30aa30)
  ) CLBLM_L_X8Y147_SLICE_X10Y147_DLUT (
.I0(CLBLM_L_X8Y150_SLICE_X10Y150_BQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_L_X8Y147_SLICE_X10Y147_DQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y147_SLICE_X10Y147_DO5),
.O6(CLBLM_L_X8Y147_SLICE_X10Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00eeeee0e0)
  ) CLBLM_L_X8Y147_SLICE_X10Y147_CLUT (
.I0(CLBLM_L_X8Y148_SLICE_X11Y148_CO6),
.I1(CLBLM_L_X8Y147_SLICE_X10Y147_CQ),
.I2(RIOB33_X105Y117_IOB_X1Y118_I),
.I3(CLBLM_L_X12Y150_SLICE_X16Y150_CQ),
.I4(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y147_SLICE_X10Y147_CO5),
.O6(CLBLM_L_X8Y147_SLICE_X10Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0aa88aa88)
  ) CLBLM_L_X8Y147_SLICE_X10Y147_BLUT (
.I0(CLBLM_L_X8Y152_SLICE_X11Y152_BO6),
.I1(CLBLM_L_X8Y147_SLICE_X10Y147_BQ),
.I2(CLBLM_L_X8Y145_SLICE_X10Y145_AQ),
.I3(CLBLM_R_X7Y145_SLICE_X8Y145_CQ),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y147_SLICE_X10Y147_BO5),
.O6(CLBLM_L_X8Y147_SLICE_X10Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffccf0ffffcca0)
  ) CLBLM_L_X8Y147_SLICE_X10Y147_ALUT (
.I0(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.I1(CLBLL_L_X4Y144_SLICE_X5Y144_A5Q),
.I2(CLBLM_L_X8Y147_SLICE_X10Y147_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y149_SLICE_X9Y149_DO6),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_L_X8Y147_SLICE_X10Y147_AO5),
.O6(CLBLM_L_X8Y147_SLICE_X10Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_L_X8Y147_SLICE_X11Y147_DLUT (
.I0(CLBLM_L_X10Y146_SLICE_X13Y146_AQ),
.I1(CLBLM_L_X10Y147_SLICE_X13Y147_BQ),
.I2(CLBLM_R_X7Y147_SLICE_X8Y147_CQ),
.I3(CLBLL_L_X4Y148_SLICE_X4Y148_CQ),
.I4(CLBLM_L_X8Y145_SLICE_X10Y145_AQ),
.I5(CLBLM_R_X5Y148_SLICE_X6Y148_BQ),
.O5(CLBLM_L_X8Y147_SLICE_X11Y147_DO5),
.O6(CLBLM_L_X8Y147_SLICE_X11Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_L_X8Y147_SLICE_X11Y147_CLUT (
.I0(CLBLM_R_X7Y146_SLICE_X9Y146_DO6),
.I1(CLBLM_R_X7Y147_SLICE_X9Y147_DO6),
.I2(CLBLM_L_X10Y146_SLICE_X12Y146_DQ),
.I3(CLBLM_L_X10Y149_SLICE_X13Y149_DQ),
.I4(CLBLM_L_X8Y147_SLICE_X11Y147_DO6),
.I5(CLBLM_L_X10Y150_SLICE_X12Y150_BQ),
.O5(CLBLM_L_X8Y147_SLICE_X11Y147_CO5),
.O6(CLBLM_L_X8Y147_SLICE_X11Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3636cccc05050505)
  ) CLBLM_L_X8Y147_SLICE_X11Y147_BLUT (
.I0(CLBLM_R_X5Y149_SLICE_X6Y149_CO6),
.I1(CLBLM_R_X7Y145_SLICE_X9Y145_BQ),
.I2(CLBLL_L_X2Y153_SLICE_X1Y153_DO6),
.I3(1'b1),
.I4(CLBLM_L_X8Y151_SLICE_X10Y151_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y147_SLICE_X11Y147_BO5),
.O6(CLBLM_L_X8Y147_SLICE_X11Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbb88888fff00000)
  ) CLBLM_L_X8Y147_SLICE_X11Y147_ALUT (
.I0(CLBLM_L_X10Y151_SLICE_X12Y151_BQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X5Y148_SLICE_X6Y148_BQ),
.I3(CLBLM_R_X7Y144_SLICE_X8Y144_BQ),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y147_SLICE_X11Y147_AO5),
.O6(CLBLM_L_X8Y147_SLICE_X11Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y148_SLICE_X10Y148_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y148_SLICE_X10Y148_AO5),
.Q(CLBLM_L_X8Y148_SLICE_X10Y148_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y148_SLICE_X10Y148_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y148_SLICE_X10Y148_AO6),
.Q(CLBLM_L_X8Y148_SLICE_X10Y148_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y148_SLICE_X10Y148_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y153_SLICE_X10Y153_CO6),
.Q(CLBLM_L_X8Y148_SLICE_X10Y148_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f1e0f0feeffeeff)
  ) CLBLM_L_X8Y148_SLICE_X10Y148_DLUT (
.I0(CLBLM_R_X7Y145_SLICE_X8Y145_BQ),
.I1(CLBLM_R_X7Y143_SLICE_X8Y143_AQ),
.I2(CLBLM_L_X8Y148_SLICE_X10Y148_AQ),
.I3(CLBLM_R_X5Y145_SLICE_X6Y145_CQ),
.I4(CLBLL_L_X4Y143_SLICE_X4Y143_BQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y148_SLICE_X10Y148_DO5),
.O6(CLBLM_L_X8Y148_SLICE_X10Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hacacacac0f0f0fff)
  ) CLBLM_L_X8Y148_SLICE_X10Y148_CLUT (
.I0(CLBLM_L_X10Y146_SLICE_X12Y146_DQ),
.I1(CLBLM_R_X11Y148_SLICE_X14Y148_BQ),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLM_L_X8Y152_SLICE_X10Y152_CQ),
.I4(CLBLM_R_X7Y147_SLICE_X8Y147_CQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y148_SLICE_X10Y148_CO5),
.O6(CLBLM_L_X8Y148_SLICE_X10Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfc0cac0ff00aa00)
  ) CLBLM_L_X8Y148_SLICE_X10Y148_BLUT (
.I0(CLBLM_R_X7Y149_SLICE_X8Y149_CQ),
.I1(CLBLM_R_X7Y146_SLICE_X9Y146_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(CLBLM_L_X8Y147_SLICE_X10Y147_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y148_SLICE_X10Y148_BO5),
.O6(CLBLM_L_X8Y148_SLICE_X10Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0e2c0e2bbbb8888)
  ) CLBLM_L_X8Y148_SLICE_X10Y148_ALUT (
.I0(CLBLM_L_X8Y148_SLICE_X10Y148_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y155_SLICE_X13Y155_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X5Y147_SLICE_X7Y147_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y148_SLICE_X10Y148_AO5),
.O6(CLBLM_L_X8Y148_SLICE_X10Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y148_SLICE_X11Y148_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y148_SLICE_X11Y148_AO6),
.Q(CLBLM_L_X8Y148_SLICE_X11Y148_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00aa00aa00aa00aa)
  ) CLBLM_L_X8Y148_SLICE_X11Y148_DLUT (
.I0(CLBLM_R_X7Y145_SLICE_X8Y145_BQ),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X7Y143_SLICE_X8Y143_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y148_SLICE_X11Y148_DO5),
.O6(CLBLM_L_X8Y148_SLICE_X11Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hebee4144eeee4444)
  ) CLBLM_L_X8Y148_SLICE_X11Y148_CLUT (
.I0(RIOB33_X105Y121_IOB_X1Y121_I),
.I1(CLBLM_L_X8Y147_SLICE_X10Y147_DQ),
.I2(CLBLL_L_X4Y143_SLICE_X4Y143_BQ),
.I3(CLBLM_R_X5Y145_SLICE_X6Y145_CQ),
.I4(CLBLM_R_X7Y147_SLICE_X8Y147_CQ),
.I5(CLBLM_L_X8Y148_SLICE_X11Y148_DO6),
.O5(CLBLM_L_X8Y148_SLICE_X11Y148_CO5),
.O6(CLBLM_L_X8Y148_SLICE_X11Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff70000ff080000)
  ) CLBLM_L_X8Y148_SLICE_X11Y148_BLUT (
.I0(CLBLM_R_X7Y143_SLICE_X8Y143_AQ),
.I1(CLBLM_L_X8Y149_SLICE_X10Y149_AO6),
.I2(CLBLM_R_X7Y145_SLICE_X8Y145_BQ),
.I3(CLBLM_R_X7Y152_SLICE_X9Y152_CQ),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(CLBLM_L_X8Y145_SLICE_X11Y145_A5Q),
.O5(CLBLM_L_X8Y148_SLICE_X11Y148_BO5),
.O6(CLBLM_L_X8Y148_SLICE_X11Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00eeeeff00e0e0)
  ) CLBLM_L_X8Y148_SLICE_X11Y148_ALUT (
.I0(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_L_X8Y148_SLICE_X11Y148_AQ),
.I3(CLBLL_L_X4Y148_SLICE_X4Y148_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X5Y148_SLICE_X7Y148_DO6),
.O5(CLBLM_L_X8Y148_SLICE_X11Y148_AO5),
.O6(CLBLM_L_X8Y148_SLICE_X11Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0f0f0f0f0e)
  ) CLBLM_L_X8Y149_SLICE_X10Y149_DLUT (
.I0(CLBLM_R_X3Y149_SLICE_X3Y149_BQ),
.I1(CLBLM_R_X7Y154_SLICE_X8Y154_CQ),
.I2(CLBLM_L_X8Y151_SLICE_X11Y151_DQ),
.I3(CLBLM_L_X8Y144_SLICE_X11Y144_CO6),
.I4(CLBLM_R_X5Y149_SLICE_X7Y149_CQ),
.I5(CLBLM_L_X8Y149_SLICE_X10Y149_BO6),
.O5(CLBLM_L_X8Y149_SLICE_X10Y149_DO5),
.O6(CLBLM_L_X8Y149_SLICE_X10Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff6aaa00006aaa)
  ) CLBLM_L_X8Y149_SLICE_X10Y149_CLUT (
.I0(CLBLM_R_X3Y149_SLICE_X3Y149_BQ),
.I1(CLBLM_L_X8Y149_SLICE_X10Y149_AO6),
.I2(CLBLM_R_X7Y143_SLICE_X8Y143_AQ),
.I3(CLBLM_R_X7Y145_SLICE_X8Y145_BQ),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(CLBLM_R_X5Y148_SLICE_X6Y148_BQ),
.O5(CLBLM_L_X8Y149_SLICE_X10Y149_CO5),
.O6(CLBLM_L_X8Y149_SLICE_X10Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_L_X8Y149_SLICE_X10Y149_BLUT (
.I0(CLBLM_L_X8Y145_SLICE_X11Y145_A5Q),
.I1(CLBLM_L_X8Y151_SLICE_X10Y151_BQ),
.I2(CLBLM_L_X8Y148_SLICE_X10Y148_AQ),
.I3(CLBLM_R_X7Y152_SLICE_X9Y152_BQ),
.I4(CLBLM_R_X7Y148_SLICE_X9Y148_AQ),
.I5(CLBLM_R_X11Y148_SLICE_X14Y148_CQ),
.O5(CLBLM_L_X8Y149_SLICE_X10Y149_BO5),
.O6(CLBLM_L_X8Y149_SLICE_X10Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h05050505f5f5f5f5)
  ) CLBLM_L_X8Y149_SLICE_X10Y149_ALUT (
.I0(CLBLL_L_X4Y143_SLICE_X4Y143_BQ),
.I1(1'b1),
.I2(CLBLM_R_X5Y145_SLICE_X6Y145_CQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y149_SLICE_X10Y149_AO5),
.O6(CLBLM_L_X8Y149_SLICE_X10Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y149_SLICE_X11Y149_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y149_SLICE_X11Y149_BO5),
.Q(CLBLM_L_X8Y149_SLICE_X11Y149_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y149_SLICE_X11Y149_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y149_SLICE_X11Y149_AO6),
.Q(CLBLM_L_X8Y149_SLICE_X11Y149_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y149_SLICE_X11Y149_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y149_SLICE_X11Y149_BO6),
.Q(CLBLM_L_X8Y149_SLICE_X11Y149_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y149_SLICE_X11Y149_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y149_SLICE_X11Y149_CO6),
.Q(CLBLM_L_X8Y149_SLICE_X11Y149_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h36c99c63c9c96363)
  ) CLBLM_L_X8Y149_SLICE_X11Y149_DLUT (
.I0(CLBLM_L_X8Y149_SLICE_X11Y149_BQ),
.I1(CLBLM_L_X8Y149_SLICE_X11Y149_AQ),
.I2(CLBLM_L_X8Y149_SLICE_X10Y149_DO6),
.I3(CLBLM_L_X8Y149_SLICE_X10Y149_AO6),
.I4(CLBLM_L_X8Y151_SLICE_X11Y151_DQ),
.I5(CLBLM_L_X8Y148_SLICE_X11Y148_DO6),
.O5(CLBLM_L_X8Y149_SLICE_X11Y149_DO5),
.O6(CLBLM_L_X8Y149_SLICE_X11Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdddf000feeef000)
  ) CLBLM_L_X8Y149_SLICE_X11Y149_CLUT (
.I0(CLBLM_L_X8Y146_SLICE_X11Y146_CO6),
.I1(CLBLM_L_X8Y149_SLICE_X11Y149_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y149_SLICE_X8Y149_BQ),
.I4(CLBLM_L_X10Y149_SLICE_X12Y149_AO5),
.I5(CLBLM_L_X8Y149_SLICE_X11Y149_DO6),
.O5(CLBLM_L_X8Y149_SLICE_X11Y149_CO5),
.O6(CLBLM_L_X8Y149_SLICE_X11Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0f3c0c0eeee2222)
  ) CLBLM_L_X8Y149_SLICE_X11Y149_BLUT (
.I0(CLBLM_R_X3Y151_SLICE_X3Y151_AO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y150_SLICE_X12Y150_DQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_L_X8Y149_SLICE_X11Y149_BQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y149_SLICE_X11Y149_BO5),
.O6(CLBLM_L_X8Y149_SLICE_X11Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000f030f030)
  ) CLBLM_L_X8Y149_SLICE_X11Y149_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_L_X8Y149_SLICE_X11Y149_AQ),
.I3(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.I4(CLBLM_L_X12Y149_SLICE_X17Y149_CQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y149_SLICE_X11Y149_AO5),
.O6(CLBLM_L_X8Y149_SLICE_X11Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y150_SLICE_X10Y150_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y150_SLICE_X10Y150_AO6),
.Q(CLBLM_L_X8Y150_SLICE_X10Y150_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y150_SLICE_X10Y150_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y150_SLICE_X10Y150_BO6),
.Q(CLBLM_L_X8Y150_SLICE_X10Y150_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y150_SLICE_X10Y150_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y150_SLICE_X10Y150_CO6),
.Q(CLBLM_L_X8Y150_SLICE_X10Y150_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcd81ccc0ccc0ccc0)
  ) CLBLM_L_X8Y150_SLICE_X10Y150_DLUT (
.I0(CLBLM_L_X8Y149_SLICE_X10Y149_AO5),
.I1(RIOB33_X105Y121_IOB_X1Y121_I),
.I2(CLBLM_R_X7Y154_SLICE_X8Y154_CQ),
.I3(CLBLM_R_X7Y149_SLICE_X8Y149_CQ),
.I4(CLBLM_R_X7Y145_SLICE_X8Y145_BQ),
.I5(CLBLM_R_X7Y143_SLICE_X8Y143_AQ),
.O5(CLBLM_L_X8Y150_SLICE_X10Y150_DO5),
.O6(CLBLM_L_X8Y150_SLICE_X10Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000005a005a)
  ) CLBLM_L_X8Y150_SLICE_X10Y150_CLUT (
.I0(CLBLM_L_X8Y152_SLICE_X11Y152_AQ),
.I1(1'b1),
.I2(CLBLM_L_X8Y148_SLICE_X10Y148_BO5),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X7Y144_SLICE_X8Y144_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y150_SLICE_X10Y150_CO5),
.O6(CLBLM_L_X8Y150_SLICE_X10Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0d1c0d1c0e2c0e2)
  ) CLBLM_L_X8Y150_SLICE_X10Y150_BLUT (
.I0(CLBLM_L_X8Y149_SLICE_X10Y149_CO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y145_SLICE_X12Y145_BQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(1'b1),
.I5(CLBLM_R_X7Y151_SLICE_X9Y151_CQ),
.O5(CLBLM_L_X8Y150_SLICE_X10Y150_BO5),
.O6(CLBLM_L_X8Y150_SLICE_X10Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfe32fe32fe32cc00)
  ) CLBLM_L_X8Y150_SLICE_X10Y150_ALUT (
.I0(CLBLM_L_X8Y149_SLICE_X10Y149_CO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X8Y150_SLICE_X10Y150_AQ),
.I3(CLBLM_L_X10Y153_SLICE_X13Y153_AQ),
.I4(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_L_X8Y150_SLICE_X10Y150_AO5),
.O6(CLBLM_L_X8Y150_SLICE_X10Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y150_SLICE_X11Y150_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y150_SLICE_X11Y150_AO6),
.Q(CLBLM_L_X8Y150_SLICE_X11Y150_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y150_SLICE_X11Y150_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y150_SLICE_X11Y150_BO6),
.Q(CLBLM_L_X8Y150_SLICE_X11Y150_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffdfdfdfd)
  ) CLBLM_L_X8Y150_SLICE_X11Y150_DLUT (
.I0(CLBLM_L_X8Y152_SLICE_X11Y152_AQ),
.I1(CLBLM_L_X10Y147_SLICE_X12Y147_CQ),
.I2(CLBLM_L_X10Y150_SLICE_X12Y150_DQ),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X7Y150_SLICE_X8Y150_CQ),
.O5(CLBLM_L_X8Y150_SLICE_X11Y150_DO5),
.O6(CLBLM_L_X8Y150_SLICE_X11Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffffef)
  ) CLBLM_L_X8Y150_SLICE_X11Y150_CLUT (
.I0(CLBLM_R_X7Y148_SLICE_X9Y148_CQ),
.I1(CLBLM_L_X8Y152_SLICE_X10Y152_DQ),
.I2(CLBLM_L_X8Y152_SLICE_X11Y152_BO5),
.I3(CLBLM_L_X10Y150_SLICE_X12Y150_CQ),
.I4(CLBLM_L_X8Y150_SLICE_X11Y150_DO6),
.I5(CLBLM_R_X7Y149_SLICE_X8Y149_BQ),
.O5(CLBLM_L_X8Y150_SLICE_X11Y150_CO5),
.O6(CLBLM_L_X8Y150_SLICE_X11Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcc00ccffaa00aa)
  ) CLBLM_L_X8Y150_SLICE_X11Y150_BLUT (
.I0(CLBLM_R_X7Y148_SLICE_X8Y148_CQ),
.I1(CLBLM_L_X8Y150_SLICE_X11Y150_BQ),
.I2(1'b1),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y149_SLICE_X13Y149_AQ),
.I5(CLBLM_L_X8Y152_SLICE_X11Y152_BO6),
.O5(CLBLM_L_X8Y150_SLICE_X11Y150_BO5),
.O6(CLBLM_L_X8Y150_SLICE_X11Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haafcaafcaa00aa00)
  ) CLBLM_L_X8Y150_SLICE_X11Y150_ALUT (
.I0(CLBLM_L_X12Y151_SLICE_X16Y151_CQ),
.I1(CLBLM_L_X10Y147_SLICE_X12Y147_CQ),
.I2(CLBLM_L_X8Y150_SLICE_X11Y150_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLM_L_X8Y152_SLICE_X11Y152_BO6),
.O5(CLBLM_L_X8Y150_SLICE_X11Y150_AO5),
.O6(CLBLM_L_X8Y150_SLICE_X11Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y151_SLICE_X10Y151_B5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y151_SLICE_X10Y151_BO5),
.Q(CLBLM_L_X8Y151_SLICE_X10Y151_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y151_SLICE_X10Y151_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y151_SLICE_X10Y151_AO6),
.Q(CLBLM_L_X8Y151_SLICE_X10Y151_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y151_SLICE_X10Y151_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y151_SLICE_X10Y151_BO6),
.Q(CLBLM_L_X8Y151_SLICE_X10Y151_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y151_SLICE_X10Y151_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y151_SLICE_X10Y151_CO6),
.Q(CLBLM_L_X8Y151_SLICE_X10Y151_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y151_SLICE_X10Y151_D_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y151_SLICE_X10Y151_DO6),
.Q(CLBLM_L_X8Y151_SLICE_X10Y151_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hbb88b888bbbbb8b8)
  ) CLBLM_L_X8Y151_SLICE_X10Y151_DLUT (
.I0(CLBLM_L_X10Y144_SLICE_X13Y144_CQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X8Y151_SLICE_X10Y151_DQ),
.I3(CLBLM_R_X11Y150_SLICE_X14Y150_BO6),
.I4(CLBLM_R_X5Y145_SLICE_X7Y145_AQ),
.I5(CLBLM_L_X8Y148_SLICE_X10Y148_A5Q),
.O5(CLBLM_L_X8Y151_SLICE_X10Y151_DO5),
.O6(CLBLM_L_X8Y151_SLICE_X10Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafff8fc0a0f080c)
  ) CLBLM_L_X8Y151_SLICE_X10Y151_CLUT (
.I0(CLBLM_R_X11Y150_SLICE_X14Y150_BO6),
.I1(CLBLM_L_X8Y151_SLICE_X10Y151_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y148_SLICE_X10Y148_A5Q),
.I4(CLBLM_R_X11Y147_SLICE_X14Y147_BQ),
.I5(CLBLM_R_X7Y152_SLICE_X9Y152_BQ),
.O5(CLBLM_L_X8Y151_SLICE_X10Y151_CO5),
.O6(CLBLM_L_X8Y151_SLICE_X10Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcacac0c0fff00f00)
  ) CLBLM_L_X8Y151_SLICE_X10Y151_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X10Y150_SLICE_X12Y150_AQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLL_L_X4Y148_SLICE_X5Y148_CQ),
.I4(CLBLM_L_X8Y151_SLICE_X10Y151_BQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y151_SLICE_X10Y151_BO5),
.O6(CLBLM_L_X8Y151_SLICE_X10Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haafcaafcaafcaa00)
  ) CLBLM_L_X8Y151_SLICE_X10Y151_ALUT (
.I0(CLBLM_L_X8Y151_SLICE_X10Y151_B5Q),
.I1(CLBLM_L_X10Y151_SLICE_X12Y151_CQ),
.I2(CLBLM_L_X8Y151_SLICE_X10Y151_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_L_X8Y151_SLICE_X10Y151_AO5),
.O6(CLBLM_L_X8Y151_SLICE_X10Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y151_SLICE_X11Y151_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y151_SLICE_X11Y151_AO6),
.Q(CLBLM_L_X8Y151_SLICE_X11Y151_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y151_SLICE_X11Y151_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y151_SLICE_X11Y151_BO6),
.Q(CLBLM_L_X8Y151_SLICE_X11Y151_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y151_SLICE_X11Y151_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y151_SLICE_X11Y151_CO6),
.Q(CLBLM_L_X8Y151_SLICE_X11Y151_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y151_SLICE_X11Y151_D_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y151_SLICE_X11Y151_DO6),
.Q(CLBLM_L_X8Y151_SLICE_X11Y151_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc00f000f0)
  ) CLBLM_L_X8Y151_SLICE_X11Y151_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X12Y152_SLICE_X16Y152_AQ),
.I2(CLBLM_L_X8Y151_SLICE_X11Y151_DQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y151_SLICE_X11Y151_DO5),
.O6(CLBLM_L_X8Y151_SLICE_X11Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000f0e4f0e4)
  ) CLBLM_L_X8Y151_SLICE_X11Y151_CLUT (
.I0(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.I1(CLBLM_L_X8Y151_SLICE_X11Y151_CQ),
.I2(CLBLM_L_X10Y151_SLICE_X13Y151_DQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_L_X8Y148_SLICE_X11Y148_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y151_SLICE_X11Y151_CO5),
.O6(CLBLM_L_X8Y151_SLICE_X11Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf1f4f0f001040000)
  ) CLBLM_L_X8Y151_SLICE_X11Y151_BLUT (
.I0(CLBLM_R_X5Y152_SLICE_X7Y152_BQ),
.I1(CLBLM_L_X8Y151_SLICE_X11Y151_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X11Y151_SLICE_X14Y151_CO6),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X7Y153_SLICE_X9Y153_A5Q),
.O5(CLBLM_L_X8Y151_SLICE_X11Y151_BO5),
.O6(CLBLM_L_X8Y151_SLICE_X11Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccfff0cccc0000)
  ) CLBLM_L_X8Y151_SLICE_X11Y151_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y145_SLICE_X6Y145_CQ),
.I2(CLBLM_L_X10Y150_SLICE_X12Y150_DQ),
.I3(CLBLM_L_X8Y151_SLICE_X11Y151_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y152_SLICE_X11Y152_BO6),
.O5(CLBLM_L_X8Y151_SLICE_X11Y151_AO5),
.O6(CLBLM_L_X8Y151_SLICE_X11Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y152_SLICE_X10Y152_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y152_SLICE_X10Y152_AO6),
.Q(CLBLM_L_X8Y152_SLICE_X10Y152_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y152_SLICE_X10Y152_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y152_SLICE_X10Y152_BO6),
.Q(CLBLM_L_X8Y152_SLICE_X10Y152_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y152_SLICE_X10Y152_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y152_SLICE_X10Y152_CO6),
.Q(CLBLM_L_X8Y152_SLICE_X10Y152_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y152_SLICE_X10Y152_D_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y152_SLICE_X10Y152_DO6),
.Q(CLBLM_L_X8Y152_SLICE_X10Y152_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0b1e4b1e4)
  ) CLBLM_L_X8Y152_SLICE_X10Y152_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y152_SLICE_X12Y152_CO5),
.I2(CLBLM_R_X7Y152_SLICE_X9Y152_AQ),
.I3(CLBLM_L_X8Y150_SLICE_X10Y150_CQ),
.I4(1'b1),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X8Y152_SLICE_X10Y152_DO5),
.O6(CLBLM_L_X8Y152_SLICE_X10Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaafcfcfc00)
  ) CLBLM_L_X8Y152_SLICE_X10Y152_CLUT (
.I0(CLBLM_L_X8Y154_SLICE_X10Y154_AQ),
.I1(CLBLM_L_X8Y152_SLICE_X10Y152_CQ),
.I2(CLBLM_L_X8Y150_SLICE_X10Y150_DO6),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y152_SLICE_X10Y152_CO5),
.O6(CLBLM_L_X8Y152_SLICE_X10Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fff000f0ccf000)
  ) CLBLM_L_X8Y152_SLICE_X10Y152_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y152_SLICE_X10Y152_BQ),
.I2(CLBLM_L_X12Y149_SLICE_X17Y149_BQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y152_SLICE_X11Y152_BO6),
.I5(CLBLM_L_X10Y150_SLICE_X12Y150_CQ),
.O5(CLBLM_L_X8Y152_SLICE_X10Y152_BO5),
.O6(CLBLM_L_X8Y152_SLICE_X10Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haafcaafcaa30aa30)
  ) CLBLM_L_X8Y152_SLICE_X10Y152_ALUT (
.I0(CLBLM_L_X10Y153_SLICE_X13Y153_DQ),
.I1(CLBLM_L_X8Y152_SLICE_X11Y152_BO6),
.I2(CLBLM_L_X8Y152_SLICE_X10Y152_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLM_L_X8Y152_SLICE_X10Y152_DQ),
.O5(CLBLM_L_X8Y152_SLICE_X10Y152_AO5),
.O6(CLBLM_L_X8Y152_SLICE_X10Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y152_SLICE_X11Y152_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y152_SLICE_X11Y152_AO6),
.Q(CLBLM_L_X8Y152_SLICE_X11Y152_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y152_SLICE_X11Y152_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y152_SLICE_X11Y152_DO5),
.O6(CLBLM_L_X8Y152_SLICE_X11Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y152_SLICE_X11Y152_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y152_SLICE_X11Y152_CO5),
.O6(CLBLM_L_X8Y152_SLICE_X11Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcff000003000300)
  ) CLBLM_L_X8Y152_SLICE_X11Y152_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y147_SLICE_X15Y147_CQ),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLM_R_X11Y146_SLICE_X14Y146_DQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y152_SLICE_X11Y152_BO5),
.O6(CLBLM_L_X8Y152_SLICE_X11Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888bb8888bb)
  ) CLBLM_L_X8Y152_SLICE_X11Y152_ALUT (
.I0(CLBLM_L_X8Y153_SLICE_X10Y153_BQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(1'b1),
.I3(CLBLM_R_X7Y149_SLICE_X8Y149_BQ),
.I4(CLBLM_L_X10Y149_SLICE_X13Y149_CO5),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X8Y152_SLICE_X11Y152_AO5),
.O6(CLBLM_L_X8Y152_SLICE_X11Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y153_SLICE_X10Y153_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y153_SLICE_X10Y153_AO6),
.Q(CLBLM_L_X8Y153_SLICE_X10Y153_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y153_SLICE_X10Y153_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y153_SLICE_X10Y153_BO6),
.Q(CLBLM_L_X8Y153_SLICE_X10Y153_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00fe0000abab)
  ) CLBLM_L_X8Y153_SLICE_X10Y153_DLUT (
.I0(CLBLM_R_X7Y155_SLICE_X8Y155_A5Q),
.I1(CLBLL_L_X4Y147_SLICE_X5Y147_B5Q),
.I2(CLBLM_R_X7Y153_SLICE_X8Y153_CQ),
.I3(CLBLM_L_X10Y156_SLICE_X12Y156_CO6),
.I4(CLBLM_R_X7Y154_SLICE_X8Y154_BQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y153_SLICE_X10Y153_DO5),
.O6(CLBLM_L_X8Y153_SLICE_X10Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaa0000cf00cf)
  ) CLBLM_L_X8Y153_SLICE_X10Y153_CLUT (
.I0(CLBLM_L_X8Y153_SLICE_X11Y153_AQ),
.I1(CLBLM_L_X8Y154_SLICE_X10Y154_BO5),
.I2(CLBLM_L_X10Y156_SLICE_X12Y156_CO6),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y150_SLICE_X12Y150_B5Q),
.I5(1'b1),
.O5(CLBLM_L_X8Y153_SLICE_X10Y153_CO5),
.O6(CLBLM_L_X8Y153_SLICE_X10Y153_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa00f0ccf0)
  ) CLBLM_L_X8Y153_SLICE_X10Y153_BLUT (
.I0(CLBLM_R_X5Y153_SLICE_X7Y153_BQ),
.I1(CLBLM_L_X8Y153_SLICE_X10Y153_BQ),
.I2(CLBLM_L_X10Y153_SLICE_X13Y153_AQ),
.I3(CLBLM_R_X5Y155_SLICE_X7Y155_CO6),
.I4(CLBLM_R_X7Y155_SLICE_X8Y155_BO5),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y153_SLICE_X10Y153_BO5),
.O6(CLBLM_L_X8Y153_SLICE_X10Y153_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaeefaee00445044)
  ) CLBLM_L_X8Y153_SLICE_X10Y153_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y153_SLICE_X10Y153_BQ),
.I2(CLBLM_L_X8Y153_SLICE_X10Y153_AQ),
.I3(CLBLM_R_X5Y155_SLICE_X7Y155_CO6),
.I4(CLBLM_R_X7Y155_SLICE_X8Y155_BO5),
.I5(CLBLM_L_X10Y146_SLICE_X13Y146_BQ),
.O5(CLBLM_L_X8Y153_SLICE_X10Y153_AO5),
.O6(CLBLM_L_X8Y153_SLICE_X10Y153_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y153_SLICE_X11Y153_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y153_SLICE_X11Y153_AO6),
.Q(CLBLM_L_X8Y153_SLICE_X11Y153_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y153_SLICE_X11Y153_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y153_SLICE_X11Y153_BO6),
.Q(CLBLM_L_X8Y153_SLICE_X11Y153_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y153_SLICE_X11Y153_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y153_SLICE_X11Y153_CO6),
.Q(CLBLM_L_X8Y153_SLICE_X11Y153_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y153_SLICE_X11Y153_D_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y153_SLICE_X11Y153_DO6),
.Q(CLBLM_L_X8Y153_SLICE_X11Y153_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0aa22aa00)
  ) CLBLM_L_X8Y153_SLICE_X11Y153_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(RIOB33_X105Y121_IOB_X1Y121_I),
.I2(CLBLM_R_X7Y153_SLICE_X9Y153_AQ),
.I3(CLBLM_L_X8Y153_SLICE_X11Y153_DQ),
.I4(CLBLM_R_X11Y146_SLICE_X14Y146_DQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y153_SLICE_X11Y153_DO5),
.O6(CLBLM_L_X8Y153_SLICE_X11Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8200ff008282ffff)
  ) CLBLM_L_X8Y153_SLICE_X11Y153_CLUT (
.I0(CLBLM_L_X8Y153_SLICE_X10Y153_DO6),
.I1(CLBLM_L_X8Y153_SLICE_X11Y153_CQ),
.I2(CLBLM_L_X8Y154_SLICE_X11Y154_CO6),
.I3(CLBLM_R_X7Y154_SLICE_X8Y154_CQ),
.I4(CLBLM_L_X8Y153_SLICE_X10Y153_CO5),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y153_SLICE_X11Y153_CO5),
.O6(CLBLM_L_X8Y153_SLICE_X11Y153_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5f0f13035f0f1303)
  ) CLBLM_L_X8Y153_SLICE_X11Y153_BLUT (
.I0(CLBLM_L_X8Y154_SLICE_X10Y154_DO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X8Y153_SLICE_X10Y153_CO5),
.I3(CLBLM_L_X8Y153_SLICE_X10Y153_DO6),
.I4(CLBLM_R_X5Y145_SLICE_X7Y145_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y153_SLICE_X11Y153_BO5),
.O6(CLBLM_L_X8Y153_SLICE_X11Y153_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00bb0000bbbbbbbb)
  ) CLBLM_L_X8Y153_SLICE_X11Y153_ALUT (
.I0(CLBLM_R_X3Y147_SLICE_X2Y147_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(1'b1),
.I3(CLBLM_L_X8Y154_SLICE_X11Y154_BO6),
.I4(CLBLM_L_X8Y153_SLICE_X10Y153_DO6),
.I5(CLBLM_L_X8Y153_SLICE_X10Y153_CO5),
.O5(CLBLM_L_X8Y153_SLICE_X11Y153_AO5),
.O6(CLBLM_L_X8Y153_SLICE_X11Y153_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y154_SLICE_X10Y154_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y154_SLICE_X10Y154_AO6),
.Q(CLBLM_L_X8Y154_SLICE_X10Y154_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa5955aaaa5955)
  ) CLBLM_L_X8Y154_SLICE_X10Y154_DLUT (
.I0(CLBLM_L_X8Y153_SLICE_X11Y153_BQ),
.I1(CLBLM_L_X10Y154_SLICE_X12Y154_CQ),
.I2(CLBLM_L_X8Y154_SLICE_X11Y154_DO6),
.I3(CLBLM_L_X8Y154_SLICE_X10Y154_CO6),
.I4(CLBLM_L_X8Y155_SLICE_X10Y155_CO6),
.I5(1'b1),
.O5(CLBLM_L_X8Y154_SLICE_X10Y154_DO5),
.O6(CLBLM_L_X8Y154_SLICE_X10Y154_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0008888811100000)
  ) CLBLM_L_X8Y154_SLICE_X10Y154_CLUT (
.I0(CLBLM_L_X8Y153_SLICE_X11Y153_AQ),
.I1(CLBLM_L_X8Y153_SLICE_X11Y153_CQ),
.I2(CLBLM_R_X7Y154_SLICE_X8Y154_BQ),
.I3(CLBLL_L_X4Y147_SLICE_X5Y147_B5Q),
.I4(CLBLM_R_X7Y153_SLICE_X8Y153_CQ),
.I5(CLBLM_L_X8Y155_SLICE_X10Y155_BQ),
.O5(CLBLM_L_X8Y154_SLICE_X10Y154_CO5),
.O6(CLBLM_L_X8Y154_SLICE_X10Y154_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8caf333350dc33cf)
  ) CLBLM_L_X8Y154_SLICE_X10Y154_BLUT (
.I0(CLBLM_R_X7Y155_SLICE_X8Y155_AQ),
.I1(CLBLM_R_X7Y153_SLICE_X8Y153_CQ),
.I2(CLBLM_R_X7Y155_SLICE_X8Y155_A5Q),
.I3(CLBLL_L_X4Y147_SLICE_X5Y147_B5Q),
.I4(CLBLM_R_X7Y154_SLICE_X8Y154_BQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y154_SLICE_X10Y154_BO5),
.O6(CLBLM_L_X8Y154_SLICE_X10Y154_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00aaf0aaf0)
  ) CLBLM_L_X8Y154_SLICE_X10Y154_ALUT (
.I0(CLBLM_L_X10Y154_SLICE_X12Y154_CQ),
.I1(1'b1),
.I2(CLBLM_R_X5Y150_SLICE_X7Y150_BQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X8Y154_SLICE_X10Y154_AO5),
.O6(CLBLM_L_X8Y154_SLICE_X10Y154_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f1f0fff0f1f0fff)
  ) CLBLM_L_X8Y154_SLICE_X11Y154_DLUT (
.I0(CLBLM_R_X7Y153_SLICE_X8Y153_CQ),
.I1(CLBLL_L_X4Y147_SLICE_X5Y147_B5Q),
.I2(CLBLM_R_X5Y155_SLICE_X7Y155_BO5),
.I3(CLBLM_L_X8Y154_SLICE_X11Y154_AO5),
.I4(CLBLM_R_X7Y153_SLICE_X9Y153_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y154_SLICE_X11Y154_DO5),
.O6(CLBLM_L_X8Y154_SLICE_X11Y154_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0b0f0f0f0f07)
  ) CLBLM_L_X8Y154_SLICE_X11Y154_CLUT (
.I0(CLBLM_L_X8Y154_SLICE_X11Y154_AO6),
.I1(CLBLM_R_X7Y154_SLICE_X8Y154_AQ),
.I2(CLBLM_L_X8Y155_SLICE_X10Y155_CO6),
.I3(CLBLM_L_X8Y153_SLICE_X11Y153_AQ),
.I4(CLBLM_L_X8Y154_SLICE_X11Y154_DO6),
.I5(CLBLM_L_X8Y155_SLICE_X10Y155_BQ),
.O5(CLBLM_L_X8Y154_SLICE_X11Y154_CO5),
.O6(CLBLM_L_X8Y154_SLICE_X11Y154_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f00f4b4b0f)
  ) CLBLM_L_X8Y154_SLICE_X11Y154_BLUT (
.I0(CLBLM_L_X8Y154_SLICE_X11Y154_DO6),
.I1(CLBLM_R_X7Y153_SLICE_X8Y153_BQ),
.I2(CLBLM_L_X8Y153_SLICE_X11Y153_AQ),
.I3(CLBLM_L_X8Y155_SLICE_X10Y155_BQ),
.I4(CLBLM_L_X8Y154_SLICE_X11Y154_AO6),
.I5(CLBLM_L_X8Y155_SLICE_X10Y155_CO6),
.O5(CLBLM_L_X8Y154_SLICE_X11Y154_BO5),
.O6(CLBLM_L_X8Y154_SLICE_X11Y154_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccc0c055000000)
  ) CLBLM_L_X8Y154_SLICE_X11Y154_ALUT (
.I0(CLBLM_R_X7Y155_SLICE_X8Y155_AQ),
.I1(CLBLM_R_X7Y153_SLICE_X8Y153_CQ),
.I2(CLBLL_L_X4Y147_SLICE_X5Y147_B5Q),
.I3(CLBLM_R_X7Y155_SLICE_X8Y155_A5Q),
.I4(CLBLM_R_X7Y154_SLICE_X8Y154_BQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y154_SLICE_X11Y154_AO5),
.O6(CLBLM_L_X8Y154_SLICE_X11Y154_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y155_SLICE_X10Y155_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y155_SLICE_X10Y155_AO6),
.Q(CLBLM_L_X8Y155_SLICE_X10Y155_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y155_SLICE_X10Y155_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y155_SLICE_X10Y155_BO6),
.Q(CLBLM_L_X8Y155_SLICE_X10Y155_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha5f0a5a5a5f0a5a5)
  ) CLBLM_L_X8Y155_SLICE_X10Y155_DLUT (
.I0(CLBLM_L_X8Y155_SLICE_X10Y155_CO6),
.I1(1'b1),
.I2(CLBLM_L_X8Y155_SLICE_X10Y155_BQ),
.I3(CLBLM_L_X8Y154_SLICE_X11Y154_DO6),
.I4(CLBLM_R_X7Y155_SLICE_X9Y155_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y155_SLICE_X10Y155_DO5),
.O6(CLBLM_L_X8Y155_SLICE_X10Y155_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h33333333fffffbff)
  ) CLBLM_L_X8Y155_SLICE_X10Y155_CLUT (
.I0(CLBLL_L_X4Y147_SLICE_X5Y147_B5Q),
.I1(CLBLM_R_X5Y155_SLICE_X7Y155_BO5),
.I2(CLBLM_R_X7Y153_SLICE_X8Y153_CQ),
.I3(CLBLM_R_X7Y154_SLICE_X8Y154_BQ),
.I4(CLBLM_R_X7Y155_SLICE_X8Y155_A5Q),
.I5(CLBLM_R_X7Y155_SLICE_X8Y155_AQ),
.O5(CLBLM_L_X8Y155_SLICE_X10Y155_CO5),
.O6(CLBLM_L_X8Y155_SLICE_X10Y155_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h4c4c5f5f0c0c0f0f)
  ) CLBLM_L_X8Y155_SLICE_X10Y155_BLUT (
.I0(CLBLM_L_X8Y155_SLICE_X10Y155_DO6),
.I1(CLBLM_L_X8Y151_SLICE_X10Y151_DQ),
.I2(CLBLM_L_X8Y153_SLICE_X10Y153_CO5),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y153_SLICE_X10Y153_DO6),
.O5(CLBLM_L_X8Y155_SLICE_X10Y155_BO5),
.O6(CLBLM_L_X8Y155_SLICE_X10Y155_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hb00bbbbb0000bbbb)
  ) CLBLM_L_X8Y155_SLICE_X10Y155_ALUT (
.I0(CLBLM_R_X5Y152_SLICE_X7Y152_BQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X8Y155_SLICE_X11Y155_AO6),
.I3(CLBLM_L_X8Y155_SLICE_X10Y155_AQ),
.I4(CLBLM_L_X8Y153_SLICE_X10Y153_CO5),
.I5(CLBLM_L_X8Y153_SLICE_X10Y153_DO6),
.O5(CLBLM_L_X8Y155_SLICE_X10Y155_AO5),
.O6(CLBLM_L_X8Y155_SLICE_X10Y155_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000010100000000)
  ) CLBLM_L_X8Y155_SLICE_X11Y155_DLUT (
.I0(CLBLM_L_X8Y153_SLICE_X11Y153_CQ),
.I1(CLBLM_L_X8Y155_SLICE_X10Y155_BQ),
.I2(CLBLM_L_X8Y153_SLICE_X11Y153_BQ),
.I3(1'b1),
.I4(CLBLM_L_X8Y153_SLICE_X11Y153_AQ),
.I5(CLBLM_L_X8Y154_SLICE_X11Y154_AO6),
.O5(CLBLM_L_X8Y155_SLICE_X11Y155_DO5),
.O6(CLBLM_L_X8Y155_SLICE_X11Y155_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0a0000002a000000)
  ) CLBLM_L_X8Y155_SLICE_X11Y155_CLUT (
.I0(CLBLM_L_X8Y153_SLICE_X11Y153_CQ),
.I1(CLBLM_R_X7Y154_SLICE_X8Y154_BQ),
.I2(CLBLM_R_X7Y153_SLICE_X8Y153_CQ),
.I3(CLBLM_L_X8Y153_SLICE_X11Y153_AQ),
.I4(CLBLM_L_X8Y155_SLICE_X10Y155_BQ),
.I5(CLBLL_L_X4Y147_SLICE_X5Y147_B5Q),
.O5(CLBLM_L_X8Y155_SLICE_X11Y155_CO5),
.O6(CLBLM_L_X8Y155_SLICE_X11Y155_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h2000000000000000)
  ) CLBLM_L_X8Y155_SLICE_X11Y155_BLUT (
.I0(CLBLM_L_X8Y155_SLICE_X10Y155_BQ),
.I1(CLBLM_L_X8Y154_SLICE_X11Y154_AO6),
.I2(CLBLM_L_X8Y153_SLICE_X11Y153_AQ),
.I3(CLBLM_L_X10Y154_SLICE_X12Y154_DQ),
.I4(CLBLM_L_X8Y153_SLICE_X11Y153_BQ),
.I5(CLBLM_L_X8Y153_SLICE_X11Y153_CQ),
.O5(CLBLM_L_X8Y155_SLICE_X11Y155_BO5),
.O6(CLBLM_L_X8Y155_SLICE_X11Y155_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0f000d0f0f)
  ) CLBLM_L_X8Y155_SLICE_X11Y155_ALUT (
.I0(CLBLM_L_X8Y155_SLICE_X11Y155_DO6),
.I1(CLBLM_L_X10Y154_SLICE_X12Y154_DQ),
.I2(CLBLM_L_X8Y155_SLICE_X10Y155_CO6),
.I3(CLBLM_L_X8Y155_SLICE_X11Y155_BO6),
.I4(CLBLM_L_X10Y154_SLICE_X12Y154_BQ),
.I5(CLBLM_L_X8Y154_SLICE_X11Y154_DO6),
.O5(CLBLM_L_X8Y155_SLICE_X11Y155_AO5),
.O6(CLBLM_L_X8Y155_SLICE_X11Y155_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y159_SLICE_X10Y159_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y159_SLICE_X10Y159_DO5),
.O6(CLBLM_L_X8Y159_SLICE_X10Y159_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y159_SLICE_X10Y159_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y159_SLICE_X10Y159_CO5),
.O6(CLBLM_L_X8Y159_SLICE_X10Y159_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y159_SLICE_X10Y159_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y159_SLICE_X10Y159_BO5),
.O6(CLBLM_L_X8Y159_SLICE_X10Y159_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555555555555555)
  ) CLBLM_L_X8Y159_SLICE_X10Y159_ALUT (
.I0(CLBLM_L_X8Y151_SLICE_X10Y151_B5Q),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y159_SLICE_X10Y159_AO5),
.O6(CLBLM_L_X8Y159_SLICE_X10Y159_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y159_SLICE_X11Y159_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y159_SLICE_X11Y159_DO5),
.O6(CLBLM_L_X8Y159_SLICE_X11Y159_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y159_SLICE_X11Y159_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y159_SLICE_X11Y159_CO5),
.O6(CLBLM_L_X8Y159_SLICE_X11Y159_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y159_SLICE_X11Y159_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y159_SLICE_X11Y159_BO5),
.O6(CLBLM_L_X8Y159_SLICE_X11Y159_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y159_SLICE_X11Y159_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y159_SLICE_X11Y159_AO5),
.O6(CLBLM_L_X8Y159_SLICE_X11Y159_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333333336333633)
  ) CLBLM_L_X10Y141_SLICE_X12Y141_DLUT (
.I0(CLBLM_L_X12Y144_SLICE_X16Y144_BQ),
.I1(CLBLM_R_X7Y142_SLICE_X8Y142_CQ),
.I2(CLBLM_L_X12Y144_SLICE_X16Y144_CQ),
.I3(CLBLM_L_X12Y144_SLICE_X16Y144_AQ),
.I4(1'b1),
.I5(CLBLM_L_X12Y145_SLICE_X16Y145_AQ),
.O5(CLBLM_L_X10Y141_SLICE_X12Y141_DO5),
.O6(CLBLM_L_X10Y141_SLICE_X12Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000cfff3000)
  ) CLBLM_L_X10Y141_SLICE_X12Y141_CLUT (
.I0(1'b1),
.I1(CLBLM_L_X12Y144_SLICE_X16Y144_CQ),
.I2(CLBLM_L_X12Y144_SLICE_X16Y144_BQ),
.I3(CLBLM_L_X12Y144_SLICE_X16Y144_AQ),
.I4(CLBLM_R_X11Y146_SLICE_X15Y146_AQ),
.I5(CLBLM_L_X12Y145_SLICE_X16Y145_AQ),
.O5(CLBLM_L_X10Y141_SLICE_X12Y141_CO5),
.O6(CLBLM_L_X10Y141_SLICE_X12Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ffffcc9ccccc)
  ) CLBLM_L_X10Y141_SLICE_X12Y141_BLUT (
.I0(CLBLM_L_X12Y144_SLICE_X16Y144_AQ),
.I1(CLBLM_R_X7Y142_SLICE_X8Y142_BQ),
.I2(CLBLM_L_X12Y144_SLICE_X16Y144_CQ),
.I3(CLBLM_L_X12Y145_SLICE_X16Y145_AQ),
.I4(CLBLM_L_X12Y144_SLICE_X16Y144_BQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y141_SLICE_X12Y141_BO5),
.O6(CLBLM_L_X10Y141_SLICE_X12Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaa9accffccff)
  ) CLBLM_L_X10Y141_SLICE_X12Y141_ALUT (
.I0(CLBLM_R_X7Y144_SLICE_X8Y144_DQ),
.I1(CLBLM_L_X12Y145_SLICE_X16Y145_AQ),
.I2(CLBLM_L_X12Y144_SLICE_X16Y144_CQ),
.I3(CLBLM_L_X12Y144_SLICE_X16Y144_AQ),
.I4(CLBLM_L_X12Y144_SLICE_X16Y144_BQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y141_SLICE_X12Y141_AO5),
.O6(CLBLM_L_X10Y141_SLICE_X12Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y141_SLICE_X13Y141_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y141_SLICE_X13Y141_DO5),
.O6(CLBLM_L_X10Y141_SLICE_X13Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y141_SLICE_X13Y141_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y141_SLICE_X13Y141_CO5),
.O6(CLBLM_L_X10Y141_SLICE_X13Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y141_SLICE_X13Y141_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y141_SLICE_X13Y141_BO5),
.O6(CLBLM_L_X10Y141_SLICE_X13Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y141_SLICE_X13Y141_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y141_SLICE_X13Y141_AO5),
.O6(CLBLM_L_X10Y141_SLICE_X13Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hef01fe1001ef10fe)
  ) CLBLM_L_X10Y142_SLICE_X12Y142_DLUT (
.I0(CLBLM_R_X5Y144_SLICE_X6Y144_DO6),
.I1(CLBLM_R_X3Y151_SLICE_X2Y151_AO6),
.I2(CLBLM_L_X10Y142_SLICE_X13Y142_BO5),
.I3(CLBLM_L_X10Y145_SLICE_X13Y145_A5Q),
.I4(CLBLM_L_X10Y141_SLICE_X12Y141_DO6),
.I5(CLBLM_L_X8Y148_SLICE_X10Y148_BQ),
.O5(CLBLM_L_X10Y142_SLICE_X12Y142_DO5),
.O6(CLBLM_L_X10Y142_SLICE_X12Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaa5500ffae5100)
  ) CLBLM_L_X10Y142_SLICE_X12Y142_CLUT (
.I0(CLBLM_R_X5Y144_SLICE_X6Y144_DO6),
.I1(CLBLM_R_X5Y143_SLICE_X7Y143_BO6),
.I2(CLBLM_R_X5Y145_SLICE_X6Y145_DO6),
.I3(CLBLM_L_X10Y141_SLICE_X12Y141_CO6),
.I4(CLBLM_R_X5Y144_SLICE_X7Y144_B5Q),
.I5(CLBLM_R_X7Y142_SLICE_X9Y142_AO6),
.O5(CLBLM_L_X10Y142_SLICE_X12Y142_CO5),
.O6(CLBLM_L_X10Y142_SLICE_X12Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_L_X10Y142_SLICE_X12Y142_BLUT (
.I0(CLBLM_L_X10Y142_SLICE_X12Y142_DO6),
.I1(CLBLM_L_X10Y142_SLICE_X13Y142_DO6),
.I2(CLBLM_L_X10Y142_SLICE_X13Y142_CO6),
.I3(CLBLM_L_X10Y143_SLICE_X13Y143_DO6),
.I4(CLBLM_L_X10Y142_SLICE_X12Y142_AO6),
.I5(CLBLM_L_X10Y142_SLICE_X12Y142_CO6),
.O5(CLBLM_L_X10Y142_SLICE_X12Y142_BO5),
.O6(CLBLM_L_X10Y142_SLICE_X12Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h33330f1b33330f0f)
  ) CLBLM_L_X10Y142_SLICE_X12Y142_ALUT (
.I0(CLBLM_R_X5Y145_SLICE_X6Y145_DO6),
.I1(CLBLM_R_X15Y151_SLICE_X20Y151_AQ),
.I2(CLBLM_L_X10Y141_SLICE_X12Y141_BO5),
.I3(CLBLM_R_X7Y142_SLICE_X9Y142_AO6),
.I4(CLBLM_R_X5Y144_SLICE_X6Y144_DO6),
.I5(CLBLM_R_X5Y143_SLICE_X7Y143_BO6),
.O5(CLBLM_L_X10Y142_SLICE_X12Y142_AO5),
.O6(CLBLM_L_X10Y142_SLICE_X12Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y142_SLICE_X13Y142_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y142_SLICE_X13Y142_AO6),
.Q(CLBLM_L_X10Y142_SLICE_X13Y142_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haab85574aa8b5547)
  ) CLBLM_L_X10Y142_SLICE_X13Y142_DLUT (
.I0(CLBLM_L_X10Y145_SLICE_X12Y145_C5Q),
.I1(CLBLM_R_X5Y144_SLICE_X6Y144_DO6),
.I2(CLBLM_L_X10Y143_SLICE_X13Y143_CO6),
.I3(CLBLM_R_X3Y151_SLICE_X2Y151_AO6),
.I4(CLBLM_R_X3Y145_SLICE_X3Y145_DQ),
.I5(CLBLM_L_X10Y141_SLICE_X12Y141_AO6),
.O5(CLBLM_L_X10Y142_SLICE_X13Y142_DO5),
.O6(CLBLM_L_X10Y142_SLICE_X13Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaa00aafbaa08)
  ) CLBLM_L_X10Y142_SLICE_X13Y142_CLUT (
.I0(CLBLM_L_X8Y145_SLICE_X11Y145_BQ),
.I1(CLBLM_R_X5Y143_SLICE_X7Y143_BO6),
.I2(CLBLM_R_X5Y145_SLICE_X6Y145_DO6),
.I3(CLBLM_R_X5Y144_SLICE_X6Y144_DO6),
.I4(CLBLM_R_X11Y143_SLICE_X14Y143_CO6),
.I5(CLBLM_R_X7Y142_SLICE_X9Y142_AO6),
.O5(CLBLM_L_X10Y142_SLICE_X13Y142_CO5),
.O6(CLBLM_L_X10Y142_SLICE_X13Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffff3f3aaaaa6aa)
  ) CLBLM_L_X10Y142_SLICE_X13Y142_BLUT (
.I0(CLBLM_L_X10Y143_SLICE_X13Y143_BQ),
.I1(CLBLM_L_X12Y145_SLICE_X16Y145_AQ),
.I2(CLBLM_L_X12Y144_SLICE_X16Y144_BQ),
.I3(CLBLM_L_X12Y144_SLICE_X16Y144_CQ),
.I4(CLBLM_L_X12Y144_SLICE_X16Y144_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y142_SLICE_X13Y142_BO5),
.O6(CLBLM_L_X10Y142_SLICE_X13Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000030303030)
  ) CLBLM_L_X10Y142_SLICE_X13Y142_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_L_X10Y142_SLICE_X13Y142_AQ),
.I3(1'b1),
.I4(CLBLM_L_X10Y145_SLICE_X12Y145_C5Q),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y142_SLICE_X13Y142_AO5),
.O6(CLBLM_L_X10Y142_SLICE_X13Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3c3cffffffff3c3c)
  ) CLBLM_L_X10Y143_SLICE_X12Y143_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y144_SLICE_X12Y144_BQ),
.I2(CLBLM_R_X5Y144_SLICE_X7Y144_B5Q),
.I3(1'b1),
.I4(CLBLM_R_X11Y148_SLICE_X15Y148_A5Q),
.I5(CLBLM_L_X8Y144_SLICE_X10Y144_BQ),
.O5(CLBLM_L_X10Y143_SLICE_X12Y143_DO5),
.O6(CLBLM_L_X10Y143_SLICE_X12Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff6f6ffffff6f6)
  ) CLBLM_L_X10Y143_SLICE_X12Y143_CLUT (
.I0(CLBLM_L_X10Y145_SLICE_X12Y145_C5Q),
.I1(CLBLM_L_X10Y145_SLICE_X12Y145_DQ),
.I2(CLBLM_L_X8Y144_SLICE_X11Y144_AQ),
.I3(1'b1),
.I4(CLBLM_L_X10Y143_SLICE_X12Y143_DO6),
.I5(CLBLM_L_X8Y145_SLICE_X11Y145_BQ),
.O5(CLBLM_L_X10Y143_SLICE_X12Y143_CO5),
.O6(CLBLM_L_X10Y143_SLICE_X12Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000f5500003c55)
  ) CLBLM_L_X10Y143_SLICE_X12Y143_BLUT (
.I0(CLBLM_R_X5Y144_SLICE_X7Y144_B5Q),
.I1(CLBLM_L_X10Y141_SLICE_X12Y141_BO6),
.I2(CLBLM_R_X11Y146_SLICE_X15Y146_AQ),
.I3(CLBLM_R_X7Y142_SLICE_X8Y142_DO6),
.I4(CLBLM_L_X10Y143_SLICE_X13Y143_AQ),
.I5(CLBLM_L_X10Y141_SLICE_X12Y141_AO5),
.O5(CLBLM_L_X10Y143_SLICE_X12Y143_BO5),
.O6(CLBLM_L_X10Y143_SLICE_X12Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h000011d10000dd1d)
  ) CLBLM_L_X10Y143_SLICE_X12Y143_ALUT (
.I0(CLBLM_R_X7Y145_SLICE_X9Y145_CQ),
.I1(CLBLM_R_X7Y142_SLICE_X8Y142_DO6),
.I2(CLBLM_L_X10Y143_SLICE_X13Y143_CO5),
.I3(CLBLM_L_X10Y141_SLICE_X12Y141_BO6),
.I4(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.I5(CLBLM_L_X10Y145_SLICE_X13Y145_CQ),
.O5(CLBLM_L_X10Y143_SLICE_X12Y143_AO5),
.O6(CLBLM_L_X10Y143_SLICE_X12Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y143_SLICE_X13Y143_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y143_SLICE_X13Y143_AO6),
.Q(CLBLM_L_X10Y143_SLICE_X13Y143_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y143_SLICE_X13Y143_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y143_SLICE_X13Y143_BO6),
.Q(CLBLM_L_X10Y143_SLICE_X13Y143_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0ff0f00f99f099)
  ) CLBLM_L_X10Y143_SLICE_X13Y143_DLUT (
.I0(CLBLM_R_X11Y144_SLICE_X15Y144_AO6),
.I1(CLBLM_R_X11Y144_SLICE_X15Y144_CO6),
.I2(CLBLM_R_X11Y148_SLICE_X15Y148_A5Q),
.I3(CLBLM_R_X5Y144_SLICE_X6Y144_DO6),
.I4(CLBLM_R_X7Y145_SLICE_X9Y145_CQ),
.I5(CLBLM_R_X3Y151_SLICE_X2Y151_AO6),
.O5(CLBLM_L_X10Y143_SLICE_X13Y143_DO5),
.O6(CLBLM_L_X10Y143_SLICE_X13Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h9ccccccc00aa00aa)
  ) CLBLM_L_X10Y143_SLICE_X13Y143_CLUT (
.I0(CLBLM_L_X12Y145_SLICE_X16Y145_AQ),
.I1(CLBLM_L_X10Y148_SLICE_X12Y148_BQ),
.I2(CLBLM_L_X12Y144_SLICE_X16Y144_CQ),
.I3(CLBLM_L_X12Y144_SLICE_X16Y144_AQ),
.I4(CLBLM_L_X12Y144_SLICE_X16Y144_BQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y143_SLICE_X13Y143_CO5),
.O6(CLBLM_L_X10Y143_SLICE_X13Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000ee00ee00)
  ) CLBLM_L_X10Y143_SLICE_X13Y143_BLUT (
.I0(CLBLM_L_X10Y145_SLICE_X13Y145_CQ),
.I1(CLBLM_L_X10Y143_SLICE_X13Y143_BQ),
.I2(1'b1),
.I3(CLBLM_R_X7Y142_SLICE_X8Y142_DO6),
.I4(CLBLM_R_X7Y143_SLICE_X9Y143_CQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y143_SLICE_X13Y143_BO5),
.O6(CLBLM_L_X10Y143_SLICE_X13Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbabbbabb10111011)
  ) CLBLM_L_X10Y143_SLICE_X13Y143_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y143_SLICE_X12Y143_BO6),
.I2(CLBLM_R_X5Y142_SLICE_X7Y142_AQ),
.I3(RIOB33_X105Y141_IOB_X1Y142_I),
.I4(1'b1),
.I5(CLBLM_L_X8Y148_SLICE_X10Y148_A5Q),
.O5(CLBLM_L_X10Y143_SLICE_X13Y143_AO5),
.O6(CLBLM_L_X10Y143_SLICE_X13Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y144_SLICE_X12Y144_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y144_SLICE_X12Y144_AO6),
.Q(CLBLM_L_X10Y144_SLICE_X12Y144_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y144_SLICE_X12Y144_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y144_SLICE_X12Y144_BO6),
.Q(CLBLM_L_X10Y144_SLICE_X12Y144_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y144_SLICE_X12Y144_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y144_SLICE_X12Y144_CO6),
.Q(CLBLM_L_X10Y144_SLICE_X12Y144_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0033003300330063)
  ) CLBLM_L_X10Y144_SLICE_X12Y144_DLUT (
.I0(CLBLM_L_X12Y145_SLICE_X16Y145_AQ),
.I1(CLBLM_R_X11Y144_SLICE_X15Y144_DO6),
.I2(CLBLM_L_X12Y144_SLICE_X16Y144_BQ),
.I3(CLBLM_L_X10Y146_SLICE_X12Y146_CQ),
.I4(CLBLM_L_X12Y144_SLICE_X16Y144_CQ),
.I5(CLBLM_L_X12Y144_SLICE_X16Y144_AQ),
.O5(CLBLM_L_X10Y144_SLICE_X12Y144_DO5),
.O6(CLBLM_L_X10Y144_SLICE_X12Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfef0fef0fff0fcf0)
  ) CLBLM_L_X10Y144_SLICE_X12Y144_CLUT (
.I0(CLBLM_R_X7Y144_SLICE_X9Y144_DO5),
.I1(CLBLM_L_X10Y144_SLICE_X12Y144_CQ),
.I2(CLBLM_R_X5Y146_SLICE_X6Y146_BO5),
.I3(CLBLM_R_X11Y151_SLICE_X15Y151_CO6),
.I4(CLBLM_L_X8Y144_SLICE_X11Y144_DO6),
.I5(CLBLM_L_X10Y142_SLICE_X12Y142_BO6),
.O5(CLBLM_L_X10Y144_SLICE_X12Y144_CO5),
.O6(CLBLM_L_X10Y144_SLICE_X12Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaafc00fc00)
  ) CLBLM_L_X10Y144_SLICE_X12Y144_BLUT (
.I0(CLBLM_R_X5Y144_SLICE_X7Y144_AQ),
.I1(CLBLM_L_X10Y144_SLICE_X12Y144_BQ),
.I2(CLBLM_R_X5Y143_SLICE_X7Y143_AQ),
.I3(CLBLM_R_X7Y142_SLICE_X8Y142_DO6),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y144_SLICE_X12Y144_BO5),
.O6(CLBLM_L_X10Y144_SLICE_X12Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heeeeecececeeecee)
  ) CLBLM_L_X10Y144_SLICE_X12Y144_ALUT (
.I0(CLBLM_R_X11Y151_SLICE_X15Y151_CO6),
.I1(CLBLM_R_X7Y151_SLICE_X8Y151_CO5),
.I2(CLBLM_L_X10Y144_SLICE_X12Y144_AQ),
.I3(CLBLM_L_X10Y142_SLICE_X12Y142_BO6),
.I4(CLBLM_R_X7Y144_SLICE_X9Y144_DO5),
.I5(CLBLM_L_X8Y147_SLICE_X11Y147_BO5),
.O5(CLBLM_L_X10Y144_SLICE_X12Y144_AO5),
.O6(CLBLM_L_X10Y144_SLICE_X12Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y144_SLICE_X13Y144_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y144_SLICE_X13Y144_AO6),
.Q(CLBLM_L_X10Y144_SLICE_X13Y144_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y144_SLICE_X13Y144_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y144_SLICE_X13Y144_BO6),
.Q(CLBLM_L_X10Y144_SLICE_X13Y144_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y144_SLICE_X13Y144_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y144_SLICE_X13Y144_CO6),
.Q(CLBLM_L_X10Y144_SLICE_X13Y144_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0c050c0503050305)
  ) CLBLM_L_X10Y144_SLICE_X13Y144_DLUT (
.I0(CLBLM_L_X10Y145_SLICE_X12Y145_C5Q),
.I1(CLBLM_L_X12Y144_SLICE_X16Y144_DO5),
.I2(CLBLM_L_X10Y144_SLICE_X13Y144_BQ),
.I3(CLBLM_R_X7Y142_SLICE_X8Y142_DO6),
.I4(1'b1),
.I5(CLBLM_L_X10Y148_SLICE_X12Y148_BQ),
.O5(CLBLM_L_X10Y144_SLICE_X13Y144_DO5),
.O6(CLBLM_L_X10Y144_SLICE_X13Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0ffc0cf000f000)
  ) CLBLM_L_X10Y144_SLICE_X13Y144_CLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y144_SLICE_X13Y144_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y147_SLICE_X12Y147_A5Q),
.I4(CLBLM_R_X11Y145_SLICE_X15Y145_AQ),
.I5(CLBLM_R_X7Y142_SLICE_X8Y142_DO6),
.O5(CLBLM_L_X10Y144_SLICE_X13Y144_CO5),
.O6(CLBLM_L_X10Y144_SLICE_X13Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0051515151)
  ) CLBLM_L_X10Y144_SLICE_X13Y144_BLUT (
.I0(CLBLM_L_X10Y144_SLICE_X13Y144_DO6),
.I1(RIOB33_X105Y141_IOB_X1Y142_I),
.I2(CLBLM_R_X5Y142_SLICE_X7Y142_AQ),
.I3(CLBLM_L_X10Y145_SLICE_X12Y145_CQ),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y144_SLICE_X13Y144_BO5),
.O6(CLBLM_L_X10Y144_SLICE_X13Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000000500050)
  ) CLBLM_L_X10Y144_SLICE_X13Y144_ALUT (
.I0(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.I1(1'b1),
.I2(CLBLM_L_X10Y144_SLICE_X13Y144_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_L_X10Y142_SLICE_X13Y142_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y144_SLICE_X13Y144_AO5),
.O6(CLBLM_L_X10Y144_SLICE_X13Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y145_SLICE_X12Y145_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y145_SLICE_X12Y145_CO5),
.Q(CLBLM_L_X10Y145_SLICE_X12Y145_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y145_SLICE_X12Y145_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y145_SLICE_X12Y145_AO6),
.Q(CLBLM_L_X10Y145_SLICE_X12Y145_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y145_SLICE_X12Y145_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y145_SLICE_X12Y145_BO6),
.Q(CLBLM_L_X10Y145_SLICE_X12Y145_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y145_SLICE_X12Y145_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y145_SLICE_X12Y145_CO6),
.Q(CLBLM_L_X10Y145_SLICE_X12Y145_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y145_SLICE_X12Y145_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y145_SLICE_X12Y145_DO6),
.Q(CLBLM_L_X10Y145_SLICE_X12Y145_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffccffc000cc00c0)
  ) CLBLM_L_X10Y145_SLICE_X12Y145_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y142_SLICE_X8Y142_DO6),
.I2(CLBLM_L_X10Y145_SLICE_X12Y145_DQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y144_SLICE_X10Y144_BQ),
.I5(CLBLM_L_X10Y151_SLICE_X13Y151_BQ),
.O5(CLBLM_L_X10Y145_SLICE_X12Y145_DO5),
.O6(CLBLM_L_X10Y145_SLICE_X12Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccf0ccf0aaffaa00)
  ) CLBLM_L_X10Y145_SLICE_X12Y145_CLUT (
.I0(CLBLM_L_X10Y144_SLICE_X13Y144_BQ),
.I1(CLBLM_R_X7Y151_SLICE_X9Y151_CQ),
.I2(CLBLM_L_X10Y149_SLICE_X12Y149_CO6),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y146_SLICE_X12Y146_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X10Y145_SLICE_X12Y145_CO5),
.O6(CLBLM_L_X10Y145_SLICE_X12Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0ffee0044)
  ) CLBLM_L_X10Y145_SLICE_X12Y145_BLUT (
.I0(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.I1(CLBLM_L_X10Y145_SLICE_X12Y145_BQ),
.I2(CLBLM_R_X7Y145_SLICE_X9Y145_BQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_R_X5Y145_SLICE_X7Y145_BQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y145_SLICE_X12Y145_BO5),
.O6(CLBLM_L_X10Y145_SLICE_X12Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffccccfcecfcec)
  ) CLBLM_L_X10Y145_SLICE_X12Y145_ALUT (
.I0(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.I1(CLBLM_L_X8Y145_SLICE_X10Y145_DO6),
.I2(CLBLM_L_X10Y145_SLICE_X12Y145_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_R_X11Y143_SLICE_X14Y143_BQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y145_SLICE_X12Y145_AO5),
.O6(CLBLM_L_X10Y145_SLICE_X12Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y145_SLICE_X13Y145_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y145_SLICE_X13Y145_AO5),
.Q(CLBLM_L_X10Y145_SLICE_X13Y145_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y145_SLICE_X13Y145_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y145_SLICE_X13Y145_AO6),
.Q(CLBLM_L_X10Y145_SLICE_X13Y145_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y145_SLICE_X13Y145_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y145_SLICE_X13Y145_BO6),
.Q(CLBLM_L_X10Y145_SLICE_X13Y145_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y145_SLICE_X13Y145_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y145_SLICE_X13Y145_CO6),
.Q(CLBLM_L_X10Y145_SLICE_X13Y145_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h010d0d0101010d0d)
  ) CLBLM_L_X10Y145_SLICE_X13Y145_DLUT (
.I0(CLBLM_L_X8Y148_SLICE_X10Y148_BQ),
.I1(CLBLM_R_X7Y142_SLICE_X8Y142_DO6),
.I2(CLBLM_R_X11Y146_SLICE_X15Y146_DQ),
.I3(CLBLM_L_X10Y142_SLICE_X13Y142_BO6),
.I4(CLBLM_L_X10Y143_SLICE_X13Y143_BQ),
.I5(CLBLM_L_X12Y144_SLICE_X16Y144_CQ),
.O5(CLBLM_L_X10Y145_SLICE_X13Y145_DO5),
.O6(CLBLM_L_X10Y145_SLICE_X13Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0f5e4a0a0f5e4)
  ) CLBLM_L_X10Y145_SLICE_X13Y145_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y145_SLICE_X13Y145_CQ),
.I2(CLBLM_L_X10Y146_SLICE_X12Y146_A5Q),
.I3(CLBLM_R_X7Y146_SLICE_X9Y146_CQ),
.I4(CLBLL_L_X4Y145_SLICE_X5Y145_DO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y145_SLICE_X13Y145_CO5),
.O6(CLBLM_L_X10Y145_SLICE_X13Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f0ccf000f0cc)
  ) CLBLM_L_X10Y145_SLICE_X13Y145_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y146_SLICE_X13Y146_AQ),
.I2(CLBLM_L_X12Y145_SLICE_X16Y145_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y145_SLICE_X13Y145_BO5),
.O6(CLBLM_L_X10Y145_SLICE_X13Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0ccf0ccffaa00aa)
  ) CLBLM_L_X10Y145_SLICE_X13Y145_ALUT (
.I0(CLBLM_L_X10Y147_SLICE_X12Y147_A5Q),
.I1(RIOB33_X105Y103_IOB_X1Y104_I),
.I2(CLBLM_R_X11Y145_SLICE_X15Y145_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLL_L_X4Y145_SLICE_X4Y145_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y145_SLICE_X13Y145_AO5),
.O6(CLBLM_L_X10Y145_SLICE_X13Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y146_SLICE_X12Y146_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y148_SLICE_X8Y148_BO6),
.Q(CLBLM_L_X10Y146_SLICE_X12Y146_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y146_SLICE_X12Y146_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y148_SLICE_X12Y148_AO6),
.Q(CLBLM_L_X10Y146_SLICE_X12Y146_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y146_SLICE_X12Y146_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y146_SLICE_X12Y146_CO5),
.Q(CLBLM_L_X10Y146_SLICE_X12Y146_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y146_SLICE_X12Y146_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y146_SLICE_X12Y146_DO5),
.Q(CLBLM_L_X10Y146_SLICE_X12Y146_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y146_SLICE_X12Y146_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y146_SLICE_X12Y146_AO6),
.Q(CLBLM_L_X10Y146_SLICE_X12Y146_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y146_SLICE_X12Y146_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y146_SLICE_X12Y146_BO6),
.Q(CLBLM_L_X10Y146_SLICE_X12Y146_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y146_SLICE_X12Y146_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y146_SLICE_X12Y146_CO6),
.Q(CLBLM_L_X10Y146_SLICE_X12Y146_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y146_SLICE_X12Y146_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y146_SLICE_X12Y146_DO6),
.Q(CLBLM_L_X10Y146_SLICE_X12Y146_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaac0c0ccccff00)
  ) CLBLM_L_X10Y146_SLICE_X12Y146_DLUT (
.I0(CLBLM_L_X8Y145_SLICE_X10Y145_BQ),
.I1(CLBLM_L_X10Y146_SLICE_X13Y146_A5Q),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X7Y148_SLICE_X8Y148_DQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y146_SLICE_X12Y146_DO5),
.O6(CLBLM_L_X10Y146_SLICE_X12Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f3c0c0ee22ee22)
  ) CLBLM_L_X10Y146_SLICE_X12Y146_CLUT (
.I0(CLBLM_R_X11Y153_SLICE_X15Y153_BQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X12Y144_SLICE_X16Y144_BQ),
.I3(CLBLM_L_X10Y144_SLICE_X12Y144_CQ),
.I4(CLBLM_L_X10Y146_SLICE_X12Y146_B5Q),
.I5(1'b1),
.O5(CLBLM_L_X10Y146_SLICE_X12Y146_CO5),
.O6(CLBLM_L_X10Y146_SLICE_X12Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff0fcf00f000c00)
  ) CLBLM_L_X10Y146_SLICE_X12Y146_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y146_SLICE_X12Y146_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y142_SLICE_X8Y142_DO6),
.I4(CLBLM_R_X11Y146_SLICE_X15Y146_AQ),
.I5(CLBLM_R_X7Y148_SLICE_X8Y148_CQ),
.O5(CLBLM_L_X10Y146_SLICE_X12Y146_BO5),
.O6(CLBLM_L_X10Y146_SLICE_X12Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaafcffffff)
  ) CLBLM_L_X10Y146_SLICE_X12Y146_ALUT (
.I0(CLBLM_L_X10Y146_SLICE_X12Y146_B5Q),
.I1(CLBLM_R_X5Y154_SLICE_X6Y154_BO6),
.I2(RIOB33_X105Y135_IOB_X1Y136_I),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(RIOB33_X105Y135_IOB_X1Y135_I),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y146_SLICE_X12Y146_AO5),
.O6(CLBLM_L_X10Y146_SLICE_X12Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y146_SLICE_X13Y146_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y146_SLICE_X13Y146_AO5),
.Q(CLBLM_L_X10Y146_SLICE_X13Y146_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y146_SLICE_X13Y146_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y146_SLICE_X13Y146_BO5),
.Q(CLBLM_L_X10Y146_SLICE_X13Y146_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y146_SLICE_X13Y146_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y146_SLICE_X13Y146_AO6),
.Q(CLBLM_L_X10Y146_SLICE_X13Y146_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y146_SLICE_X13Y146_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y146_SLICE_X13Y146_BO6),
.Q(CLBLM_L_X10Y146_SLICE_X13Y146_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y146_SLICE_X13Y146_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y146_SLICE_X13Y146_CO6),
.Q(CLBLM_L_X10Y146_SLICE_X13Y146_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffeeffee)
  ) CLBLM_L_X10Y146_SLICE_X13Y146_DLUT (
.I0(CLBLM_L_X10Y148_SLICE_X13Y148_BQ),
.I1(CLBLM_L_X10Y146_SLICE_X13Y146_CQ),
.I2(1'b1),
.I3(CLBLM_L_X10Y146_SLICE_X13Y146_A5Q),
.I4(1'b1),
.I5(CLBLM_L_X10Y145_SLICE_X13Y145_BQ),
.O5(CLBLM_L_X10Y146_SLICE_X13Y146_DO5),
.O6(CLBLM_L_X10Y146_SLICE_X13Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hbb11aa00bb11aa00)
  ) CLBLM_L_X10Y146_SLICE_X13Y146_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(1'b1),
.I3(CLBLM_R_X11Y148_SLICE_X15Y148_A5Q),
.I4(CLBLM_L_X10Y147_SLICE_X13Y147_BQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y146_SLICE_X13Y146_CO5),
.O6(CLBLM_L_X10Y146_SLICE_X13Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccf0ccf0ff440044)
  ) CLBLM_L_X10Y146_SLICE_X13Y146_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X10Y145_SLICE_X13Y145_BQ),
.I2(RIOB33_X105Y103_IOB_X1Y103_I),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y147_SLICE_X12Y147_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y146_SLICE_X13Y146_BO5),
.O6(CLBLM_L_X10Y146_SLICE_X13Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0f00ff000a0a)
  ) CLBLM_L_X10Y146_SLICE_X13Y146_ALUT (
.I0(CLBLM_R_X7Y149_SLICE_X8Y149_CQ),
.I1(CLBLM_R_X11Y149_SLICE_X14Y149_CQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_L_X10Y146_SLICE_X13Y146_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y146_SLICE_X13Y146_AO5),
.O6(CLBLM_L_X10Y146_SLICE_X13Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y147_SLICE_X12Y147_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y152_SLICE_X12Y152_CO6),
.Q(CLBLM_L_X10Y147_SLICE_X12Y147_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y147_SLICE_X12Y147_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y147_SLICE_X12Y147_AO6),
.Q(CLBLM_L_X10Y147_SLICE_X12Y147_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y147_SLICE_X12Y147_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y147_SLICE_X12Y147_CO6),
.Q(CLBLM_L_X10Y147_SLICE_X12Y147_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbb88888fff00000)
  ) CLBLM_L_X10Y147_SLICE_X12Y147_DLUT (
.I0(CLBLM_R_X3Y143_SLICE_X2Y143_BQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y146_SLICE_X13Y146_AQ),
.I3(CLBLM_R_X11Y147_SLICE_X15Y147_BQ),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y147_SLICE_X12Y147_DO5),
.O6(CLBLM_L_X10Y147_SLICE_X12Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc05cc50cc05cc50)
  ) CLBLM_L_X10Y147_SLICE_X12Y147_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X11Y146_SLICE_X14Y146_DQ),
.I2(CLBLM_L_X10Y150_SLICE_X12Y150_DQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y147_SLICE_X12Y147_BO5),
.I5(1'b1),
.O5(CLBLM_L_X10Y147_SLICE_X12Y147_CO5),
.O6(CLBLM_L_X10Y147_SLICE_X12Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcf80c08cc88cc88)
  ) CLBLM_L_X10Y147_SLICE_X12Y147_BLUT (
.I0(CLBLM_R_X11Y148_SLICE_X15Y148_CQ),
.I1(RIOB33_X105Y121_IOB_X1Y121_I),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y146_SLICE_X13Y146_B5Q),
.I4(CLBLM_L_X10Y145_SLICE_X13Y145_CQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y147_SLICE_X12Y147_BO5),
.O6(CLBLM_L_X10Y147_SLICE_X12Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaabefa00001450)
  ) CLBLM_L_X10Y147_SLICE_X12Y147_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X11Y147_SLICE_X14Y147_BQ),
.I2(CLBLM_L_X10Y147_SLICE_X12Y147_AQ),
.I3(CLBLL_L_X4Y146_SLICE_X4Y146_DO6),
.I4(CLBLM_R_X11Y146_SLICE_X14Y146_AQ),
.I5(CLBLM_L_X10Y148_SLICE_X13Y148_AQ),
.O5(CLBLM_L_X10Y147_SLICE_X12Y147_AO5),
.O6(CLBLM_L_X10Y147_SLICE_X12Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y147_SLICE_X13Y147_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y147_SLICE_X13Y147_AO6),
.Q(CLBLM_L_X10Y147_SLICE_X13Y147_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y147_SLICE_X13Y147_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y147_SLICE_X13Y147_BO6),
.Q(CLBLM_L_X10Y147_SLICE_X13Y147_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf00ff30cf00ff30c)
  ) CLBLM_L_X10Y147_SLICE_X13Y147_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y147_SLICE_X11Y147_CO6),
.I2(CLBLM_L_X10Y149_SLICE_X13Y149_DQ),
.I3(CLBLM_L_X10Y146_SLICE_X13Y146_CQ),
.I4(CLBLM_L_X10Y147_SLICE_X13Y147_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y147_SLICE_X13Y147_DO5),
.O6(CLBLM_L_X10Y147_SLICE_X13Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffdc10ffffdc10)
  ) CLBLM_L_X10Y147_SLICE_X13Y147_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X10Y144_SLICE_X13Y144_AQ),
.I2(CLBLM_R_X3Y151_SLICE_X3Y151_AO6),
.I3(CLBLM_R_X5Y145_SLICE_X6Y145_BO5),
.I4(CLBLM_R_X5Y144_SLICE_X7Y144_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y147_SLICE_X13Y147_CO5),
.O6(CLBLM_L_X10Y147_SLICE_X13Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'he2e2c0c0e2e2c0c0)
  ) CLBLM_L_X10Y147_SLICE_X13Y147_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X8Y146_SLICE_X11Y146_BQ),
.I3(1'b1),
.I4(CLBLM_L_X8Y145_SLICE_X10Y145_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y147_SLICE_X13Y147_BO5),
.O6(CLBLM_L_X10Y147_SLICE_X13Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff01ff6800010068)
  ) CLBLM_L_X10Y147_SLICE_X13Y147_ALUT (
.I0(CLBLM_L_X10Y147_SLICE_X13Y147_DO6),
.I1(CLBLM_L_X10Y147_SLICE_X13Y147_BQ),
.I2(CLBLM_L_X10Y147_SLICE_X13Y147_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_L_X8Y145_SLICE_X11Y145_A5Q),
.O5(CLBLM_L_X10Y147_SLICE_X13Y147_AO5),
.O6(CLBLM_L_X10Y147_SLICE_X13Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y148_SLICE_X12Y148_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y148_SLICE_X12Y148_BO6),
.Q(CLBLM_L_X10Y148_SLICE_X12Y148_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y148_SLICE_X12Y148_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y148_SLICE_X12Y148_CO6),
.Q(CLBLM_L_X10Y148_SLICE_X12Y148_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h313331333f3f3f3f)
  ) CLBLM_L_X10Y148_SLICE_X12Y148_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X10Y148_SLICE_X13Y148_CO6),
.I2(CLBLM_R_X5Y144_SLICE_X7Y144_AQ),
.I3(CLBLL_L_X2Y151_SLICE_X1Y151_BO6),
.I4(1'b1),
.I5(CLBLM_L_X10Y144_SLICE_X13Y144_AQ),
.O5(CLBLM_L_X10Y148_SLICE_X12Y148_DO5),
.O6(CLBLM_L_X10Y148_SLICE_X12Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'he4e4f5f5e4a0f5a0)
  ) CLBLM_L_X10Y148_SLICE_X12Y148_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y148_SLICE_X12Y148_CQ),
.I2(CLBLM_L_X10Y148_SLICE_X12Y148_BQ),
.I3(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.I4(CLBLM_L_X10Y148_SLICE_X12Y148_DO6),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_L_X10Y148_SLICE_X12Y148_CO5),
.O6(CLBLM_L_X10Y148_SLICE_X12Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff54ff5400540054)
  ) CLBLM_L_X10Y148_SLICE_X12Y148_BLUT (
.I0(CLBLL_L_X4Y145_SLICE_X5Y145_DO6),
.I1(CLBLM_L_X10Y148_SLICE_X12Y148_BQ),
.I2(CLBLM_L_X10Y146_SLICE_X12Y146_BQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLM_L_X8Y151_SLICE_X10Y151_CQ),
.O5(CLBLM_L_X10Y148_SLICE_X12Y148_BO5),
.O6(CLBLM_L_X10Y148_SLICE_X12Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbb88888fff00000)
  ) CLBLM_L_X10Y148_SLICE_X12Y148_ALUT (
.I0(CLBLM_L_X10Y149_SLICE_X13Y149_DQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLL_L_X4Y146_SLICE_X5Y146_A5Q),
.I3(CLBLM_L_X10Y148_SLICE_X12Y148_CQ),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y148_SLICE_X12Y148_AO5),
.O6(CLBLM_L_X10Y148_SLICE_X12Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y148_SLICE_X13Y148_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y148_SLICE_X13Y148_AO6),
.Q(CLBLM_L_X10Y148_SLICE_X13Y148_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y148_SLICE_X13Y148_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y148_SLICE_X13Y148_BO6),
.Q(CLBLM_L_X10Y148_SLICE_X13Y148_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5545000055550055)
  ) CLBLM_L_X10Y148_SLICE_X13Y148_DLUT (
.I0(CLBLM_L_X8Y145_SLICE_X10Y145_CO5),
.I1(CLBLM_R_X3Y151_SLICE_X3Y151_AO6),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X5Y144_SLICE_X7Y144_AQ),
.I4(CLBLM_L_X10Y148_SLICE_X13Y148_CO5),
.I5(CLBLM_L_X10Y144_SLICE_X13Y144_AQ),
.O5(CLBLM_L_X10Y148_SLICE_X13Y148_DO5),
.O6(CLBLM_L_X10Y148_SLICE_X13Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaa0000f0f0cccc)
  ) CLBLM_L_X10Y148_SLICE_X13Y148_CLUT (
.I0(CLBLL_L_X4Y146_SLICE_X5Y146_A5Q),
.I1(CLBLM_L_X10Y148_SLICE_X13Y148_AQ),
.I2(CLBLM_R_X7Y152_SLICE_X9Y152_CQ),
.I3(CLBLM_L_X8Y149_SLICE_X11Y149_CQ),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y148_SLICE_X13Y148_CO5),
.O6(CLBLM_L_X10Y148_SLICE_X13Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcfcccc03030000)
  ) CLBLM_L_X10Y148_SLICE_X13Y148_BLUT (
.I0(1'b1),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(1'b1),
.I4(CLBLL_L_X4Y148_SLICE_X4Y148_CQ),
.I5(CLBLM_L_X10Y150_SLICE_X13Y150_A5Q),
.O5(CLBLM_L_X10Y148_SLICE_X13Y148_BO5),
.O6(CLBLM_L_X10Y148_SLICE_X13Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff550055ff740074)
  ) CLBLM_L_X10Y148_SLICE_X13Y148_ALUT (
.I0(CLBLM_L_X8Y148_SLICE_X10Y148_DO6),
.I1(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.I2(CLBLM_L_X10Y148_SLICE_X13Y148_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y150_SLICE_X13Y150_AQ),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_L_X10Y148_SLICE_X13Y148_AO5),
.O6(CLBLM_L_X10Y148_SLICE_X13Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y149_SLICE_X12Y149_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y77_IOB_X0Y77_I),
.D(CLBLM_L_X8Y144_SLICE_X10Y144_CQ),
.Q(CLBLM_L_X10Y149_SLICE_X12Y149_AQ),
.R(CLBLM_R_X11Y151_SLICE_X15Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0c0e0c0e0f0f0f0f)
  ) CLBLM_L_X10Y149_SLICE_X12Y149_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X5Y144_SLICE_X7Y144_AQ),
.I2(CLBLM_L_X10Y150_SLICE_X13Y150_A5Q),
.I3(CLBLL_L_X4Y154_SLICE_X4Y154_CO6),
.I4(1'b1),
.I5(CLBLM_L_X10Y144_SLICE_X13Y144_AQ),
.O5(CLBLM_L_X10Y149_SLICE_X12Y149_DO5),
.O6(CLBLM_L_X10Y149_SLICE_X12Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0099660000669900)
  ) CLBLM_L_X10Y149_SLICE_X12Y149_CLUT (
.I0(CLBLM_R_X5Y151_SLICE_X6Y151_BQ),
.I1(CLBLM_L_X10Y150_SLICE_X13Y150_CQ),
.I2(1'b1),
.I3(CLBLM_L_X10Y145_SLICE_X12Y145_CQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_L_X10Y149_SLICE_X13Y149_BQ),
.O5(CLBLM_L_X10Y149_SLICE_X12Y149_CO5),
.O6(CLBLM_L_X10Y149_SLICE_X12Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'heeec2220aaa0aaa0)
  ) CLBLM_L_X10Y149_SLICE_X12Y149_BLUT (
.I0(RIOB33_X105Y121_IOB_X1Y121_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X7Y145_SLICE_X9Y145_C5Q),
.I3(CLBLM_L_X8Y148_SLICE_X11Y148_AQ),
.I4(CLBLM_L_X10Y146_SLICE_X12Y146_BQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y149_SLICE_X12Y149_BO5),
.O6(CLBLM_L_X10Y149_SLICE_X12Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0010100000fcfc)
  ) CLBLM_L_X10Y149_SLICE_X12Y149_ALUT (
.I0(CLBLM_L_X10Y149_SLICE_X12Y149_DO6),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.I3(CLBLM_R_X11Y147_SLICE_X15Y147_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y149_SLICE_X12Y149_AO5),
.O6(CLBLM_L_X10Y149_SLICE_X12Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y149_SLICE_X13Y149_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y149_SLICE_X13Y149_CO6),
.Q(CLBLM_L_X10Y149_SLICE_X13Y149_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y149_SLICE_X13Y149_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y149_SLICE_X13Y149_AO6),
.Q(CLBLM_L_X10Y149_SLICE_X13Y149_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y149_SLICE_X13Y149_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y149_SLICE_X13Y149_BO6),
.Q(CLBLM_L_X10Y149_SLICE_X13Y149_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y149_SLICE_X13Y149_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y149_SLICE_X13Y149_DO6),
.Q(CLBLM_L_X10Y149_SLICE_X13Y149_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hdcdcdcdc10101010)
  ) CLBLM_L_X10Y149_SLICE_X13Y149_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLL_L_X4Y146_SLICE_X5Y146_A5Q),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X11Y153_SLICE_X15Y153_AQ),
.O5(CLBLM_L_X10Y149_SLICE_X13Y149_DO5),
.O6(CLBLM_L_X10Y149_SLICE_X13Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3c0e2c000ff55ff)
  ) CLBLM_L_X10Y149_SLICE_X13Y149_CLUT (
.I0(CLBLL_L_X4Y148_SLICE_X4Y148_CQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X12Y148_SLICE_X16Y148_AQ),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(CLBLM_R_X11Y147_SLICE_X15Y147_DQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y149_SLICE_X13Y149_CO5),
.O6(CLBLM_L_X10Y149_SLICE_X13Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0f3c0c0f3c0)
  ) CLBLM_L_X10Y149_SLICE_X13Y149_BLUT (
.I0(1'b1),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X7Y145_SLICE_X9Y145_C5Q),
.I3(CLBLM_L_X10Y150_SLICE_X13Y150_CQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_L_X10Y148_SLICE_X13Y148_CO6),
.O5(CLBLM_L_X10Y149_SLICE_X13Y149_BO5),
.O6(CLBLM_L_X10Y149_SLICE_X13Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdecddcc31201100)
  ) CLBLM_L_X10Y149_SLICE_X13Y149_ALUT (
.I0(CLBLM_R_X11Y147_SLICE_X14Y147_CO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y149_SLICE_X13Y149_AQ),
.I3(CLBLM_R_X11Y150_SLICE_X15Y150_AQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_L_X8Y149_SLICE_X11Y149_CQ),
.O5(CLBLM_L_X10Y149_SLICE_X13Y149_AO5),
.O6(CLBLM_L_X10Y149_SLICE_X13Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y150_SLICE_X12Y150_A5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y149_SLICE_X12Y149_BO6),
.Q(CLBLM_L_X10Y150_SLICE_X12Y150_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y150_SLICE_X12Y150_B5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y147_SLICE_X12Y147_DO6),
.Q(CLBLM_L_X10Y150_SLICE_X12Y150_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y150_SLICE_X12Y150_C5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y147_SLICE_X11Y147_AO6),
.Q(CLBLM_L_X10Y150_SLICE_X12Y150_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y150_SLICE_X12Y150_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y150_SLICE_X12Y150_AO6),
.Q(CLBLM_L_X10Y150_SLICE_X12Y150_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y150_SLICE_X12Y150_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y150_SLICE_X12Y150_BO6),
.Q(CLBLM_L_X10Y150_SLICE_X12Y150_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y150_SLICE_X12Y150_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y150_SLICE_X12Y150_CO6),
.Q(CLBLM_L_X10Y150_SLICE_X12Y150_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y150_SLICE_X12Y150_D_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y150_SLICE_X12Y150_DO6),
.Q(CLBLM_L_X10Y150_SLICE_X12Y150_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0006060606)
  ) CLBLM_L_X10Y150_SLICE_X12Y150_DLUT (
.I0(CLBLM_L_X10Y147_SLICE_X12Y147_DO5),
.I1(CLBLM_R_X7Y148_SLICE_X8Y148_CQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_L_X12Y152_SLICE_X16Y152_BQ),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y150_SLICE_X12Y150_DO5),
.O6(CLBLM_L_X10Y150_SLICE_X12Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0d1c0d1d1c0d1c0)
  ) CLBLM_L_X10Y150_SLICE_X12Y150_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y149_SLICE_X13Y149_A5Q),
.I3(CLBLM_L_X10Y147_SLICE_X12Y147_CQ),
.I4(1'b1),
.I5(CLBLM_L_X10Y149_SLICE_X12Y149_BO5),
.O5(CLBLM_L_X10Y150_SLICE_X12Y150_CO5),
.O6(CLBLM_L_X10Y150_SLICE_X12Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff000000f0f0)
  ) CLBLM_L_X10Y150_SLICE_X12Y150_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X5Y148_SLICE_X6Y148_BQ),
.I3(CLBLM_L_X10Y150_SLICE_X13Y150_BQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y150_SLICE_X12Y150_BO5),
.O6(CLBLM_L_X10Y150_SLICE_X12Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaf0aa00aaccaacc)
  ) CLBLM_L_X10Y150_SLICE_X12Y150_ALUT (
.I0(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.I1(CLBLM_R_X11Y149_SLICE_X14Y149_BQ),
.I2(CLBLM_L_X10Y150_SLICE_X12Y150_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X11Y147_SLICE_X14Y147_CO6),
.O5(CLBLM_L_X10Y150_SLICE_X12Y150_AO5),
.O6(CLBLM_L_X10Y150_SLICE_X12Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y150_SLICE_X13Y150_A5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y149_SLICE_X12Y149_AO6),
.Q(CLBLM_L_X10Y150_SLICE_X13Y150_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y150_SLICE_X13Y150_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y150_SLICE_X13Y150_AO6),
.Q(CLBLM_L_X10Y150_SLICE_X13Y150_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y150_SLICE_X13Y150_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y150_SLICE_X13Y150_BO6),
.Q(CLBLM_L_X10Y150_SLICE_X13Y150_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y150_SLICE_X13Y150_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y150_SLICE_X13Y150_CO6),
.Q(CLBLM_L_X10Y150_SLICE_X13Y150_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333222233303330)
  ) CLBLM_L_X10Y150_SLICE_X13Y150_DLUT (
.I0(CLBLL_L_X4Y149_SLICE_X5Y149_A5Q),
.I1(CLBLM_L_X8Y146_SLICE_X10Y146_BQ),
.I2(CLBLM_R_X5Y144_SLICE_X7Y144_CQ),
.I3(CLBLM_L_X10Y150_SLICE_X13Y150_A5Q),
.I4(CLBLM_L_X10Y150_SLICE_X13Y150_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y150_SLICE_X13Y150_DO5),
.O6(CLBLM_L_X10Y150_SLICE_X13Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hab01ae04ab01ae04)
  ) CLBLM_L_X10Y150_SLICE_X13Y150_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y145_SLICE_X6Y145_AQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X11Y151_SLICE_X15Y151_A5Q),
.I4(CLBLM_L_X10Y148_SLICE_X13Y148_CO5),
.I5(1'b1),
.O5(CLBLM_L_X10Y150_SLICE_X13Y150_CO5),
.O6(CLBLM_L_X10Y150_SLICE_X13Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000088f088f0)
  ) CLBLM_L_X10Y150_SLICE_X13Y150_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X10Y150_SLICE_X13Y150_BQ),
.I2(CLBLM_L_X12Y149_SLICE_X17Y149_BQ),
.I3(CLBLM_R_X11Y147_SLICE_X14Y147_CO6),
.I4(CLBLM_L_X8Y147_SLICE_X10Y147_BQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y150_SLICE_X13Y150_BO5),
.O6(CLBLM_L_X10Y150_SLICE_X13Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffccaaffffcca0)
  ) CLBLM_L_X10Y150_SLICE_X13Y150_ALUT (
.I0(CLBLM_L_X10Y150_SLICE_X13Y150_AQ),
.I1(CLBLM_R_X11Y152_SLICE_X15Y152_BQ),
.I2(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y149_SLICE_X9Y149_DO6),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_L_X10Y150_SLICE_X13Y150_AO5),
.O6(CLBLM_L_X10Y150_SLICE_X13Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y151_SLICE_X12Y151_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y151_SLICE_X12Y151_AO6),
.Q(CLBLM_L_X10Y151_SLICE_X12Y151_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y151_SLICE_X12Y151_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y151_SLICE_X12Y151_BO6),
.Q(CLBLM_L_X10Y151_SLICE_X12Y151_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y151_SLICE_X12Y151_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y151_SLICE_X12Y151_CO6),
.Q(CLBLM_L_X10Y151_SLICE_X12Y151_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y151_SLICE_X12Y151_D_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y151_SLICE_X12Y151_DO6),
.Q(CLBLM_L_X10Y151_SLICE_X12Y151_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccf0a0ccccffaa)
  ) CLBLM_L_X10Y151_SLICE_X12Y151_DLUT (
.I0(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.I1(CLBLM_R_X3Y150_SLICE_X3Y150_A5Q),
.I2(CLBLM_L_X10Y151_SLICE_X12Y151_DQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X10Y148_SLICE_X12Y148_DO6),
.O5(CLBLM_L_X10Y151_SLICE_X12Y151_DO5),
.O6(CLBLM_L_X10Y151_SLICE_X12Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f000aa0088)
  ) CLBLM_L_X10Y151_SLICE_X12Y151_CLUT (
.I0(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.I1(CLBLM_L_X10Y144_SLICE_X12Y144_CQ),
.I2(CLBLM_L_X10Y151_SLICE_X12Y151_DQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_L_X10Y151_SLICE_X12Y151_CQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y151_SLICE_X12Y151_CO5),
.O6(CLBLM_L_X10Y151_SLICE_X12Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff88fff0008800f0)
  ) CLBLM_L_X10Y151_SLICE_X12Y151_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X10Y151_SLICE_X12Y151_BQ),
.I2(CLBLM_L_X10Y150_SLICE_X12Y150_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X11Y147_SLICE_X14Y147_CO6),
.I5(CLBLM_L_X8Y153_SLICE_X11Y153_CQ),
.O5(CLBLM_L_X10Y151_SLICE_X12Y151_BO5),
.O6(CLBLM_L_X10Y151_SLICE_X12Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hee22ee22ee22fc30)
  ) CLBLM_L_X10Y151_SLICE_X12Y151_ALUT (
.I0(CLBLM_R_X7Y151_SLICE_X8Y151_BQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y151_SLICE_X12Y151_AQ),
.I3(CLBLM_L_X10Y154_SLICE_X13Y154_BQ),
.I4(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_L_X10Y151_SLICE_X12Y151_AO5),
.O6(CLBLM_L_X10Y151_SLICE_X12Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y151_SLICE_X13Y151_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y151_SLICE_X13Y151_AO6),
.Q(CLBLM_L_X10Y151_SLICE_X13Y151_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y151_SLICE_X13Y151_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y151_SLICE_X13Y151_BO6),
.Q(CLBLM_L_X10Y151_SLICE_X13Y151_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y151_SLICE_X13Y151_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y151_SLICE_X13Y151_CO6),
.Q(CLBLM_L_X10Y151_SLICE_X13Y151_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y151_SLICE_X13Y151_D_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y151_SLICE_X13Y151_DO6),
.Q(CLBLM_L_X10Y151_SLICE_X13Y151_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff222000002220)
  ) CLBLM_L_X10Y151_SLICE_X13Y151_DLUT (
.I0(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_L_X10Y151_SLICE_X13Y151_DQ),
.I3(CLBLM_R_X11Y149_SLICE_X14Y149_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X11Y152_SLICE_X14Y152_BQ),
.O5(CLBLM_L_X10Y151_SLICE_X13Y151_DO5),
.O6(CLBLM_L_X10Y151_SLICE_X13Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa0f00cfc0)
  ) CLBLM_L_X10Y151_SLICE_X13Y151_CLUT (
.I0(CLBLM_R_X5Y150_SLICE_X6Y150_DQ),
.I1(CLBLM_L_X10Y151_SLICE_X13Y151_CQ),
.I2(CLBLM_R_X11Y153_SLICE_X14Y153_BO5),
.I3(CLBLM_R_X11Y152_SLICE_X14Y152_CQ),
.I4(CLBLM_R_X11Y154_SLICE_X15Y154_CO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y151_SLICE_X13Y151_CO5),
.O6(CLBLM_L_X10Y151_SLICE_X13Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f011004400)
  ) CLBLM_L_X10Y151_SLICE_X13Y151_BLUT (
.I0(CLBLM_R_X5Y152_SLICE_X7Y152_BQ),
.I1(CLBLM_L_X10Y151_SLICE_X13Y151_BQ),
.I2(CLBLM_R_X7Y143_SLICE_X8Y143_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X11Y151_SLICE_X14Y151_CO5),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y151_SLICE_X13Y151_BO5),
.O6(CLBLM_L_X10Y151_SLICE_X13Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hddccdccc11001000)
  ) CLBLM_L_X10Y151_SLICE_X13Y151_ALUT (
.I0(CLBLM_R_X5Y152_SLICE_X7Y152_BQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y151_SLICE_X13Y151_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X11Y151_SLICE_X14Y151_BO6),
.I5(CLBLM_L_X10Y151_SLICE_X12Y151_CQ),
.O5(CLBLM_L_X10Y151_SLICE_X13Y151_AO5),
.O6(CLBLM_L_X10Y151_SLICE_X13Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y152_SLICE_X12Y152_D5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y152_SLICE_X12Y152_DO5),
.Q(CLBLM_L_X10Y152_SLICE_X12Y152_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y152_SLICE_X12Y152_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y152_SLICE_X12Y152_AO6),
.Q(CLBLM_L_X10Y152_SLICE_X12Y152_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y152_SLICE_X12Y152_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y152_SLICE_X12Y152_BO6),
.Q(CLBLM_L_X10Y152_SLICE_X12Y152_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y152_SLICE_X12Y152_D_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y152_SLICE_X12Y152_DO6),
.Q(CLBLM_L_X10Y152_SLICE_X12Y152_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hee22ee22f3f3c0c0)
  ) CLBLM_L_X10Y152_SLICE_X12Y152_DLUT (
.I0(CLBLM_L_X10Y153_SLICE_X12Y153_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y150_SLICE_X12Y150_CQ),
.I3(CLBLM_R_X11Y144_SLICE_X14Y144_BQ),
.I4(CLBLM_R_X7Y154_SLICE_X9Y154_BQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y152_SLICE_X12Y152_DO5),
.O6(CLBLM_L_X10Y152_SLICE_X12Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffc800c8c8c8c8c8)
  ) CLBLM_L_X10Y152_SLICE_X12Y152_CLUT (
.I0(CLBLM_L_X10Y146_SLICE_X12Y146_DQ),
.I1(RIOB33_X105Y121_IOB_X1Y121_I),
.I2(CLBLM_L_X10Y152_SLICE_X12Y152_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y152_SLICE_X12Y152_D5Q),
.I5(1'b1),
.O5(CLBLM_L_X10Y152_SLICE_X12Y152_CO5),
.O6(CLBLM_L_X10Y152_SLICE_X12Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc00aaf0f0)
  ) CLBLM_L_X10Y152_SLICE_X12Y152_BLUT (
.I0(CLBLM_L_X10Y152_SLICE_X12Y152_BQ),
.I1(CLBLM_L_X10Y150_SLICE_X12Y150_BQ),
.I2(CLBLM_L_X10Y153_SLICE_X12Y153_BQ),
.I3(CLBLM_R_X11Y154_SLICE_X15Y154_CO6),
.I4(CLBLM_R_X11Y153_SLICE_X14Y153_BO5),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y152_SLICE_X12Y152_BO5),
.O6(CLBLM_L_X10Y152_SLICE_X12Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfebafebafebaeeaa)
  ) CLBLM_L_X10Y152_SLICE_X12Y152_ALUT (
.I0(CLBLM_L_X8Y145_SLICE_X10Y145_DO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y152_SLICE_X12Y152_AQ),
.I3(CLBLM_R_X7Y152_SLICE_X8Y152_AQ),
.I4(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_L_X10Y152_SLICE_X12Y152_AO5),
.O6(CLBLM_L_X10Y152_SLICE_X12Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y152_SLICE_X13Y152_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y152_SLICE_X13Y152_AO6),
.Q(CLBLM_L_X10Y152_SLICE_X13Y152_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y152_SLICE_X13Y152_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y152_SLICE_X13Y152_BO6),
.Q(CLBLM_L_X10Y152_SLICE_X13Y152_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccffffffff)
  ) CLBLM_L_X10Y152_SLICE_X13Y152_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y153_SLICE_X14Y153_BO5),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X10Y154_SLICE_X13Y154_BQ),
.O5(CLBLM_L_X10Y152_SLICE_X13Y152_DO5),
.O6(CLBLM_L_X10Y152_SLICE_X13Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00f000ee00ee)
  ) CLBLM_L_X10Y152_SLICE_X13Y152_CLUT (
.I0(CLBLM_L_X10Y145_SLICE_X12Y145_AQ),
.I1(CLBLM_L_X10Y152_SLICE_X13Y152_AQ),
.I2(CLBLM_L_X10Y153_SLICE_X13Y153_DQ),
.I3(CLBLM_L_X8Y146_SLICE_X10Y146_BQ),
.I4(CLBLM_R_X7Y144_SLICE_X8Y144_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y152_SLICE_X13Y152_CO5),
.O6(CLBLM_L_X10Y152_SLICE_X13Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0e4a0e4f5f5a0a0)
  ) CLBLM_L_X10Y152_SLICE_X13Y152_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y152_SLICE_X13Y152_BQ),
.I2(CLBLM_L_X10Y152_SLICE_X13Y152_AQ),
.I3(CLBLM_R_X11Y154_SLICE_X15Y154_CO6),
.I4(CLBLM_R_X11Y152_SLICE_X14Y152_AQ),
.I5(CLBLM_R_X11Y153_SLICE_X14Y153_BO5),
.O5(CLBLM_L_X10Y152_SLICE_X13Y152_BO5),
.O6(CLBLM_L_X10Y152_SLICE_X13Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00fe32cc00)
  ) CLBLM_L_X10Y152_SLICE_X13Y152_ALUT (
.I0(CLBLM_L_X10Y147_SLICE_X13Y147_CO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y152_SLICE_X13Y152_AQ),
.I3(CLBLM_L_X8Y151_SLICE_X11Y151_AQ),
.I4(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_L_X10Y152_SLICE_X13Y152_AO5),
.O6(CLBLM_L_X10Y152_SLICE_X13Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y153_SLICE_X12Y153_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y153_SLICE_X12Y153_AO6),
.Q(CLBLM_L_X10Y153_SLICE_X12Y153_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y153_SLICE_X12Y153_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y153_SLICE_X12Y153_BO6),
.Q(CLBLM_L_X10Y153_SLICE_X12Y153_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y153_SLICE_X12Y153_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y153_SLICE_X12Y153_CO6),
.Q(CLBLM_L_X10Y153_SLICE_X12Y153_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y153_SLICE_X12Y153_D_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y153_SLICE_X12Y153_DO6),
.Q(CLBLM_L_X10Y153_SLICE_X12Y153_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaa00feff000000)
  ) CLBLM_L_X10Y153_SLICE_X12Y153_DLUT (
.I0(CLBLM_R_X11Y154_SLICE_X15Y154_AQ),
.I1(CLBLM_R_X11Y154_SLICE_X14Y154_AQ),
.I2(CLBLM_R_X11Y154_SLICE_X15Y154_BQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y153_SLICE_X13Y153_BQ),
.I5(CLBLM_R_X7Y148_SLICE_X9Y148_BQ),
.O5(CLBLM_L_X10Y153_SLICE_X12Y153_DO5),
.O6(CLBLM_L_X10Y153_SLICE_X12Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff005555ff000101)
  ) CLBLM_L_X10Y153_SLICE_X12Y153_CLUT (
.I0(CLBLM_R_X11Y154_SLICE_X15Y154_AQ),
.I1(CLBLM_R_X11Y154_SLICE_X14Y154_AQ),
.I2(CLBLM_R_X11Y154_SLICE_X15Y154_BQ),
.I3(CLBLM_L_X10Y153_SLICE_X13Y153_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X10Y153_SLICE_X13Y153_BQ),
.O5(CLBLM_L_X10Y153_SLICE_X12Y153_CO5),
.O6(CLBLM_L_X10Y153_SLICE_X12Y153_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaffffaaaa0f0c)
  ) CLBLM_L_X10Y153_SLICE_X12Y153_BLUT (
.I0(CLBLM_L_X8Y153_SLICE_X11Y153_DQ),
.I1(CLBLM_L_X10Y153_SLICE_X12Y153_BQ),
.I2(CLBLM_R_X11Y153_SLICE_X14Y153_BO5),
.I3(CLBLM_L_X10Y154_SLICE_X13Y154_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X11Y154_SLICE_X15Y154_CO6),
.O5(CLBLM_L_X10Y153_SLICE_X12Y153_BO5),
.O6(CLBLM_L_X10Y153_SLICE_X12Y153_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcfcfcfcfcfcacf)
  ) CLBLM_L_X10Y153_SLICE_X12Y153_ALUT (
.I0(RIOB33_X105Y135_IOB_X1Y136_I),
.I1(CLBLM_L_X10Y150_SLICE_X12Y150_C5Q),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y135_IOB_X1Y135_I),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(CLBLM_R_X5Y154_SLICE_X6Y154_BO6),
.O5(CLBLM_L_X10Y153_SLICE_X12Y153_AO5),
.O6(CLBLM_L_X10Y153_SLICE_X12Y153_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y153_SLICE_X13Y153_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y153_SLICE_X13Y153_AO6),
.Q(CLBLM_L_X10Y153_SLICE_X13Y153_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y153_SLICE_X13Y153_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y153_SLICE_X13Y153_BO6),
.Q(CLBLM_L_X10Y153_SLICE_X13Y153_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y153_SLICE_X13Y153_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y153_SLICE_X13Y153_CO6),
.Q(CLBLM_L_X10Y153_SLICE_X13Y153_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y153_SLICE_X13Y153_D_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y153_SLICE_X13Y153_DO6),
.Q(CLBLM_L_X10Y153_SLICE_X13Y153_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff00c8000000c8)
  ) CLBLM_L_X10Y153_SLICE_X13Y153_DLUT (
.I0(CLBLM_R_X7Y149_SLICE_X9Y149_CO6),
.I1(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.I2(CLBLM_L_X10Y153_SLICE_X13Y153_DQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X10Y155_SLICE_X13Y155_BQ),
.O5(CLBLM_L_X10Y153_SLICE_X13Y153_DO5),
.O6(CLBLM_L_X10Y153_SLICE_X13Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0afa0a3a0aca0a3)
  ) CLBLM_L_X10Y153_SLICE_X13Y153_CLUT (
.I0(CLBLM_L_X10Y152_SLICE_X12Y152_AQ),
.I1(CLBLM_L_X10Y153_SLICE_X13Y153_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(CLBLM_L_X10Y152_SLICE_X13Y152_DO6),
.I5(CLBLM_R_X11Y153_SLICE_X14Y153_AO5),
.O5(CLBLM_L_X10Y153_SLICE_X13Y153_CO5),
.O6(CLBLM_L_X10Y153_SLICE_X13Y153_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f01144f0f01111)
  ) CLBLM_L_X10Y153_SLICE_X13Y153_BLUT (
.I0(RIOB33_X105Y121_IOB_X1Y121_I),
.I1(CLBLM_L_X10Y153_SLICE_X13Y153_BQ),
.I2(CLBLL_L_X4Y151_SLICE_X5Y151_AQ),
.I3(CLBLM_R_X11Y154_SLICE_X14Y154_BO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X11Y153_SLICE_X14Y153_BO6),
.O5(CLBLM_L_X10Y153_SLICE_X13Y153_BO5),
.O6(CLBLM_L_X10Y153_SLICE_X13Y153_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdcff1033dccc1000)
  ) CLBLM_L_X10Y153_SLICE_X13Y153_ALUT (
.I0(CLBLM_R_X7Y155_SLICE_X8Y155_BO5),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y153_SLICE_X13Y153_AQ),
.I3(CLBLM_R_X5Y155_SLICE_X7Y155_CO6),
.I4(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.I5(CLBLM_L_X10Y154_SLICE_X12Y154_BQ),
.O5(CLBLM_L_X10Y153_SLICE_X13Y153_AO5),
.O6(CLBLM_L_X10Y153_SLICE_X13Y153_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y154_SLICE_X12Y154_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y154_SLICE_X12Y154_AO6),
.Q(CLBLM_L_X10Y154_SLICE_X12Y154_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y154_SLICE_X12Y154_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y154_SLICE_X12Y154_BO6),
.Q(CLBLM_L_X10Y154_SLICE_X12Y154_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y154_SLICE_X12Y154_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y154_SLICE_X12Y154_CO6),
.Q(CLBLM_L_X10Y154_SLICE_X12Y154_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y154_SLICE_X12Y154_D_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y154_SLICE_X12Y154_DO6),
.Q(CLBLM_L_X10Y154_SLICE_X12Y154_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0cffc0ff04554055)
  ) CLBLM_L_X10Y154_SLICE_X12Y154_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y153_SLICE_X10Y153_DO6),
.I2(CLBLM_L_X10Y154_SLICE_X12Y154_DQ),
.I3(CLBLM_L_X8Y153_SLICE_X10Y153_CO5),
.I4(CLBLM_L_X10Y155_SLICE_X12Y155_DO6),
.I5(CLBLM_L_X10Y148_SLICE_X12Y148_CQ),
.O5(CLBLM_L_X10Y154_SLICE_X12Y154_DO5),
.O6(CLBLM_L_X10Y154_SLICE_X12Y154_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0f5e4f5a0a0e4a0)
  ) CLBLM_L_X10Y154_SLICE_X12Y154_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y154_SLICE_X12Y154_CQ),
.I2(CLBLM_L_X8Y145_SLICE_X11Y145_CQ),
.I3(CLBLM_R_X5Y155_SLICE_X7Y155_CO6),
.I4(CLBLM_R_X7Y155_SLICE_X8Y155_BO5),
.I5(CLBLM_R_X7Y154_SLICE_X8Y154_AQ),
.O5(CLBLM_L_X10Y154_SLICE_X12Y154_CO5),
.O6(CLBLM_L_X10Y154_SLICE_X12Y154_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000044f044f0)
  ) CLBLM_L_X10Y154_SLICE_X12Y154_BLUT (
.I0(CLBLM_R_X7Y155_SLICE_X8Y155_BO5),
.I1(CLBLM_L_X10Y154_SLICE_X12Y154_BQ),
.I2(CLBLM_L_X10Y154_SLICE_X12Y154_AQ),
.I3(CLBLM_R_X5Y155_SLICE_X7Y155_CO6),
.I4(CLBLM_R_X7Y145_SLICE_X8Y145_C5Q),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y154_SLICE_X12Y154_BO5),
.O6(CLBLM_L_X10Y154_SLICE_X12Y154_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000073407340)
  ) CLBLM_L_X10Y154_SLICE_X12Y154_ALUT (
.I0(CLBLM_R_X7Y155_SLICE_X8Y155_BO5),
.I1(CLBLM_R_X5Y155_SLICE_X7Y155_CO6),
.I2(CLBLM_L_X10Y154_SLICE_X12Y154_AQ),
.I3(CLBLM_L_X10Y154_SLICE_X12Y154_CQ),
.I4(CLBLM_L_X8Y147_SLICE_X10Y147_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y154_SLICE_X12Y154_AO5),
.O6(CLBLM_L_X10Y154_SLICE_X12Y154_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y154_SLICE_X13Y154_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y154_SLICE_X13Y154_AO6),
.Q(CLBLM_L_X10Y154_SLICE_X13Y154_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y154_SLICE_X13Y154_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y154_SLICE_X13Y154_BO6),
.Q(CLBLM_L_X10Y154_SLICE_X13Y154_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000ff000000)
  ) CLBLM_L_X10Y154_SLICE_X13Y154_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_L_X10Y150_SLICE_X12Y150_B5Q),
.I4(CLBLM_L_X10Y154_SLICE_X13Y154_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y154_SLICE_X13Y154_DO5),
.O6(CLBLM_L_X10Y154_SLICE_X13Y154_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00c001c1fa3a5414)
  ) CLBLM_L_X10Y154_SLICE_X13Y154_CLUT (
.I0(CLBLM_R_X11Y154_SLICE_X14Y154_AQ),
.I1(CLBLM_L_X10Y153_SLICE_X13Y153_BQ),
.I2(CLBLM_R_X11Y154_SLICE_X15Y154_AQ),
.I3(CLBLM_L_X10Y153_SLICE_X13Y153_CQ),
.I4(CLBLM_R_X11Y154_SLICE_X15Y154_BQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y154_SLICE_X13Y154_CO5),
.O6(CLBLM_L_X10Y154_SLICE_X13Y154_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8ddd88d88d8d8888)
  ) CLBLM_L_X10Y154_SLICE_X13Y154_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y154_SLICE_X8Y154_AQ),
.I2(CLBLM_R_X11Y153_SLICE_X14Y153_BO5),
.I3(CLBLM_R_X11Y154_SLICE_X15Y154_CO6),
.I4(CLBLM_L_X10Y151_SLICE_X13Y151_CQ),
.I5(CLBLM_L_X10Y154_SLICE_X13Y154_BQ),
.O5(CLBLM_L_X10Y154_SLICE_X13Y154_BO5),
.O6(CLBLM_L_X10Y154_SLICE_X13Y154_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffcca0ccffccaa)
  ) CLBLM_L_X10Y154_SLICE_X13Y154_ALUT (
.I0(CLBLM_L_X10Y154_SLICE_X13Y154_AQ),
.I1(CLBLM_R_X5Y153_SLICE_X6Y153_BQ),
.I2(CLBLM_R_X11Y154_SLICE_X15Y154_CO5),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X11Y154_SLICE_X14Y154_BO6),
.I5(CLBLM_L_X10Y154_SLICE_X13Y154_CO6),
.O5(CLBLM_L_X10Y154_SLICE_X13Y154_AO5),
.O6(CLBLM_L_X10Y154_SLICE_X13Y154_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y155_SLICE_X12Y155_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y155_SLICE_X12Y155_AO6),
.Q(CLBLM_L_X10Y155_SLICE_X12Y155_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaafefaaaaa)
  ) CLBLM_L_X10Y155_SLICE_X12Y155_DLUT (
.I0(CLBLM_L_X8Y155_SLICE_X10Y155_CO6),
.I1(CLBLM_L_X8Y153_SLICE_X11Y153_BQ),
.I2(CLBLM_L_X8Y155_SLICE_X11Y155_DO6),
.I3(CLBLM_L_X8Y155_SLICE_X11Y155_CO6),
.I4(CLBLM_L_X10Y154_SLICE_X12Y154_AQ),
.I5(CLBLM_L_X8Y154_SLICE_X11Y154_DO6),
.O5(CLBLM_L_X10Y155_SLICE_X12Y155_DO5),
.O6(CLBLM_L_X10Y155_SLICE_X12Y155_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555151555551155)
  ) CLBLM_L_X10Y155_SLICE_X12Y155_CLUT (
.I0(CLBLM_L_X8Y155_SLICE_X10Y155_CO6),
.I1(CLBLM_L_X8Y153_SLICE_X10Y153_BQ),
.I2(CLBLM_L_X10Y155_SLICE_X13Y155_DO6),
.I3(CLBLM_L_X10Y156_SLICE_X12Y156_AO5),
.I4(CLBLM_L_X8Y154_SLICE_X11Y154_DO6),
.I5(CLBLM_L_X10Y155_SLICE_X13Y155_BQ),
.O5(CLBLM_L_X10Y155_SLICE_X12Y155_CO5),
.O6(CLBLM_L_X10Y155_SLICE_X12Y155_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0000ffff00e01f)
  ) CLBLM_L_X10Y155_SLICE_X12Y155_BLUT (
.I0(CLBLM_L_X10Y156_SLICE_X12Y156_AO5),
.I1(CLBLM_L_X10Y155_SLICE_X13Y155_DO6),
.I2(CLBLM_L_X10Y153_SLICE_X13Y153_AQ),
.I3(CLBLM_L_X10Y155_SLICE_X13Y155_BQ),
.I4(CLBLM_L_X8Y155_SLICE_X10Y155_CO6),
.I5(CLBLM_L_X8Y154_SLICE_X11Y154_DO6),
.O5(CLBLM_L_X10Y155_SLICE_X12Y155_BO5),
.O6(CLBLM_L_X10Y155_SLICE_X12Y155_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0aaa0fff0a0a0f0f)
  ) CLBLM_L_X10Y155_SLICE_X12Y155_ALUT (
.I0(CLBLM_L_X10Y150_SLICE_X12Y150_B5Q),
.I1(1'b1),
.I2(CLBLM_L_X8Y153_SLICE_X10Y153_CO5),
.I3(CLBLM_L_X10Y156_SLICE_X12Y156_BO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y153_SLICE_X10Y153_DO6),
.O5(CLBLM_L_X10Y155_SLICE_X12Y155_AO5),
.O6(CLBLM_L_X10Y155_SLICE_X12Y155_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y155_SLICE_X13Y155_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y155_SLICE_X13Y155_AO6),
.Q(CLBLM_L_X10Y155_SLICE_X13Y155_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y155_SLICE_X13Y155_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y155_SLICE_X13Y155_BO6),
.Q(CLBLM_L_X10Y155_SLICE_X13Y155_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y155_SLICE_X13Y155_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y155_SLICE_X13Y155_CO6),
.Q(CLBLM_L_X10Y155_SLICE_X13Y155_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hc000c00000000000)
  ) CLBLM_L_X10Y155_SLICE_X13Y155_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y154_SLICE_X12Y154_DQ),
.I2(CLBLM_L_X8Y153_SLICE_X11Y153_BQ),
.I3(CLBLM_L_X8Y155_SLICE_X10Y155_AQ),
.I4(1'b1),
.I5(CLBLM_L_X8Y155_SLICE_X11Y155_CO6),
.O5(CLBLM_L_X10Y155_SLICE_X13Y155_DO5),
.O6(CLBLM_L_X10Y155_SLICE_X13Y155_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hd0507050dd557755)
  ) CLBLM_L_X10Y155_SLICE_X13Y155_CLUT (
.I0(CLBLM_L_X8Y153_SLICE_X10Y153_CO5),
.I1(CLBLM_L_X10Y155_SLICE_X12Y155_CO6),
.I2(CLBLM_R_X11Y148_SLICE_X15Y148_CQ),
.I3(CLBLM_L_X8Y153_SLICE_X10Y153_DO6),
.I4(CLBLM_L_X10Y155_SLICE_X13Y155_CQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y155_SLICE_X13Y155_CO5),
.O6(CLBLM_L_X10Y155_SLICE_X13Y155_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3033f0ff0000f0ff)
  ) CLBLM_L_X10Y155_SLICE_X13Y155_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y155_SLICE_X12Y155_BO6),
.I2(CLBLM_L_X10Y154_SLICE_X13Y154_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y153_SLICE_X10Y153_CO5),
.I5(CLBLM_L_X8Y153_SLICE_X10Y153_DO6),
.O5(CLBLM_L_X10Y155_SLICE_X13Y155_BO5),
.O6(CLBLM_L_X10Y155_SLICE_X13Y155_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hb8b8b8b8bbb8bbb8)
  ) CLBLM_L_X10Y155_SLICE_X13Y155_ALUT (
.I0(CLBLM_L_X10Y155_SLICE_X13Y155_CQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y155_SLICE_X13Y155_AQ),
.I3(RIOB33_X105Y141_IOB_X1Y142_I),
.I4(1'b1),
.I5(CLBLM_R_X5Y142_SLICE_X7Y142_AQ),
.O5(CLBLM_L_X10Y155_SLICE_X13Y155_AO5),
.O6(CLBLM_L_X10Y155_SLICE_X13Y155_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_L_X10Y156_SLICE_X12Y156_DLUT (
.I0(CLBLM_L_X8Y155_SLICE_X11Y155_CO6),
.I1(CLBLM_L_X10Y154_SLICE_X12Y154_DQ),
.I2(CLBLM_L_X8Y153_SLICE_X11Y153_BQ),
.I3(CLBLM_L_X10Y155_SLICE_X13Y155_CQ),
.I4(CLBLM_L_X8Y155_SLICE_X10Y155_AQ),
.I5(CLBLM_L_X10Y155_SLICE_X13Y155_BQ),
.O5(CLBLM_L_X10Y156_SLICE_X12Y156_DO5),
.O6(CLBLM_L_X10Y156_SLICE_X12Y156_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0c000a0a00000a0a)
  ) CLBLM_L_X10Y156_SLICE_X12Y156_CLUT (
.I0(CLBLM_L_X10Y156_SLICE_X12Y156_AO6),
.I1(CLBLM_L_X10Y155_SLICE_X13Y155_CQ),
.I2(CLBLM_L_X8Y154_SLICE_X11Y154_DO6),
.I3(CLBLM_L_X10Y155_SLICE_X13Y155_DO6),
.I4(CLBLM_L_X10Y155_SLICE_X12Y155_AQ),
.I5(CLBLM_L_X10Y155_SLICE_X13Y155_BQ),
.O5(CLBLM_L_X10Y156_SLICE_X12Y156_CO5),
.O6(CLBLM_L_X10Y156_SLICE_X12Y156_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc3ccc39cc33cc33)
  ) CLBLM_L_X10Y156_SLICE_X12Y156_BLUT (
.I0(CLBLM_L_X10Y156_SLICE_X12Y156_DO6),
.I1(CLBLM_L_X10Y155_SLICE_X12Y155_AQ),
.I2(CLBLM_L_X8Y154_SLICE_X11Y154_DO6),
.I3(CLBLM_L_X8Y155_SLICE_X10Y155_CO6),
.I4(CLBLM_L_X10Y156_SLICE_X12Y156_AO6),
.I5(CLBLM_L_X8Y153_SLICE_X10Y153_AQ),
.O5(CLBLM_L_X10Y156_SLICE_X12Y156_BO5),
.O6(CLBLM_L_X10Y156_SLICE_X12Y156_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000202020202)
  ) CLBLM_L_X10Y156_SLICE_X12Y156_ALUT (
.I0(CLBLM_L_X8Y155_SLICE_X11Y155_DO6),
.I1(CLBLM_L_X8Y155_SLICE_X10Y155_AQ),
.I2(CLBLM_L_X10Y154_SLICE_X12Y154_DQ),
.I3(CLBLM_L_X10Y155_SLICE_X13Y155_BQ),
.I4(CLBLM_L_X10Y155_SLICE_X13Y155_CQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y156_SLICE_X12Y156_AO5),
.O6(CLBLM_L_X10Y156_SLICE_X12Y156_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y156_SLICE_X13Y156_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y156_SLICE_X13Y156_DO5),
.O6(CLBLM_L_X10Y156_SLICE_X13Y156_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y156_SLICE_X13Y156_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y156_SLICE_X13Y156_CO5),
.O6(CLBLM_L_X10Y156_SLICE_X13Y156_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y156_SLICE_X13Y156_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y156_SLICE_X13Y156_BO5),
.O6(CLBLM_L_X10Y156_SLICE_X13Y156_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y156_SLICE_X13Y156_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y156_SLICE_X13Y156_AO5),
.O6(CLBLM_L_X10Y156_SLICE_X13Y156_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y144_SLICE_X16Y144_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y144_SLICE_X16Y144_AO6),
.Q(CLBLM_L_X12Y144_SLICE_X16Y144_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y144_SLICE_X16Y144_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y144_SLICE_X16Y144_BO6),
.Q(CLBLM_L_X12Y144_SLICE_X16Y144_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y144_SLICE_X16Y144_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y144_SLICE_X16Y144_CO6),
.Q(CLBLM_L_X12Y144_SLICE_X16Y144_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8f0fffff44000000)
  ) CLBLM_L_X12Y144_SLICE_X16Y144_DLUT (
.I0(CLBLM_L_X12Y145_SLICE_X16Y145_AQ),
.I1(CLBLM_L_X12Y144_SLICE_X16Y144_CQ),
.I2(CLBLM_R_X7Y142_SLICE_X8Y142_DO6),
.I3(CLBLM_L_X12Y144_SLICE_X16Y144_AQ),
.I4(CLBLM_L_X12Y144_SLICE_X16Y144_BQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y144_SLICE_X16Y144_DO5),
.O6(CLBLM_L_X12Y144_SLICE_X16Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff40ff1000400010)
  ) CLBLM_L_X12Y144_SLICE_X16Y144_CLUT (
.I0(CLBLM_L_X10Y152_SLICE_X12Y152_DQ),
.I1(CLBLM_L_X12Y144_SLICE_X16Y144_CQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X12Y144_SLICE_X16Y144_DO6),
.I5(CLBLM_L_X12Y154_SLICE_X16Y154_AQ),
.O5(CLBLM_L_X12Y144_SLICE_X16Y144_CO5),
.O6(CLBLM_L_X12Y144_SLICE_X16Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffa8a8a8ff000000)
  ) CLBLM_L_X12Y144_SLICE_X16Y144_BLUT (
.I0(CLBLM_L_X12Y144_SLICE_X16Y144_DO6),
.I1(CLBLM_L_X12Y144_SLICE_X16Y144_BQ),
.I2(CLBLM_R_X7Y142_SLICE_X8Y142_DO6),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y144_SLICE_X12Y144_AQ),
.I5(CLBLM_L_X12Y144_SLICE_X16Y144_AO5),
.O5(CLBLM_L_X12Y144_SLICE_X16Y144_BO5),
.O6(CLBLM_L_X12Y144_SLICE_X16Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a3a003000300)
  ) CLBLM_L_X12Y144_SLICE_X16Y144_ALUT (
.I0(CLBLM_R_X3Y145_SLICE_X2Y145_AQ),
.I1(CLBLM_L_X10Y152_SLICE_X12Y152_DQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_L_X12Y145_SLICE_X16Y145_CO5),
.I5(1'b1),
.O5(CLBLM_L_X12Y144_SLICE_X16Y144_AO5),
.O6(CLBLM_L_X12Y144_SLICE_X16Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y144_SLICE_X17Y144_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y144_SLICE_X17Y144_DO5),
.O6(CLBLM_L_X12Y144_SLICE_X17Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y144_SLICE_X17Y144_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y144_SLICE_X17Y144_CO5),
.O6(CLBLM_L_X12Y144_SLICE_X17Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y144_SLICE_X17Y144_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y144_SLICE_X17Y144_BO5),
.O6(CLBLM_L_X12Y144_SLICE_X17Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y144_SLICE_X17Y144_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y144_SLICE_X17Y144_AO5),
.O6(CLBLM_L_X12Y144_SLICE_X17Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y145_SLICE_X16Y145_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y145_SLICE_X16Y145_AO6),
.Q(CLBLM_L_X12Y145_SLICE_X16Y145_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y145_SLICE_X16Y145_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y145_SLICE_X16Y145_BO6),
.Q(CLBLM_L_X12Y145_SLICE_X16Y145_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y145_SLICE_X16Y145_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y145_SLICE_X16Y145_DO5),
.O6(CLBLM_L_X12Y145_SLICE_X16Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h2000000020005fff)
  ) CLBLM_L_X12Y145_SLICE_X16Y145_CLUT (
.I0(CLBLM_L_X12Y144_SLICE_X16Y144_BQ),
.I1(CLBLM_L_X12Y145_SLICE_X16Y145_AQ),
.I2(CLBLM_R_X7Y142_SLICE_X8Y142_DO6),
.I3(CLBLM_L_X12Y144_SLICE_X16Y144_CQ),
.I4(CLBLM_L_X12Y144_SLICE_X16Y144_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y145_SLICE_X16Y145_CO5),
.O6(CLBLM_L_X12Y145_SLICE_X16Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf055f044f055f044)
  ) CLBLM_L_X12Y145_SLICE_X16Y145_BLUT (
.I0(CLBLL_L_X4Y145_SLICE_X5Y145_DO6),
.I1(CLBLM_L_X12Y145_SLICE_X16Y145_BQ),
.I2(CLBLM_R_X11Y152_SLICE_X14Y152_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X11Y145_SLICE_X14Y145_BQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y145_SLICE_X16Y145_BO5),
.O6(CLBLM_L_X12Y145_SLICE_X16Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00ee44aa00ea40)
  ) CLBLM_L_X12Y145_SLICE_X16Y145_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_L_X12Y145_SLICE_X16Y145_AQ),
.I3(CLBLM_R_X7Y142_SLICE_X8Y142_BQ),
.I4(CLBLM_L_X10Y152_SLICE_X12Y152_DQ),
.I5(CLBLM_L_X12Y145_SLICE_X16Y145_CO6),
.O5(CLBLM_L_X12Y145_SLICE_X16Y145_AO5),
.O6(CLBLM_L_X12Y145_SLICE_X16Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y145_SLICE_X17Y145_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y145_SLICE_X17Y145_DO5),
.O6(CLBLM_L_X12Y145_SLICE_X17Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y145_SLICE_X17Y145_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y145_SLICE_X17Y145_CO5),
.O6(CLBLM_L_X12Y145_SLICE_X17Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y145_SLICE_X17Y145_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y145_SLICE_X17Y145_BO5),
.O6(CLBLM_L_X12Y145_SLICE_X17Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y145_SLICE_X17Y145_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y145_SLICE_X17Y145_AO5),
.O6(CLBLM_L_X12Y145_SLICE_X17Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y146_SLICE_X16Y146_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y146_SLICE_X16Y146_AO6),
.Q(CLBLM_L_X12Y146_SLICE_X16Y146_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y146_SLICE_X16Y146_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y146_SLICE_X16Y146_DO5),
.O6(CLBLM_L_X12Y146_SLICE_X16Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y146_SLICE_X16Y146_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y146_SLICE_X16Y146_CO5),
.O6(CLBLM_L_X12Y146_SLICE_X16Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y146_SLICE_X16Y146_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y146_SLICE_X16Y146_BO5),
.O6(CLBLM_L_X12Y146_SLICE_X16Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa33003000)
  ) CLBLM_L_X12Y146_SLICE_X16Y146_ALUT (
.I0(CLBLM_R_X11Y146_SLICE_X15Y146_CQ),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_L_X12Y146_SLICE_X16Y146_AQ),
.I3(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.I4(CLBLM_L_X10Y143_SLICE_X13Y143_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X12Y146_SLICE_X16Y146_AO5),
.O6(CLBLM_L_X12Y146_SLICE_X16Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y146_SLICE_X17Y146_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y146_SLICE_X17Y146_DO5),
.O6(CLBLM_L_X12Y146_SLICE_X17Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y146_SLICE_X17Y146_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y146_SLICE_X17Y146_CO5),
.O6(CLBLM_L_X12Y146_SLICE_X17Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y146_SLICE_X17Y146_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y146_SLICE_X17Y146_BO5),
.O6(CLBLM_L_X12Y146_SLICE_X17Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y146_SLICE_X17Y146_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y146_SLICE_X17Y146_AO5),
.O6(CLBLM_L_X12Y146_SLICE_X17Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y147_SLICE_X16Y147_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y147_SLICE_X16Y147_AO6),
.Q(CLBLM_L_X12Y147_SLICE_X16Y147_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y147_SLICE_X16Y147_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y147_SLICE_X16Y147_DO5),
.O6(CLBLM_L_X12Y147_SLICE_X16Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y147_SLICE_X16Y147_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y147_SLICE_X16Y147_CO5),
.O6(CLBLM_L_X12Y147_SLICE_X16Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y147_SLICE_X16Y147_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y147_SLICE_X16Y147_BO5),
.O6(CLBLM_L_X12Y147_SLICE_X16Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hddddddd8888888d8)
  ) CLBLM_L_X12Y147_SLICE_X16Y147_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y151_SLICE_X13Y151_CQ),
.I2(CLBLM_L_X12Y147_SLICE_X16Y147_AQ),
.I3(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLM_L_X12Y146_SLICE_X16Y146_AQ),
.O5(CLBLM_L_X12Y147_SLICE_X16Y147_AO5),
.O6(CLBLM_L_X12Y147_SLICE_X16Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y147_SLICE_X17Y147_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y147_SLICE_X17Y147_DO5),
.O6(CLBLM_L_X12Y147_SLICE_X17Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y147_SLICE_X17Y147_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y147_SLICE_X17Y147_CO5),
.O6(CLBLM_L_X12Y147_SLICE_X17Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y147_SLICE_X17Y147_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y147_SLICE_X17Y147_BO5),
.O6(CLBLM_L_X12Y147_SLICE_X17Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y147_SLICE_X17Y147_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y147_SLICE_X17Y147_AO5),
.O6(CLBLM_L_X12Y147_SLICE_X17Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y148_SLICE_X16Y148_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y148_SLICE_X16Y148_AO6),
.Q(CLBLM_L_X12Y148_SLICE_X16Y148_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y148_SLICE_X16Y148_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y148_SLICE_X16Y148_BO6),
.Q(CLBLM_L_X12Y148_SLICE_X16Y148_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y148_SLICE_X16Y148_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y148_SLICE_X16Y148_DO5),
.O6(CLBLM_L_X12Y148_SLICE_X16Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h55aaaa55aa5555aa)
  ) CLBLM_L_X12Y148_SLICE_X16Y148_CLUT (
.I0(CLBLM_L_X8Y144_SLICE_X10Y144_AQ),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_L_X8Y151_SLICE_X11Y151_CQ),
.I4(CLBLM_L_X10Y145_SLICE_X12Y145_BQ),
.I5(CLBLL_L_X4Y148_SLICE_X5Y148_BQ),
.O5(CLBLM_L_X12Y148_SLICE_X16Y148_CO5),
.O6(CLBLM_L_X12Y148_SLICE_X16Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'he4f5e4a0a0f5a0a0)
  ) CLBLM_L_X12Y148_SLICE_X16Y148_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X12Y148_SLICE_X16Y148_BQ),
.I2(CLBLM_L_X12Y150_SLICE_X16Y150_AQ),
.I3(CLBLM_R_X11Y147_SLICE_X14Y147_CO6),
.I4(CLBLM_L_X12Y149_SLICE_X16Y149_AQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X12Y148_SLICE_X16Y148_BO5),
.O6(CLBLM_L_X12Y148_SLICE_X16Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccf0cc00ccaaccaa)
  ) CLBLM_L_X12Y148_SLICE_X16Y148_ALUT (
.I0(CLBLM_L_X10Y151_SLICE_X12Y151_BQ),
.I1(CLBLM_L_X10Y152_SLICE_X12Y152_DQ),
.I2(CLBLM_L_X12Y148_SLICE_X16Y148_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X11Y147_SLICE_X14Y147_CO6),
.O5(CLBLM_L_X12Y148_SLICE_X16Y148_AO5),
.O6(CLBLM_L_X12Y148_SLICE_X16Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y148_SLICE_X17Y148_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y148_SLICE_X17Y148_DO5),
.O6(CLBLM_L_X12Y148_SLICE_X17Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y148_SLICE_X17Y148_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y148_SLICE_X17Y148_CO5),
.O6(CLBLM_L_X12Y148_SLICE_X17Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y148_SLICE_X17Y148_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y148_SLICE_X17Y148_BO5),
.O6(CLBLM_L_X12Y148_SLICE_X17Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y148_SLICE_X17Y148_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y148_SLICE_X17Y148_AO5),
.O6(CLBLM_L_X12Y148_SLICE_X17Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y149_SLICE_X16Y149_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y149_SLICE_X16Y149_AO6),
.Q(CLBLM_L_X12Y149_SLICE_X16Y149_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7dbe7dbe7dbe7dbe)
  ) CLBLM_L_X12Y149_SLICE_X16Y149_DLUT (
.I0(CLBLM_R_X7Y146_SLICE_X9Y146_BQ),
.I1(CLBLL_L_X4Y148_SLICE_X5Y148_BQ),
.I2(CLBLM_L_X10Y151_SLICE_X12Y151_BQ),
.I3(CLBLM_L_X12Y149_SLICE_X17Y149_CQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y149_SLICE_X16Y149_DO5),
.O6(CLBLM_L_X12Y149_SLICE_X16Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5ff55ff5affaaffa)
  ) CLBLM_L_X12Y149_SLICE_X16Y149_CLUT (
.I0(CLBLM_L_X12Y150_SLICE_X16Y150_BQ),
.I1(1'b1),
.I2(CLBLM_L_X8Y151_SLICE_X11Y151_CQ),
.I3(CLBLM_L_X10Y150_SLICE_X12Y150_AQ),
.I4(1'b1),
.I5(CLBLM_L_X8Y144_SLICE_X10Y144_AQ),
.O5(CLBLM_L_X12Y149_SLICE_X16Y149_CO5),
.O6(CLBLM_L_X12Y149_SLICE_X16Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffaaffffaa)
  ) CLBLM_L_X12Y149_SLICE_X16Y149_BLUT (
.I0(CLBLM_L_X12Y149_SLICE_X16Y149_DO6),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X11Y149_SLICE_X14Y149_AQ),
.I4(CLBLM_L_X10Y145_SLICE_X12Y145_BQ),
.I5(CLBLM_L_X12Y149_SLICE_X16Y149_CO6),
.O5(CLBLM_L_X12Y149_SLICE_X16Y149_BO5),
.O6(CLBLM_L_X12Y149_SLICE_X16Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaf3aa33aac0aa00)
  ) CLBLM_L_X12Y149_SLICE_X16Y149_ALUT (
.I0(CLBLL_L_X4Y143_SLICE_X4Y143_BQ),
.I1(CLBLM_R_X11Y147_SLICE_X14Y147_CO6),
.I2(CLBLM_L_X12Y149_SLICE_X16Y149_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_L_X12Y149_SLICE_X17Y149_CQ),
.O5(CLBLM_L_X12Y149_SLICE_X16Y149_AO5),
.O6(CLBLM_L_X12Y149_SLICE_X16Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y149_SLICE_X17Y149_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y149_SLICE_X17Y149_AO6),
.Q(CLBLM_L_X12Y149_SLICE_X17Y149_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y149_SLICE_X17Y149_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y149_SLICE_X17Y149_BO6),
.Q(CLBLM_L_X12Y149_SLICE_X17Y149_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y149_SLICE_X17Y149_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y149_SLICE_X17Y149_CO6),
.Q(CLBLM_L_X12Y149_SLICE_X17Y149_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y149_SLICE_X17Y149_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y149_SLICE_X17Y149_DO5),
.O6(CLBLM_L_X12Y149_SLICE_X17Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc0cf000fa0afa0a)
  ) CLBLM_L_X12Y149_SLICE_X17Y149_CLUT (
.I0(CLBLM_L_X12Y150_SLICE_X16Y150_BQ),
.I1(CLBLM_L_X12Y149_SLICE_X17Y149_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y151_SLICE_X9Y151_AQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X11Y147_SLICE_X14Y147_CO6),
.O5(CLBLM_L_X12Y149_SLICE_X17Y149_CO5),
.O6(CLBLM_L_X12Y149_SLICE_X17Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hacafa0afaca0a0a0)
  ) CLBLM_L_X12Y149_SLICE_X17Y149_BLUT (
.I0(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.I1(CLBLM_L_X12Y149_SLICE_X17Y149_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X11Y147_SLICE_X14Y147_CO6),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_L_X12Y149_SLICE_X17Y149_AQ),
.O5(CLBLM_L_X12Y149_SLICE_X17Y149_BO5),
.O6(CLBLM_L_X12Y149_SLICE_X17Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hafa0acaca0a0acac)
  ) CLBLM_L_X12Y149_SLICE_X17Y149_ALUT (
.I0(CLBLM_R_X11Y152_SLICE_X14Y152_DQ),
.I1(CLBLM_L_X12Y148_SLICE_X16Y148_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X11Y147_SLICE_X14Y147_CO6),
.I5(CLBLM_L_X12Y149_SLICE_X17Y149_AQ),
.O5(CLBLM_L_X12Y149_SLICE_X17Y149_AO5),
.O6(CLBLM_L_X12Y149_SLICE_X17Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y150_SLICE_X16Y150_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X12Y150_SLICE_X16Y150_AO6),
.Q(CLBLM_L_X12Y150_SLICE_X16Y150_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y150_SLICE_X16Y150_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X12Y150_SLICE_X16Y150_BO6),
.Q(CLBLM_L_X12Y150_SLICE_X16Y150_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y150_SLICE_X16Y150_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X12Y150_SLICE_X16Y150_CO6),
.Q(CLBLM_L_X12Y150_SLICE_X16Y150_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0aaf0aa03030000)
  ) CLBLM_L_X12Y150_SLICE_X16Y150_DLUT (
.I0(CLBLM_L_X10Y149_SLICE_X13Y149_A5Q),
.I1(CLBLM_R_X11Y151_SLICE_X15Y151_A5Q),
.I2(CLBLM_L_X12Y151_SLICE_X16Y151_BQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y147_SLICE_X9Y147_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y150_SLICE_X16Y150_DO5),
.O6(CLBLM_L_X12Y150_SLICE_X16Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa03aa00aa0caa0c)
  ) CLBLM_L_X12Y150_SLICE_X16Y150_CLUT (
.I0(CLBLM_R_X11Y150_SLICE_X15Y150_CQ),
.I1(CLBLM_L_X12Y150_SLICE_X16Y150_CQ),
.I2(CLBLM_R_X11Y154_SLICE_X15Y154_CO6),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X12Y151_SLICE_X16Y151_CQ),
.I5(CLBLM_L_X12Y150_SLICE_X16Y150_DO5),
.O5(CLBLM_L_X12Y150_SLICE_X16Y150_CO5),
.O6(CLBLM_L_X12Y150_SLICE_X16Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hee44aa00fa50fa50)
  ) CLBLM_L_X12Y150_SLICE_X16Y150_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X12Y150_SLICE_X16Y150_BQ),
.I2(CLBLM_L_X12Y148_SLICE_X16Y148_AQ),
.I3(CLBLM_L_X12Y152_SLICE_X17Y152_BQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X11Y147_SLICE_X14Y147_CO6),
.O5(CLBLM_L_X12Y150_SLICE_X16Y150_BO5),
.O6(CLBLM_L_X12Y150_SLICE_X16Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00ccccd8d8)
  ) CLBLM_L_X12Y150_SLICE_X16Y150_ALUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_R_X11Y150_SLICE_X15Y150_CQ),
.I2(CLBLM_L_X12Y150_SLICE_X16Y150_AQ),
.I3(CLBLM_L_X12Y151_SLICE_X16Y151_AQ),
.I4(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X12Y150_SLICE_X16Y150_AO5),
.O6(CLBLM_L_X12Y150_SLICE_X16Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y150_SLICE_X17Y150_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y150_SLICE_X17Y150_DO5),
.O6(CLBLM_L_X12Y150_SLICE_X17Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y150_SLICE_X17Y150_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y150_SLICE_X17Y150_CO5),
.O6(CLBLM_L_X12Y150_SLICE_X17Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y150_SLICE_X17Y150_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y150_SLICE_X17Y150_BO5),
.O6(CLBLM_L_X12Y150_SLICE_X17Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y150_SLICE_X17Y150_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y150_SLICE_X17Y150_AO5),
.O6(CLBLM_L_X12Y150_SLICE_X17Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y151_SLICE_X16Y151_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X12Y151_SLICE_X16Y151_AO6),
.Q(CLBLM_L_X12Y151_SLICE_X16Y151_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y151_SLICE_X16Y151_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X12Y151_SLICE_X16Y151_BO6),
.Q(CLBLM_L_X12Y151_SLICE_X16Y151_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y151_SLICE_X16Y151_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X12Y151_SLICE_X16Y151_CO6),
.Q(CLBLM_L_X12Y151_SLICE_X16Y151_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0010001000000010)
  ) CLBLM_L_X12Y151_SLICE_X16Y151_DLUT (
.I0(CLBLM_L_X12Y151_SLICE_X16Y151_BQ),
.I1(CLBLM_R_X11Y151_SLICE_X15Y151_A5Q),
.I2(CLBLM_R_X7Y147_SLICE_X9Y147_AQ),
.I3(CLBLM_L_X12Y150_SLICE_X16Y150_CQ),
.I4(CLBLM_L_X12Y151_SLICE_X16Y151_CQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y151_SLICE_X16Y151_DO5),
.O6(CLBLM_L_X12Y151_SLICE_X16Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaf3f3fcfc)
  ) CLBLM_L_X12Y151_SLICE_X16Y151_CLUT (
.I0(CLBLL_L_X4Y149_SLICE_X4Y149_AQ),
.I1(CLBLM_L_X12Y151_SLICE_X16Y151_CQ),
.I2(CLBLM_R_X11Y154_SLICE_X15Y154_CO6),
.I3(1'b1),
.I4(CLBLM_L_X12Y151_SLICE_X16Y151_DO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X12Y151_SLICE_X16Y151_CO5),
.O6(CLBLM_L_X12Y151_SLICE_X16Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f000110044)
  ) CLBLM_L_X12Y151_SLICE_X16Y151_BLUT (
.I0(CLBLM_R_X11Y154_SLICE_X15Y154_CO6),
.I1(CLBLM_R_X11Y151_SLICE_X14Y151_AO5),
.I2(CLBLM_R_X11Y151_SLICE_X14Y151_BQ),
.I3(CLBLM_L_X12Y151_SLICE_X16Y151_DO5),
.I4(CLBLM_L_X12Y151_SLICE_X16Y151_BQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X12Y151_SLICE_X16Y151_BO5),
.O6(CLBLM_L_X12Y151_SLICE_X16Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff0fffa00f000fa)
  ) CLBLM_L_X12Y151_SLICE_X16Y151_ALUT (
.I0(RIOB33_X105Y141_IOB_X1Y142_I),
.I1(1'b1),
.I2(CLBLM_L_X12Y151_SLICE_X16Y151_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X5Y142_SLICE_X7Y142_AQ),
.I5(CLBLM_L_X8Y152_SLICE_X10Y152_CQ),
.O5(CLBLM_L_X12Y151_SLICE_X16Y151_AO5),
.O6(CLBLM_L_X12Y151_SLICE_X16Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000010001)
  ) CLBLM_L_X12Y151_SLICE_X17Y151_DLUT (
.I0(CLBLM_L_X12Y154_SLICE_X16Y154_AQ),
.I1(CLBLM_L_X12Y152_SLICE_X16Y152_AQ),
.I2(CLBLM_L_X12Y153_SLICE_X17Y153_DO6),
.I3(CLBLM_L_X12Y153_SLICE_X16Y153_AQ),
.I4(1'b1),
.I5(CLBLM_L_X12Y152_SLICE_X17Y152_BQ),
.O5(CLBLM_L_X12Y151_SLICE_X17Y151_DO5),
.O6(CLBLM_L_X12Y151_SLICE_X17Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h4b5a5a5a4b5a4b5a)
  ) CLBLM_L_X12Y151_SLICE_X17Y151_CLUT (
.I0(CLBLM_L_X12Y153_SLICE_X16Y153_DO6),
.I1(CLBLM_R_X11Y153_SLICE_X14Y153_CO5),
.I2(CLBLM_L_X12Y152_SLICE_X17Y152_CQ),
.I3(CLBLM_L_X10Y151_SLICE_X13Y151_CQ),
.I4(CLBLM_L_X12Y151_SLICE_X17Y151_DO6),
.I5(CLBLM_R_X13Y151_SLICE_X18Y151_CO6),
.O5(CLBLM_L_X12Y151_SLICE_X17Y151_CO5),
.O6(CLBLM_L_X12Y151_SLICE_X17Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h33333333c9ccc3cc)
  ) CLBLM_L_X12Y151_SLICE_X17Y151_BLUT (
.I0(CLBLM_R_X13Y151_SLICE_X18Y151_AO6),
.I1(CLBLM_L_X12Y152_SLICE_X17Y152_BQ),
.I2(CLBLM_R_X11Y153_SLICE_X14Y153_CO5),
.I3(CLBLM_R_X11Y152_SLICE_X14Y152_BQ),
.I4(CLBLM_R_X13Y151_SLICE_X18Y151_BO6),
.I5(CLBLM_L_X12Y153_SLICE_X16Y153_DO6),
.O5(CLBLM_L_X12Y151_SLICE_X17Y151_BO5),
.O6(CLBLM_L_X12Y151_SLICE_X17Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3332303233333333)
  ) CLBLM_L_X12Y151_SLICE_X17Y151_ALUT (
.I0(CLBLM_R_X13Y151_SLICE_X18Y151_AO6),
.I1(CLBLM_L_X12Y153_SLICE_X16Y153_DO6),
.I2(CLBLM_R_X11Y153_SLICE_X14Y153_CO5),
.I3(CLBLM_L_X12Y152_SLICE_X17Y152_BQ),
.I4(CLBLM_R_X13Y151_SLICE_X18Y151_BO6),
.I5(CLBLM_R_X11Y152_SLICE_X14Y152_CQ),
.O5(CLBLM_L_X12Y151_SLICE_X17Y151_AO5),
.O6(CLBLM_L_X12Y151_SLICE_X17Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y152_SLICE_X16Y152_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X12Y152_SLICE_X16Y152_AO6),
.Q(CLBLM_L_X12Y152_SLICE_X16Y152_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y152_SLICE_X16Y152_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X12Y152_SLICE_X16Y152_BO6),
.Q(CLBLM_L_X12Y152_SLICE_X16Y152_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h55aa55aa45ba15ea)
  ) CLBLM_L_X12Y152_SLICE_X16Y152_DLUT (
.I0(CLBLM_L_X12Y153_SLICE_X16Y153_DO6),
.I1(CLBLM_R_X11Y153_SLICE_X15Y153_AQ),
.I2(CLBLM_L_X10Y152_SLICE_X12Y152_BQ),
.I3(CLBLM_L_X12Y152_SLICE_X16Y152_BQ),
.I4(CLBLM_L_X12Y154_SLICE_X16Y154_BO5),
.I5(CLBLM_R_X11Y153_SLICE_X14Y153_CO5),
.O5(CLBLM_L_X12Y152_SLICE_X16Y152_DO5),
.O6(CLBLM_L_X12Y152_SLICE_X16Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5554445455555555)
  ) CLBLM_L_X12Y152_SLICE_X16Y152_CLUT (
.I0(CLBLM_L_X12Y153_SLICE_X16Y153_DO6),
.I1(CLBLM_R_X11Y153_SLICE_X14Y153_CO5),
.I2(CLBLM_L_X12Y153_SLICE_X17Y153_DO6),
.I3(CLBLM_L_X12Y153_SLICE_X16Y153_AQ),
.I4(CLBLM_L_X12Y153_SLICE_X17Y153_CO6),
.I5(CLBLM_L_X10Y152_SLICE_X13Y152_BQ),
.O5(CLBLM_L_X12Y152_SLICE_X16Y152_CO5),
.O6(CLBLM_L_X12Y152_SLICE_X16Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff32ff3200320032)
  ) CLBLM_L_X12Y152_SLICE_X16Y152_BLUT (
.I0(CLBLM_L_X12Y152_SLICE_X16Y152_DO6),
.I1(CLBLM_R_X11Y154_SLICE_X15Y154_CO5),
.I2(CLBLM_L_X10Y154_SLICE_X13Y154_CO5),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLM_R_X11Y147_SLICE_X15Y147_CQ),
.O5(CLBLM_L_X12Y152_SLICE_X16Y152_BO5),
.O6(CLBLM_L_X12Y152_SLICE_X16Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00fe54ef45)
  ) CLBLM_L_X12Y152_SLICE_X16Y152_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y154_SLICE_X13Y154_CO5),
.I2(CLBLM_L_X12Y152_SLICE_X16Y152_AQ),
.I3(CLBLM_R_X7Y152_SLICE_X9Y152_CQ),
.I4(CLBLM_L_X12Y151_SLICE_X17Y151_AO6),
.I5(CLBLM_R_X11Y154_SLICE_X15Y154_CO5),
.O5(CLBLM_L_X12Y152_SLICE_X16Y152_AO5),
.O6(CLBLM_L_X12Y152_SLICE_X16Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y152_SLICE_X17Y152_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X12Y152_SLICE_X17Y152_AO6),
.Q(CLBLM_L_X12Y152_SLICE_X17Y152_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y152_SLICE_X17Y152_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X12Y152_SLICE_X17Y152_BO6),
.Q(CLBLM_L_X12Y152_SLICE_X17Y152_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y152_SLICE_X17Y152_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X12Y152_SLICE_X17Y152_CO6),
.Q(CLBLM_L_X12Y152_SLICE_X17Y152_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555555551555515)
  ) CLBLM_L_X12Y152_SLICE_X17Y152_DLUT (
.I0(CLBLM_L_X12Y153_SLICE_X16Y153_DO6),
.I1(CLBLM_R_X11Y152_SLICE_X14Y152_DQ),
.I2(CLBLM_L_X12Y154_SLICE_X16Y154_BO5),
.I3(CLBLM_R_X11Y153_SLICE_X15Y153_AQ),
.I4(CLBLM_L_X12Y152_SLICE_X16Y152_BQ),
.I5(CLBLM_R_X11Y153_SLICE_X14Y153_CO5),
.O5(CLBLM_L_X12Y152_SLICE_X17Y152_DO5),
.O6(CLBLM_L_X12Y152_SLICE_X17Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0ff000ff0fa000a)
  ) CLBLM_L_X12Y152_SLICE_X17Y152_CLUT (
.I0(CLBLM_L_X10Y154_SLICE_X13Y154_CO5),
.I1(1'b1),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X11Y154_SLICE_X15Y154_CO5),
.I4(CLBLM_R_X11Y148_SLICE_X14Y148_DQ),
.I5(CLBLM_L_X12Y151_SLICE_X17Y151_CO6),
.O5(CLBLM_L_X12Y152_SLICE_X17Y152_CO5),
.O6(CLBLM_L_X12Y152_SLICE_X17Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5f5f005050500)
  ) CLBLM_L_X12Y152_SLICE_X17Y152_BLUT (
.I0(CLBLM_R_X11Y154_SLICE_X15Y154_CO5),
.I1(1'b1),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X12Y151_SLICE_X17Y151_BO6),
.I4(CLBLM_L_X10Y154_SLICE_X13Y154_CO5),
.I5(CLBLM_R_X7Y144_SLICE_X8Y144_CQ),
.O5(CLBLM_L_X12Y152_SLICE_X17Y152_BO5),
.O6(CLBLM_L_X12Y152_SLICE_X17Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5a0f5f5f5a0f5a0)
  ) CLBLM_L_X12Y152_SLICE_X17Y152_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(1'b1),
.I2(CLBLM_L_X12Y152_SLICE_X17Y152_CQ),
.I3(CLBLM_L_X12Y152_SLICE_X17Y152_AQ),
.I4(CLBLM_R_X5Y142_SLICE_X7Y142_AQ),
.I5(RIOB33_X105Y141_IOB_X1Y142_I),
.O5(CLBLM_L_X12Y152_SLICE_X17Y152_AO5),
.O6(CLBLM_L_X12Y152_SLICE_X17Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y153_SLICE_X16Y153_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X12Y153_SLICE_X16Y153_AO6),
.Q(CLBLM_L_X12Y153_SLICE_X16Y153_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7777777577777777)
  ) CLBLM_L_X12Y153_SLICE_X16Y153_DLUT (
.I0(CLBLM_L_X12Y151_SLICE_X16Y151_DO5),
.I1(CLBLM_L_X10Y153_SLICE_X13Y153_CQ),
.I2(CLBLM_L_X10Y153_SLICE_X13Y153_BQ),
.I3(CLBLM_R_X11Y154_SLICE_X15Y154_BQ),
.I4(CLBLM_R_X11Y154_SLICE_X14Y154_AQ),
.I5(CLBLM_R_X11Y154_SLICE_X15Y154_AQ),
.O5(CLBLM_L_X12Y153_SLICE_X16Y153_DO5),
.O6(CLBLM_L_X12Y153_SLICE_X16Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3b3ffffffffcfdf)
  ) CLBLM_L_X12Y153_SLICE_X16Y153_CLUT (
.I0(CLBLM_R_X11Y154_SLICE_X15Y154_AQ),
.I1(CLBLM_R_X11Y152_SLICE_X15Y152_AQ),
.I2(CLBLM_R_X11Y154_SLICE_X14Y154_AQ),
.I3(CLBLM_R_X11Y154_SLICE_X15Y154_BQ),
.I4(CLBLM_R_X11Y153_SLICE_X15Y153_AQ),
.I5(CLBLM_L_X12Y152_SLICE_X16Y152_BQ),
.O5(CLBLM_L_X12Y153_SLICE_X16Y153_CO5),
.O6(CLBLM_L_X12Y153_SLICE_X16Y153_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hdededededecfdede)
  ) CLBLM_L_X12Y153_SLICE_X16Y153_BLUT (
.I0(CLBLM_L_X12Y153_SLICE_X16Y153_DO6),
.I1(CLBLM_L_X10Y154_SLICE_X13Y154_CO5),
.I2(CLBLM_L_X12Y153_SLICE_X16Y153_AQ),
.I3(CLBLM_R_X11Y153_SLICE_X14Y153_CO5),
.I4(CLBLM_R_X11Y152_SLICE_X14Y152_AQ),
.I5(CLBLM_L_X12Y153_SLICE_X16Y153_CO6),
.O5(CLBLM_L_X12Y153_SLICE_X16Y153_BO5),
.O6(CLBLM_L_X12Y153_SLICE_X16Y153_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888bb88bb88)
  ) CLBLM_L_X12Y153_SLICE_X16Y153_ALUT (
.I0(CLBLM_R_X7Y154_SLICE_X9Y154_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(1'b1),
.I3(CLBLM_L_X12Y153_SLICE_X16Y153_BO6),
.I4(1'b1),
.I5(CLBLM_R_X11Y154_SLICE_X15Y154_CO5),
.O5(CLBLM_L_X12Y153_SLICE_X16Y153_AO5),
.O6(CLBLM_L_X12Y153_SLICE_X16Y153_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y153_SLICE_X17Y153_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X12Y153_SLICE_X17Y153_AO6),
.Q(CLBLM_L_X12Y153_SLICE_X17Y153_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffff57)
  ) CLBLM_L_X12Y153_SLICE_X17Y153_DLUT (
.I0(CLBLM_R_X11Y154_SLICE_X14Y154_AQ),
.I1(CLBLM_R_X11Y154_SLICE_X15Y154_AQ),
.I2(CLBLM_R_X11Y154_SLICE_X15Y154_BQ),
.I3(CLBLM_R_X11Y152_SLICE_X15Y152_AQ),
.I4(CLBLM_R_X11Y153_SLICE_X15Y153_AQ),
.I5(CLBLM_L_X12Y152_SLICE_X16Y152_BQ),
.O5(CLBLM_L_X12Y153_SLICE_X17Y153_DO5),
.O6(CLBLM_L_X12Y153_SLICE_X17Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3b3ffffffffffff)
  ) CLBLM_L_X12Y153_SLICE_X17Y153_CLUT (
.I0(CLBLM_R_X11Y154_SLICE_X15Y154_AQ),
.I1(CLBLM_R_X11Y153_SLICE_X15Y153_AQ),
.I2(CLBLM_R_X11Y154_SLICE_X14Y154_AQ),
.I3(CLBLM_R_X11Y154_SLICE_X15Y154_BQ),
.I4(CLBLM_R_X11Y152_SLICE_X15Y152_AQ),
.I5(CLBLM_L_X12Y152_SLICE_X16Y152_BQ),
.O5(CLBLM_L_X12Y153_SLICE_X17Y153_CO5),
.O6(CLBLM_L_X12Y153_SLICE_X17Y153_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5599559a55aa55aa)
  ) CLBLM_L_X12Y153_SLICE_X17Y153_BLUT (
.I0(CLBLM_L_X12Y153_SLICE_X17Y153_AQ),
.I1(CLBLM_R_X11Y153_SLICE_X14Y153_CO5),
.I2(CLBLM_R_X13Y152_SLICE_X18Y152_AO6),
.I3(CLBLM_L_X12Y153_SLICE_X16Y153_DO6),
.I4(CLBLM_R_X13Y152_SLICE_X18Y152_BO6),
.I5(CLBLM_L_X10Y154_SLICE_X13Y154_BQ),
.O5(CLBLM_L_X12Y153_SLICE_X17Y153_BO5),
.O6(CLBLM_L_X12Y153_SLICE_X17Y153_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdddd1111ddcc1100)
  ) CLBLM_L_X12Y153_SLICE_X17Y153_ALUT (
.I0(CLBLM_R_X11Y154_SLICE_X15Y154_CO5),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(1'b1),
.I3(CLBLM_L_X12Y153_SLICE_X17Y153_BO6),
.I4(CLBLM_R_X11Y154_SLICE_X15Y154_AQ),
.I5(CLBLM_L_X10Y154_SLICE_X13Y154_CO5),
.O5(CLBLM_L_X12Y153_SLICE_X17Y153_AO5),
.O6(CLBLM_L_X12Y153_SLICE_X17Y153_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y154_SLICE_X16Y154_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X12Y154_SLICE_X16Y154_AO6),
.Q(CLBLM_L_X12Y154_SLICE_X16Y154_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y154_SLICE_X16Y154_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y154_SLICE_X16Y154_DO5),
.O6(CLBLM_L_X12Y154_SLICE_X16Y154_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y154_SLICE_X16Y154_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y154_SLICE_X16Y154_CO5),
.O6(CLBLM_L_X12Y154_SLICE_X16Y154_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hd00fd0dfff00f000)
  ) CLBLM_L_X12Y154_SLICE_X16Y154_BLUT (
.I0(CLBLM_L_X10Y153_SLICE_X13Y153_BQ),
.I1(CLBLM_L_X10Y153_SLICE_X13Y153_CQ),
.I2(CLBLM_R_X11Y154_SLICE_X15Y154_AQ),
.I3(CLBLM_R_X11Y154_SLICE_X14Y154_AQ),
.I4(CLBLM_R_X11Y154_SLICE_X15Y154_BQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y154_SLICE_X16Y154_BO5),
.O6(CLBLM_L_X12Y154_SLICE_X16Y154_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00ccfacc00ccaf)
  ) CLBLM_L_X12Y154_SLICE_X16Y154_ALUT (
.I0(CLBLM_L_X10Y154_SLICE_X13Y154_CO5),
.I1(CLBLL_L_X4Y150_SLICE_X5Y150_AQ),
.I2(CLBLM_L_X12Y154_SLICE_X16Y154_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X11Y154_SLICE_X15Y154_CO5),
.I5(CLBLM_L_X12Y152_SLICE_X16Y152_CO6),
.O5(CLBLM_L_X12Y154_SLICE_X16Y154_AO5),
.O6(CLBLM_L_X12Y154_SLICE_X16Y154_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y154_SLICE_X17Y154_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y154_SLICE_X17Y154_DO5),
.O6(CLBLM_L_X12Y154_SLICE_X17Y154_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y154_SLICE_X17Y154_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y154_SLICE_X17Y154_CO5),
.O6(CLBLM_L_X12Y154_SLICE_X17Y154_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y154_SLICE_X17Y154_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y154_SLICE_X17Y154_BO5),
.O6(CLBLM_L_X12Y154_SLICE_X17Y154_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y154_SLICE_X17Y154_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y154_SLICE_X17Y154_AO5),
.O6(CLBLM_L_X12Y154_SLICE_X17Y154_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y155_SLICE_X16Y155_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y155_SLICE_X16Y155_DO5),
.O6(CLBLM_L_X12Y155_SLICE_X16Y155_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y155_SLICE_X16Y155_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y155_SLICE_X16Y155_CO5),
.O6(CLBLM_L_X12Y155_SLICE_X16Y155_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y155_SLICE_X16Y155_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y155_SLICE_X16Y155_BO5),
.O6(CLBLM_L_X12Y155_SLICE_X16Y155_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y155_SLICE_X16Y155_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y155_SLICE_X16Y155_AO5),
.O6(CLBLM_L_X12Y155_SLICE_X16Y155_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y155_SLICE_X17Y155_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X12Y155_SLICE_X17Y155_AO6),
.Q(CLBLM_L_X12Y155_SLICE_X17Y155_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y155_SLICE_X17Y155_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y155_SLICE_X17Y155_DO5),
.O6(CLBLM_L_X12Y155_SLICE_X17Y155_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y155_SLICE_X17Y155_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y155_SLICE_X17Y155_CO5),
.O6(CLBLM_L_X12Y155_SLICE_X17Y155_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y155_SLICE_X17Y155_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y155_SLICE_X17Y155_BO5),
.O6(CLBLM_L_X12Y155_SLICE_X17Y155_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccf0ccfaccf0ccfa)
  ) CLBLM_L_X12Y155_SLICE_X17Y155_ALUT (
.I0(RIOB33_X105Y141_IOB_X1Y142_I),
.I1(CLBLM_R_X7Y155_SLICE_X9Y155_AQ),
.I2(CLBLM_L_X12Y155_SLICE_X17Y155_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X5Y142_SLICE_X7Y142_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y155_SLICE_X17Y155_AO5),
.O6(CLBLM_L_X12Y155_SLICE_X17Y155_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y158_SLICE_X22Y158_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y158_SLICE_X22Y158_DO5),
.O6(CLBLM_L_X16Y158_SLICE_X22Y158_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y158_SLICE_X22Y158_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y158_SLICE_X22Y158_CO5),
.O6(CLBLM_L_X16Y158_SLICE_X22Y158_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y158_SLICE_X22Y158_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y158_SLICE_X22Y158_BO5),
.O6(CLBLM_L_X16Y158_SLICE_X22Y158_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffff0ff55ff55)
  ) CLBLM_L_X16Y158_SLICE_X22Y158_ALUT (
.I0(RIOB33_X105Y137_IOB_X1Y137_I),
.I1(1'b1),
.I2(RIOB33_X105Y127_IOB_X1Y128_I),
.I3(RIOB33_X105Y129_IOB_X1Y129_I),
.I4(RIOB33_X105Y129_IOB_X1Y130_I),
.I5(1'b1),
.O5(CLBLM_L_X16Y158_SLICE_X22Y158_AO5),
.O6(CLBLM_L_X16Y158_SLICE_X22Y158_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y158_SLICE_X23Y158_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y158_SLICE_X23Y158_DO5),
.O6(CLBLM_L_X16Y158_SLICE_X23Y158_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y158_SLICE_X23Y158_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y158_SLICE_X23Y158_CO5),
.O6(CLBLM_L_X16Y158_SLICE_X23Y158_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y158_SLICE_X23Y158_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y158_SLICE_X23Y158_BO5),
.O6(CLBLM_L_X16Y158_SLICE_X23Y158_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y158_SLICE_X23Y158_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y158_SLICE_X23Y158_AO5),
.O6(CLBLM_L_X16Y158_SLICE_X23Y158_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y141_SLICE_X2Y141_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y141_SLICE_X2Y141_DO5),
.O6(CLBLM_R_X3Y141_SLICE_X2Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y141_SLICE_X2Y141_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y141_SLICE_X2Y141_CO5),
.O6(CLBLM_R_X3Y141_SLICE_X2Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfaf0aa00fefceecc)
  ) CLBLM_R_X3Y141_SLICE_X2Y141_BLUT (
.I0(CLBLM_R_X3Y144_SLICE_X3Y144_BO5),
.I1(CLBLM_R_X3Y150_SLICE_X2Y150_BO6),
.I2(CLBLM_R_X3Y151_SLICE_X3Y151_AO6),
.I3(CLBLM_R_X3Y152_SLICE_X3Y152_CO6),
.I4(LIOB33_X0Y53_IOB_X0Y53_I),
.I5(CLBLL_L_X4Y142_SLICE_X5Y142_AO5),
.O5(CLBLM_R_X3Y141_SLICE_X2Y141_BO5),
.O6(CLBLM_R_X3Y141_SLICE_X2Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_R_X3Y141_SLICE_X2Y141_ALUT (
.I0(CLBLM_R_X3Y143_SLICE_X3Y143_A5Q),
.I1(CLBLM_R_X3Y142_SLICE_X2Y142_BQ),
.I2(CLBLM_R_X3Y142_SLICE_X2Y142_AQ),
.I3(CLBLM_R_X3Y143_SLICE_X3Y143_BQ),
.I4(CLBLL_L_X2Y145_SLICE_X1Y145_AQ),
.I5(CLBLM_R_X3Y143_SLICE_X2Y143_CQ),
.O5(CLBLM_R_X3Y141_SLICE_X2Y141_AO5),
.O6(CLBLM_R_X3Y141_SLICE_X2Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y141_SLICE_X3Y141_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y141_SLICE_X3Y141_DO5),
.O6(CLBLM_R_X3Y141_SLICE_X3Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y141_SLICE_X3Y141_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y141_SLICE_X3Y141_CO5),
.O6(CLBLM_R_X3Y141_SLICE_X3Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y141_SLICE_X3Y141_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y141_SLICE_X3Y141_BO5),
.O6(CLBLM_R_X3Y141_SLICE_X3Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y141_SLICE_X3Y141_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y141_SLICE_X3Y141_AO5),
.O6(CLBLM_R_X3Y141_SLICE_X3Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y142_SLICE_X2Y142_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y142_SLICE_X2Y142_AO6),
.Q(CLBLM_R_X3Y142_SLICE_X2Y142_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y142_SLICE_X2Y142_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y142_SLICE_X2Y142_BO6),
.Q(CLBLM_R_X3Y142_SLICE_X2Y142_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y142_SLICE_X2Y142_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y142_SLICE_X2Y142_CO6),
.Q(CLBLM_R_X3Y142_SLICE_X2Y142_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h80000000c0000000)
  ) CLBLM_R_X3Y142_SLICE_X2Y142_DLUT (
.I0(CLBLM_R_X3Y142_SLICE_X2Y142_AQ),
.I1(CLBLM_R_X3Y143_SLICE_X2Y143_CQ),
.I2(CLBLM_R_X3Y143_SLICE_X3Y143_A5Q),
.I3(CLBLM_R_X3Y142_SLICE_X2Y142_BQ),
.I4(CLBLL_L_X2Y145_SLICE_X1Y145_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y142_SLICE_X2Y142_DO5),
.O6(CLBLM_R_X3Y142_SLICE_X2Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00be14aa00)
  ) CLBLM_R_X3Y142_SLICE_X2Y142_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X3Y142_SLICE_X2Y142_CQ),
.I2(CLBLM_R_X3Y143_SLICE_X3Y143_DO5),
.I3(CLBLM_R_X3Y148_SLICE_X3Y148_BQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X3Y145_SLICE_X3Y145_D5Q),
.O5(CLBLM_R_X3Y142_SLICE_X2Y142_CO5),
.O6(CLBLM_R_X3Y142_SLICE_X2Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff006060ff00c0c0)
  ) CLBLM_R_X3Y142_SLICE_X2Y142_BLUT (
.I0(CLBLM_R_X3Y143_SLICE_X3Y143_A5Q),
.I1(CLBLM_R_X3Y142_SLICE_X2Y142_BQ),
.I2(CLBLM_R_X3Y143_SLICE_X3Y143_CO5),
.I3(CLBLL_L_X2Y145_SLICE_X1Y145_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X3Y143_SLICE_X2Y143_CQ),
.O5(CLBLM_R_X3Y142_SLICE_X2Y142_BO5),
.O6(CLBLM_R_X3Y142_SLICE_X2Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff022000000220)
  ) CLBLM_R_X3Y142_SLICE_X2Y142_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X3Y145_SLICE_X3Y145_D5Q),
.I2(CLBLM_R_X3Y142_SLICE_X2Y142_AQ),
.I3(CLBLM_R_X3Y142_SLICE_X2Y142_DO5),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X5Y149_SLICE_X6Y149_AQ),
.O5(CLBLM_R_X3Y142_SLICE_X2Y142_AO5),
.O6(CLBLM_R_X3Y142_SLICE_X2Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y142_SLICE_X3Y142_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y142_SLICE_X3Y142_DO5),
.O6(CLBLM_R_X3Y142_SLICE_X3Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y142_SLICE_X3Y142_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y142_SLICE_X3Y142_CO5),
.O6(CLBLM_R_X3Y142_SLICE_X3Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y142_SLICE_X3Y142_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y142_SLICE_X3Y142_BO5),
.O6(CLBLM_R_X3Y142_SLICE_X3Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y142_SLICE_X3Y142_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y142_SLICE_X3Y142_AO5),
.O6(CLBLM_R_X3Y142_SLICE_X3Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y143_SLICE_X2Y143_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y143_SLICE_X2Y143_AO6),
.Q(CLBLM_R_X3Y143_SLICE_X2Y143_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y143_SLICE_X2Y143_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y143_SLICE_X2Y143_BO6),
.Q(CLBLM_R_X3Y143_SLICE_X2Y143_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y143_SLICE_X2Y143_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y143_SLICE_X2Y143_CO6),
.Q(CLBLM_R_X3Y143_SLICE_X2Y143_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y143_SLICE_X2Y143_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y143_SLICE_X2Y143_DO6),
.Q(CLBLM_R_X3Y143_SLICE_X2Y143_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccf0fff000)
  ) CLBLM_R_X3Y143_SLICE_X2Y143_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y143_SLICE_X2Y143_CQ),
.I2(CLBLM_R_X3Y143_SLICE_X2Y143_DQ),
.I3(CLBLM_R_X3Y144_SLICE_X2Y144_CO6),
.I4(CLBLM_R_X3Y144_SLICE_X2Y144_A5Q),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X3Y143_SLICE_X2Y143_DO5),
.O6(CLBLM_R_X3Y143_SLICE_X2Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00ba10ea40)
  ) CLBLM_R_X3Y143_SLICE_X2Y143_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X3Y143_SLICE_X2Y143_CQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X5Y143_SLICE_X6Y143_AQ),
.I4(CLBLM_R_X3Y143_SLICE_X3Y143_A5Q),
.I5(CLBLM_R_X3Y145_SLICE_X3Y145_D5Q),
.O5(CLBLM_R_X3Y143_SLICE_X2Y143_CO5),
.O6(CLBLM_R_X3Y143_SLICE_X2Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa3fc0aaaaff00)
  ) CLBLM_R_X3Y143_SLICE_X2Y143_BLUT (
.I0(CLBLL_L_X4Y145_SLICE_X4Y145_CQ),
.I1(CLBLM_R_X3Y143_SLICE_X3Y143_DO5),
.I2(CLBLM_R_X3Y143_SLICE_X2Y143_AQ),
.I3(CLBLM_R_X3Y145_SLICE_X3Y145_D5Q),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X3Y142_SLICE_X2Y142_CQ),
.O5(CLBLM_R_X3Y143_SLICE_X2Y143_BO5),
.O6(CLBLM_R_X3Y143_SLICE_X2Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa30c0aaaaf000)
  ) CLBLM_R_X3Y143_SLICE_X2Y143_ALUT (
.I0(CLBLM_R_X3Y144_SLICE_X2Y144_A5Q),
.I1(CLBLM_R_X3Y143_SLICE_X3Y143_DO5),
.I2(CLBLM_R_X3Y143_SLICE_X3Y143_CO5),
.I3(CLBLM_R_X3Y143_SLICE_X2Y143_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X3Y142_SLICE_X2Y142_CQ),
.O5(CLBLM_R_X3Y143_SLICE_X2Y143_AO5),
.O6(CLBLM_R_X3Y143_SLICE_X2Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y143_SLICE_X3Y143_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y143_SLICE_X3Y143_CO6),
.Q(CLBLM_R_X3Y143_SLICE_X3Y143_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y143_SLICE_X3Y143_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y143_SLICE_X3Y143_DO6),
.Q(CLBLM_R_X3Y143_SLICE_X3Y143_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y143_SLICE_X3Y143_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y143_SLICE_X3Y143_AO6),
.Q(CLBLM_R_X3Y143_SLICE_X3Y143_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y143_SLICE_X3Y143_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y143_SLICE_X3Y143_BO6),
.Q(CLBLM_R_X3Y143_SLICE_X3Y143_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hbb88bb88a0a00000)
  ) CLBLM_R_X3Y143_SLICE_X3Y143_DLUT (
.I0(CLBLM_R_X3Y143_SLICE_X3Y143_BQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X3Y142_SLICE_X2Y142_DO6),
.I3(CLBLM_R_X3Y146_SLICE_X3Y146_CQ),
.I4(CLBLM_R_X3Y143_SLICE_X3Y143_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y143_SLICE_X3Y143_DO5),
.O6(CLBLM_R_X3Y143_SLICE_X3Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0b1a0a033330000)
  ) CLBLM_R_X3Y143_SLICE_X3Y143_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X3Y145_SLICE_X3Y145_D5Q),
.I2(CLBLM_R_X5Y155_SLICE_X7Y155_AQ),
.I3(CLBLM_R_X3Y143_SLICE_X3Y143_A5Q),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y143_SLICE_X3Y143_CO5),
.O6(CLBLM_R_X3Y143_SLICE_X3Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccdcccec00100020)
  ) CLBLM_R_X3Y143_SLICE_X3Y143_BLUT (
.I0(CLBLM_R_X3Y142_SLICE_X2Y142_DO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X3Y145_SLICE_X3Y145_D5Q),
.I4(CLBLM_R_X3Y143_SLICE_X3Y143_BQ),
.I5(CLBLM_L_X8Y145_SLICE_X10Y145_A5Q),
.O5(CLBLM_R_X3Y143_SLICE_X3Y143_BO5),
.O6(CLBLM_R_X3Y143_SLICE_X3Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa03aa30aa00aa00)
  ) CLBLM_R_X3Y143_SLICE_X3Y143_ALUT (
.I0(CLBLM_L_X8Y155_SLICE_X10Y155_AQ),
.I1(CLBLM_R_X3Y145_SLICE_X3Y145_D5Q),
.I2(CLBLM_R_X3Y143_SLICE_X3Y143_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X3Y141_SLICE_X2Y141_AO6),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X3Y143_SLICE_X3Y143_AO5),
.O6(CLBLM_R_X3Y143_SLICE_X3Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y144_SLICE_X2Y144_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y144_SLICE_X2Y144_AO5),
.Q(CLBLM_R_X3Y144_SLICE_X2Y144_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y144_SLICE_X2Y144_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y144_SLICE_X2Y144_BO5),
.Q(CLBLM_R_X3Y144_SLICE_X2Y144_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y144_SLICE_X2Y144_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y144_SLICE_X2Y144_AO6),
.Q(CLBLM_R_X3Y144_SLICE_X2Y144_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y144_SLICE_X2Y144_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y144_SLICE_X2Y144_BO6),
.Q(CLBLM_R_X3Y144_SLICE_X2Y144_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffff7fffffffff)
  ) CLBLM_R_X3Y144_SLICE_X2Y144_DLUT (
.I0(CLBLM_R_X3Y144_SLICE_X3Y144_AQ),
.I1(CLBLL_L_X4Y143_SLICE_X4Y143_CO6),
.I2(CLBLL_L_X2Y146_SLICE_X1Y146_CQ),
.I3(CLBLM_R_X7Y142_SLICE_X8Y142_DO6),
.I4(CLBLM_L_X8Y144_SLICE_X11Y144_BO6),
.I5(CLBLL_L_X2Y146_SLICE_X1Y146_AQ),
.O5(CLBLM_R_X3Y144_SLICE_X2Y144_DO5),
.O6(CLBLM_R_X3Y144_SLICE_X2Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000004000000cc)
  ) CLBLM_R_X3Y144_SLICE_X2Y144_CLUT (
.I0(CLBLM_R_X3Y148_SLICE_X3Y148_BQ),
.I1(CLBLL_L_X4Y143_SLICE_X4Y143_CO6),
.I2(CLBLM_R_X3Y144_SLICE_X3Y144_BO5),
.I3(CLBLM_R_X7Y142_SLICE_X8Y142_DO6),
.I4(CLBLM_L_X8Y144_SLICE_X11Y144_BO6),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X3Y144_SLICE_X2Y144_CO5),
.O6(CLBLM_R_X3Y144_SLICE_X2Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff33cc00f3f3c0c0)
  ) CLBLM_R_X3Y144_SLICE_X2Y144_BLUT (
.I0(1'b1),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X3Y146_SLICE_X3Y146_AQ),
.I3(CLBLM_R_X3Y146_SLICE_X2Y146_BQ),
.I4(RIOB33_X105Y127_IOB_X1Y127_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y144_SLICE_X2Y144_BO5),
.O6(CLBLM_R_X3Y144_SLICE_X2Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaccaaccfff000f0)
  ) CLBLM_R_X3Y144_SLICE_X2Y144_ALUT (
.I0(CLBLM_R_X3Y144_SLICE_X2Y144_B5Q),
.I1(CLBLM_R_X3Y145_SLICE_X2Y145_BQ),
.I2(CLBLL_L_X4Y144_SLICE_X4Y144_BQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X3Y147_SLICE_X3Y147_DQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y144_SLICE_X2Y144_AO5),
.O6(CLBLM_R_X3Y144_SLICE_X2Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y144_SLICE_X3Y144_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y144_SLICE_X3Y144_AO6),
.Q(CLBLM_R_X3Y144_SLICE_X3Y144_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y144_SLICE_X3Y144_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y144_SLICE_X3Y144_DO5),
.O6(CLBLM_R_X3Y144_SLICE_X3Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h07ff07ff77ff77ff)
  ) CLBLM_R_X3Y144_SLICE_X3Y144_CLUT (
.I0(CLBLM_R_X3Y146_SLICE_X2Y146_AQ),
.I1(CLBLM_R_X3Y146_SLICE_X2Y146_BQ),
.I2(CLBLL_L_X4Y144_SLICE_X4Y144_BQ),
.I3(CLBLM_R_X3Y146_SLICE_X3Y146_CQ),
.I4(1'b1),
.I5(CLBLL_L_X4Y144_SLICE_X4Y144_AQ),
.O5(CLBLM_R_X3Y144_SLICE_X3Y144_CO5),
.O6(CLBLM_R_X3Y144_SLICE_X3Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hdc00ff0050505050)
  ) CLBLM_R_X3Y144_SLICE_X3Y144_BLUT (
.I0(CLBLM_R_X5Y147_SLICE_X7Y147_D5Q),
.I1(CLBLM_R_X3Y148_SLICE_X3Y148_BQ),
.I2(CLBLL_L_X2Y147_SLICE_X1Y147_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_L_X8Y145_SLICE_X11Y145_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y144_SLICE_X3Y144_BO5),
.O6(CLBLM_R_X3Y144_SLICE_X3Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa3c00f000)
  ) CLBLM_R_X3Y144_SLICE_X3Y144_ALUT (
.I0(CLBLM_R_X11Y146_SLICE_X15Y146_AQ),
.I1(CLBLM_R_X7Y144_SLICE_X9Y144_DO6),
.I2(CLBLM_R_X3Y144_SLICE_X3Y144_AQ),
.I3(CLBLM_R_X3Y144_SLICE_X3Y144_BO6),
.I4(CLBLL_L_X2Y146_SLICE_X1Y146_CQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X3Y144_SLICE_X3Y144_AO5),
.O6(CLBLM_R_X3Y144_SLICE_X3Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y145_SLICE_X2Y145_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y145_SLICE_X2Y145_CO6),
.Q(CLBLM_R_X3Y145_SLICE_X2Y145_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y145_SLICE_X2Y145_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y145_SLICE_X2Y145_AO6),
.Q(CLBLM_R_X3Y145_SLICE_X2Y145_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y145_SLICE_X2Y145_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y145_SLICE_X2Y145_BO6),
.Q(CLBLM_R_X3Y145_SLICE_X2Y145_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_R_X3Y145_SLICE_X2Y145_DLUT (
.I0(CLBLL_L_X4Y144_SLICE_X4Y144_BQ),
.I1(CLBLM_R_X5Y144_SLICE_X6Y144_AQ),
.I2(CLBLM_R_X3Y145_SLICE_X2Y145_A5Q),
.I3(CLBLM_R_X3Y145_SLICE_X3Y145_CQ),
.I4(CLBLM_R_X3Y145_SLICE_X2Y145_BQ),
.I5(CLBLL_L_X4Y144_SLICE_X4Y144_AQ),
.O5(CLBLM_R_X3Y145_SLICE_X2Y145_DO5),
.O6(CLBLM_R_X3Y145_SLICE_X2Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hdffd1331f000f000)
  ) CLBLM_R_X3Y145_SLICE_X2Y145_CLUT (
.I0(CLBLM_R_X5Y144_SLICE_X6Y144_BO5),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X5Y144_SLICE_X6Y144_AQ),
.I3(CLBLM_R_X3Y145_SLICE_X2Y145_A5Q),
.I4(CLBLM_L_X12Y147_SLICE_X16Y147_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y145_SLICE_X2Y145_CO5),
.O6(CLBLM_R_X3Y145_SLICE_X2Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf202f808f808f808)
  ) CLBLM_R_X3Y145_SLICE_X2Y145_BLUT (
.I0(CLBLM_R_X5Y144_SLICE_X6Y144_BO5),
.I1(CLBLM_R_X3Y145_SLICE_X2Y145_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X5Y148_SLICE_X7Y148_CQ),
.I4(CLBLM_R_X3Y145_SLICE_X2Y145_CO5),
.I5(CLBLM_R_X3Y145_SLICE_X3Y145_CQ),
.O5(CLBLM_R_X3Y145_SLICE_X2Y145_BO5),
.O6(CLBLM_R_X3Y145_SLICE_X2Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heeaaeeaaeca0eca0)
  ) CLBLM_R_X3Y145_SLICE_X2Y145_ALUT (
.I0(CLBLM_R_X5Y152_SLICE_X7Y152_DO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X3Y145_SLICE_X2Y145_AQ),
.I3(CLBLL_L_X2Y145_SLICE_X1Y145_AQ),
.I4(1'b1),
.I5(CLBLM_R_X5Y152_SLICE_X6Y152_A5Q),
.O5(CLBLM_R_X3Y145_SLICE_X2Y145_AO5),
.O6(CLBLM_R_X3Y145_SLICE_X2Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y145_SLICE_X3Y145_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y145_SLICE_X3Y145_AO5),
.Q(CLBLM_R_X3Y145_SLICE_X3Y145_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y145_SLICE_X3Y145_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y145_SLICE_X3Y145_DO5),
.Q(CLBLM_R_X3Y145_SLICE_X3Y145_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y145_SLICE_X3Y145_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y145_SLICE_X3Y145_AO6),
.Q(CLBLM_R_X3Y145_SLICE_X3Y145_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y145_SLICE_X3Y145_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y145_SLICE_X3Y145_BO6),
.Q(CLBLM_R_X3Y145_SLICE_X3Y145_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y145_SLICE_X3Y145_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y145_SLICE_X3Y145_CO6),
.Q(CLBLM_R_X3Y145_SLICE_X3Y145_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y145_SLICE_X3Y145_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y145_SLICE_X3Y145_DO6),
.Q(CLBLM_R_X3Y145_SLICE_X3Y145_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hee44ee44fafa5050)
  ) CLBLM_R_X3Y145_SLICE_X3Y145_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLL_L_X4Y146_SLICE_X4Y146_A5Q),
.I2(CLBLM_R_X11Y146_SLICE_X14Y146_AQ),
.I3(CLBLM_R_X3Y145_SLICE_X3Y145_BQ),
.I4(CLBLL_L_X2Y147_SLICE_X1Y147_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y145_SLICE_X3Y145_DO5),
.O6(CLBLM_R_X3Y145_SLICE_X3Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hb3ecececa0a0a0a0)
  ) CLBLM_R_X3Y145_SLICE_X3Y145_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X3Y145_SLICE_X3Y145_CQ),
.I2(CLBLL_L_X4Y146_SLICE_X4Y146_AQ),
.I3(CLBLM_R_X5Y144_SLICE_X6Y144_AQ),
.I4(CLBLM_R_X3Y145_SLICE_X2Y145_A5Q),
.I5(CLBLM_R_X5Y144_SLICE_X6Y144_BO6),
.O5(CLBLM_R_X3Y145_SLICE_X3Y145_CO5),
.O6(CLBLM_R_X3Y145_SLICE_X3Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ffee000000ee)
  ) CLBLM_R_X3Y145_SLICE_X3Y145_BLUT (
.I0(CLBLM_R_X5Y147_SLICE_X7Y147_CQ),
.I1(CLBLM_R_X3Y145_SLICE_X3Y145_BQ),
.I2(1'b1),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X5Y152_SLICE_X7Y152_DO6),
.I5(CLBLM_R_X3Y142_SLICE_X2Y142_CQ),
.O5(CLBLM_R_X3Y145_SLICE_X3Y145_BO5),
.O6(CLBLM_R_X3Y145_SLICE_X3Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaccccff00aaaa)
  ) CLBLM_R_X3Y145_SLICE_X3Y145_ALUT (
.I0(CLBLM_R_X5Y144_SLICE_X6Y144_AQ),
.I1(CLBLL_L_X4Y154_SLICE_X4Y154_CO6),
.I2(1'b1),
.I3(CLBLM_R_X3Y145_SLICE_X3Y145_D5Q),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y145_SLICE_X3Y145_AO5),
.O6(CLBLM_R_X3Y145_SLICE_X3Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y146_SLICE_X2Y146_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y146_SLICE_X2Y146_AO6),
.Q(CLBLM_R_X3Y146_SLICE_X2Y146_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y146_SLICE_X2Y146_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y146_SLICE_X2Y146_BO6),
.Q(CLBLM_R_X3Y146_SLICE_X2Y146_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f00000000000)
  ) CLBLM_R_X3Y146_SLICE_X2Y146_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X11Y147_SLICE_X14Y147_BQ),
.I3(CLBLL_L_X4Y146_SLICE_X4Y146_DO6),
.I4(1'b1),
.I5(CLBLM_L_X10Y147_SLICE_X12Y147_AQ),
.O5(CLBLM_R_X3Y146_SLICE_X2Y146_DO5),
.O6(CLBLM_R_X3Y146_SLICE_X2Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hc000c000c000c000)
  ) CLBLM_R_X3Y146_SLICE_X2Y146_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y146_SLICE_X2Y146_AQ),
.I2(CLBLM_R_X3Y146_SLICE_X2Y146_BQ),
.I3(CLBLM_R_X3Y145_SLICE_X2Y145_DO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y146_SLICE_X2Y146_CO5),
.O6(CLBLM_R_X3Y146_SLICE_X2Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hbeaa3c00eeaacc00)
  ) CLBLM_R_X3Y146_SLICE_X2Y146_BLUT (
.I0(CLBLM_R_X5Y148_SLICE_X6Y148_AQ),
.I1(CLBLM_R_X3Y146_SLICE_X2Y146_BQ),
.I2(CLBLM_R_X3Y146_SLICE_X2Y146_AQ),
.I3(CLBLM_R_X5Y144_SLICE_X6Y144_BO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X3Y145_SLICE_X2Y145_DO6),
.O5(CLBLM_R_X3Y146_SLICE_X2Y146_BO5),
.O6(CLBLM_R_X3Y146_SLICE_X2Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8f888f88f888f888)
  ) CLBLM_R_X3Y146_SLICE_X2Y146_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X3Y149_SLICE_X2Y149_BQ),
.I2(CLBLM_R_X3Y146_SLICE_X2Y146_AQ),
.I3(CLBLM_R_X5Y144_SLICE_X6Y144_BO6),
.I4(1'b1),
.I5(CLBLM_R_X3Y145_SLICE_X2Y145_DO6),
.O5(CLBLM_R_X3Y146_SLICE_X2Y146_AO5),
.O6(CLBLM_R_X3Y146_SLICE_X2Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y146_SLICE_X3Y146_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y146_SLICE_X3Y146_AO6),
.Q(CLBLM_R_X3Y146_SLICE_X3Y146_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y146_SLICE_X3Y146_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y146_SLICE_X3Y146_BO6),
.Q(CLBLM_R_X3Y146_SLICE_X3Y146_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y146_SLICE_X3Y146_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y146_SLICE_X3Y146_CO6),
.Q(CLBLM_R_X3Y146_SLICE_X3Y146_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h80000000c0000000)
  ) CLBLM_R_X3Y146_SLICE_X3Y146_DLUT (
.I0(CLBLL_L_X4Y147_SLICE_X5Y147_BQ),
.I1(CLBLM_L_X10Y147_SLICE_X12Y147_AQ),
.I2(CLBLM_R_X3Y146_SLICE_X3Y146_BQ),
.I3(CLBLL_L_X4Y146_SLICE_X4Y146_DO6),
.I4(CLBLM_R_X11Y147_SLICE_X14Y147_BQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y146_SLICE_X3Y146_DO5),
.O6(CLBLM_R_X3Y146_SLICE_X3Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff22ff8822228888)
  ) CLBLM_R_X3Y146_SLICE_X3Y146_CLUT (
.I0(CLBLM_R_X5Y144_SLICE_X6Y144_BO6),
.I1(CLBLM_R_X3Y146_SLICE_X2Y146_CO6),
.I2(1'b1),
.I3(CLBLM_R_X3Y147_SLICE_X3Y147_BQ),
.I4(CLBLM_R_X3Y146_SLICE_X3Y146_CQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X3Y146_SLICE_X3Y146_CO5),
.O6(CLBLM_R_X3Y146_SLICE_X3Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h888b888b888b8888)
  ) CLBLM_R_X3Y146_SLICE_X3Y146_BLUT (
.I0(CLBLM_L_X8Y149_SLICE_X11Y149_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X11Y146_SLICE_X14Y146_AQ),
.I3(CLBLM_R_X3Y146_SLICE_X3Y146_DO5),
.I4(CLBLM_R_X3Y146_SLICE_X2Y146_DO6),
.I5(CLBLM_R_X3Y146_SLICE_X3Y146_BQ),
.O5(CLBLM_R_X3Y146_SLICE_X3Y146_BO5),
.O6(CLBLM_R_X3Y146_SLICE_X3Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff5f005fff4c004c)
  ) CLBLM_R_X3Y146_SLICE_X3Y146_ALUT (
.I0(CLBLM_L_X8Y149_SLICE_X11Y149_AQ),
.I1(CLBLM_R_X3Y146_SLICE_X3Y146_BQ),
.I2(CLBLL_L_X4Y151_SLICE_X4Y151_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLL_L_X4Y143_SLICE_X4Y143_AQ),
.I5(CLBLM_R_X3Y146_SLICE_X3Y146_AQ),
.O5(CLBLM_R_X3Y146_SLICE_X3Y146_AO5),
.O6(CLBLM_R_X3Y146_SLICE_X3Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y147_SLICE_X2Y147_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y147_SLICE_X2Y147_BO6),
.Q(CLBLM_R_X3Y147_SLICE_X2Y147_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y147_SLICE_X2Y147_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y147_SLICE_X2Y147_AO6),
.Q(CLBLM_R_X3Y147_SLICE_X2Y147_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y147_SLICE_X2Y147_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y147_SLICE_X2Y147_CO6),
.Q(CLBLM_R_X3Y147_SLICE_X2Y147_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y147_SLICE_X2Y147_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y147_SLICE_X2Y147_DO6),
.Q(CLBLM_R_X3Y147_SLICE_X2Y147_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbeafbea51405140)
  ) CLBLM_R_X3Y147_SLICE_X2Y147_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y152_SLICE_X11Y152_BO6),
.I2(CLBLM_R_X3Y147_SLICE_X2Y147_DQ),
.I3(CLBLM_R_X5Y146_SLICE_X6Y146_CQ),
.I4(1'b1),
.I5(CLBLM_R_X3Y148_SLICE_X2Y148_AQ),
.O5(CLBLM_R_X3Y147_SLICE_X2Y147_DO5),
.O6(CLBLM_R_X3Y147_SLICE_X2Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfd0dff0ff808f000)
  ) CLBLM_R_X3Y147_SLICE_X2Y147_CLUT (
.I0(CLBLL_L_X4Y151_SLICE_X4Y151_AQ),
.I1(CLBLM_R_X3Y147_SLICE_X2Y147_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLL_L_X4Y146_SLICE_X4Y146_A5Q),
.I4(CLBLM_L_X8Y149_SLICE_X11Y149_AQ),
.I5(CLBLM_R_X11Y147_SLICE_X14Y147_BQ),
.O5(CLBLM_R_X3Y147_SLICE_X2Y147_CO5),
.O6(CLBLM_R_X3Y147_SLICE_X2Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc00a05f5f5f5f)
  ) CLBLM_R_X3Y147_SLICE_X2Y147_BLUT (
.I0(CLBLM_L_X8Y149_SLICE_X11Y149_AQ),
.I1(CLBLM_R_X3Y147_SLICE_X3Y147_AQ),
.I2(CLBLL_L_X4Y151_SLICE_X4Y151_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y147_SLICE_X2Y147_BO5),
.O6(CLBLM_R_X3Y147_SLICE_X2Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccfff0ccccfff0)
  ) CLBLM_R_X3Y147_SLICE_X2Y147_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y79_IOB_X0Y79_I),
.I2(CLBLM_R_X3Y147_SLICE_X2Y147_AQ),
.I3(CLBLM_R_X5Y152_SLICE_X7Y152_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y147_SLICE_X2Y147_AO5),
.O6(CLBLM_R_X3Y147_SLICE_X2Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y147_SLICE_X3Y147_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y147_SLICE_X3Y147_CO5),
.Q(CLBLM_R_X3Y147_SLICE_X3Y147_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y147_SLICE_X3Y147_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y147_SLICE_X3Y147_AO6),
.Q(CLBLM_R_X3Y147_SLICE_X3Y147_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y147_SLICE_X3Y147_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y147_SLICE_X3Y147_BO6),
.Q(CLBLM_R_X3Y147_SLICE_X3Y147_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y147_SLICE_X3Y147_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y147_SLICE_X3Y147_CO6),
.Q(CLBLM_R_X3Y147_SLICE_X3Y147_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y147_SLICE_X3Y147_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y147_SLICE_X3Y147_DO6),
.Q(CLBLM_R_X3Y147_SLICE_X3Y147_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000fa32fa32)
  ) CLBLM_R_X3Y147_SLICE_X3Y147_DLUT (
.I0(CLBLL_L_X4Y147_SLICE_X5Y147_BQ),
.I1(CLBLM_L_X8Y148_SLICE_X10Y148_A5Q),
.I2(CLBLM_R_X3Y147_SLICE_X3Y147_DQ),
.I3(CLBLM_R_X11Y150_SLICE_X14Y150_BO6),
.I4(CLBLM_R_X5Y142_SLICE_X7Y142_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X3Y147_SLICE_X3Y147_DO5),
.O6(CLBLM_R_X3Y147_SLICE_X3Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccaaaaff00aaaa)
  ) CLBLM_R_X3Y147_SLICE_X3Y147_CLUT (
.I0(RIOB33_X105Y101_IOB_X1Y102_I),
.I1(CLBLL_L_X4Y147_SLICE_X4Y147_BQ),
.I2(1'b1),
.I3(CLBLM_R_X3Y147_SLICE_X2Y147_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y147_SLICE_X3Y147_CO5),
.O6(CLBLM_R_X3Y147_SLICE_X3Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a3a0a3a0aca0ac)
  ) CLBLM_R_X3Y147_SLICE_X3Y147_BLUT (
.I0(CLBLM_R_X3Y147_SLICE_X2Y147_DQ),
.I1(CLBLM_R_X3Y147_SLICE_X3Y147_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X11Y146_SLICE_X14Y146_AQ),
.I4(1'b1),
.I5(CLBLM_R_X3Y146_SLICE_X3Y146_DO6),
.O5(CLBLM_R_X3Y147_SLICE_X3Y147_BO5),
.O6(CLBLM_R_X3Y147_SLICE_X3Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heeeeeaeaccccc0c0)
  ) CLBLM_R_X3Y147_SLICE_X3Y147_ALUT (
.I0(CLBLL_L_X4Y144_SLICE_X5Y144_AQ),
.I1(CLBLM_R_X5Y152_SLICE_X7Y152_DO6),
.I2(CLBLM_R_X3Y147_SLICE_X3Y147_AQ),
.I3(1'b1),
.I4(CLBLM_R_X3Y150_SLICE_X3Y150_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X3Y147_SLICE_X3Y147_AO5),
.O6(CLBLM_R_X3Y147_SLICE_X3Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y148_SLICE_X2Y148_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y148_SLICE_X2Y148_AO6),
.Q(CLBLM_R_X3Y148_SLICE_X2Y148_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y148_SLICE_X2Y148_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y148_SLICE_X2Y148_BO6),
.Q(CLBLM_R_X3Y148_SLICE_X2Y148_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y148_SLICE_X2Y148_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y148_SLICE_X2Y148_CO6),
.Q(CLBLM_R_X3Y148_SLICE_X2Y148_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y148_SLICE_X2Y148_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y148_SLICE_X2Y148_DO6),
.Q(CLBLM_R_X3Y148_SLICE_X2Y148_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffcff00fcfc0000)
  ) CLBLM_R_X3Y148_SLICE_X2Y148_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y145_SLICE_X12Y145_CQ),
.I2(CLBLM_R_X3Y148_SLICE_X2Y148_DQ),
.I3(CLBLM_R_X3Y147_SLICE_X3Y147_CQ),
.I4(CLBLM_R_X5Y152_SLICE_X7Y152_DO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X3Y148_SLICE_X2Y148_DO5),
.O6(CLBLM_R_X3Y148_SLICE_X2Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf2f8f2f802080208)
  ) CLBLM_R_X3Y148_SLICE_X2Y148_CLUT (
.I0(CLBLL_L_X2Y147_SLICE_X1Y147_AO6),
.I1(CLBLM_R_X3Y148_SLICE_X2Y148_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X3Y148_SLICE_X2Y148_AO5),
.I4(1'b1),
.I5(CLBLM_R_X7Y144_SLICE_X9Y144_CQ),
.O5(CLBLM_R_X3Y148_SLICE_X2Y148_CO5),
.O6(CLBLM_R_X3Y148_SLICE_X2Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa30c0aaaac0c0)
  ) CLBLM_R_X3Y148_SLICE_X2Y148_BLUT (
.I0(CLBLM_L_X8Y150_SLICE_X11Y150_AQ),
.I1(CLBLM_R_X3Y148_SLICE_X2Y148_BQ),
.I2(CLBLL_L_X2Y147_SLICE_X1Y147_AO6),
.I3(CLBLM_R_X3Y148_SLICE_X2Y148_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X3Y148_SLICE_X2Y148_AO5),
.O5(CLBLM_R_X3Y148_SLICE_X2Y148_BO5),
.O6(CLBLM_R_X3Y148_SLICE_X2Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8888f88f00f000f0)
  ) CLBLM_R_X3Y148_SLICE_X2Y148_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLL_L_X4Y148_SLICE_X4Y148_C5Q),
.I2(CLBLM_R_X3Y148_SLICE_X2Y148_AQ),
.I3(CLBLM_R_X11Y150_SLICE_X14Y150_BO6),
.I4(CLBLL_L_X2Y148_SLICE_X1Y148_BO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y148_SLICE_X2Y148_AO5),
.O6(CLBLM_R_X3Y148_SLICE_X2Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y148_SLICE_X3Y148_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y148_SLICE_X3Y148_BO5),
.Q(CLBLM_R_X3Y148_SLICE_X3Y148_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y148_SLICE_X3Y148_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y148_SLICE_X3Y148_AO6),
.Q(CLBLM_R_X3Y148_SLICE_X3Y148_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y148_SLICE_X3Y148_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y148_SLICE_X3Y148_BO6),
.Q(CLBLM_R_X3Y148_SLICE_X3Y148_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y148_SLICE_X3Y148_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y148_SLICE_X3Y148_CO6),
.Q(CLBLM_R_X3Y148_SLICE_X3Y148_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3133020033330000)
  ) CLBLM_R_X3Y148_SLICE_X3Y148_DLUT (
.I0(CLBLM_R_X3Y148_SLICE_X2Y148_AQ),
.I1(CLBLL_L_X2Y148_SLICE_X1Y148_BO6),
.I2(CLBLM_R_X11Y150_SLICE_X14Y150_BO6),
.I3(CLBLM_R_X3Y148_SLICE_X2Y148_CQ),
.I4(CLBLM_R_X3Y148_SLICE_X3Y148_B5Q),
.I5(CLBLM_R_X3Y148_SLICE_X2Y148_BQ),
.O5(CLBLM_R_X3Y148_SLICE_X3Y148_DO5),
.O6(CLBLM_R_X3Y148_SLICE_X3Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00cacaff00caca)
  ) CLBLM_R_X3Y148_SLICE_X3Y148_CLUT (
.I0(CLBLL_L_X4Y148_SLICE_X4Y148_C5Q),
.I1(CLBLM_R_X3Y148_SLICE_X3Y148_CQ),
.I2(CLBLM_R_X3Y144_SLICE_X2Y144_CO6),
.I3(CLBLL_L_X4Y146_SLICE_X5Y146_A5Q),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y148_SLICE_X3Y148_CO5),
.O6(CLBLM_R_X3Y148_SLICE_X3Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfc3030ff88ff88)
  ) CLBLM_R_X3Y148_SLICE_X3Y148_BLUT (
.I0(CLBLL_L_X4Y149_SLICE_X4Y149_CQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLL_L_X4Y144_SLICE_X4Y144_DO6),
.I3(CLBLM_R_X3Y148_SLICE_X3Y148_DO6),
.I4(CLBLM_R_X7Y149_SLICE_X8Y149_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y148_SLICE_X3Y148_BO5),
.O6(CLBLM_R_X3Y148_SLICE_X3Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf808f000f000f000)
  ) CLBLM_R_X3Y148_SLICE_X3Y148_ALUT (
.I0(CLBLM_R_X3Y148_SLICE_X3Y148_B5Q),
.I1(CLBLM_R_X3Y148_SLICE_X2Y148_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X5Y148_SLICE_X7Y148_C5Q),
.I4(CLBLM_R_X3Y148_SLICE_X2Y148_AQ),
.I5(CLBLM_R_X3Y148_SLICE_X2Y148_BQ),
.O5(CLBLM_R_X3Y148_SLICE_X3Y148_AO5),
.O6(CLBLM_R_X3Y148_SLICE_X3Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y149_SLICE_X2Y149_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y149_SLICE_X2Y149_AO6),
.Q(CLBLM_R_X3Y149_SLICE_X2Y149_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y149_SLICE_X2Y149_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y149_SLICE_X2Y149_BO6),
.Q(CLBLM_R_X3Y149_SLICE_X2Y149_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y149_SLICE_X2Y149_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y149_SLICE_X2Y149_CO6),
.Q(CLBLM_R_X3Y149_SLICE_X2Y149_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ff00aaaaffaa)
  ) CLBLM_R_X3Y149_SLICE_X2Y149_DLUT (
.I0(CLBLM_R_X7Y145_SLICE_X9Y145_AQ),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X3Y147_SLICE_X2Y147_CQ),
.I4(CLBLL_L_X2Y152_SLICE_X1Y152_BO6),
.I5(CLBLL_L_X4Y152_SLICE_X5Y152_AO6),
.O5(CLBLM_R_X3Y149_SLICE_X2Y149_DO5),
.O6(CLBLM_R_X3Y149_SLICE_X2Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hafafacaca0a0acac)
  ) CLBLM_R_X3Y149_SLICE_X2Y149_CLUT (
.I0(CLBLM_R_X7Y150_SLICE_X9Y150_A5Q),
.I1(CLBLM_R_X5Y152_SLICE_X7Y152_B5Q),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(CLBLM_R_X3Y144_SLICE_X2Y144_CO6),
.I5(CLBLM_R_X3Y149_SLICE_X2Y149_CQ),
.O5(CLBLM_R_X3Y149_SLICE_X2Y149_CO5),
.O6(CLBLM_R_X3Y149_SLICE_X2Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hacacafa0acacafa0)
  ) CLBLM_R_X3Y149_SLICE_X2Y149_BLUT (
.I0(CLBLM_R_X5Y150_SLICE_X7Y150_AQ),
.I1(CLBLM_R_X3Y149_SLICE_X2Y149_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y150_SLICE_X9Y150_A5Q),
.I4(CLBLM_L_X8Y152_SLICE_X11Y152_BO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y149_SLICE_X2Y149_BO5),
.O6(CLBLM_R_X3Y149_SLICE_X2Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaf3c0ff00)
  ) CLBLM_R_X3Y149_SLICE_X2Y149_ALUT (
.I0(CLBLM_R_X3Y148_SLICE_X2Y148_DQ),
.I1(CLBLL_L_X4Y151_SLICE_X4Y151_AQ),
.I2(CLBLM_R_X3Y149_SLICE_X2Y149_AQ),
.I3(CLBLL_L_X4Y145_SLICE_X4Y145_CQ),
.I4(CLBLM_L_X8Y149_SLICE_X11Y149_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X3Y149_SLICE_X2Y149_AO5),
.O6(CLBLM_R_X3Y149_SLICE_X2Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y149_SLICE_X3Y149_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y149_SLICE_X3Y149_BO5),
.Q(CLBLM_R_X3Y149_SLICE_X3Y149_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y149_SLICE_X3Y149_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y149_SLICE_X3Y149_AO6),
.Q(CLBLM_R_X3Y149_SLICE_X3Y149_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y149_SLICE_X3Y149_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y149_SLICE_X3Y149_BO6),
.Q(CLBLM_R_X3Y149_SLICE_X3Y149_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y149_SLICE_X3Y149_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y149_SLICE_X3Y149_CO6),
.Q(CLBLM_R_X3Y149_SLICE_X3Y149_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y149_SLICE_X3Y149_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y149_SLICE_X3Y149_DO6),
.Q(CLBLM_R_X3Y149_SLICE_X3Y149_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaafcffaaaa3000)
  ) CLBLM_R_X3Y149_SLICE_X3Y149_DLUT (
.I0(CLBLM_R_X5Y153_SLICE_X6Y153_A5Q),
.I1(CLBLM_R_X11Y150_SLICE_X14Y150_BO6),
.I2(CLBLM_R_X3Y149_SLICE_X3Y149_DQ),
.I3(CLBLM_L_X8Y148_SLICE_X10Y148_A5Q),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y145_SLICE_X8Y145_AQ),
.O5(CLBLM_R_X3Y149_SLICE_X3Y149_DO5),
.O6(CLBLM_R_X3Y149_SLICE_X3Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfaeefafa50445050)
  ) CLBLM_R_X3Y149_SLICE_X3Y149_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X3Y149_SLICE_X3Y149_CQ),
.I2(CLBLL_L_X4Y145_SLICE_X4Y145_CQ),
.I3(CLBLM_R_X11Y150_SLICE_X14Y150_BO6),
.I4(CLBLM_L_X8Y148_SLICE_X10Y148_A5Q),
.I5(CLBLM_R_X11Y150_SLICE_X15Y150_AQ),
.O5(CLBLM_R_X3Y149_SLICE_X3Y149_CO5),
.O6(CLBLM_R_X3Y149_SLICE_X3Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaee0044d8d8d8d8)
  ) CLBLM_R_X3Y149_SLICE_X3Y149_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X3Y149_SLICE_X3Y149_BQ),
.I2(CLBLM_R_X3Y146_SLICE_X2Y146_BQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X3Y149_SLICE_X2Y149_CQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y149_SLICE_X3Y149_BO5),
.O6(CLBLM_R_X3Y149_SLICE_X3Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heeecaaa0eeecaaa0)
  ) CLBLM_R_X3Y149_SLICE_X3Y149_ALUT (
.I0(CLBLM_R_X5Y152_SLICE_X7Y152_DO6),
.I1(CLBLM_R_X11Y148_SLICE_X15Y148_B5Q),
.I2(CLBLM_R_X7Y149_SLICE_X8Y149_AQ),
.I3(CLBLM_R_X3Y149_SLICE_X3Y149_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y149_SLICE_X3Y149_AO5),
.O6(CLBLM_R_X3Y149_SLICE_X3Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000aaaaf0f0fafa)
  ) CLBLM_R_X3Y150_SLICE_X2Y150_DLUT (
.I0(CLBLM_R_X3Y149_SLICE_X2Y149_BQ),
.I1(1'b1),
.I2(CLBLM_R_X7Y150_SLICE_X8Y150_AQ),
.I3(1'b1),
.I4(CLBLL_L_X4Y152_SLICE_X5Y152_AO6),
.I5(CLBLL_L_X2Y152_SLICE_X1Y152_BO6),
.O5(CLBLM_R_X3Y150_SLICE_X2Y150_DO5),
.O6(CLBLM_R_X3Y150_SLICE_X2Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h1010331000000000)
  ) CLBLM_R_X3Y150_SLICE_X2Y150_CLUT (
.I0(CLBLM_R_X3Y156_SLICE_X2Y156_AO6),
.I1(CLBLL_L_X2Y155_SLICE_X1Y155_DO6),
.I2(CLBLM_R_X3Y147_SLICE_X2Y147_DQ),
.I3(CLBLM_L_X10Y146_SLICE_X12Y146_C5Q),
.I4(CLBLL_L_X2Y150_SLICE_X0Y150_AO6),
.I5(RIOB33_X105Y131_IOB_X1Y131_I),
.O5(CLBLM_R_X3Y150_SLICE_X2Y150_CO5),
.O6(CLBLM_R_X3Y150_SLICE_X2Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_R_X3Y150_SLICE_X2Y150_BLUT (
.I0(CLBLM_R_X3Y151_SLICE_X2Y151_DO6),
.I1(CLBLL_L_X4Y150_SLICE_X4Y150_DO6),
.I2(CLBLM_R_X3Y149_SLICE_X2Y149_DO6),
.I3(CLBLL_L_X2Y150_SLICE_X1Y150_AO6),
.I4(CLBLM_R_X3Y155_SLICE_X2Y155_DO6),
.I5(CLBLL_L_X4Y150_SLICE_X5Y150_DO6),
.O5(CLBLM_R_X3Y150_SLICE_X2Y150_BO5),
.O6(CLBLM_R_X3Y150_SLICE_X2Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000005004544)
  ) CLBLM_R_X3Y150_SLICE_X2Y150_ALUT (
.I0(CLBLL_L_X2Y155_SLICE_X1Y155_DO6),
.I1(CLBLM_L_X8Y153_SLICE_X11Y153_DQ),
.I2(CLBLM_R_X3Y156_SLICE_X2Y156_AO6),
.I3(CLBLM_L_X8Y150_SLICE_X11Y150_AQ),
.I4(CLBLL_L_X2Y150_SLICE_X0Y150_AO6),
.I5(RIOB33_X105Y131_IOB_X1Y131_I),
.O5(CLBLM_R_X3Y150_SLICE_X2Y150_AO5),
.O6(CLBLM_R_X3Y150_SLICE_X2Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y150_SLICE_X3Y150_A5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X3Y150_SLICE_X3Y150_AO5),
.Q(CLBLM_R_X3Y150_SLICE_X3Y150_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y150_SLICE_X3Y150_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.Q(CLBLM_R_X3Y150_SLICE_X3Y150_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y150_SLICE_X3Y150_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X3Y150_SLICE_X3Y150_BO6),
.Q(CLBLM_R_X3Y150_SLICE_X3Y150_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000003202)
  ) CLBLM_R_X3Y150_SLICE_X3Y150_DLUT (
.I0(CLBLL_L_X4Y145_SLICE_X4Y145_AQ),
.I1(CLBLL_L_X4Y155_SLICE_X4Y155_AO5),
.I2(RIOB33_X105Y135_IOB_X1Y136_I),
.I3(CLBLM_R_X3Y147_SLICE_X3Y147_DQ),
.I4(CLBLL_L_X2Y151_SLICE_X0Y151_CO5),
.I5(RIOB33_X105Y135_IOB_X1Y135_I),
.O5(CLBLM_R_X3Y150_SLICE_X3Y150_DO5),
.O6(CLBLM_R_X3Y150_SLICE_X3Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffceceffffffce)
  ) CLBLM_R_X3Y150_SLICE_X3Y150_CLUT (
.I0(RIOB33_X105Y109_IOB_X1Y110_I),
.I1(CLBLL_L_X2Y150_SLICE_X1Y150_DO6),
.I2(CLBLL_L_X2Y154_SLICE_X1Y154_BO6),
.I3(CLBLL_L_X4Y149_SLICE_X4Y149_AQ),
.I4(CLBLL_L_X2Y149_SLICE_X1Y149_DO6),
.I5(CLBLL_L_X4Y152_SLICE_X4Y152_AO6),
.O5(CLBLM_R_X3Y150_SLICE_X3Y150_CO5),
.O6(CLBLM_R_X3Y150_SLICE_X3Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hafaeafae05040504)
  ) CLBLM_R_X3Y150_SLICE_X3Y150_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X3Y150_SLICE_X3Y150_BQ),
.I2(CLBLM_R_X3Y144_SLICE_X2Y144_CO6),
.I3(CLBLM_R_X3Y143_SLICE_X3Y143_B5Q),
.I4(1'b1),
.I5(CLBLM_R_X5Y150_SLICE_X6Y150_A5Q),
.O5(CLBLM_R_X3Y150_SLICE_X3Y150_BO5),
.O6(CLBLM_R_X3Y150_SLICE_X3Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0acaccfc0cfc0)
  ) CLBLM_R_X3Y150_SLICE_X3Y150_ALUT (
.I0(CLBLL_L_X4Y151_SLICE_X4Y151_A5Q),
.I1(CLBLM_R_X5Y152_SLICE_X6Y152_A5Q),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X3Y147_SLICE_X2Y147_A5Q),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y150_SLICE_X3Y150_AO5),
.O6(CLBLM_R_X3Y150_SLICE_X3Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff3f0fffff3300)
  ) CLBLM_R_X3Y151_SLICE_X2Y151_DLUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y155_SLICE_X5Y155_AO5),
.I2(CLBLL_L_X2Y152_SLICE_X1Y152_BO5),
.I3(CLBLM_R_X7Y151_SLICE_X8Y151_AQ),
.I4(CLBLM_R_X5Y152_SLICE_X6Y152_DO6),
.I5(CLBLM_R_X3Y148_SLICE_X2Y148_BQ),
.O5(CLBLM_R_X3Y151_SLICE_X2Y151_DO5),
.O6(CLBLM_R_X3Y151_SLICE_X2Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffff0ace)
  ) CLBLM_R_X3Y151_SLICE_X2Y151_CLUT (
.I0(CLBLM_R_X3Y148_SLICE_X2Y148_CQ),
.I1(CLBLL_L_X4Y148_SLICE_X4Y148_AQ),
.I2(CLBLL_L_X2Y152_SLICE_X1Y152_BO5),
.I3(CLBLL_L_X4Y155_SLICE_X5Y155_AO5),
.I4(CLBLM_R_X3Y152_SLICE_X2Y152_CO6),
.I5(CLBLM_R_X3Y151_SLICE_X2Y151_BO6),
.O5(CLBLM_R_X3Y151_SLICE_X2Y151_CO5),
.O6(CLBLM_R_X3Y151_SLICE_X2Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00cc00dc50)
  ) CLBLM_R_X3Y151_SLICE_X2Y151_BLUT (
.I0(CLBLL_L_X2Y151_SLICE_X1Y151_AO5),
.I1(CLBLM_L_X8Y149_SLICE_X11Y149_B5Q),
.I2(CLBLM_R_X7Y151_SLICE_X8Y151_A5Q),
.I3(CLBLM_L_X16Y158_SLICE_X22Y158_AO5),
.I4(RIOB33_X105Y131_IOB_X1Y132_I),
.I5(CLBLL_L_X2Y152_SLICE_X1Y152_AO5),
.O5(CLBLM_R_X3Y151_SLICE_X2Y151_BO5),
.O6(CLBLM_R_X3Y151_SLICE_X2Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000004)
  ) CLBLM_R_X3Y151_SLICE_X2Y151_ALUT (
.I0(CLBLL_L_X2Y151_SLICE_X1Y151_BO6),
.I1(CLBLM_R_X3Y153_SLICE_X2Y153_AO6),
.I2(CLBLM_R_X3Y151_SLICE_X3Y151_AO6),
.I3(CLBLM_R_X3Y154_SLICE_X3Y154_AO6),
.I4(CLBLM_R_X3Y150_SLICE_X2Y150_BO6),
.I5(CLBLM_R_X3Y152_SLICE_X3Y152_CO6),
.O5(CLBLM_R_X3Y151_SLICE_X2Y151_AO5),
.O6(CLBLM_R_X3Y151_SLICE_X2Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff3bff3bff0aff0a)
  ) CLBLM_R_X3Y151_SLICE_X3Y151_DLUT (
.I0(CLBLM_R_X3Y147_SLICE_X3Y147_AQ),
.I1(CLBLL_L_X4Y155_SLICE_X5Y155_AO5),
.I2(CLBLM_R_X3Y152_SLICE_X2Y152_AO5),
.I3(CLBLM_R_X3Y151_SLICE_X3Y151_CO6),
.I4(1'b1),
.I5(CLBLM_R_X5Y147_SLICE_X6Y147_BQ),
.O5(CLBLM_R_X3Y151_SLICE_X3Y151_DO5),
.O6(CLBLM_R_X3Y151_SLICE_X3Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000003f0f3300)
  ) CLBLM_R_X3Y151_SLICE_X3Y151_CLUT (
.I0(1'b1),
.I1(CLBLL_L_X2Y151_SLICE_X0Y151_CO5),
.I2(CLBLL_L_X2Y154_SLICE_X1Y154_BO5),
.I3(CLBLM_R_X3Y149_SLICE_X3Y149_AQ),
.I4(CLBLM_R_X5Y150_SLICE_X6Y150_DQ),
.I5(CLBLL_L_X2Y155_SLICE_X1Y155_DO6),
.O5(CLBLM_R_X3Y151_SLICE_X3Y151_CO5),
.O6(CLBLM_R_X3Y151_SLICE_X3Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0fcfafef00ccaaee)
  ) CLBLM_R_X3Y151_SLICE_X3Y151_BLUT (
.I0(CLBLL_L_X4Y149_SLICE_X4Y149_CQ),
.I1(CLBLM_L_X8Y151_SLICE_X10Y151_DQ),
.I2(CLBLL_L_X2Y154_SLICE_X1Y154_BO6),
.I3(CLBLL_L_X4Y152_SLICE_X4Y152_AO6),
.I4(CLBLL_L_X4Y155_SLICE_X5Y155_AO6),
.I5(RIOB33_X105Y107_IOB_X1Y107_I),
.O5(CLBLM_R_X3Y151_SLICE_X3Y151_BO5),
.O6(CLBLM_R_X3Y151_SLICE_X3Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_R_X3Y151_SLICE_X3Y151_ALUT (
.I0(CLBLM_R_X3Y152_SLICE_X2Y152_DO6),
.I1(CLBLL_L_X4Y150_SLICE_X4Y150_CO6),
.I2(CLBLM_R_X3Y151_SLICE_X2Y151_CO6),
.I3(CLBLM_R_X3Y151_SLICE_X3Y151_BO6),
.I4(CLBLM_R_X3Y155_SLICE_X2Y155_DO6),
.I5(CLBLL_L_X4Y151_SLICE_X4Y151_BO6),
.O5(CLBLM_R_X3Y151_SLICE_X3Y151_AO5),
.O6(CLBLM_R_X3Y151_SLICE_X3Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h75ff757530ff3030)
  ) CLBLM_R_X3Y152_SLICE_X2Y152_DLUT (
.I0(CLBLM_R_X3Y152_SLICE_X2Y152_AO6),
.I1(CLBLL_L_X2Y151_SLICE_X0Y151_BO6),
.I2(LIOB33_X0Y61_IOB_X0Y61_I),
.I3(CLBLM_R_X3Y152_SLICE_X2Y152_AO5),
.I4(CLBLM_R_X5Y154_SLICE_X6Y154_AQ),
.I5(CLBLM_R_X5Y147_SLICE_X6Y147_AQ),
.O5(CLBLM_R_X3Y152_SLICE_X2Y152_DO5),
.O6(CLBLM_R_X3Y152_SLICE_X2Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000002000)
  ) CLBLM_R_X3Y152_SLICE_X2Y152_CLUT (
.I0(RIOB33_X105Y133_IOB_X1Y133_I),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(RIOB33_X105Y115_IOB_X1Y115_I),
.I3(RIOB33_X105Y131_IOB_X1Y132_I),
.I4(RIOB33_X105Y133_IOB_X1Y134_I),
.I5(CLBLL_L_X2Y152_SLICE_X1Y152_AO6),
.O5(CLBLM_R_X3Y152_SLICE_X2Y152_CO5),
.O6(CLBLM_R_X3Y152_SLICE_X2Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffafcc0ccc0c)
  ) CLBLM_R_X3Y152_SLICE_X2Y152_BLUT (
.I0(RIOB33_X105Y127_IOB_X1Y128_I),
.I1(CLBLL_L_X4Y151_SLICE_X5Y151_BQ),
.I2(RIOB33_X105Y137_IOB_X1Y137_I),
.I3(RIOB33_X105Y129_IOB_X1Y129_I),
.I4(CLBLM_R_X5Y145_SLICE_X6Y145_DO5),
.I5(1'b1),
.O5(CLBLM_R_X3Y152_SLICE_X2Y152_BO5),
.O6(CLBLM_R_X3Y152_SLICE_X2Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffdfffffdff)
  ) CLBLM_R_X3Y152_SLICE_X2Y152_ALUT (
.I0(RIOB33_X105Y133_IOB_X1Y134_I),
.I1(CLBLL_L_X2Y155_SLICE_X1Y155_DO6),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(RIOB33_X105Y133_IOB_X1Y133_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y152_SLICE_X2Y152_AO5),
.O6(CLBLM_R_X3Y152_SLICE_X2Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000050445044)
  ) CLBLM_R_X3Y152_SLICE_X3Y152_DLUT (
.I0(CLBLL_L_X4Y154_SLICE_X5Y154_CO5),
.I1(CLBLM_R_X3Y149_SLICE_X3Y149_DQ),
.I2(CLBLM_R_X3Y148_SLICE_X2Y148_AQ),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(1'b1),
.I5(CLBLL_L_X2Y152_SLICE_X1Y152_AO6),
.O5(CLBLM_R_X3Y152_SLICE_X3Y152_DO5),
.O6(CLBLM_R_X3Y152_SLICE_X3Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffefffefffffffe)
  ) CLBLM_R_X3Y152_SLICE_X3Y152_CLUT (
.I0(CLBLL_L_X4Y153_SLICE_X5Y153_CO6),
.I1(CLBLM_R_X3Y151_SLICE_X3Y151_DO6),
.I2(CLBLL_L_X4Y152_SLICE_X4Y152_DO6),
.I3(CLBLM_R_X3Y150_SLICE_X3Y150_CO6),
.I4(CLBLM_R_X3Y155_SLICE_X3Y155_AO5),
.I5(CLBLL_L_X2Y155_SLICE_X1Y155_BO6),
.O5(CLBLM_R_X3Y152_SLICE_X3Y152_CO5),
.O6(CLBLM_R_X3Y152_SLICE_X3Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffafffffffe)
  ) CLBLM_R_X3Y152_SLICE_X3Y152_BLUT (
.I0(CLBLM_R_X3Y152_SLICE_X3Y152_DO6),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(CLBLL_L_X4Y152_SLICE_X4Y152_CO6),
.I3(CLBLL_L_X4Y152_SLICE_X5Y152_CO6),
.I4(CLBLM_R_X3Y152_SLICE_X3Y152_AO6),
.I5(CLBLL_L_X2Y154_SLICE_X1Y154_BO6),
.O5(CLBLM_R_X3Y152_SLICE_X3Y152_BO5),
.O6(CLBLM_R_X3Y152_SLICE_X3Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0055307500003030)
  ) CLBLM_R_X3Y152_SLICE_X3Y152_ALUT (
.I0(CLBLL_L_X4Y155_SLICE_X4Y155_BO6),
.I1(CLBLL_L_X2Y152_SLICE_X1Y152_AO6),
.I2(RIOB33_X105Y113_IOB_X1Y114_I),
.I3(CLBLL_L_X2Y155_SLICE_X1Y155_DO6),
.I4(CLBLL_L_X2Y151_SLICE_X1Y151_AO6),
.I5(CLBLM_R_X7Y152_SLICE_X8Y152_DQ),
.O5(CLBLM_R_X3Y152_SLICE_X3Y152_AO5),
.O6(CLBLM_R_X3Y152_SLICE_X3Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffff1fff1)
  ) CLBLM_R_X3Y153_SLICE_X2Y153_DLUT (
.I0(CLBLL_L_X2Y155_SLICE_X1Y155_AO6),
.I1(CLBLM_R_X3Y156_SLICE_X2Y156_CO6),
.I2(CLBLM_R_X3Y154_SLICE_X3Y154_DO6),
.I3(CLBLL_L_X4Y153_SLICE_X5Y153_DO6),
.I4(1'b1),
.I5(CLBLM_R_X3Y153_SLICE_X2Y153_BO6),
.O5(CLBLM_R_X3Y153_SLICE_X2Y153_DO5),
.O6(CLBLM_R_X3Y153_SLICE_X2Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0010000000000000)
  ) CLBLM_R_X3Y153_SLICE_X2Y153_CLUT (
.I0(RIOB33_X105Y133_IOB_X1Y134_I),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(RIOB33_X105Y133_IOB_X1Y133_I),
.I3(CLBLL_L_X2Y155_SLICE_X1Y155_DO6),
.I4(RIOB33_X105Y131_IOB_X1Y132_I),
.I5(CLBLM_R_X3Y148_SLICE_X2Y148_DQ),
.O5(CLBLM_R_X3Y153_SLICE_X2Y153_CO5),
.O6(CLBLM_R_X3Y153_SLICE_X2Y153_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffff7f3f5f0)
  ) CLBLM_R_X3Y153_SLICE_X2Y153_BLUT (
.I0(CLBLL_L_X2Y151_SLICE_X0Y151_AO6),
.I1(CLBLM_R_X3Y152_SLICE_X2Y152_AO5),
.I2(CLBLM_R_X3Y153_SLICE_X3Y153_CO6),
.I3(CLBLM_R_X5Y152_SLICE_X7Y152_CQ),
.I4(CLBLM_R_X3Y145_SLICE_X2Y145_AQ),
.I5(CLBLM_R_X3Y153_SLICE_X2Y153_CO6),
.O5(CLBLM_R_X3Y153_SLICE_X2Y153_BO5),
.O6(CLBLM_R_X3Y153_SLICE_X2Y153_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0003000100030000)
  ) CLBLM_R_X3Y153_SLICE_X2Y153_ALUT (
.I0(CLBLL_L_X2Y152_SLICE_X1Y152_BO5),
.I1(CLBLL_L_X4Y151_SLICE_X5Y151_CO6),
.I2(CLBLM_R_X3Y153_SLICE_X3Y153_AO6),
.I3(CLBLL_L_X2Y153_SLICE_X1Y153_AO6),
.I4(CLBLL_L_X2Y155_SLICE_X1Y155_AO6),
.I5(CLBLM_R_X3Y156_SLICE_X2Y156_CO6),
.O5(CLBLM_R_X3Y153_SLICE_X2Y153_AO5),
.O6(CLBLM_R_X3Y153_SLICE_X2Y153_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0044004400ff0044)
  ) CLBLM_R_X3Y153_SLICE_X3Y153_DLUT (
.I0(CLBLL_L_X2Y151_SLICE_X1Y151_AO6),
.I1(CLBLM_R_X3Y148_SLICE_X2Y148_DQ),
.I2(1'b1),
.I3(CLBLL_L_X2Y155_SLICE_X1Y155_DO6),
.I4(CLBLM_R_X3Y145_SLICE_X2Y145_AQ),
.I5(CLBLL_L_X4Y155_SLICE_X4Y155_BO6),
.O5(CLBLM_R_X3Y153_SLICE_X3Y153_DO5),
.O6(CLBLM_R_X3Y153_SLICE_X3Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccee0c0c0cae)
  ) CLBLM_R_X3Y153_SLICE_X3Y153_CLUT (
.I0(LIOB33_X0Y65_IOB_X0Y66_I),
.I1(CLBLL_L_X4Y151_SLICE_X5Y151_BQ),
.I2(RIOB33_X105Y137_IOB_X1Y137_I),
.I3(CLBLL_L_X2Y152_SLICE_X1Y152_AO5),
.I4(CLBLL_L_X2Y154_SLICE_X1Y154_BO5),
.I5(RIOB33_X105Y129_IOB_X1Y129_I),
.O5(CLBLM_R_X3Y153_SLICE_X3Y153_CO5),
.O6(CLBLM_R_X3Y153_SLICE_X3Y153_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff005d000c)
  ) CLBLM_R_X3Y153_SLICE_X3Y153_BLUT (
.I0(CLBLL_L_X2Y154_SLICE_X1Y154_BO5),
.I1(CLBLM_R_X5Y152_SLICE_X7Y152_CQ),
.I2(CLBLL_L_X2Y151_SLICE_X0Y151_CO5),
.I3(CLBLL_L_X2Y152_SLICE_X1Y152_AO5),
.I4(LIOB33_X0Y65_IOB_X0Y66_I),
.I5(CLBLM_R_X3Y152_SLICE_X2Y152_BO5),
.O5(CLBLM_R_X3Y153_SLICE_X3Y153_BO5),
.O6(CLBLM_R_X3Y153_SLICE_X3Y153_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_R_X3Y153_SLICE_X3Y153_ALUT (
.I0(CLBLM_R_X3Y153_SLICE_X3Y153_DO6),
.I1(CLBLM_R_X3Y155_SLICE_X3Y155_BO6),
.I2(CLBLL_L_X4Y154_SLICE_X5Y154_DO6),
.I3(CLBLM_R_X3Y153_SLICE_X3Y153_BO6),
.I4(CLBLL_L_X4Y153_SLICE_X4Y153_BO6),
.I5(CLBLM_R_X3Y150_SLICE_X3Y150_DO6),
.O5(CLBLM_R_X3Y153_SLICE_X3Y153_AO5),
.O6(CLBLM_R_X3Y153_SLICE_X3Y153_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaeeaaeefafefafe)
  ) CLBLM_R_X3Y154_SLICE_X2Y154_DLUT (
.I0(CLBLL_L_X4Y151_SLICE_X4Y151_DO6),
.I1(RIOB33_X105Y113_IOB_X1Y113_I),
.I2(CLBLM_R_X3Y149_SLICE_X3Y149_CQ),
.I3(CLBLL_L_X2Y154_SLICE_X1Y154_BO6),
.I4(1'b1),
.I5(CLBLL_L_X2Y152_SLICE_X1Y152_BO5),
.O5(CLBLM_R_X3Y154_SLICE_X2Y154_DO5),
.O6(CLBLM_R_X3Y154_SLICE_X2Y154_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff3030ffffbaba)
  ) CLBLM_R_X3Y154_SLICE_X2Y154_CLUT (
.I0(LIOB33_X0Y67_IOB_X0Y68_I),
.I1(CLBLL_L_X2Y154_SLICE_X1Y154_AO5),
.I2(CLBLM_R_X3Y149_SLICE_X2Y149_AQ),
.I3(1'b1),
.I4(CLBLL_L_X4Y155_SLICE_X4Y155_DO6),
.I5(CLBLL_L_X2Y151_SLICE_X0Y151_BO6),
.O5(CLBLM_R_X3Y154_SLICE_X2Y154_CO5),
.O6(CLBLM_R_X3Y154_SLICE_X2Y154_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffafefaaee)
  ) CLBLM_R_X3Y154_SLICE_X2Y154_BLUT (
.I0(CLBLM_R_X3Y154_SLICE_X2Y154_DO6),
.I1(CLBLM_R_X3Y155_SLICE_X2Y155_BO6),
.I2(CLBLL_L_X4Y152_SLICE_X5Y152_AO6),
.I3(CLBLM_R_X3Y156_SLICE_X2Y156_BO6),
.I4(CLBLM_R_X7Y153_SLICE_X9Y153_BQ),
.I5(CLBLM_R_X3Y154_SLICE_X2Y154_CO6),
.O5(CLBLM_R_X3Y154_SLICE_X2Y154_BO5),
.O6(CLBLM_R_X3Y154_SLICE_X2Y154_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000004000000)
  ) CLBLM_R_X3Y154_SLICE_X2Y154_ALUT (
.I0(RIOB33_X105Y133_IOB_X1Y134_I),
.I1(RIOB33_X105Y133_IOB_X1Y133_I),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(CLBLM_R_X7Y153_SLICE_X9Y153_BQ),
.I5(CLBLL_L_X2Y155_SLICE_X1Y155_DO6),
.O5(CLBLM_R_X3Y154_SLICE_X2Y154_AO5),
.O6(CLBLM_R_X3Y154_SLICE_X2Y154_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbbbffbbaaaaffaa)
  ) CLBLM_R_X3Y154_SLICE_X3Y154_DLUT (
.I0(CLBLM_R_X3Y150_SLICE_X3Y150_DO6),
.I1(CLBLL_L_X2Y154_SLICE_X1Y154_BO6),
.I2(1'b1),
.I3(CLBLL_L_X4Y150_SLICE_X5Y150_BQ),
.I4(CLBLL_L_X4Y155_SLICE_X5Y155_AO6),
.I5(RIOB33_X105Y111_IOB_X1Y111_I),
.O5(CLBLM_R_X3Y154_SLICE_X3Y154_DO5),
.O6(CLBLM_R_X3Y154_SLICE_X3Y154_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000077553300)
  ) CLBLM_R_X3Y154_SLICE_X3Y154_CLUT (
.I0(CLBLL_L_X2Y154_SLICE_X1Y154_BO5),
.I1(CLBLL_L_X4Y155_SLICE_X4Y155_BO6),
.I2(1'b1),
.I3(CLBLM_R_X3Y149_SLICE_X3Y149_CQ),
.I4(RIOB33_X105Y113_IOB_X1Y113_I),
.I5(CLBLL_L_X2Y152_SLICE_X1Y152_AO6),
.O5(CLBLM_R_X3Y154_SLICE_X3Y154_CO5),
.O6(CLBLM_R_X3Y154_SLICE_X3Y154_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffbfa)
  ) CLBLM_R_X3Y154_SLICE_X3Y154_BLUT (
.I0(CLBLL_L_X4Y155_SLICE_X4Y155_CO6),
.I1(CLBLL_L_X2Y154_SLICE_X1Y154_AO5),
.I2(CLBLM_R_X3Y154_SLICE_X2Y154_AO6),
.I3(CLBLM_R_X3Y149_SLICE_X2Y149_AQ),
.I4(CLBLM_R_X3Y154_SLICE_X3Y154_CO6),
.I5(CLBLL_L_X4Y151_SLICE_X4Y151_DO6),
.O5(CLBLM_R_X3Y154_SLICE_X3Y154_BO5),
.O6(CLBLM_R_X3Y154_SLICE_X3Y154_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_R_X3Y154_SLICE_X3Y154_ALUT (
.I0(CLBLL_L_X2Y150_SLICE_X1Y150_CO6),
.I1(CLBLM_R_X5Y154_SLICE_X7Y154_DO6),
.I2(CLBLM_R_X3Y155_SLICE_X2Y155_DO6),
.I3(CLBLM_R_X3Y154_SLICE_X3Y154_BO6),
.I4(CLBLL_L_X4Y154_SLICE_X4Y154_BO6),
.I5(CLBLM_R_X3Y155_SLICE_X2Y155_AO6),
.O5(CLBLM_R_X3Y154_SLICE_X3Y154_AO5),
.O6(CLBLM_R_X3Y154_SLICE_X3Y154_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000002000000000)
  ) CLBLM_R_X3Y155_SLICE_X2Y155_DLUT (
.I0(CLBLL_L_X2Y152_SLICE_X1Y152_BO5),
.I1(CLBLM_R_X3Y155_SLICE_X3Y155_CO6),
.I2(CLBLL_L_X2Y154_SLICE_X1Y154_AO6),
.I3(CLBLM_R_X3Y155_SLICE_X2Y155_CO6),
.I4(CLBLL_L_X2Y154_SLICE_X1Y154_CO6),
.I5(CLBLL_L_X4Y154_SLICE_X5Y154_CO6),
.O5(CLBLM_R_X3Y155_SLICE_X2Y155_DO5),
.O6(CLBLM_R_X3Y155_SLICE_X2Y155_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000001ab0101)
  ) CLBLM_R_X3Y155_SLICE_X2Y155_CLUT (
.I0(RIOB33_X105Y135_IOB_X1Y136_I),
.I1(CLBLL_L_X2Y150_SLICE_X0Y150_AO6),
.I2(RIOB33_X105Y135_IOB_X1Y135_I),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(CLBLM_R_X3Y156_SLICE_X2Y156_AO5),
.I5(CLBLL_L_X4Y155_SLICE_X4Y155_AO5),
.O5(CLBLM_R_X3Y155_SLICE_X2Y155_CO5),
.O6(CLBLM_R_X3Y155_SLICE_X2Y155_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h1000000000000000)
  ) CLBLM_R_X3Y155_SLICE_X2Y155_BLUT (
.I0(CLBLL_L_X2Y154_SLICE_X1Y154_CO6),
.I1(RIOB33_X105Y129_IOB_X1Y129_I),
.I2(CLBLM_R_X3Y155_SLICE_X3Y155_AO6),
.I3(RIOB33_X105Y137_IOB_X1Y137_I),
.I4(CLBLL_L_X2Y154_SLICE_X1Y154_CO5),
.I5(CLBLL_L_X4Y154_SLICE_X5Y154_CO6),
.O5(CLBLM_R_X3Y155_SLICE_X2Y155_BO5),
.O6(CLBLM_R_X3Y155_SLICE_X2Y155_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000001000000)
  ) CLBLM_R_X3Y155_SLICE_X2Y155_ALUT (
.I0(CLBLM_R_X3Y156_SLICE_X2Y156_CO6),
.I1(CLBLL_L_X4Y155_SLICE_X4Y155_BO5),
.I2(CLBLM_R_X3Y155_SLICE_X3Y155_CO6),
.I3(CLBLL_L_X4Y154_SLICE_X5Y154_CO6),
.I4(CLBLL_L_X2Y152_SLICE_X1Y152_BO5),
.I5(CLBLL_L_X2Y154_SLICE_X1Y154_CO6),
.O5(CLBLM_R_X3Y155_SLICE_X2Y155_AO5),
.O6(CLBLM_R_X3Y155_SLICE_X2Y155_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00ffffffff)
  ) CLBLM_R_X3Y155_SLICE_X3Y155_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(RIOB33_X105Y133_IOB_X1Y134_I),
.I4(1'b1),
.I5(RIOB33_X105Y133_IOB_X1Y133_I),
.O5(CLBLM_R_X3Y155_SLICE_X3Y155_DO5),
.O6(CLBLM_R_X3Y155_SLICE_X3Y155_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff05ff00ff27)
  ) CLBLM_R_X3Y155_SLICE_X3Y155_CLUT (
.I0(RIOB33_X105Y131_IOB_X1Y132_I),
.I1(CLBLL_L_X2Y152_SLICE_X1Y152_AO5),
.I2(CLBLL_L_X2Y155_SLICE_X1Y155_DO6),
.I3(CLBLM_L_X16Y158_SLICE_X22Y158_AO5),
.I4(CLBLM_R_X3Y155_SLICE_X3Y155_DO6),
.I5(RIOB33_X105Y131_IOB_X1Y131_I),
.O5(CLBLM_R_X3Y155_SLICE_X3Y155_CO5),
.O6(CLBLM_R_X3Y155_SLICE_X3Y155_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000000c000a)
  ) CLBLM_R_X3Y155_SLICE_X3Y155_BLUT (
.I0(CLBLL_L_X4Y150_SLICE_X5Y150_BQ),
.I1(RIOB33_X105Y111_IOB_X1Y111_I),
.I2(CLBLL_L_X2Y154_SLICE_X1Y154_BO5),
.I3(CLBLL_L_X4Y155_SLICE_X4Y155_AO5),
.I4(RIOB33_X105Y135_IOB_X1Y136_I),
.I5(RIOB33_X105Y135_IOB_X1Y135_I),
.O5(CLBLM_R_X3Y155_SLICE_X3Y155_BO5),
.O6(CLBLM_R_X3Y155_SLICE_X3Y155_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffbfffbffefffef)
  ) CLBLM_R_X3Y155_SLICE_X3Y155_ALUT (
.I0(RIOB33_X105Y133_IOB_X1Y134_I),
.I1(RIOB33_X105Y133_IOB_X1Y133_I),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(CLBLL_L_X2Y155_SLICE_X1Y155_DO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y155_SLICE_X3Y155_AO5),
.O6(CLBLM_R_X3Y155_SLICE_X3Y155_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y156_SLICE_X2Y156_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y156_SLICE_X2Y156_DO5),
.O6(CLBLM_R_X3Y156_SLICE_X2Y156_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000002000)
  ) CLBLM_R_X3Y156_SLICE_X2Y156_CLUT (
.I0(RIOB33_X105Y135_IOB_X1Y136_I),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(RIOB33_X105Y135_IOB_X1Y135_I),
.I3(CLBLM_R_X3Y156_SLICE_X2Y156_AO5),
.I4(CLBLM_L_X16Y158_SLICE_X22Y158_AO5),
.I5(RIOB33_X105Y129_IOB_X1Y130_I),
.O5(CLBLM_R_X3Y156_SLICE_X2Y156_CO5),
.O6(CLBLM_R_X3Y156_SLICE_X2Y156_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf4f4f1f0f0f0f0f0)
  ) CLBLM_R_X3Y156_SLICE_X2Y156_BLUT (
.I0(CLBLL_L_X2Y152_SLICE_X1Y152_AO6),
.I1(RIOB33_X105Y133_IOB_X1Y133_I),
.I2(CLBLM_R_X3Y156_SLICE_X2Y156_CO6),
.I3(RIOB33_X105Y133_IOB_X1Y134_I),
.I4(RIOB33_X105Y131_IOB_X1Y132_I),
.I5(RIOB33_X105Y131_IOB_X1Y131_I),
.O5(CLBLM_R_X3Y156_SLICE_X2Y156_BO5),
.O6(CLBLM_R_X3Y156_SLICE_X2Y156_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff3fff300c000c0)
  ) CLBLM_R_X3Y156_SLICE_X2Y156_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y133_IOB_X1Y133_I),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(RIOB33_X105Y133_IOB_X1Y134_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y156_SLICE_X2Y156_AO5),
.O6(CLBLM_R_X3Y156_SLICE_X2Y156_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y156_SLICE_X3Y156_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y156_SLICE_X3Y156_DO5),
.O6(CLBLM_R_X3Y156_SLICE_X3Y156_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y156_SLICE_X3Y156_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y156_SLICE_X3Y156_CO5),
.O6(CLBLM_R_X3Y156_SLICE_X3Y156_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y156_SLICE_X3Y156_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y156_SLICE_X3Y156_BO5),
.O6(CLBLM_R_X3Y156_SLICE_X3Y156_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y156_SLICE_X3Y156_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y156_SLICE_X3Y156_AO5),
.O6(CLBLM_R_X3Y156_SLICE_X3Y156_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y142_SLICE_X6Y142_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y142_SLICE_X6Y142_DO5),
.O6(CLBLM_R_X5Y142_SLICE_X6Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y142_SLICE_X6Y142_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y142_SLICE_X6Y142_CO5),
.O6(CLBLM_R_X5Y142_SLICE_X6Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y142_SLICE_X6Y142_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y142_SLICE_X6Y142_BO5),
.O6(CLBLM_R_X5Y142_SLICE_X6Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y142_SLICE_X6Y142_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y142_SLICE_X6Y142_AO5),
.O6(CLBLM_R_X5Y142_SLICE_X6Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y142_SLICE_X7Y142_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y142_SLICE_X8Y142_AO6),
.Q(CLBLM_R_X5Y142_SLICE_X7Y142_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y142_SLICE_X7Y142_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y142_SLICE_X7Y142_DO5),
.O6(CLBLM_R_X5Y142_SLICE_X7Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y142_SLICE_X7Y142_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y142_SLICE_X7Y142_CO5),
.O6(CLBLM_R_X5Y142_SLICE_X7Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y142_SLICE_X7Y142_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y142_SLICE_X7Y142_BO5),
.O6(CLBLM_R_X5Y142_SLICE_X7Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y142_SLICE_X7Y142_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y142_SLICE_X7Y142_AO5),
.O6(CLBLM_R_X5Y142_SLICE_X7Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y143_SLICE_X6Y143_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y143_SLICE_X6Y143_AO6),
.Q(CLBLM_R_X5Y143_SLICE_X6Y143_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y143_SLICE_X6Y143_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y143_SLICE_X6Y143_DO5),
.O6(CLBLM_R_X5Y143_SLICE_X6Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y143_SLICE_X6Y143_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y143_SLICE_X6Y143_CO5),
.O6(CLBLM_R_X5Y143_SLICE_X6Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y143_SLICE_X6Y143_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y143_SLICE_X6Y143_BO5),
.O6(CLBLM_R_X5Y143_SLICE_X6Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffc000000fc00)
  ) CLBLM_R_X5Y143_SLICE_X6Y143_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y143_SLICE_X14Y143_AQ),
.I2(CLBLM_R_X5Y143_SLICE_X6Y143_AQ),
.I3(CLBLM_R_X7Y142_SLICE_X8Y142_DO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLL_L_X4Y145_SLICE_X4Y145_A5Q),
.O5(CLBLM_R_X5Y143_SLICE_X6Y143_AO5),
.O6(CLBLM_R_X5Y143_SLICE_X6Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y143_SLICE_X7Y143_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y143_SLICE_X7Y143_AO6),
.Q(CLBLM_R_X5Y143_SLICE_X7Y143_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y143_SLICE_X7Y143_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y143_SLICE_X7Y143_DO5),
.O6(CLBLM_R_X5Y143_SLICE_X7Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffff01ffffff00)
  ) CLBLM_R_X5Y143_SLICE_X7Y143_CLUT (
.I0(CLBLM_R_X3Y152_SLICE_X3Y152_CO6),
.I1(CLBLL_L_X2Y151_SLICE_X1Y151_BO6),
.I2(CLBLM_R_X5Y145_SLICE_X6Y145_DO6),
.I3(CLBLM_R_X5Y152_SLICE_X7Y152_B5Q),
.I4(CLBLL_L_X4Y144_SLICE_X5Y144_DO6),
.I5(CLBLM_R_X5Y143_SLICE_X7Y143_BO6),
.O5(CLBLM_R_X5Y143_SLICE_X7Y143_CO5),
.O6(CLBLM_R_X5Y143_SLICE_X7Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0001000103330fff)
  ) CLBLM_R_X5Y143_SLICE_X7Y143_BLUT (
.I0(CLBLL_L_X4Y154_SLICE_X4Y154_CO6),
.I1(CLBLM_R_X3Y153_SLICE_X2Y153_DO6),
.I2(CLBLL_L_X2Y153_SLICE_X1Y153_DO6),
.I3(CLBLM_R_X3Y154_SLICE_X2Y154_BO6),
.I4(CLBLM_R_X3Y152_SLICE_X3Y152_CO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y143_SLICE_X7Y143_BO5),
.O6(CLBLM_R_X5Y143_SLICE_X7Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0000ccccfff0)
  ) CLBLM_R_X5Y143_SLICE_X7Y143_ALUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y144_SLICE_X4Y144_BQ),
.I2(CLBLM_R_X5Y143_SLICE_X7Y143_AQ),
.I3(CLBLM_L_X8Y143_SLICE_X11Y143_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X5Y143_SLICE_X7Y143_CO6),
.O5(CLBLM_R_X5Y143_SLICE_X7Y143_AO5),
.O6(CLBLM_R_X5Y143_SLICE_X7Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y144_SLICE_X6Y144_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y144_SLICE_X6Y144_AO6),
.Q(CLBLM_R_X5Y144_SLICE_X6Y144_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffaffffffff)
  ) CLBLM_R_X5Y144_SLICE_X6Y144_DLUT (
.I0(CLBLL_L_X4Y148_SLICE_X4Y148_C5Q),
.I1(1'b1),
.I2(CLBLM_R_X5Y152_SLICE_X7Y152_B5Q),
.I3(CLBLM_R_X5Y144_SLICE_X6Y144_CO6),
.I4(CLBLM_R_X3Y145_SLICE_X3Y145_A5Q),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X5Y144_SLICE_X6Y144_DO5),
.O6(CLBLM_R_X5Y144_SLICE_X6Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_R_X5Y144_SLICE_X6Y144_CLUT (
.I0(CLBLM_R_X3Y149_SLICE_X3Y149_B5Q),
.I1(CLBLL_L_X4Y145_SLICE_X4Y145_A5Q),
.I2(CLBLM_R_X3Y144_SLICE_X2Y144_AQ),
.I3(CLBLM_R_X7Y145_SLICE_X8Y145_C5Q),
.I4(CLBLM_R_X3Y144_SLICE_X2Y144_A5Q),
.I5(CLBLM_R_X3Y143_SLICE_X3Y143_B5Q),
.O5(CLBLM_R_X5Y144_SLICE_X6Y144_CO5),
.O6(CLBLM_R_X5Y144_SLICE_X6Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000808080808080)
  ) CLBLM_R_X5Y144_SLICE_X6Y144_BLUT (
.I0(CLBLM_R_X7Y147_SLICE_X8Y147_B5Q),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X7Y147_SLICE_X8Y147_C5Q),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y144_SLICE_X6Y144_BO5),
.O6(CLBLM_R_X5Y144_SLICE_X6Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc5fffccccffff)
  ) CLBLM_R_X5Y144_SLICE_X6Y144_ALUT (
.I0(CLBLM_R_X7Y147_SLICE_X8Y147_B5Q),
.I1(CLBLM_R_X5Y147_SLICE_X7Y147_AQ),
.I2(CLBLM_R_X5Y144_SLICE_X6Y144_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y147_SLICE_X8Y147_C5Q),
.O5(CLBLM_R_X5Y144_SLICE_X6Y144_AO5),
.O6(CLBLM_R_X5Y144_SLICE_X6Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y144_SLICE_X7Y144_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y144_SLICE_X7Y144_BO5),
.Q(CLBLM_R_X5Y144_SLICE_X7Y144_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y144_SLICE_X7Y144_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y144_SLICE_X7Y144_AO6),
.Q(CLBLM_R_X5Y144_SLICE_X7Y144_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y144_SLICE_X7Y144_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y144_SLICE_X7Y144_BO6),
.Q(CLBLM_R_X5Y144_SLICE_X7Y144_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y144_SLICE_X7Y144_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y144_SLICE_X7Y144_CO6),
.Q(CLBLM_R_X5Y144_SLICE_X7Y144_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0500050100000101)
  ) CLBLM_R_X5Y144_SLICE_X7Y144_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y144_SLICE_X13Y144_AQ),
.I2(CLBLM_L_X8Y145_SLICE_X10Y145_CO6),
.I3(CLBLM_R_X5Y146_SLICE_X7Y146_AO5),
.I4(CLBLM_R_X5Y144_SLICE_X7Y144_AQ),
.I5(CLBLM_R_X3Y150_SLICE_X2Y150_BO6),
.O5(CLBLM_R_X5Y144_SLICE_X7Y144_DO5),
.O6(CLBLM_R_X5Y144_SLICE_X7Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaaf0aaccaac0)
  ) CLBLM_R_X5Y144_SLICE_X7Y144_CLUT (
.I0(CLBLM_R_X7Y143_SLICE_X8Y143_B5Q),
.I1(CLBLM_R_X5Y144_SLICE_X7Y144_CQ),
.I2(RIOB33_X105Y117_IOB_X1Y118_I),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.I5(CLBLM_R_X5Y146_SLICE_X7Y146_DO6),
.O5(CLBLM_R_X5Y144_SLICE_X7Y144_CO5),
.O6(CLBLM_R_X5Y144_SLICE_X7Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hacacacacfafa0a0a)
  ) CLBLM_R_X5Y144_SLICE_X7Y144_BLUT (
.I0(CLBLM_R_X7Y144_SLICE_X9Y144_A5Q),
.I1(CLBLM_R_X3Y148_SLICE_X3Y148_AQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(CLBLM_R_X5Y152_SLICE_X7Y152_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y144_SLICE_X7Y144_BO5),
.O6(CLBLM_R_X5Y144_SLICE_X7Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffef0f20f0e0002)
  ) CLBLM_R_X5Y144_SLICE_X7Y144_ALUT (
.I0(CLBLM_R_X5Y144_SLICE_X7Y144_AQ),
.I1(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_R_X11Y146_SLICE_X14Y146_AQ),
.I5(CLBLM_R_X3Y143_SLICE_X3Y143_A5Q),
.O5(CLBLM_R_X5Y144_SLICE_X7Y144_AO5),
.O6(CLBLM_R_X5Y144_SLICE_X7Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y145_SLICE_X6Y145_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y145_SLICE_X6Y145_BO6),
.Q(CLBLM_R_X5Y145_SLICE_X6Y145_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y145_SLICE_X6Y145_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y145_SLICE_X6Y145_AO6),
.Q(CLBLM_R_X5Y145_SLICE_X6Y145_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y145_SLICE_X6Y145_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y145_SLICE_X6Y145_CO6),
.Q(CLBLM_R_X5Y145_SLICE_X6Y145_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaaffaa69969669)
  ) CLBLM_R_X5Y145_SLICE_X6Y145_DLUT (
.I0(CLBLM_R_X3Y151_SLICE_X3Y151_AO6),
.I1(CLBLL_L_X2Y151_SLICE_X1Y151_BO6),
.I2(CLBLM_R_X3Y154_SLICE_X2Y154_BO6),
.I3(CLBLM_R_X3Y150_SLICE_X2Y150_BO6),
.I4(CLBLM_R_X5Y147_SLICE_X6Y147_DO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y145_SLICE_X6Y145_DO5),
.O6(CLBLM_R_X5Y145_SLICE_X6Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hae04aa00ae04aa00)
  ) CLBLM_R_X5Y145_SLICE_X6Y145_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y145_SLICE_X6Y145_CQ),
.I2(CLBLM_R_X5Y148_SLICE_X7Y148_CQ),
.I3(CLBLM_R_X5Y147_SLICE_X7Y147_CQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y145_SLICE_X6Y145_CO5),
.O6(CLBLM_R_X5Y145_SLICE_X6Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff00f00aaaa8888)
  ) CLBLM_R_X5Y145_SLICE_X6Y145_BLUT (
.I0(RIOB33_X105Y121_IOB_X1Y121_I),
.I1(CLBLM_L_X10Y146_SLICE_X13Y146_AQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLL_L_X4Y145_SLICE_X5Y145_AQ),
.I4(CLBLL_L_X4Y145_SLICE_X4Y145_BQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y145_SLICE_X6Y145_BO5),
.O6(CLBLM_R_X5Y145_SLICE_X6Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f6f600000606)
  ) CLBLM_R_X5Y145_SLICE_X6Y145_ALUT (
.I0(CLBLM_R_X5Y146_SLICE_X7Y146_AO5),
.I1(CLBLM_R_X5Y145_SLICE_X7Y145_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X5Y145_SLICE_X6Y145_A5Q),
.O5(CLBLM_R_X5Y145_SLICE_X6Y145_AO5),
.O6(CLBLM_R_X5Y145_SLICE_X6Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y145_SLICE_X7Y145_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y145_SLICE_X7Y145_AO6),
.Q(CLBLM_R_X5Y145_SLICE_X7Y145_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y145_SLICE_X7Y145_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y145_SLICE_X7Y145_BO6),
.Q(CLBLM_R_X5Y145_SLICE_X7Y145_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y145_SLICE_X7Y145_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y145_SLICE_X7Y145_CO6),
.Q(CLBLM_R_X5Y145_SLICE_X7Y145_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h404000003f3f3f3f)
  ) CLBLM_R_X5Y145_SLICE_X7Y145_DLUT (
.I0(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.I1(CLBLM_R_X7Y147_SLICE_X8Y147_AQ),
.I2(CLBLL_L_X4Y145_SLICE_X4Y145_CQ),
.I3(1'b1),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y145_SLICE_X7Y145_DO5),
.O6(CLBLM_R_X5Y145_SLICE_X7Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0b1e4a0a0b1e4)
  ) CLBLM_R_X5Y145_SLICE_X7Y145_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y148_SLICE_X10Y148_CO6),
.I2(CLBLM_R_X5Y145_SLICE_X7Y145_BQ),
.I3(CLBLM_R_X5Y147_SLICE_X7Y147_CQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y145_SLICE_X7Y145_CO5),
.O6(CLBLM_R_X5Y145_SLICE_X7Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf505f000f404f000)
  ) CLBLM_R_X5Y145_SLICE_X7Y145_BLUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_R_X5Y145_SLICE_X7Y145_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X5Y147_SLICE_X7Y147_D5Q),
.I4(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.I5(CLBLM_R_X11Y145_SLICE_X14Y145_AQ),
.O5(CLBLM_R_X5Y145_SLICE_X7Y145_BO5),
.O6(CLBLM_R_X5Y145_SLICE_X7Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc005a00f0)
  ) CLBLM_R_X5Y145_SLICE_X7Y145_ALUT (
.I0(CLBLM_R_X5Y145_SLICE_X7Y145_DO6),
.I1(CLBLM_R_X5Y148_SLICE_X6Y148_BQ),
.I2(CLBLM_R_X5Y145_SLICE_X7Y145_AQ),
.I3(CLBLM_R_X11Y146_SLICE_X14Y146_AQ),
.I4(CLBLM_R_X7Y145_SLICE_X8Y145_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X5Y145_SLICE_X7Y145_AO5),
.O6(CLBLM_R_X5Y145_SLICE_X7Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y146_SLICE_X6Y146_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y146_SLICE_X6Y146_BO6),
.Q(CLBLM_R_X5Y146_SLICE_X6Y146_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y146_SLICE_X6Y146_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y146_SLICE_X6Y146_AO6),
.Q(CLBLM_R_X5Y146_SLICE_X6Y146_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y146_SLICE_X6Y146_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y146_SLICE_X6Y146_CO6),
.Q(CLBLM_R_X5Y146_SLICE_X6Y146_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y146_SLICE_X6Y146_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y146_SLICE_X6Y146_DO6),
.Q(CLBLM_R_X5Y146_SLICE_X6Y146_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haeaeabab04040101)
  ) CLBLM_R_X5Y146_SLICE_X6Y146_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y146_SLICE_X7Y146_AO6),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(1'b1),
.I4(CLBLM_R_X7Y146_SLICE_X9Y146_AQ),
.I5(CLBLM_R_X5Y151_SLICE_X7Y151_AQ),
.O5(CLBLM_R_X5Y146_SLICE_X6Y146_DO5),
.O6(CLBLM_R_X5Y146_SLICE_X6Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hab01ae04ab01ae04)
  ) CLBLM_R_X5Y146_SLICE_X6Y146_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y146_SLICE_X8Y146_BO5),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X5Y150_SLICE_X6Y150_BQ),
.I4(CLBLM_L_X8Y146_SLICE_X10Y146_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y146_SLICE_X6Y146_CO5),
.O6(CLBLM_R_X5Y146_SLICE_X6Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fc00ccaaaa0000)
  ) CLBLM_R_X5Y146_SLICE_X6Y146_BLUT (
.I0(CLBLM_L_X10Y146_SLICE_X12Y146_CQ),
.I1(CLBLM_R_X5Y146_SLICE_X6Y146_A5Q),
.I2(CLBLM_R_X5Y150_SLICE_X6Y150_AQ),
.I3(CLBLL_L_X4Y145_SLICE_X5Y145_CO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y146_SLICE_X6Y146_BO5),
.O6(CLBLM_R_X5Y146_SLICE_X6Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0072725050)
  ) CLBLM_R_X5Y146_SLICE_X6Y146_ALUT (
.I0(CLBLL_L_X4Y149_SLICE_X5Y149_BO5),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X5Y146_SLICE_X6Y146_AQ),
.I3(CLBLM_R_X7Y146_SLICE_X9Y146_CQ),
.I4(CLBLM_R_X3Y151_SLICE_X3Y151_AO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X5Y146_SLICE_X6Y146_AO5),
.O6(CLBLM_R_X5Y146_SLICE_X6Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h55dd550055ff5500)
  ) CLBLM_R_X5Y146_SLICE_X7Y146_DLUT (
.I0(CLBLM_R_X5Y146_SLICE_X7Y146_AO6),
.I1(CLBLM_R_X3Y153_SLICE_X2Y153_DO6),
.I2(1'b1),
.I3(CLBLM_R_X5Y144_SLICE_X7Y144_AQ),
.I4(CLBLM_L_X10Y144_SLICE_X13Y144_AQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X5Y146_SLICE_X7Y146_DO5),
.O6(CLBLM_R_X5Y146_SLICE_X7Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h55ff7fff00003f3f)
  ) CLBLM_R_X5Y146_SLICE_X7Y146_CLUT (
.I0(CLBLM_R_X5Y145_SLICE_X7Y145_AQ),
.I1(CLBLM_L_X10Y147_SLICE_X12Y147_AQ),
.I2(CLBLM_R_X11Y147_SLICE_X14Y147_BQ),
.I3(CLBLM_R_X7Y145_SLICE_X8Y145_AQ),
.I4(CLBLL_L_X4Y146_SLICE_X5Y146_BO5),
.I5(CLBLM_R_X5Y145_SLICE_X7Y145_DO5),
.O5(CLBLM_R_X5Y146_SLICE_X7Y146_CO5),
.O6(CLBLM_R_X5Y146_SLICE_X7Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haabf0000bfbf0000)
  ) CLBLM_R_X5Y146_SLICE_X7Y146_BLUT (
.I0(CLBLM_R_X5Y143_SLICE_X7Y143_BO5),
.I1(CLBLL_L_X2Y151_SLICE_X1Y151_BO6),
.I2(CLBLM_R_X3Y151_SLICE_X3Y151_AO6),
.I3(CLBLM_R_X3Y150_SLICE_X2Y150_BO6),
.I4(CLBLM_R_X5Y146_SLICE_X7Y146_CO6),
.I5(CLBLL_L_X4Y154_SLICE_X4Y154_CO6),
.O5(CLBLM_R_X5Y146_SLICE_X7Y146_BO5),
.O6(CLBLM_R_X5Y146_SLICE_X7Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0fff8f8f8f8f)
  ) CLBLM_R_X5Y146_SLICE_X7Y146_ALUT (
.I0(CLBLL_L_X4Y149_SLICE_X5Y149_DQ),
.I1(CLBLM_R_X5Y148_SLICE_X6Y148_BQ),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.I4(CLBLL_L_X4Y148_SLICE_X4Y148_CQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y146_SLICE_X7Y146_AO5),
.O6(CLBLM_R_X5Y146_SLICE_X7Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y147_SLICE_X6Y147_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y147_SLICE_X6Y147_AO6),
.Q(CLBLM_R_X5Y147_SLICE_X6Y147_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y147_SLICE_X6Y147_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y147_SLICE_X6Y147_BO6),
.Q(CLBLM_R_X5Y147_SLICE_X6Y147_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y147_SLICE_X6Y147_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y147_SLICE_X6Y147_CO6),
.Q(CLBLM_R_X5Y147_SLICE_X6Y147_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h4bb4b44bb44b4bb4)
  ) CLBLM_R_X5Y147_SLICE_X6Y147_DLUT (
.I0(CLBLM_R_X7Y157_SLICE_X8Y157_AQ),
.I1(CLBLM_L_X16Y158_SLICE_X22Y158_AO5),
.I2(CLBLM_R_X3Y152_SLICE_X3Y152_CO6),
.I3(CLBLL_L_X4Y154_SLICE_X4Y154_CO6),
.I4(CLBLL_L_X2Y153_SLICE_X1Y153_DO6),
.I5(CLBLM_R_X3Y153_SLICE_X2Y153_DO6),
.O5(CLBLM_R_X5Y147_SLICE_X6Y147_DO5),
.O6(CLBLM_R_X5Y147_SLICE_X6Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h888d88d8888d88d8)
  ) CLBLM_R_X5Y147_SLICE_X6Y147_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y147_SLICE_X8Y147_B5Q),
.I2(CLBLM_R_X5Y145_SLICE_X6Y145_BO5),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLL_L_X4Y148_SLICE_X4Y148_BQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y147_SLICE_X6Y147_CO5),
.O6(CLBLM_R_X5Y147_SLICE_X6Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0ccffcc00)
  ) CLBLM_R_X5Y147_SLICE_X6Y147_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y147_SLICE_X6Y147_BQ),
.I2(CLBLM_L_X12Y144_SLICE_X16Y144_AQ),
.I3(CLBLM_R_X5Y152_SLICE_X7Y152_DO5),
.I4(CLBLL_L_X4Y148_SLICE_X4Y148_BQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X5Y147_SLICE_X6Y147_BO5),
.O6(CLBLM_R_X5Y147_SLICE_X6Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefcaa00fefcaa00)
  ) CLBLM_R_X5Y147_SLICE_X6Y147_ALUT (
.I0(CLBLM_L_X10Y147_SLICE_X13Y147_BQ),
.I1(CLBLM_R_X7Y151_SLICE_X9Y151_CQ),
.I2(CLBLM_R_X5Y147_SLICE_X6Y147_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X5Y152_SLICE_X7Y152_DO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y147_SLICE_X6Y147_AO5),
.O6(CLBLM_R_X5Y147_SLICE_X6Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y147_SLICE_X7Y147_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y147_SLICE_X7Y147_DO5),
.Q(CLBLM_R_X5Y147_SLICE_X7Y147_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y147_SLICE_X7Y147_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y147_SLICE_X7Y147_AO6),
.Q(CLBLM_R_X5Y147_SLICE_X7Y147_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y147_SLICE_X7Y147_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y147_SLICE_X7Y147_BO6),
.Q(CLBLM_R_X5Y147_SLICE_X7Y147_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y147_SLICE_X7Y147_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y147_SLICE_X7Y147_CO6),
.Q(CLBLM_R_X5Y147_SLICE_X7Y147_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y147_SLICE_X7Y147_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y147_SLICE_X7Y147_DO6),
.Q(CLBLM_R_X5Y147_SLICE_X7Y147_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff000f0aaccaacc)
  ) CLBLM_R_X5Y147_SLICE_X7Y147_DLUT (
.I0(CLBLM_R_X7Y157_SLICE_X8Y157_AQ),
.I1(CLBLL_L_X2Y147_SLICE_X1Y147_AQ),
.I2(CLBLM_R_X7Y148_SLICE_X8Y148_D5Q),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y153_SLICE_X10Y153_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y147_SLICE_X7Y147_DO5),
.O6(CLBLM_R_X5Y147_SLICE_X7Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888d8d8888d8d8)
  ) CLBLM_R_X5Y147_SLICE_X7Y147_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y146_SLICE_X10Y146_BQ),
.I2(CLBLM_R_X5Y146_SLICE_X6Y146_DQ),
.I3(1'b1),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X7Y147_SLICE_X9Y147_CO5),
.O5(CLBLM_R_X5Y147_SLICE_X7Y147_CO5),
.O6(CLBLM_R_X5Y147_SLICE_X7Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfef40e04fef40e04)
  ) CLBLM_R_X5Y147_SLICE_X7Y147_BLUT (
.I0(CLBLM_R_X5Y152_SLICE_X7Y152_DO5),
.I1(CLBLM_R_X5Y147_SLICE_X7Y147_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLL_L_X4Y147_SLICE_X4Y147_CQ),
.I4(CLBLM_L_X8Y143_SLICE_X11Y143_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y147_SLICE_X7Y147_BO5),
.O6(CLBLM_R_X5Y147_SLICE_X7Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccf505ccccf5f5)
  ) CLBLM_R_X5Y147_SLICE_X7Y147_ALUT (
.I0(CLBLL_L_X4Y150_SLICE_X4Y150_B5Q),
.I1(CLBLM_R_X15Y151_SLICE_X20Y151_AQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X5Y144_SLICE_X7Y144_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X3Y148_SLICE_X3Y148_AQ),
.O5(CLBLM_R_X5Y147_SLICE_X7Y147_AO5),
.O6(CLBLM_R_X5Y147_SLICE_X7Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y148_SLICE_X6Y148_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y148_SLICE_X6Y148_AO6),
.Q(CLBLM_R_X5Y148_SLICE_X6Y148_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y148_SLICE_X6Y148_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y148_SLICE_X6Y148_BO6),
.Q(CLBLM_R_X5Y148_SLICE_X6Y148_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffeeee)
  ) CLBLM_R_X5Y148_SLICE_X6Y148_DLUT (
.I0(CLBLL_L_X4Y148_SLICE_X4Y148_BQ),
.I1(CLBLM_R_X5Y145_SLICE_X7Y145_CQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X5Y147_SLICE_X7Y147_CQ),
.I5(CLBLM_R_X5Y149_SLICE_X7Y149_BQ),
.O5(CLBLM_R_X5Y148_SLICE_X6Y148_DO5),
.O6(CLBLM_R_X5Y148_SLICE_X6Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf7ffffffffffffff)
  ) CLBLM_R_X5Y148_SLICE_X6Y148_CLUT (
.I0(CLBLM_R_X7Y146_SLICE_X9Y146_AQ),
.I1(CLBLM_R_X5Y148_SLICE_X6Y148_AQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X5Y147_SLICE_X6Y147_CQ),
.I4(CLBLM_R_X5Y146_SLICE_X6Y146_DQ),
.I5(CLBLM_R_X5Y151_SLICE_X6Y151_CQ),
.O5(CLBLM_R_X5Y148_SLICE_X6Y148_CO5),
.O6(CLBLM_R_X5Y148_SLICE_X6Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000c0c0c0c0)
  ) CLBLM_R_X5Y148_SLICE_X6Y148_BLUT (
.I0(1'b1),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X5Y148_SLICE_X7Y148_C5Q),
.I3(1'b1),
.I4(CLBLM_R_X5Y150_SLICE_X6Y150_CQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X5Y148_SLICE_X6Y148_BO5),
.O6(CLBLM_R_X5Y148_SLICE_X6Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0000cccc55aa)
  ) CLBLM_R_X5Y148_SLICE_X6Y148_ALUT (
.I0(CLBLM_R_X7Y147_SLICE_X9Y147_CO6),
.I1(CLBLM_R_X5Y151_SLICE_X6Y151_CQ),
.I2(1'b1),
.I3(CLBLM_R_X5Y149_SLICE_X7Y149_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X5Y148_SLICE_X6Y148_AO5),
.O6(CLBLM_R_X5Y148_SLICE_X6Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y148_SLICE_X7Y148_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y148_SLICE_X7Y148_CO5),
.Q(CLBLM_R_X5Y148_SLICE_X7Y148_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y148_SLICE_X7Y148_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y148_SLICE_X7Y148_AO6),
.Q(CLBLM_R_X5Y148_SLICE_X7Y148_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y148_SLICE_X7Y148_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y148_SLICE_X7Y148_BO6),
.Q(CLBLM_R_X5Y148_SLICE_X7Y148_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y148_SLICE_X7Y148_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y148_SLICE_X7Y148_CO6),
.Q(CLBLM_R_X5Y148_SLICE_X7Y148_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffddff11ffccff00)
  ) CLBLM_R_X5Y148_SLICE_X7Y148_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X10Y144_SLICE_X13Y144_AQ),
.I2(1'b1),
.I3(CLBLM_R_X5Y144_SLICE_X7Y144_AQ),
.I4(CLBLM_R_X7Y147_SLICE_X9Y147_CO6),
.I5(CLBLM_R_X3Y154_SLICE_X2Y154_BO6),
.O5(CLBLM_R_X5Y148_SLICE_X7Y148_DO5),
.O6(CLBLM_R_X5Y148_SLICE_X7Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'he2e2e2e2cc00fc30)
  ) CLBLM_R_X5Y148_SLICE_X7Y148_CLUT (
.I0(CLBLM_R_X7Y148_SLICE_X8Y148_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y146_SLICE_X12Y146_DQ),
.I3(CLBLL_L_X4Y150_SLICE_X5Y150_BQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y148_SLICE_X7Y148_CO5),
.O6(CLBLM_R_X5Y148_SLICE_X7Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ffcc000000cc)
  ) CLBLM_R_X5Y148_SLICE_X7Y148_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y147_SLICE_X8Y147_CQ),
.I2(1'b1),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X5Y155_SLICE_X6Y155_BQ),
.O5(CLBLM_R_X5Y148_SLICE_X7Y148_BO5),
.O6(CLBLM_R_X5Y148_SLICE_X7Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff3333ccfc0030)
  ) CLBLM_R_X5Y148_SLICE_X7Y148_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X5Y148_SLICE_X7Y148_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X7Y148_SLICE_X8Y148_AQ),
.I5(CLBLM_R_X5Y150_SLICE_X7Y150_CO6),
.O5(CLBLM_R_X5Y148_SLICE_X7Y148_AO5),
.O6(CLBLM_R_X5Y148_SLICE_X7Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y149_SLICE_X6Y149_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y149_SLICE_X6Y149_AO6),
.Q(CLBLM_R_X5Y149_SLICE_X6Y149_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y149_SLICE_X6Y149_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y149_SLICE_X6Y149_BO6),
.Q(CLBLM_R_X5Y149_SLICE_X6Y149_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000008000000000)
  ) CLBLM_R_X5Y149_SLICE_X6Y149_DLUT (
.I0(CLBLM_R_X5Y145_SLICE_X6Y145_AQ),
.I1(CLBLM_L_X10Y150_SLICE_X13Y150_CQ),
.I2(CLBLM_L_X10Y145_SLICE_X12Y145_CQ),
.I3(CLBLM_R_X5Y148_SLICE_X6Y148_DO6),
.I4(CLBLM_R_X7Y151_SLICE_X8Y151_DO6),
.I5(CLBLM_R_X5Y151_SLICE_X6Y151_BQ),
.O5(CLBLM_R_X5Y149_SLICE_X6Y149_DO5),
.O6(CLBLM_R_X5Y149_SLICE_X6Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h000011000fff0fff)
  ) CLBLM_R_X5Y149_SLICE_X6Y149_CLUT (
.I0(RIOB33_X105Y135_IOB_X1Y136_I),
.I1(CLBLM_R_X5Y154_SLICE_X6Y154_BO6),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(RIOB33_X105Y135_IOB_X1Y135_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y149_SLICE_X6Y149_CO5),
.O6(CLBLM_R_X5Y149_SLICE_X6Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaf0ccf0cc)
  ) CLBLM_R_X5Y149_SLICE_X6Y149_BLUT (
.I0(CLBLM_L_X10Y148_SLICE_X13Y148_BQ),
.I1(CLBLM_R_X5Y149_SLICE_X6Y149_BQ),
.I2(CLBLM_L_X10Y149_SLICE_X13Y149_BQ),
.I3(CLBLM_R_X5Y152_SLICE_X7Y152_DO5),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X5Y149_SLICE_X6Y149_BO5),
.O6(CLBLM_R_X5Y149_SLICE_X6Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc00f0ccccaafa)
  ) CLBLM_R_X5Y149_SLICE_X6Y149_ALUT (
.I0(CLBLM_R_X5Y149_SLICE_X6Y149_DO6),
.I1(CLBLM_L_X10Y151_SLICE_X13Y151_AQ),
.I2(CLBLM_R_X5Y149_SLICE_X6Y149_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X5Y148_SLICE_X6Y148_CO6),
.O5(CLBLM_R_X5Y149_SLICE_X6Y149_AO5),
.O6(CLBLM_R_X5Y149_SLICE_X6Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y149_SLICE_X7Y149_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y149_SLICE_X7Y149_AO6),
.Q(CLBLM_R_X5Y149_SLICE_X7Y149_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y149_SLICE_X7Y149_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y149_SLICE_X7Y149_BO6),
.Q(CLBLM_R_X5Y149_SLICE_X7Y149_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y149_SLICE_X7Y149_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y149_SLICE_X7Y149_CO6),
.Q(CLBLM_R_X5Y149_SLICE_X7Y149_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0505050505050101)
  ) CLBLM_R_X5Y149_SLICE_X7Y149_DLUT (
.I0(CLBLL_L_X4Y149_SLICE_X5Y149_A5Q),
.I1(CLBLM_R_X3Y150_SLICE_X2Y150_BO6),
.I2(CLBLM_R_X5Y144_SLICE_X7Y144_AQ),
.I3(1'b1),
.I4(CLBLM_L_X10Y144_SLICE_X13Y144_AQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X5Y149_SLICE_X7Y149_DO5),
.O6(CLBLM_R_X5Y149_SLICE_X7Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0e4e4e4e4)
  ) CLBLM_R_X5Y149_SLICE_X7Y149_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y149_SLICE_X7Y149_CQ),
.I2(CLBLM_R_X7Y149_SLICE_X8Y149_DQ),
.I3(1'b1),
.I4(1'b1),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X5Y149_SLICE_X7Y149_CO5),
.O6(CLBLM_R_X5Y149_SLICE_X7Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc00aa0055)
  ) CLBLM_R_X5Y149_SLICE_X7Y149_BLUT (
.I0(CLBLL_L_X4Y146_SLICE_X4Y146_CO5),
.I1(CLBLM_R_X5Y151_SLICE_X7Y151_BQ),
.I2(1'b1),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X5Y147_SLICE_X6Y147_CQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X5Y149_SLICE_X7Y149_BO5),
.O6(CLBLM_R_X5Y149_SLICE_X7Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff001111ff004444)
  ) CLBLM_R_X5Y149_SLICE_X7Y149_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X7Y149_SLICE_X9Y149_BO6),
.I2(1'b1),
.I3(CLBLL_L_X4Y148_SLICE_X5Y148_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLL_L_X4Y147_SLICE_X4Y147_BQ),
.O5(CLBLM_R_X5Y149_SLICE_X7Y149_AO5),
.O6(CLBLM_R_X5Y149_SLICE_X7Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y150_SLICE_X6Y150_A5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y150_SLICE_X6Y150_AO5),
.Q(CLBLM_R_X5Y150_SLICE_X6Y150_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y150_SLICE_X6Y150_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y150_SLICE_X6Y150_AO6),
.Q(CLBLM_R_X5Y150_SLICE_X6Y150_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y150_SLICE_X6Y150_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y150_SLICE_X6Y150_BO6),
.Q(CLBLM_R_X5Y150_SLICE_X6Y150_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y150_SLICE_X6Y150_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y150_SLICE_X6Y150_CO6),
.Q(CLBLM_R_X5Y150_SLICE_X6Y150_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y150_SLICE_X6Y150_D_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y150_SLICE_X6Y150_DO6),
.Q(CLBLM_R_X5Y150_SLICE_X6Y150_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffaff00fafa0000)
  ) CLBLM_R_X5Y150_SLICE_X6Y150_DLUT (
.I0(CLBLM_R_X5Y145_SLICE_X6Y145_AQ),
.I1(1'b1),
.I2(CLBLM_R_X5Y150_SLICE_X6Y150_DQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X5Y152_SLICE_X7Y152_DO6),
.I5(CLBLM_R_X5Y147_SLICE_X6Y147_AQ),
.O5(CLBLM_R_X5Y150_SLICE_X6Y150_DO5),
.O6(CLBLM_R_X5Y150_SLICE_X6Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000ff00aaaa)
  ) CLBLM_R_X5Y150_SLICE_X6Y150_CLUT (
.I0(CLBLM_R_X5Y150_SLICE_X7Y150_AQ),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X7Y142_SLICE_X8Y142_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y153_SLICE_X10Y153_DO5),
.O5(CLBLM_R_X5Y150_SLICE_X6Y150_CO5),
.O6(CLBLM_R_X5Y150_SLICE_X6Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fe000efefe0e0e)
  ) CLBLM_R_X5Y150_SLICE_X6Y150_BLUT (
.I0(CLBLM_R_X5Y150_SLICE_X6Y150_BQ),
.I1(CLBLM_R_X3Y147_SLICE_X3Y147_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y148_SLICE_X10Y148_A5Q),
.I4(CLBLM_R_X5Y149_SLICE_X7Y149_CQ),
.I5(CLBLM_R_X11Y150_SLICE_X14Y150_AO6),
.O5(CLBLM_R_X5Y150_SLICE_X6Y150_BO5),
.O6(CLBLM_R_X5Y150_SLICE_X6Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcc00ccaaf0aaf0)
  ) CLBLM_R_X5Y150_SLICE_X6Y150_ALUT (
.I0(CLBLM_R_X7Y153_SLICE_X8Y153_BQ),
.I1(CLBLM_R_X3Y150_SLICE_X2Y150_BO6),
.I2(CLBLM_R_X3Y152_SLICE_X3Y152_CO6),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y144_SLICE_X13Y144_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y150_SLICE_X6Y150_AO5),
.O6(CLBLM_R_X5Y150_SLICE_X6Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y150_SLICE_X7Y150_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y150_SLICE_X7Y150_AO6),
.Q(CLBLM_R_X5Y150_SLICE_X7Y150_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y150_SLICE_X7Y150_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y150_SLICE_X7Y150_BO6),
.Q(CLBLM_R_X5Y150_SLICE_X7Y150_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbffffffffffffff)
  ) CLBLM_R_X5Y150_SLICE_X7Y150_DLUT (
.I0(CLBLM_R_X5Y149_SLICE_X7Y149_AQ),
.I1(CLBLM_R_X7Y151_SLICE_X9Y151_CQ),
.I2(1'b1),
.I3(CLBLM_R_X7Y153_SLICE_X9Y153_DQ),
.I4(CLBLM_R_X7Y149_SLICE_X8Y149_AQ),
.I5(CLBLL_L_X4Y147_SLICE_X4Y147_CQ),
.O5(CLBLM_R_X5Y150_SLICE_X7Y150_DO5),
.O6(CLBLM_R_X5Y150_SLICE_X7Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000050)
  ) CLBLM_R_X5Y150_SLICE_X7Y150_CLUT (
.I0(CLBLM_R_X3Y150_SLICE_X3Y150_AQ),
.I1(1'b1),
.I2(CLBLL_L_X4Y150_SLICE_X5Y150_CO6),
.I3(CLBLM_R_X7Y153_SLICE_X9Y153_A5Q),
.I4(CLBLM_R_X7Y152_SLICE_X9Y152_DO6),
.I5(CLBLM_R_X5Y150_SLICE_X7Y150_DO6),
.O5(CLBLM_R_X5Y150_SLICE_X7Y150_CO5),
.O6(CLBLM_R_X5Y150_SLICE_X7Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0055550000)
  ) CLBLM_R_X5Y150_SLICE_X7Y150_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X7Y147_SLICE_X8Y147_C5Q),
.I4(CLBLM_R_X3Y150_SLICE_X3Y150_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X5Y150_SLICE_X7Y150_BO5),
.O6(CLBLM_R_X5Y150_SLICE_X7Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbbbb8b8bbbbb8b8)
  ) CLBLM_R_X5Y150_SLICE_X7Y150_ALUT (
.I0(CLBLM_L_X8Y149_SLICE_X11Y149_B5Q),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X8Y153_SLICE_X10Y153_DO5),
.I3(1'b1),
.I4(CLBLM_R_X5Y152_SLICE_X6Y152_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y150_SLICE_X7Y150_AO5),
.O6(CLBLM_R_X5Y150_SLICE_X7Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y151_SLICE_X6Y151_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y151_SLICE_X6Y151_AO6),
.Q(CLBLM_R_X5Y151_SLICE_X6Y151_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y151_SLICE_X6Y151_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y151_SLICE_X6Y151_BO6),
.Q(CLBLM_R_X5Y151_SLICE_X6Y151_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y151_SLICE_X6Y151_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y151_SLICE_X6Y151_CO6),
.Q(CLBLM_R_X5Y151_SLICE_X6Y151_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y151_SLICE_X6Y151_D_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y151_SLICE_X6Y151_DO6),
.Q(CLBLM_R_X5Y151_SLICE_X6Y151_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00fa50ee44fa50)
  ) CLBLM_R_X5Y151_SLICE_X6Y151_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLL_L_X2Y151_SLICE_X1Y151_BO6),
.I2(CLBLM_R_X5Y151_SLICE_X6Y151_DQ),
.I3(CLBLM_L_X8Y151_SLICE_X11Y151_BQ),
.I4(CLBLL_L_X4Y149_SLICE_X5Y149_BO5),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X5Y151_SLICE_X6Y151_DO5),
.O6(CLBLM_R_X5Y151_SLICE_X6Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00ff55aa00)
  ) CLBLM_R_X5Y151_SLICE_X6Y151_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X5Y151_SLICE_X7Y151_CQ),
.I4(CLBLM_L_X10Y149_SLICE_X13Y149_BQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X5Y151_SLICE_X6Y151_CO5),
.O6(CLBLM_R_X5Y151_SLICE_X6Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000000aa00aa)
  ) CLBLM_R_X5Y151_SLICE_X6Y151_BLUT (
.I0(CLBLM_R_X5Y151_SLICE_X6Y151_CQ),
.I1(1'b1),
.I2(1'b1),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLL_L_X4Y148_SLICE_X5Y148_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X5Y151_SLICE_X6Y151_BO5),
.O6(CLBLM_R_X5Y151_SLICE_X6Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccfff0cccc00f0)
  ) CLBLM_R_X5Y151_SLICE_X6Y151_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y147_SLICE_X6Y147_BQ),
.I2(CLBLM_R_X5Y151_SLICE_X6Y151_AQ),
.I3(CLBLM_R_X5Y152_SLICE_X7Y152_DO5),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X5Y146_SLICE_X6Y146_DQ),
.O5(CLBLM_R_X5Y151_SLICE_X6Y151_AO5),
.O6(CLBLM_R_X5Y151_SLICE_X6Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y151_SLICE_X7Y151_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y151_SLICE_X7Y151_AO6),
.Q(CLBLM_R_X5Y151_SLICE_X7Y151_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y151_SLICE_X7Y151_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y151_SLICE_X7Y151_BO6),
.Q(CLBLM_R_X5Y151_SLICE_X7Y151_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y151_SLICE_X7Y151_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y151_SLICE_X7Y151_CO6),
.Q(CLBLM_R_X5Y151_SLICE_X7Y151_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00300030cece0202)
  ) CLBLM_R_X5Y151_SLICE_X7Y151_DLUT (
.I0(CLBLM_R_X5Y149_SLICE_X7Y149_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X5Y152_SLICE_X7Y152_BQ),
.I4(CLBLL_L_X4Y150_SLICE_X4Y150_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y151_SLICE_X7Y151_DO5),
.O6(CLBLM_R_X5Y151_SLICE_X7Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hafaaeeee05004444)
  ) CLBLM_R_X5Y151_SLICE_X7Y151_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y151_SLICE_X7Y151_CQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLL_L_X4Y154_SLICE_X4Y154_CO6),
.I4(CLBLL_L_X4Y149_SLICE_X5Y149_BO5),
.I5(CLBLM_R_X5Y145_SLICE_X7Y145_CQ),
.O5(CLBLM_R_X5Y151_SLICE_X7Y151_CO5),
.O6(CLBLM_R_X5Y151_SLICE_X7Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffcf0fc0f0c000c)
  ) CLBLM_R_X5Y151_SLICE_X7Y151_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y151_SLICE_X7Y151_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X5Y152_SLICE_X7Y152_DO5),
.I4(CLBLL_L_X4Y147_SLICE_X4Y147_BQ),
.I5(CLBLM_R_X7Y153_SLICE_X8Y153_AQ),
.O5(CLBLM_R_X5Y151_SLICE_X7Y151_BO5),
.O6(CLBLM_R_X5Y151_SLICE_X7Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa33ff30f0)
  ) CLBLM_R_X5Y151_SLICE_X7Y151_ALUT (
.I0(CLBLM_L_X10Y155_SLICE_X12Y155_AQ),
.I1(CLBLL_L_X4Y151_SLICE_X4Y151_AQ),
.I2(CLBLM_R_X5Y151_SLICE_X7Y151_AQ),
.I3(CLBLM_L_X8Y149_SLICE_X11Y149_AQ),
.I4(CLBLM_R_X7Y147_SLICE_X8Y147_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X5Y151_SLICE_X7Y151_AO5),
.O6(CLBLM_R_X5Y151_SLICE_X7Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y152_SLICE_X6Y152_A5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y151_SLICE_X7Y151_DO5),
.Q(CLBLM_R_X5Y152_SLICE_X6Y152_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y152_SLICE_X6Y152_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y152_SLICE_X6Y152_AO6),
.Q(CLBLM_R_X5Y152_SLICE_X6Y152_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y152_SLICE_X6Y152_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y152_SLICE_X6Y152_BO6),
.Q(CLBLM_R_X5Y152_SLICE_X6Y152_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y152_SLICE_X6Y152_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y152_SLICE_X6Y152_CO6),
.Q(CLBLM_R_X5Y152_SLICE_X6Y152_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h1110111000100010)
  ) CLBLM_R_X5Y152_SLICE_X6Y152_DLUT (
.I0(CLBLL_L_X4Y154_SLICE_X5Y154_CO5),
.I1(CLBLL_L_X2Y155_SLICE_X1Y155_DO6),
.I2(CLBLM_R_X7Y152_SLICE_X8Y152_CQ),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(1'b1),
.I5(CLBLM_R_X7Y152_SLICE_X8Y152_BQ),
.O5(CLBLM_R_X5Y152_SLICE_X6Y152_DO5),
.O6(CLBLM_R_X5Y152_SLICE_X6Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaccfcaaaa0000)
  ) CLBLM_R_X5Y152_SLICE_X6Y152_CLUT (
.I0(CLBLM_R_X5Y146_SLICE_X6Y146_AQ),
.I1(CLBLM_R_X5Y152_SLICE_X6Y152_CQ),
.I2(CLBLM_R_X11Y146_SLICE_X14Y146_DQ),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X5Y152_SLICE_X6Y152_CO5),
.O6(CLBLM_R_X5Y152_SLICE_X6Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccffcc00003300)
  ) CLBLM_R_X5Y152_SLICE_X6Y152_BLUT (
.I0(1'b1),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(1'b1),
.I3(CLBLM_R_X5Y150_SLICE_X6Y150_CQ),
.I4(CLBLM_L_X8Y153_SLICE_X10Y153_DO5),
.I5(CLBLM_L_X8Y152_SLICE_X10Y152_BQ),
.O5(CLBLM_R_X5Y152_SLICE_X6Y152_BO5),
.O6(CLBLM_R_X5Y152_SLICE_X6Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00fc30fc30)
  ) CLBLM_R_X5Y152_SLICE_X6Y152_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X7Y152_SLICE_X9Y152_AQ),
.I3(CLBLM_R_X3Y150_SLICE_X3Y150_BQ),
.I4(1'b1),
.I5(CLBLM_L_X8Y153_SLICE_X10Y153_DO5),
.O5(CLBLM_R_X5Y152_SLICE_X6Y152_AO5),
.O6(CLBLM_R_X5Y152_SLICE_X6Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y152_SLICE_X7Y152_B5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y152_SLICE_X7Y152_BO5),
.Q(CLBLM_R_X5Y152_SLICE_X7Y152_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y152_SLICE_X7Y152_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y152_SLICE_X7Y152_AO6),
.Q(CLBLM_R_X5Y152_SLICE_X7Y152_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y152_SLICE_X7Y152_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y152_SLICE_X7Y152_BO6),
.Q(CLBLM_R_X5Y152_SLICE_X7Y152_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y152_SLICE_X7Y152_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y152_SLICE_X7Y152_CO6),
.Q(CLBLM_R_X5Y152_SLICE_X7Y152_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h50405050f0c0f0f0)
  ) CLBLM_R_X5Y152_SLICE_X7Y152_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y121_IOB_X1Y121_I),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X5Y152_SLICE_X6Y152_CQ),
.I4(CLBLM_R_X11Y146_SLICE_X14Y146_DQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y152_SLICE_X7Y152_DO5),
.O6(CLBLM_R_X5Y152_SLICE_X7Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0f5f5e4e4)
  ) CLBLM_R_X5Y152_SLICE_X7Y152_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y152_SLICE_X7Y152_CQ),
.I2(CLBLM_L_X10Y153_SLICE_X12Y153_BQ),
.I3(1'b1),
.I4(CLBLM_R_X3Y149_SLICE_X3Y149_B5Q),
.I5(CLBLM_R_X3Y144_SLICE_X2Y144_CO6),
.O5(CLBLM_R_X5Y152_SLICE_X7Y152_CO5),
.O6(CLBLM_R_X5Y152_SLICE_X7Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0aaf0aaffcc00cc)
  ) CLBLM_R_X5Y152_SLICE_X7Y152_BLUT (
.I0(CLBLM_R_X7Y153_SLICE_X8Y153_AQ),
.I1(CLBLM_R_X3Y145_SLICE_X3Y145_CQ),
.I2(CLBLM_R_X7Y154_SLICE_X8Y154_BQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y143_SLICE_X8Y143_CQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y152_SLICE_X7Y152_BO5),
.O6(CLBLM_R_X5Y152_SLICE_X7Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heeecaaa0eeecaaa0)
  ) CLBLM_R_X5Y152_SLICE_X7Y152_ALUT (
.I0(CLBLM_R_X5Y152_SLICE_X7Y152_DO6),
.I1(CLBLM_R_X5Y144_SLICE_X7Y144_CQ),
.I2(CLBLM_R_X5Y152_SLICE_X7Y152_AQ),
.I3(CLBLM_R_X5Y149_SLICE_X7Y149_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y152_SLICE_X7Y152_AO5),
.O6(CLBLM_R_X5Y152_SLICE_X7Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y153_SLICE_X6Y153_A5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y153_SLICE_X6Y153_CO5),
.Q(CLBLM_R_X5Y153_SLICE_X6Y153_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y153_SLICE_X6Y153_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y153_SLICE_X6Y153_AO6),
.Q(CLBLM_R_X5Y153_SLICE_X6Y153_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y153_SLICE_X6Y153_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y153_SLICE_X6Y153_BO6),
.Q(CLBLM_R_X5Y153_SLICE_X6Y153_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfffcfcfefffefe)
  ) CLBLM_R_X5Y153_SLICE_X6Y153_DLUT (
.I0(CLBLM_R_X7Y152_SLICE_X8Y152_AQ),
.I1(CLBLM_R_X5Y153_SLICE_X7Y153_CO6),
.I2(CLBLM_R_X5Y153_SLICE_X7Y153_DO6),
.I3(CLBLL_L_X2Y154_SLICE_X1Y154_AO5),
.I4(CLBLM_R_X5Y151_SLICE_X6Y151_DQ),
.I5(CLBLM_R_X5Y154_SLICE_X7Y154_AO6),
.O5(CLBLM_R_X5Y153_SLICE_X6Y153_DO5),
.O6(CLBLM_R_X5Y153_SLICE_X6Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hafafafafbbaa3300)
  ) CLBLM_R_X5Y153_SLICE_X6Y153_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLL_L_X4Y145_SLICE_X5Y145_CO6),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLM_R_X5Y153_SLICE_X6Y153_A5Q),
.I4(CLBLM_L_X10Y154_SLICE_X12Y154_BQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y153_SLICE_X6Y153_CO5),
.O6(CLBLM_R_X5Y153_SLICE_X6Y153_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaf0aaccaaf0aacc)
  ) CLBLM_R_X5Y153_SLICE_X6Y153_BLUT (
.I0(CLBLM_R_X3Y145_SLICE_X3Y145_DQ),
.I1(CLBLM_R_X5Y153_SLICE_X6Y153_BQ),
.I2(CLBLM_L_X10Y150_SLICE_X13Y150_CQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X5Y152_SLICE_X7Y152_DO5),
.I5(1'b1),
.O5(CLBLM_R_X5Y153_SLICE_X6Y153_BO5),
.O6(CLBLM_R_X5Y153_SLICE_X6Y153_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffaff5000fa0050)
  ) CLBLM_R_X5Y153_SLICE_X6Y153_ALUT (
.I0(CLBLM_L_X8Y152_SLICE_X11Y152_BO6),
.I1(1'b1),
.I2(CLBLM_R_X5Y153_SLICE_X6Y153_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y146_SLICE_X10Y146_AQ),
.I5(CLBLM_R_X3Y145_SLICE_X3Y145_CQ),
.O5(CLBLM_R_X5Y153_SLICE_X6Y153_AO5),
.O6(CLBLM_R_X5Y153_SLICE_X6Y153_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y153_SLICE_X7Y153_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y153_SLICE_X7Y153_AO6),
.Q(CLBLM_R_X5Y153_SLICE_X7Y153_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y153_SLICE_X7Y153_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y153_SLICE_X7Y153_BO6),
.Q(CLBLM_R_X5Y153_SLICE_X7Y153_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000040)
  ) CLBLM_R_X5Y153_SLICE_X7Y153_DLUT (
.I0(RIOB33_X105Y133_IOB_X1Y133_I),
.I1(CLBLM_R_X11Y147_SLICE_X15Y147_CQ),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(CLBLL_L_X2Y155_SLICE_X1Y155_DO6),
.I4(RIOB33_X105Y133_IOB_X1Y134_I),
.I5(RIOB33_X105Y131_IOB_X1Y131_I),
.O5(CLBLM_R_X5Y153_SLICE_X7Y153_DO5),
.O6(CLBLM_R_X5Y153_SLICE_X7Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000080)
  ) CLBLM_R_X5Y153_SLICE_X7Y153_CLUT (
.I0(CLBLM_R_X7Y150_SLICE_X9Y150_AQ),
.I1(RIOB33_X105Y131_IOB_X1Y132_I),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(CLBLL_L_X2Y155_SLICE_X1Y155_DO6),
.I4(RIOB33_X105Y133_IOB_X1Y134_I),
.I5(RIOB33_X105Y133_IOB_X1Y133_I),
.O5(CLBLM_R_X5Y153_SLICE_X7Y153_CO5),
.O6(CLBLM_R_X5Y153_SLICE_X7Y153_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf505f505f404f404)
  ) CLBLM_R_X5Y153_SLICE_X7Y153_BLUT (
.I0(CLBLM_R_X3Y144_SLICE_X2Y144_CO6),
.I1(CLBLM_R_X5Y153_SLICE_X7Y153_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y154_SLICE_X9Y154_BQ),
.I4(1'b1),
.I5(CLBLM_R_X3Y145_SLICE_X3Y145_A5Q),
.O5(CLBLM_R_X5Y153_SLICE_X7Y153_BO5),
.O6(CLBLM_R_X5Y153_SLICE_X7Y153_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0f3c0f3c0c0c0d1)
  ) CLBLM_R_X5Y153_SLICE_X7Y153_ALUT (
.I0(CLBLM_R_X7Y153_SLICE_X8Y153_CQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLL_L_X4Y142_SLICE_X5Y142_AQ),
.I3(CLBLM_R_X7Y154_SLICE_X8Y154_BQ),
.I4(CLBLL_L_X4Y147_SLICE_X5Y147_B5Q),
.I5(CLBLM_R_X7Y155_SLICE_X8Y155_A5Q),
.O5(CLBLM_R_X5Y153_SLICE_X7Y153_AO5),
.O6(CLBLM_R_X5Y153_SLICE_X7Y153_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y154_SLICE_X6Y154_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y154_SLICE_X6Y154_AO6),
.Q(CLBLM_R_X5Y154_SLICE_X6Y154_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y154_SLICE_X6Y154_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y154_SLICE_X6Y154_DO5),
.O6(CLBLM_R_X5Y154_SLICE_X6Y154_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y154_SLICE_X6Y154_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y154_SLICE_X6Y154_CO5),
.O6(CLBLM_R_X5Y154_SLICE_X6Y154_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_R_X5Y154_SLICE_X6Y154_BLUT (
.I0(RIOB33_X105Y127_IOB_X1Y128_I),
.I1(RIOB33_X105Y129_IOB_X1Y130_I),
.I2(RIOB33_X105Y137_IOB_X1Y137_I),
.I3(RIOB33_X105Y133_IOB_X1Y134_I),
.I4(RIOB33_X105Y131_IOB_X1Y132_I),
.I5(RIOB33_X105Y133_IOB_X1Y133_I),
.O5(CLBLM_R_X5Y154_SLICE_X6Y154_BO5),
.O6(CLBLM_R_X5Y154_SLICE_X6Y154_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00e4e4e4e4)
  ) CLBLM_R_X5Y154_SLICE_X6Y154_ALUT (
.I0(CLBLM_R_X5Y152_SLICE_X7Y152_DO5),
.I1(CLBLM_R_X7Y154_SLICE_X9Y154_AQ),
.I2(CLBLM_R_X5Y154_SLICE_X6Y154_AQ),
.I3(CLBLM_R_X5Y149_SLICE_X7Y149_BQ),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X5Y154_SLICE_X6Y154_AO5),
.O6(CLBLM_R_X5Y154_SLICE_X6Y154_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff44f444f4)
  ) CLBLM_R_X5Y154_SLICE_X7Y154_DLUT (
.I0(CLBLM_R_X5Y154_SLICE_X7Y154_AO6),
.I1(CLBLM_L_X8Y151_SLICE_X11Y151_AQ),
.I2(CLBLM_L_X10Y153_SLICE_X12Y153_CQ),
.I3(CLBLM_R_X5Y154_SLICE_X7Y154_AO5),
.I4(1'b1),
.I5(CLBLM_R_X5Y154_SLICE_X7Y154_BO6),
.O5(CLBLM_R_X5Y154_SLICE_X7Y154_DO5),
.O6(CLBLM_R_X5Y154_SLICE_X7Y154_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffbffffff)
  ) CLBLM_R_X5Y154_SLICE_X7Y154_CLUT (
.I0(RIOB33_X105Y135_IOB_X1Y135_I),
.I1(RIOB33_X105Y135_IOB_X1Y136_I),
.I2(RIOB33_X105Y129_IOB_X1Y129_I),
.I3(RIOB33_X105Y137_IOB_X1Y137_I),
.I4(RIOB33_X105Y131_IOB_X1Y132_I),
.I5(RIOB33_X105Y129_IOB_X1Y130_I),
.O5(CLBLM_R_X5Y154_SLICE_X7Y154_CO5),
.O6(CLBLM_R_X5Y154_SLICE_X7Y154_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000088800800)
  ) CLBLM_R_X5Y154_SLICE_X7Y154_BLUT (
.I0(RIOB33_X105Y133_IOB_X1Y133_I),
.I1(RIOB33_X105Y133_IOB_X1Y134_I),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(CLBLL_L_X4Y148_SLICE_X5Y148_AQ),
.I4(CLBLM_R_X5Y151_SLICE_X7Y151_CQ),
.I5(CLBLM_R_X5Y154_SLICE_X7Y154_CO6),
.O5(CLBLM_R_X5Y154_SLICE_X7Y154_BO5),
.O6(CLBLM_R_X5Y154_SLICE_X7Y154_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffdfffeffff)
  ) CLBLM_R_X5Y154_SLICE_X7Y154_ALUT (
.I0(RIOB33_X105Y133_IOB_X1Y133_I),
.I1(RIOB33_X105Y133_IOB_X1Y134_I),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(CLBLL_L_X2Y155_SLICE_X1Y155_DO6),
.I4(RIOB33_X105Y131_IOB_X1Y132_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y154_SLICE_X7Y154_AO5),
.O6(CLBLM_R_X5Y154_SLICE_X7Y154_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y155_SLICE_X6Y155_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y155_SLICE_X6Y155_AO6),
.Q(CLBLM_R_X5Y155_SLICE_X6Y155_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y155_SLICE_X6Y155_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y155_SLICE_X6Y155_BO6),
.Q(CLBLM_R_X5Y155_SLICE_X6Y155_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y155_SLICE_X6Y155_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y155_SLICE_X6Y155_DO5),
.O6(CLBLM_R_X5Y155_SLICE_X6Y155_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y155_SLICE_X6Y155_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y155_SLICE_X6Y155_CO5),
.O6(CLBLM_R_X5Y155_SLICE_X6Y155_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf303f000fc0cf000)
  ) CLBLM_R_X5Y155_SLICE_X6Y155_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y155_SLICE_X6Y155_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X5Y154_SLICE_X6Y154_AQ),
.I4(CLBLM_R_X5Y155_SLICE_X7Y155_BO6),
.I5(CLBLM_R_X5Y152_SLICE_X6Y152_AQ),
.O5(CLBLM_R_X5Y155_SLICE_X6Y155_BO5),
.O6(CLBLM_R_X5Y155_SLICE_X6Y155_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hebfaaaaa41500000)
  ) CLBLM_R_X5Y155_SLICE_X6Y155_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y155_SLICE_X6Y155_BQ),
.I2(CLBLM_R_X5Y155_SLICE_X6Y155_AQ),
.I3(CLBLM_R_X5Y152_SLICE_X6Y152_AQ),
.I4(CLBLM_R_X5Y155_SLICE_X7Y155_BO6),
.I5(CLBLM_R_X7Y152_SLICE_X8Y152_BQ),
.O5(CLBLM_R_X5Y155_SLICE_X6Y155_AO5),
.O6(CLBLM_R_X5Y155_SLICE_X6Y155_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y155_SLICE_X7Y155_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y155_SLICE_X7Y155_AO6),
.Q(CLBLM_R_X5Y155_SLICE_X7Y155_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000044444444)
  ) CLBLM_R_X5Y155_SLICE_X7Y155_DLUT (
.I0(CLBLM_R_X5Y155_SLICE_X6Y155_AQ),
.I1(CLBLM_R_X5Y152_SLICE_X6Y152_AQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X5Y155_SLICE_X6Y155_BQ),
.O5(CLBLM_R_X5Y155_SLICE_X7Y155_DO5),
.O6(CLBLM_R_X5Y155_SLICE_X7Y155_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000040)
  ) CLBLM_R_X5Y155_SLICE_X7Y155_CLUT (
.I0(CLBLM_R_X5Y155_SLICE_X6Y155_AQ),
.I1(CLBLM_R_X5Y152_SLICE_X6Y152_AQ),
.I2(CLBLM_R_X7Y155_SLICE_X8Y155_AQ),
.I3(CLBLM_R_X7Y155_SLICE_X8Y155_A5Q),
.I4(CLBLM_R_X5Y155_SLICE_X7Y155_AQ),
.I5(CLBLM_R_X5Y155_SLICE_X6Y155_BQ),
.O5(CLBLM_R_X5Y155_SLICE_X7Y155_CO5),
.O6(CLBLM_R_X5Y155_SLICE_X7Y155_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h555555510000000c)
  ) CLBLM_R_X5Y155_SLICE_X7Y155_BLUT (
.I0(CLBLM_R_X7Y155_SLICE_X8Y155_BO5),
.I1(CLBLM_R_X5Y152_SLICE_X6Y152_AQ),
.I2(CLBLM_R_X5Y155_SLICE_X7Y155_AQ),
.I3(CLBLM_R_X5Y155_SLICE_X6Y155_BQ),
.I4(CLBLM_R_X5Y155_SLICE_X6Y155_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y155_SLICE_X7Y155_BO5),
.O6(CLBLM_R_X5Y155_SLICE_X7Y155_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff50f05fffa0f0a)
  ) CLBLM_R_X5Y155_SLICE_X7Y155_ALUT (
.I0(CLBLM_R_X5Y155_SLICE_X7Y155_DO6),
.I1(1'b1),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y155_SLICE_X8Y155_BO5),
.I4(CLBLM_R_X5Y149_SLICE_X7Y149_AQ),
.I5(CLBLM_R_X5Y155_SLICE_X7Y155_AQ),
.O5(CLBLM_R_X5Y155_SLICE_X7Y155_AO5),
.O6(CLBLM_R_X5Y155_SLICE_X7Y155_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y142_SLICE_X8Y142_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y142_SLICE_X8Y142_BO6),
.Q(CLBLM_R_X7Y142_SLICE_X8Y142_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y142_SLICE_X8Y142_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y142_SLICE_X8Y142_CO6),
.Q(CLBLM_R_X7Y142_SLICE_X8Y142_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ffef0000ffef)
  ) CLBLM_R_X7Y142_SLICE_X8Y142_DLUT (
.I0(CLBLM_R_X3Y152_SLICE_X3Y152_CO6),
.I1(CLBLM_R_X5Y145_SLICE_X6Y145_DO6),
.I2(CLBLM_R_X5Y143_SLICE_X7Y143_BO6),
.I3(CLBLL_L_X2Y151_SLICE_X1Y151_BO6),
.I4(CLBLM_R_X5Y144_SLICE_X6Y144_DO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y142_SLICE_X8Y142_DO5),
.O6(CLBLM_R_X7Y142_SLICE_X8Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hafaca0a0afaca0a0)
  ) CLBLM_R_X7Y142_SLICE_X8Y142_CLUT (
.I0(CLBLM_R_X3Y148_SLICE_X3Y148_AQ),
.I1(CLBLM_R_X7Y142_SLICE_X8Y142_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y142_SLICE_X8Y142_BQ),
.I4(CLBLM_R_X7Y142_SLICE_X8Y142_DO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y142_SLICE_X8Y142_CO5),
.O6(CLBLM_R_X7Y142_SLICE_X8Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfc0cfc0cac0cac0)
  ) CLBLM_R_X7Y142_SLICE_X8Y142_BLUT (
.I0(CLBLM_R_X7Y144_SLICE_X8Y144_DQ),
.I1(CLBLM_L_X8Y142_SLICE_X10Y142_AQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y142_SLICE_X8Y142_DO6),
.I4(1'b1),
.I5(CLBLM_R_X7Y142_SLICE_X8Y142_BQ),
.O5(CLBLM_R_X7Y142_SLICE_X8Y142_BO5),
.O6(CLBLM_R_X7Y142_SLICE_X8Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaf3aa0033330000)
  ) CLBLM_R_X7Y142_SLICE_X8Y142_ALUT (
.I0(CLBLM_R_X7Y144_SLICE_X8Y144_DQ),
.I1(RIOB33_X105Y141_IOB_X1Y142_I),
.I2(CLBLM_R_X5Y142_SLICE_X7Y142_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y147_SLICE_X8Y147_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X7Y142_SLICE_X8Y142_AO5),
.O6(CLBLM_R_X7Y142_SLICE_X8Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y142_SLICE_X9Y142_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y142_SLICE_X9Y142_DO5),
.O6(CLBLM_R_X7Y142_SLICE_X9Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y142_SLICE_X9Y142_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y142_SLICE_X9Y142_CO5),
.O6(CLBLM_R_X7Y142_SLICE_X9Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y142_SLICE_X9Y142_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y142_SLICE_X9Y142_BO5),
.O6(CLBLM_R_X7Y142_SLICE_X9Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafafafafafafafa)
  ) CLBLM_R_X7Y142_SLICE_X9Y142_ALUT (
.I0(CLBLL_L_X2Y151_SLICE_X1Y151_BO6),
.I1(1'b1),
.I2(CLBLM_R_X3Y152_SLICE_X3Y152_CO6),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y142_SLICE_X9Y142_AO5),
.O6(CLBLM_R_X7Y142_SLICE_X9Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y143_SLICE_X8Y143_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y143_SLICE_X8Y143_BO5),
.Q(CLBLM_R_X7Y143_SLICE_X8Y143_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y143_SLICE_X8Y143_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y143_SLICE_X8Y143_AO6),
.Q(CLBLM_R_X7Y143_SLICE_X8Y143_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y143_SLICE_X8Y143_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y143_SLICE_X8Y143_BO6),
.Q(CLBLM_R_X7Y143_SLICE_X8Y143_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y143_SLICE_X8Y143_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y143_SLICE_X8Y143_CO6),
.Q(CLBLM_R_X7Y143_SLICE_X8Y143_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0011223302132031)
  ) CLBLM_R_X7Y143_SLICE_X8Y143_DLUT (
.I0(CLBLM_R_X7Y142_SLICE_X8Y142_DO6),
.I1(CLBLM_R_X7Y143_SLICE_X8Y143_CQ),
.I2(CLBLM_L_X12Y144_SLICE_X16Y144_CQ),
.I3(CLBLM_L_X8Y145_SLICE_X11Y145_BQ),
.I4(CLBLM_R_X7Y146_SLICE_X9Y146_CQ),
.I5(CLBLM_L_X10Y142_SLICE_X13Y142_BO6),
.O5(CLBLM_R_X7Y143_SLICE_X8Y143_DO5),
.O6(CLBLM_R_X7Y143_SLICE_X8Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f00000aaff)
  ) CLBLM_R_X7Y143_SLICE_X8Y143_CLUT (
.I0(CLBLM_R_X5Y142_SLICE_X7Y142_AQ),
.I1(1'b1),
.I2(CLBLM_R_X7Y145_SLICE_X8Y145_CQ),
.I3(RIOB33_X105Y141_IOB_X1Y142_I),
.I4(CLBLM_R_X7Y143_SLICE_X8Y143_DO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X7Y143_SLICE_X8Y143_CO5),
.O6(CLBLM_R_X7Y143_SLICE_X8Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccf0f0aaaaf0f0)
  ) CLBLM_R_X7Y143_SLICE_X8Y143_BLUT (
.I0(CLBLL_L_X4Y148_SLICE_X4Y148_AQ),
.I1(CLBLM_R_X7Y144_SLICE_X9Y144_BQ),
.I2(RIOB33_X105Y101_IOB_X1Y101_I),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y143_SLICE_X8Y143_BO5),
.O6(CLBLM_R_X7Y143_SLICE_X8Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa30003000)
  ) CLBLM_R_X7Y143_SLICE_X8Y143_ALUT (
.I0(CLBLM_L_X8Y147_SLICE_X10Y147_DQ),
.I1(CLBLM_R_X5Y148_SLICE_X7Y148_CQ),
.I2(CLBLM_R_X7Y143_SLICE_X8Y143_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X7Y143_SLICE_X8Y143_AO5),
.O6(CLBLM_R_X7Y143_SLICE_X8Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y143_SLICE_X9Y143_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y143_SLICE_X9Y143_AO6),
.Q(CLBLM_R_X7Y143_SLICE_X9Y143_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y143_SLICE_X9Y143_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y143_SLICE_X9Y143_BO6),
.Q(CLBLM_R_X7Y143_SLICE_X9Y143_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y143_SLICE_X9Y143_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y143_SLICE_X9Y143_CO6),
.Q(CLBLM_R_X7Y143_SLICE_X9Y143_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffefffefffefffe)
  ) CLBLM_R_X7Y143_SLICE_X9Y143_DLUT (
.I0(CLBLM_L_X8Y143_SLICE_X11Y143_AQ),
.I1(CLBLM_R_X5Y143_SLICE_X7Y143_AQ),
.I2(CLBLM_R_X7Y143_SLICE_X9Y143_BQ),
.I3(CLBLM_R_X7Y143_SLICE_X9Y143_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y143_SLICE_X9Y143_DO5),
.O6(CLBLM_R_X7Y143_SLICE_X9Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaaee00550044)
  ) CLBLM_R_X7Y143_SLICE_X9Y143_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y143_SLICE_X9Y143_CQ),
.I2(1'b1),
.I3(CLBLM_R_X5Y143_SLICE_X7Y143_CO6),
.I4(CLBLM_R_X7Y143_SLICE_X9Y143_AQ),
.I5(CLBLM_R_X7Y143_SLICE_X8Y143_BQ),
.O5(CLBLM_R_X7Y143_SLICE_X9Y143_CO5),
.O6(CLBLM_R_X7Y143_SLICE_X9Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0f0faaaa0c0c)
  ) CLBLM_R_X7Y143_SLICE_X9Y143_BLUT (
.I0(CLBLM_R_X3Y149_SLICE_X3Y149_B5Q),
.I1(CLBLM_R_X7Y143_SLICE_X9Y143_BQ),
.I2(CLBLM_R_X5Y143_SLICE_X7Y143_CO6),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y143_SLICE_X10Y143_BQ),
.O5(CLBLM_R_X7Y143_SLICE_X9Y143_BO5),
.O6(CLBLM_R_X7Y143_SLICE_X9Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000fffc00fc)
  ) CLBLM_R_X7Y143_SLICE_X9Y143_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y143_SLICE_X9Y143_BQ),
.I2(CLBLM_R_X7Y143_SLICE_X9Y143_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y144_SLICE_X9Y144_AQ),
.I5(CLBLM_R_X5Y143_SLICE_X7Y143_CO6),
.O5(CLBLM_R_X7Y143_SLICE_X9Y143_AO5),
.O6(CLBLM_R_X7Y143_SLICE_X9Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y144_SLICE_X8Y144_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y144_SLICE_X8Y144_AO6),
.Q(CLBLM_R_X7Y144_SLICE_X8Y144_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y144_SLICE_X8Y144_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y144_SLICE_X8Y144_BO6),
.Q(CLBLM_R_X7Y144_SLICE_X8Y144_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y144_SLICE_X8Y144_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y144_SLICE_X8Y144_CO6),
.Q(CLBLM_R_X7Y144_SLICE_X8Y144_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y144_SLICE_X8Y144_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y144_SLICE_X8Y144_DO6),
.Q(CLBLM_R_X7Y144_SLICE_X8Y144_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000fa00fa00)
  ) CLBLM_R_X7Y144_SLICE_X8Y144_DLUT (
.I0(CLBLM_R_X11Y144_SLICE_X15Y144_DO6),
.I1(1'b1),
.I2(CLBLM_R_X7Y144_SLICE_X8Y144_DQ),
.I3(CLBLM_R_X7Y142_SLICE_X8Y142_DO6),
.I4(CLBLM_R_X3Y145_SLICE_X2Y145_A5Q),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X7Y144_SLICE_X8Y144_DO5),
.O6(CLBLM_R_X7Y144_SLICE_X8Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f0aaf000f088)
  ) CLBLM_R_X7Y144_SLICE_X8Y144_CLUT (
.I0(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.I1(CLBLM_R_X7Y144_SLICE_X8Y144_CQ),
.I2(CLBLM_R_X3Y145_SLICE_X3Y145_A5Q),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLM_L_X10Y144_SLICE_X13Y144_BQ),
.O5(CLBLM_R_X7Y144_SLICE_X8Y144_CO5),
.O6(CLBLM_R_X7Y144_SLICE_X8Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffeeffeaaaeeaaea)
  ) CLBLM_R_X7Y144_SLICE_X8Y144_BLUT (
.I0(CLBLM_R_X5Y144_SLICE_X7Y144_DO6),
.I1(CLBLM_R_X7Y144_SLICE_X8Y144_BQ),
.I2(RIOB33_X105Y117_IOB_X1Y118_I),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.I5(CLBLL_L_X4Y148_SLICE_X4Y148_CQ),
.O5(CLBLM_R_X7Y144_SLICE_X8Y144_BO5),
.O6(CLBLM_R_X7Y144_SLICE_X8Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heefaeefaeefaeeaa)
  ) CLBLM_R_X7Y144_SLICE_X8Y144_ALUT (
.I0(CLBLM_R_X5Y144_SLICE_X7Y144_DO6),
.I1(CLBLM_R_X3Y144_SLICE_X2Y144_BQ),
.I2(CLBLM_R_X7Y144_SLICE_X8Y144_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_R_X7Y144_SLICE_X8Y144_AO5),
.O6(CLBLM_R_X7Y144_SLICE_X8Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y144_SLICE_X9Y144_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y148_SLICE_X10Y148_BO6),
.Q(CLBLM_R_X7Y144_SLICE_X9Y144_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y144_SLICE_X9Y144_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y144_SLICE_X9Y144_AO6),
.Q(CLBLM_R_X7Y144_SLICE_X9Y144_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y144_SLICE_X9Y144_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y144_SLICE_X9Y144_BO6),
.Q(CLBLM_R_X7Y144_SLICE_X9Y144_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y144_SLICE_X9Y144_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y144_SLICE_X9Y144_CO6),
.Q(CLBLM_R_X7Y144_SLICE_X9Y144_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00002020ff00ffff)
  ) CLBLM_R_X7Y144_SLICE_X9Y144_DLUT (
.I0(CLBLL_L_X2Y146_SLICE_X1Y146_AQ),
.I1(CLBLM_L_X8Y144_SLICE_X11Y144_BO6),
.I2(CLBLL_L_X4Y143_SLICE_X4Y143_CO6),
.I3(CLBLM_L_X10Y144_SLICE_X12Y144_DO6),
.I4(CLBLM_R_X7Y142_SLICE_X8Y142_DO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y144_SLICE_X9Y144_DO5),
.O6(CLBLM_R_X7Y144_SLICE_X9Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f0ccf000f0cc)
  ) CLBLM_R_X7Y144_SLICE_X9Y144_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y144_SLICE_X9Y144_CQ),
.I2(CLBLM_R_X5Y144_SLICE_X7Y144_B5Q),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y144_SLICE_X9Y144_CO5),
.O6(CLBLM_R_X7Y144_SLICE_X9Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0050504040)
  ) CLBLM_R_X7Y144_SLICE_X9Y144_BLUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_R_X7Y144_SLICE_X9Y144_BQ),
.I2(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.I3(CLBLM_L_X8Y150_SLICE_X10Y150_AQ),
.I4(CLBLM_L_X10Y144_SLICE_X12Y144_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X7Y144_SLICE_X9Y144_BO5),
.O6(CLBLM_R_X7Y144_SLICE_X9Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccfe0032cccc0000)
  ) CLBLM_R_X7Y144_SLICE_X9Y144_ALUT (
.I0(CLBLM_R_X7Y144_SLICE_X9Y144_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_R_X3Y150_SLICE_X3Y150_AQ),
.I5(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.O5(CLBLM_R_X7Y144_SLICE_X9Y144_AO5),
.O6(CLBLM_R_X7Y144_SLICE_X9Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y145_SLICE_X8Y145_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y145_SLICE_X8Y145_CO5),
.Q(CLBLM_R_X7Y145_SLICE_X8Y145_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y145_SLICE_X8Y145_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y145_SLICE_X8Y145_AO6),
.Q(CLBLM_R_X7Y145_SLICE_X8Y145_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y145_SLICE_X8Y145_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y145_SLICE_X8Y145_BO6),
.Q(CLBLM_R_X7Y145_SLICE_X8Y145_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y145_SLICE_X8Y145_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y145_SLICE_X8Y145_CO6),
.Q(CLBLM_R_X7Y145_SLICE_X8Y145_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000033336333)
  ) CLBLM_R_X7Y145_SLICE_X8Y145_DLUT (
.I0(CLBLM_R_X7Y143_SLICE_X8Y143_AQ),
.I1(CLBLM_R_X11Y148_SLICE_X14Y148_CQ),
.I2(CLBLL_L_X4Y143_SLICE_X4Y143_BQ),
.I3(CLBLM_R_X5Y145_SLICE_X6Y145_CQ),
.I4(CLBLM_R_X7Y145_SLICE_X8Y145_BQ),
.I5(CLBLL_L_X4Y145_SLICE_X4Y145_BQ),
.O5(CLBLM_R_X7Y145_SLICE_X8Y145_DO5),
.O6(CLBLM_R_X7Y145_SLICE_X8Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc00f0f0f0aaaa)
  ) CLBLM_R_X7Y145_SLICE_X8Y145_CLUT (
.I0(CLBLM_R_X3Y145_SLICE_X2Y145_A5Q),
.I1(CLBLM_R_X5Y147_SLICE_X6Y147_CQ),
.I2(CLBLM_R_X7Y148_SLICE_X9Y148_CQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y145_SLICE_X8Y145_CO5),
.O6(CLBLM_R_X7Y145_SLICE_X8Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf202f202f000f000)
  ) CLBLM_R_X7Y145_SLICE_X8Y145_BLUT (
.I0(CLBLM_R_X7Y145_SLICE_X8Y145_BQ),
.I1(CLBLM_R_X5Y148_SLICE_X7Y148_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y147_SLICE_X8Y147_BQ),
.I4(1'b1),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X7Y145_SLICE_X8Y145_BO5),
.O6(CLBLM_R_X7Y145_SLICE_X8Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc005a005a)
  ) CLBLM_R_X7Y145_SLICE_X8Y145_ALUT (
.I0(CLBLM_R_X5Y145_SLICE_X7Y145_DO6),
.I1(CLBLM_L_X12Y145_SLICE_X16Y145_BQ),
.I2(CLBLM_R_X7Y145_SLICE_X8Y145_AQ),
.I3(CLBLM_R_X11Y146_SLICE_X14Y146_AQ),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X7Y145_SLICE_X8Y145_AO5),
.O6(CLBLM_R_X7Y145_SLICE_X8Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y145_SLICE_X9Y145_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y145_SLICE_X9Y145_CO5),
.Q(CLBLM_R_X7Y145_SLICE_X9Y145_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y145_SLICE_X9Y145_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y145_SLICE_X9Y145_AO6),
.Q(CLBLM_R_X7Y145_SLICE_X9Y145_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y145_SLICE_X9Y145_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y145_SLICE_X9Y145_BO6),
.Q(CLBLM_R_X7Y145_SLICE_X9Y145_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y145_SLICE_X9Y145_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y145_SLICE_X9Y145_CO6),
.Q(CLBLM_R_X7Y145_SLICE_X9Y145_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffdfdf)
  ) CLBLM_R_X7Y145_SLICE_X9Y145_DLUT (
.I0(CLBLM_R_X7Y153_SLICE_X9Y153_CO5),
.I1(CLBLL_L_X2Y151_SLICE_X1Y151_BO6),
.I2(CLBLL_L_X4Y154_SLICE_X4Y154_CO6),
.I3(1'b1),
.I4(CLBLM_R_X5Y149_SLICE_X6Y149_CO6),
.I5(CLBLM_R_X5Y145_SLICE_X6Y145_DO6),
.O5(CLBLM_R_X7Y145_SLICE_X9Y145_DO5),
.O6(CLBLM_R_X7Y145_SLICE_X9Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5a0a0ea40ea40)
  ) CLBLM_R_X7Y145_SLICE_X9Y145_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X7Y147_SLICE_X8Y147_DQ),
.I3(CLBLM_L_X12Y149_SLICE_X16Y149_AQ),
.I4(CLBLM_L_X8Y145_SLICE_X10Y145_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X7Y145_SLICE_X9Y145_CO5),
.O6(CLBLM_R_X7Y145_SLICE_X9Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffac80000fac8)
  ) CLBLM_R_X7Y145_SLICE_X9Y145_BLUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_R_X7Y145_SLICE_X9Y145_BQ),
.I2(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.I3(CLBLM_R_X7Y144_SLICE_X9Y144_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X3Y144_SLICE_X2Y144_AQ),
.O5(CLBLM_R_X7Y145_SLICE_X9Y145_BO5),
.O6(CLBLM_R_X7Y145_SLICE_X9Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffc8ffc800c800c8)
  ) CLBLM_R_X7Y145_SLICE_X9Y145_ALUT (
.I0(CLBLM_R_X7Y148_SLICE_X9Y148_CQ),
.I1(CLBLM_L_X8Y152_SLICE_X11Y152_BO6),
.I2(CLBLM_R_X7Y145_SLICE_X9Y145_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLM_L_X8Y145_SLICE_X11Y145_BQ),
.O5(CLBLM_R_X7Y145_SLICE_X9Y145_AO5),
.O6(CLBLM_R_X7Y145_SLICE_X9Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y146_SLICE_X8Y146_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y146_SLICE_X8Y146_CO5),
.Q(CLBLM_R_X7Y146_SLICE_X8Y146_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y146_SLICE_X8Y146_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y146_SLICE_X8Y146_AO6),
.Q(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y146_SLICE_X8Y146_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y146_SLICE_X8Y146_CO6),
.Q(CLBLM_R_X7Y146_SLICE_X8Y146_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y146_SLICE_X8Y146_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y146_SLICE_X8Y146_DO6),
.Q(CLBLM_R_X7Y146_SLICE_X8Y146_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa0000ff00)
  ) CLBLM_R_X7Y146_SLICE_X8Y146_DLUT (
.I0(CLBLM_L_X8Y145_SLICE_X11Y145_AQ),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X7Y152_SLICE_X9Y152_CQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X7Y146_SLICE_X8Y146_DO5),
.O6(CLBLM_R_X7Y146_SLICE_X8Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff330033f044f044)
  ) CLBLM_R_X7Y146_SLICE_X8Y146_CLUT (
.I0(CLBLM_R_X7Y146_SLICE_X8Y146_C5Q),
.I1(RIOB33_X105Y119_IOB_X1Y119_I),
.I2(CLBLM_L_X10Y146_SLICE_X13Y146_B5Q),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X5Y146_SLICE_X6Y146_DQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y146_SLICE_X8Y146_CO5),
.O6(CLBLM_R_X7Y146_SLICE_X8Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hbb88b888ff00f000)
  ) CLBLM_R_X7Y146_SLICE_X8Y146_BLUT (
.I0(CLBLM_R_X11Y146_SLICE_X15Y146_DQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X11Y148_SLICE_X15Y148_AQ),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(CLBLM_R_X7Y152_SLICE_X9Y152_CQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y146_SLICE_X8Y146_BO5),
.O6(CLBLM_R_X7Y146_SLICE_X8Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccce00000002)
  ) CLBLM_R_X7Y146_SLICE_X8Y146_ALUT (
.I0(RIOB33_X105Y119_IOB_X1Y119_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.I3(CLBLM_R_X7Y146_SLICE_X8Y146_CQ),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLL_L_X4Y149_SLICE_X5Y149_CQ),
.O5(CLBLM_R_X7Y146_SLICE_X8Y146_AO5),
.O6(CLBLM_R_X7Y146_SLICE_X8Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y146_SLICE_X9Y146_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y146_SLICE_X9Y146_AO6),
.Q(CLBLM_R_X7Y146_SLICE_X9Y146_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y146_SLICE_X9Y146_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y146_SLICE_X9Y146_BO6),
.Q(CLBLM_R_X7Y146_SLICE_X9Y146_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y146_SLICE_X9Y146_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y146_SLICE_X9Y146_CO6),
.Q(CLBLM_R_X7Y146_SLICE_X9Y146_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_R_X7Y146_SLICE_X9Y146_DLUT (
.I0(CLBLM_R_X7Y145_SLICE_X9Y145_C5Q),
.I1(CLBLM_R_X7Y152_SLICE_X9Y152_CQ),
.I2(CLBLM_R_X7Y147_SLICE_X8Y147_DQ),
.I3(CLBLM_R_X7Y149_SLICE_X8Y149_CQ),
.I4(CLBLM_R_X7Y146_SLICE_X8Y146_DQ),
.I5(CLBLL_L_X4Y146_SLICE_X5Y146_A5Q),
.O5(CLBLM_R_X7Y146_SLICE_X9Y146_DO5),
.O6(CLBLM_R_X7Y146_SLICE_X9Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa0000fcfc)
  ) CLBLM_R_X7Y146_SLICE_X9Y146_CLUT (
.I0(CLBLM_R_X5Y148_SLICE_X7Y148_AQ),
.I1(CLBLM_R_X7Y146_SLICE_X9Y146_CQ),
.I2(CLBLM_L_X10Y148_SLICE_X12Y148_BQ),
.I3(1'b1),
.I4(CLBLL_L_X4Y145_SLICE_X5Y145_DO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X7Y146_SLICE_X9Y146_CO5),
.O6(CLBLM_R_X7Y146_SLICE_X9Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0aaaaaacc)
  ) CLBLM_R_X7Y146_SLICE_X9Y146_BLUT (
.I0(CLBLL_L_X4Y146_SLICE_X4Y146_BQ),
.I1(CLBLM_R_X7Y146_SLICE_X9Y146_BQ),
.I2(CLBLM_R_X7Y147_SLICE_X9Y147_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X7Y146_SLICE_X9Y146_BO5),
.O6(CLBLM_R_X7Y146_SLICE_X9Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc00a5cccc00a5)
  ) CLBLM_R_X7Y146_SLICE_X9Y146_ALUT (
.I0(CLBLM_R_X5Y148_SLICE_X6Y148_AQ),
.I1(CLBLM_R_X7Y143_SLICE_X9Y143_AQ),
.I2(CLBLM_L_X8Y148_SLICE_X10Y148_CO5),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y146_SLICE_X9Y146_AO5),
.O6(CLBLM_R_X7Y146_SLICE_X9Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y147_SLICE_X8Y147_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y147_SLICE_X8Y147_BO5),
.Q(CLBLM_R_X7Y147_SLICE_X8Y147_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y147_SLICE_X8Y147_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y147_SLICE_X8Y147_CO5),
.Q(CLBLM_R_X7Y147_SLICE_X8Y147_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y147_SLICE_X8Y147_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y147_SLICE_X8Y147_AO6),
.Q(CLBLM_R_X7Y147_SLICE_X8Y147_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y147_SLICE_X8Y147_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y147_SLICE_X8Y147_BO6),
.Q(CLBLM_R_X7Y147_SLICE_X8Y147_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y147_SLICE_X8Y147_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y147_SLICE_X8Y147_CO6),
.Q(CLBLM_R_X7Y147_SLICE_X8Y147_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y147_SLICE_X8Y147_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y147_SLICE_X8Y147_DO6),
.Q(CLBLM_R_X7Y147_SLICE_X8Y147_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc55cc55cc00cc00)
  ) CLBLM_R_X7Y147_SLICE_X8Y147_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X5Y152_SLICE_X7Y152_CQ),
.I2(1'b1),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLM_L_X10Y146_SLICE_X13Y146_B5Q),
.O5(CLBLM_R_X7Y147_SLICE_X8Y147_DO5),
.O6(CLBLM_R_X7Y147_SLICE_X8Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf404f404cfcfc0c0)
  ) CLBLM_R_X7Y147_SLICE_X8Y147_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X7Y147_SLICE_X9Y147_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y153_SLICE_X8Y153_CQ),
.I4(CLBLM_R_X7Y147_SLICE_X8Y147_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X7Y147_SLICE_X8Y147_CO5),
.O6(CLBLM_R_X7Y147_SLICE_X8Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0c000caaffaa00)
  ) CLBLM_R_X7Y147_SLICE_X8Y147_BLUT (
.I0(CLBLM_R_X7Y147_SLICE_X8Y147_CQ),
.I1(CLBLM_R_X7Y153_SLICE_X8Y153_DQ),
.I2(CLBLM_R_X11Y153_SLICE_X14Y153_AO6),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X5Y147_SLICE_X7Y147_DQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y147_SLICE_X8Y147_BO5),
.O6(CLBLM_R_X7Y147_SLICE_X8Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffccffccf0cc5a)
  ) CLBLM_R_X7Y147_SLICE_X8Y147_ALUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_L_X8Y150_SLICE_X10Y150_CQ),
.I2(CLBLM_R_X7Y147_SLICE_X8Y147_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.I5(CLBLM_R_X11Y146_SLICE_X14Y146_AQ),
.O5(CLBLM_R_X7Y147_SLICE_X8Y147_AO5),
.O6(CLBLM_R_X7Y147_SLICE_X8Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y147_SLICE_X9Y147_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y147_SLICE_X9Y147_AO6),
.Q(CLBLM_R_X7Y147_SLICE_X9Y147_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y147_SLICE_X9Y147_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y147_SLICE_X9Y147_BO6),
.Q(CLBLM_R_X7Y147_SLICE_X9Y147_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffefffffffe)
  ) CLBLM_R_X7Y147_SLICE_X9Y147_DLUT (
.I0(CLBLM_R_X5Y148_SLICE_X7Y148_C5Q),
.I1(CLBLM_L_X10Y146_SLICE_X13Y146_B5Q),
.I2(CLBLM_R_X7Y147_SLICE_X9Y147_BQ),
.I3(CLBLM_R_X5Y148_SLICE_X7Y148_BQ),
.I4(CLBLM_L_X10Y146_SLICE_X13Y146_DO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y147_SLICE_X9Y147_DO5),
.O6(CLBLM_R_X7Y147_SLICE_X9Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hee00ee00ff00f000)
  ) CLBLM_R_X7Y147_SLICE_X9Y147_CLUT (
.I0(CLBLM_R_X7Y145_SLICE_X9Y145_C5Q),
.I1(CLBLL_L_X4Y147_SLICE_X4Y147_AQ),
.I2(CLBLM_R_X7Y149_SLICE_X8Y149_CQ),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(CLBLM_L_X8Y150_SLICE_X10Y150_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y147_SLICE_X9Y147_CO5),
.O6(CLBLM_R_X7Y147_SLICE_X9Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0f3c0c0c0f3c0c0)
  ) CLBLM_R_X7Y147_SLICE_X9Y147_BLUT (
.I0(1'b1),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y151_SLICE_X12Y151_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X7Y145_SLICE_X9Y145_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X7Y147_SLICE_X9Y147_BO5),
.O6(CLBLM_R_X7Y147_SLICE_X9Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0f3c0c0c0f3c0)
  ) CLBLM_R_X7Y147_SLICE_X9Y147_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X8Y146_SLICE_X10Y146_AQ),
.I3(CLBLM_R_X7Y147_SLICE_X8Y147_BQ),
.I4(CLBLM_R_X11Y153_SLICE_X14Y153_AO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y147_SLICE_X9Y147_AO5),
.O6(CLBLM_R_X7Y147_SLICE_X9Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y148_SLICE_X8Y148_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y148_SLICE_X8Y148_DO5),
.Q(CLBLM_R_X7Y148_SLICE_X8Y148_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y148_SLICE_X8Y148_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y148_SLICE_X8Y148_AO6),
.Q(CLBLM_R_X7Y148_SLICE_X8Y148_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y148_SLICE_X8Y148_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y148_SLICE_X8Y148_CO6),
.Q(CLBLM_R_X7Y148_SLICE_X8Y148_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y148_SLICE_X8Y148_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y148_SLICE_X8Y148_DO6),
.Q(CLBLM_R_X7Y148_SLICE_X8Y148_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5a0a0dddd8888)
  ) CLBLM_R_X7Y148_SLICE_X8Y148_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y154_SLICE_X12Y154_DQ),
.I2(CLBLL_L_X2Y146_SLICE_X1Y146_AQ),
.I3(1'b1),
.I4(RIOB33_X105Y143_IOB_X1Y144_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y148_SLICE_X8Y148_DO5),
.O6(CLBLM_R_X7Y148_SLICE_X8Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f0f3f003000300)
  ) CLBLM_R_X7Y148_SLICE_X8Y148_CLUT (
.I0(1'b1),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y150_SLICE_X8Y150_CQ),
.I4(1'b1),
.I5(CLBLM_R_X5Y147_SLICE_X7Y147_BQ),
.O5(CLBLM_R_X7Y148_SLICE_X8Y148_CO5),
.O6(CLBLM_R_X7Y148_SLICE_X8Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00c8c8c8c8c8c8)
  ) CLBLM_R_X7Y148_SLICE_X8Y148_BLUT (
.I0(CLBLM_R_X7Y148_SLICE_X9Y148_DQ),
.I1(RIOB33_X105Y121_IOB_X1Y121_I),
.I2(CLBLM_R_X7Y147_SLICE_X8Y147_CQ),
.I3(CLBLM_R_X5Y146_SLICE_X6Y146_A5Q),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y148_SLICE_X8Y148_BO5),
.O6(CLBLM_R_X7Y148_SLICE_X8Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff3333ffef3323)
  ) CLBLM_R_X7Y148_SLICE_X8Y148_ALUT (
.I0(CLBLM_R_X5Y154_SLICE_X6Y154_BO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(RIOB33_X105Y135_IOB_X1Y136_I),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(CLBLM_R_X7Y148_SLICE_X9Y148_AQ),
.I5(RIOB33_X105Y135_IOB_X1Y135_I),
.O5(CLBLM_R_X7Y148_SLICE_X8Y148_AO5),
.O6(CLBLM_R_X7Y148_SLICE_X8Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y148_SLICE_X9Y148_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y148_SLICE_X9Y148_AO6),
.Q(CLBLM_R_X7Y148_SLICE_X9Y148_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y148_SLICE_X9Y148_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y148_SLICE_X9Y148_BO6),
.Q(CLBLM_R_X7Y148_SLICE_X9Y148_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y148_SLICE_X9Y148_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y148_SLICE_X9Y148_CO6),
.Q(CLBLM_R_X7Y148_SLICE_X9Y148_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y148_SLICE_X9Y148_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y148_SLICE_X9Y148_DO6),
.Q(CLBLM_R_X7Y148_SLICE_X9Y148_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hddddd8d8dd88d888)
  ) CLBLM_R_X7Y148_SLICE_X9Y148_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y145_SLICE_X8Y145_AQ),
.I2(CLBLM_R_X7Y148_SLICE_X9Y148_DQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_L_X8Y146_SLICE_X10Y146_DO6),
.I5(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.O5(CLBLM_R_X7Y148_SLICE_X9Y148_DO5),
.O6(CLBLM_R_X7Y148_SLICE_X9Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0b1e4a0a0b1e4)
  ) CLBLM_R_X7Y148_SLICE_X9Y148_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y148_SLICE_X12Y148_AO5),
.I2(CLBLM_R_X7Y148_SLICE_X9Y148_BQ),
.I3(CLBLM_R_X5Y146_SLICE_X6Y146_CQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y148_SLICE_X9Y148_CO5),
.O6(CLBLM_R_X7Y148_SLICE_X9Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hddddd8d8ddddd8d8)
  ) CLBLM_R_X7Y148_SLICE_X9Y148_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLL_L_X4Y150_SLICE_X4Y150_B5Q),
.I2(CLBLM_R_X11Y153_SLICE_X14Y153_AO6),
.I3(1'b1),
.I4(CLBLM_R_X7Y147_SLICE_X9Y147_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y148_SLICE_X9Y148_BO5),
.O6(CLBLM_R_X7Y148_SLICE_X9Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafa5050aaaa0000)
  ) CLBLM_R_X7Y148_SLICE_X9Y148_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(1'b1),
.I2(CLBLM_R_X7Y148_SLICE_X9Y148_AQ),
.I3(1'b1),
.I4(CLBLM_R_X7Y148_SLICE_X9Y148_DQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X7Y148_SLICE_X9Y148_AO5),
.O6(CLBLM_R_X7Y148_SLICE_X9Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y149_SLICE_X8Y149_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y149_SLICE_X8Y149_AO6),
.Q(CLBLM_R_X7Y149_SLICE_X8Y149_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y149_SLICE_X8Y149_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y149_SLICE_X8Y149_BO6),
.Q(CLBLM_R_X7Y149_SLICE_X8Y149_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y149_SLICE_X8Y149_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y149_SLICE_X8Y149_CO6),
.Q(CLBLM_R_X7Y149_SLICE_X8Y149_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y149_SLICE_X8Y149_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y149_SLICE_X8Y149_DO6),
.Q(CLBLM_R_X7Y149_SLICE_X8Y149_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff228800002288)
  ) CLBLM_R_X7Y149_SLICE_X8Y149_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X7Y150_SLICE_X8Y150_DO6),
.I2(1'b1),
.I3(CLBLM_L_X8Y146_SLICE_X11Y146_CO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X5Y148_SLICE_X7Y148_BQ),
.O5(CLBLM_R_X7Y149_SLICE_X8Y149_DO5),
.O6(CLBLM_R_X7Y149_SLICE_X8Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5a0a0a0f5a0a0a0)
  ) CLBLM_R_X7Y149_SLICE_X8Y149_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(1'b1),
.I2(CLBLM_R_X3Y149_SLICE_X2Y149_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_L_X10Y148_SLICE_X13Y148_BQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y149_SLICE_X8Y149_CO5),
.O6(CLBLM_R_X7Y149_SLICE_X8Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff001111ff002222)
  ) CLBLM_R_X7Y149_SLICE_X8Y149_BLUT (
.I0(CLBLM_R_X7Y148_SLICE_X8Y148_BO5),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(1'b1),
.I3(CLBLL_L_X4Y149_SLICE_X4Y149_DQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X10Y150_SLICE_X12Y150_CQ),
.O5(CLBLM_R_X7Y149_SLICE_X8Y149_BO5),
.O6(CLBLM_R_X7Y149_SLICE_X8Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h888888888dd88dd8)
  ) CLBLM_R_X7Y149_SLICE_X8Y149_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y149_SLICE_X13Y149_BQ),
.I2(CLBLM_R_X7Y149_SLICE_X8Y149_DQ),
.I3(CLBLM_L_X8Y148_SLICE_X11Y148_CO6),
.I4(1'b1),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X7Y149_SLICE_X8Y149_AO5),
.O6(CLBLM_R_X7Y149_SLICE_X8Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y149_SLICE_X9Y149_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y149_SLICE_X9Y149_AO6),
.Q(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc04cc04c000c000)
  ) CLBLM_R_X7Y149_SLICE_X9Y149_DLUT (
.I0(CLBLM_R_X7Y153_SLICE_X9Y153_CO5),
.I1(CLBLM_L_X10Y149_SLICE_X12Y149_AO5),
.I2(CLBLM_R_X5Y144_SLICE_X7Y144_AQ),
.I3(CLBLM_R_X7Y147_SLICE_X9Y147_CO5),
.I4(1'b1),
.I5(CLBLM_L_X10Y144_SLICE_X13Y144_AQ),
.O5(CLBLM_R_X7Y149_SLICE_X9Y149_DO5),
.O6(CLBLM_R_X7Y149_SLICE_X9Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff3fffff0f0f0f0)
  ) CLBLM_R_X7Y149_SLICE_X9Y149_CLUT (
.I0(1'b1),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X5Y144_SLICE_X7Y144_AQ),
.I3(CLBLL_L_X2Y151_SLICE_X1Y151_BO6),
.I4(CLBLL_L_X4Y146_SLICE_X4Y146_CO5),
.I5(CLBLM_L_X10Y144_SLICE_X13Y144_AQ),
.O5(CLBLM_R_X7Y149_SLICE_X9Y149_CO5),
.O6(CLBLM_R_X7Y149_SLICE_X9Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfeffcccc00000500)
  ) CLBLM_R_X7Y149_SLICE_X9Y149_BLUT (
.I0(CLBLM_L_X8Y149_SLICE_X10Y149_AO5),
.I1(CLBLL_L_X4Y146_SLICE_X5Y146_A5Q),
.I2(CLBLM_R_X7Y143_SLICE_X8Y143_AQ),
.I3(CLBLM_R_X7Y145_SLICE_X8Y145_BQ),
.I4(CLBLM_R_X7Y152_SLICE_X9Y152_BQ),
.I5(RIOB33_X105Y121_IOB_X1Y121_I),
.O5(CLBLM_R_X7Y149_SLICE_X9Y149_BO5),
.O6(CLBLM_R_X7Y149_SLICE_X9Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaffccaaaaf0c0)
  ) CLBLM_R_X7Y149_SLICE_X9Y149_ALUT (
.I0(CLBLM_R_X3Y143_SLICE_X3Y143_B5Q),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_R_X7Y150_SLICE_X9Y150_DO6),
.I3(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.O5(CLBLM_R_X7Y149_SLICE_X9Y149_AO5),
.O6(CLBLM_R_X7Y149_SLICE_X9Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y150_SLICE_X8Y150_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y150_SLICE_X8Y150_AO6),
.Q(CLBLM_R_X7Y150_SLICE_X8Y150_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y150_SLICE_X8Y150_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y150_SLICE_X8Y150_BO6),
.Q(CLBLM_R_X7Y150_SLICE_X8Y150_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y150_SLICE_X8Y150_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y150_SLICE_X8Y150_CO6),
.Q(CLBLM_R_X7Y150_SLICE_X8Y150_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6666999999996666)
  ) CLBLM_R_X7Y150_SLICE_X8Y150_DLUT (
.I0(CLBLM_L_X8Y154_SLICE_X10Y154_AQ),
.I1(CLBLM_R_X7Y153_SLICE_X9Y153_A5Q),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X7Y149_SLICE_X8Y149_DQ),
.I5(CLBLM_R_X5Y150_SLICE_X7Y150_BQ),
.O5(CLBLM_R_X7Y150_SLICE_X8Y150_DO5),
.O6(CLBLM_R_X7Y150_SLICE_X8Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0b1e4a0a0a0b1e4)
  ) CLBLM_R_X7Y150_SLICE_X8Y150_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y150_SLICE_X8Y150_CQ),
.I2(CLBLM_R_X7Y148_SLICE_X8Y148_DQ),
.I3(CLBLM_R_X7Y148_SLICE_X9Y148_CQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X7Y150_SLICE_X9Y150_CO5),
.O5(CLBLM_R_X7Y150_SLICE_X8Y150_CO5),
.O6(CLBLM_R_X7Y150_SLICE_X8Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0ccf0ccf0aaf0aa)
  ) CLBLM_R_X7Y150_SLICE_X8Y150_BLUT (
.I0(CLBLM_L_X8Y150_SLICE_X10Y150_CQ),
.I1(CLBLM_R_X7Y150_SLICE_X8Y150_BQ),
.I2(CLBLM_R_X7Y149_SLICE_X8Y149_CQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLM_L_X8Y152_SLICE_X11Y152_BO6),
.O5(CLBLM_R_X7Y150_SLICE_X8Y150_BO5),
.O6(CLBLM_R_X7Y150_SLICE_X8Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hb8bbbbbbb8888888)
  ) CLBLM_R_X7Y150_SLICE_X8Y150_ALUT (
.I0(CLBLM_L_X8Y151_SLICE_X11Y151_DQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X7Y150_SLICE_X8Y150_AQ),
.I3(CLBLL_L_X4Y151_SLICE_X4Y151_AQ),
.I4(CLBLM_L_X8Y149_SLICE_X11Y149_AQ),
.I5(CLBLM_R_X7Y145_SLICE_X8Y145_AQ),
.O5(CLBLM_R_X7Y150_SLICE_X8Y150_AO5),
.O6(CLBLM_R_X7Y150_SLICE_X8Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y150_SLICE_X9Y150_A5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y150_SLICE_X9Y150_BO6),
.Q(CLBLM_R_X7Y150_SLICE_X9Y150_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y150_SLICE_X9Y150_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y150_SLICE_X9Y150_AO6),
.Q(CLBLM_R_X7Y150_SLICE_X9Y150_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaa0a8b1aaa0aaa0)
  ) CLBLM_R_X7Y150_SLICE_X9Y150_DLUT (
.I0(RIOB33_X105Y121_IOB_X1Y121_I),
.I1(CLBLM_L_X8Y149_SLICE_X10Y149_AO5),
.I2(CLBLM_L_X10Y146_SLICE_X12Y146_DQ),
.I3(CLBLM_R_X5Y149_SLICE_X7Y149_CQ),
.I4(CLBLM_R_X7Y145_SLICE_X8Y145_BQ),
.I5(CLBLM_R_X7Y143_SLICE_X8Y143_AQ),
.O5(CLBLM_R_X7Y150_SLICE_X9Y150_DO5),
.O6(CLBLM_R_X7Y150_SLICE_X9Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000020033cc33cc)
  ) CLBLM_R_X7Y150_SLICE_X9Y150_CLUT (
.I0(CLBLM_R_X7Y148_SLICE_X8Y148_CQ),
.I1(CLBLM_R_X5Y146_SLICE_X6Y146_CQ),
.I2(CLBLM_L_X8Y146_SLICE_X10Y146_AQ),
.I3(CLBLM_R_X7Y150_SLICE_X9Y150_A5Q),
.I4(CLBLM_R_X7Y150_SLICE_X9Y150_BO5),
.I5(1'b1),
.O5(CLBLM_R_X7Y150_SLICE_X9Y150_CO5),
.O6(CLBLM_R_X7Y150_SLICE_X9Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000fc0cfffff7f7)
  ) CLBLM_R_X7Y150_SLICE_X9Y150_BLUT (
.I0(CLBLM_L_X8Y150_SLICE_X10Y150_CQ),
.I1(CLBLM_R_X7Y145_SLICE_X8Y145_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X11Y153_SLICE_X14Y153_BQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y150_SLICE_X9Y150_BO5),
.O6(CLBLM_R_X7Y150_SLICE_X9Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff33b3b3ff00a0a0)
  ) CLBLM_R_X7Y150_SLICE_X9Y150_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X8Y150_SLICE_X11Y150_CO6),
.I2(CLBLM_R_X7Y150_SLICE_X9Y150_AQ),
.I3(CLBLM_L_X8Y143_SLICE_X10Y143_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y150_SLICE_X9Y150_CO6),
.O5(CLBLM_R_X7Y150_SLICE_X9Y150_AO5),
.O6(CLBLM_R_X7Y150_SLICE_X9Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y151_SLICE_X8Y151_A5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y151_SLICE_X8Y151_CO6),
.Q(CLBLM_R_X7Y151_SLICE_X8Y151_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y151_SLICE_X8Y151_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y151_SLICE_X8Y151_AO6),
.Q(CLBLM_R_X7Y151_SLICE_X8Y151_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y151_SLICE_X8Y151_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y151_SLICE_X8Y151_BO6),
.Q(CLBLM_R_X7Y151_SLICE_X8Y151_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffeeffff33330000)
  ) CLBLM_R_X7Y151_SLICE_X8Y151_DLUT (
.I0(CLBLM_L_X10Y149_SLICE_X13Y149_BQ),
.I1(RIOB33_X105Y121_IOB_X1Y121_I),
.I2(1'b1),
.I3(CLBLM_R_X5Y152_SLICE_X6Y152_CQ),
.I4(CLBLM_R_X11Y146_SLICE_X14Y146_DQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y151_SLICE_X8Y151_DO5),
.O6(CLBLM_R_X7Y151_SLICE_X8Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbaa3300f0f00000)
  ) CLBLM_R_X7Y151_SLICE_X8Y151_CLUT (
.I0(CLBLM_R_X7Y151_SLICE_X8Y151_BQ),
.I1(CLBLL_L_X4Y145_SLICE_X5Y145_CO6),
.I2(CLBLM_L_X10Y153_SLICE_X12Y153_CQ),
.I3(CLBLM_R_X7Y151_SLICE_X8Y151_A5Q),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y151_SLICE_X8Y151_CO5),
.O6(CLBLM_R_X7Y151_SLICE_X8Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa00f0aaaa00c0)
  ) CLBLM_R_X7Y151_SLICE_X8Y151_BLUT (
.I0(CLBLM_R_X3Y149_SLICE_X3Y149_AQ),
.I1(CLBLM_R_X7Y151_SLICE_X8Y151_BQ),
.I2(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y143_SLICE_X8Y143_CQ),
.O5(CLBLM_R_X7Y151_SLICE_X8Y151_BO5),
.O6(CLBLM_R_X7Y151_SLICE_X8Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc5550cccc5550)
  ) CLBLM_R_X7Y151_SLICE_X8Y151_ALUT (
.I0(CLBLM_R_X5Y152_SLICE_X7Y152_DO5),
.I1(CLBLM_L_X10Y149_SLICE_X12Y149_AQ),
.I2(CLBLM_R_X7Y151_SLICE_X8Y151_AQ),
.I3(CLBLM_R_X5Y149_SLICE_X7Y149_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y151_SLICE_X8Y151_AO5),
.O6(CLBLM_R_X7Y151_SLICE_X8Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y151_SLICE_X9Y151_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y151_SLICE_X9Y151_AO6),
.Q(CLBLM_R_X7Y151_SLICE_X9Y151_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y151_SLICE_X9Y151_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y151_SLICE_X9Y151_BO6),
.Q(CLBLM_R_X7Y151_SLICE_X9Y151_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y151_SLICE_X9Y151_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y151_SLICE_X9Y151_CO6),
.Q(CLBLM_R_X7Y151_SLICE_X9Y151_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff00f0011551155)
  ) CLBLM_R_X7Y151_SLICE_X9Y151_DLUT (
.I0(CLBLM_L_X8Y146_SLICE_X10Y146_BQ),
.I1(CLBLM_R_X3Y147_SLICE_X3Y147_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLL_L_X2Y151_SLICE_X1Y151_BO6),
.I4(CLBLM_L_X8Y151_SLICE_X11Y151_CQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y151_SLICE_X9Y151_DO5),
.O6(CLBLM_R_X7Y151_SLICE_X9Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccfccfc00030030)
  ) CLBLM_R_X7Y151_SLICE_X9Y151_CLUT (
.I0(1'b1),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X7Y153_SLICE_X9Y153_DQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X7Y150_SLICE_X9Y150_DO6),
.I5(CLBLM_L_X8Y151_SLICE_X10Y151_AQ),
.O5(CLBLM_R_X7Y151_SLICE_X9Y151_CO5),
.O6(CLBLM_R_X7Y151_SLICE_X9Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0afafafa0acacac)
  ) CLBLM_R_X7Y151_SLICE_X9Y151_BLUT (
.I0(CLBLM_L_X10Y152_SLICE_X13Y152_BQ),
.I1(CLBLM_R_X7Y151_SLICE_X9Y151_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLL_L_X4Y151_SLICE_X4Y151_AQ),
.I4(CLBLM_L_X8Y149_SLICE_X11Y149_AQ),
.I5(CLBLM_R_X3Y147_SLICE_X3Y147_BQ),
.O5(CLBLM_R_X7Y151_SLICE_X9Y151_BO5),
.O6(CLBLM_R_X7Y151_SLICE_X9Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff007070f8f8)
  ) CLBLM_R_X7Y151_SLICE_X9Y151_ALUT (
.I0(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_R_X7Y151_SLICE_X9Y151_AQ),
.I3(CLBLL_L_X4Y151_SLICE_X4Y151_AQ),
.I4(CLBLM_R_X7Y153_SLICE_X9Y153_CO5),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X7Y151_SLICE_X9Y151_AO5),
.O6(CLBLM_R_X7Y151_SLICE_X9Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y152_SLICE_X8Y152_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y152_SLICE_X8Y152_AO6),
.Q(CLBLM_R_X7Y152_SLICE_X8Y152_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y152_SLICE_X8Y152_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y152_SLICE_X8Y152_BO6),
.Q(CLBLM_R_X7Y152_SLICE_X8Y152_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y152_SLICE_X8Y152_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y152_SLICE_X8Y152_CO6),
.Q(CLBLM_R_X7Y152_SLICE_X8Y152_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y152_SLICE_X8Y152_D_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y152_SLICE_X8Y152_DO6),
.Q(CLBLM_R_X7Y152_SLICE_X8Y152_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hee44ee44fa50fa50)
  ) CLBLM_R_X7Y152_SLICE_X8Y152_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y153_SLICE_X9Y153_A5Q),
.I2(CLBLM_R_X7Y152_SLICE_X8Y152_DQ),
.I3(CLBLM_L_X10Y150_SLICE_X13Y150_CQ),
.I4(1'b1),
.I5(CLBLM_R_X5Y152_SLICE_X7Y152_DO5),
.O5(CLBLM_R_X7Y152_SLICE_X8Y152_DO5),
.O6(CLBLM_R_X7Y152_SLICE_X8Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafa5050eeee4444)
  ) CLBLM_R_X7Y152_SLICE_X8Y152_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y152_SLICE_X8Y152_CQ),
.I2(CLBLM_R_X7Y153_SLICE_X9Y153_DQ),
.I3(1'b1),
.I4(CLBLM_R_X7Y155_SLICE_X8Y155_A5Q),
.I5(CLBLM_R_X5Y152_SLICE_X7Y152_DO5),
.O5(CLBLM_R_X7Y152_SLICE_X8Y152_CO5),
.O6(CLBLM_R_X7Y152_SLICE_X8Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcacfcacfcac0cac0)
  ) CLBLM_R_X7Y152_SLICE_X8Y152_BLUT (
.I0(CLBLM_L_X8Y154_SLICE_X10Y154_AQ),
.I1(CLBLM_L_X10Y151_SLICE_X13Y151_DQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X5Y152_SLICE_X7Y152_DO5),
.I4(1'b1),
.I5(CLBLM_R_X7Y152_SLICE_X8Y152_BQ),
.O5(CLBLM_R_X7Y152_SLICE_X8Y152_BO5),
.O6(CLBLM_R_X7Y152_SLICE_X8Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ccccff00c0c0)
  ) CLBLM_R_X7Y152_SLICE_X8Y152_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y152_SLICE_X11Y152_BO6),
.I2(CLBLM_R_X7Y152_SLICE_X8Y152_AQ),
.I3(CLBLM_R_X5Y151_SLICE_X6Y151_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y149_SLICE_X8Y149_BQ),
.O5(CLBLM_R_X7Y152_SLICE_X8Y152_AO5),
.O6(CLBLM_R_X7Y152_SLICE_X8Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y152_SLICE_X9Y152_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y152_SLICE_X9Y152_AO6),
.Q(CLBLM_R_X7Y152_SLICE_X9Y152_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y152_SLICE_X9Y152_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y152_SLICE_X9Y152_BO6),
.Q(CLBLM_R_X7Y152_SLICE_X9Y152_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y152_SLICE_X9Y152_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y152_SLICE_X9Y152_CO6),
.Q(CLBLM_R_X7Y152_SLICE_X9Y152_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffefffffffffff)
  ) CLBLM_R_X7Y152_SLICE_X9Y152_DLUT (
.I0(CLBLM_L_X8Y150_SLICE_X10Y150_BQ),
.I1(CLBLM_R_X5Y152_SLICE_X6Y152_CQ),
.I2(CLBLM_L_X8Y154_SLICE_X10Y154_AQ),
.I3(CLBLM_R_X7Y154_SLICE_X9Y154_AQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X7Y151_SLICE_X8Y151_DO5),
.O5(CLBLM_R_X7Y152_SLICE_X9Y152_DO5),
.O6(CLBLM_R_X7Y152_SLICE_X9Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haac0aac0aac0aac0)
  ) CLBLM_R_X7Y152_SLICE_X9Y152_CLUT (
.I0(CLBLM_R_X7Y150_SLICE_X9Y150_AQ),
.I1(CLBLM_L_X10Y150_SLICE_X12Y150_BQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y152_SLICE_X9Y152_CO5),
.O6(CLBLM_R_X7Y152_SLICE_X9Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0c0c00000c0c)
  ) CLBLM_R_X7Y152_SLICE_X9Y152_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y152_SLICE_X9Y152_BQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y152_SLICE_X8Y152_CQ),
.O5(CLBLM_R_X7Y152_SLICE_X9Y152_BO5),
.O6(CLBLM_R_X7Y152_SLICE_X9Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f00300f3f00300)
  ) CLBLM_R_X7Y152_SLICE_X9Y152_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y153_SLICE_X10Y153_DO5),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X5Y152_SLICE_X6Y152_BQ),
.I4(CLBLM_L_X10Y152_SLICE_X12Y152_BQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y152_SLICE_X9Y152_AO5),
.O6(CLBLM_R_X7Y152_SLICE_X9Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y153_SLICE_X8Y153_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y153_SLICE_X8Y153_AO6),
.Q(CLBLM_R_X7Y153_SLICE_X8Y153_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y153_SLICE_X8Y153_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y153_SLICE_X8Y153_BO6),
.Q(CLBLM_R_X7Y153_SLICE_X8Y153_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y153_SLICE_X8Y153_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y153_SLICE_X8Y153_CO6),
.Q(CLBLM_R_X7Y153_SLICE_X8Y153_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y153_SLICE_X8Y153_D_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y153_SLICE_X8Y153_DO6),
.Q(CLBLM_R_X7Y153_SLICE_X8Y153_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hae04ae04ae04ae04)
  ) CLBLM_R_X7Y153_SLICE_X8Y153_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y153_SLICE_X12Y153_DQ),
.I2(CLBLM_R_X11Y153_SLICE_X14Y153_AO6),
.I3(CLBLL_L_X4Y151_SLICE_X5Y151_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y153_SLICE_X8Y153_DO5),
.O6(CLBLM_R_X7Y153_SLICE_X8Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f05544f0f00044)
  ) CLBLM_R_X7Y153_SLICE_X8Y153_CLUT (
.I0(RIOB33_X105Y121_IOB_X1Y121_I),
.I1(CLBLM_R_X7Y153_SLICE_X8Y153_CQ),
.I2(CLBLM_R_X3Y143_SLICE_X3Y143_AQ),
.I3(CLBLM_L_X10Y156_SLICE_X12Y156_CO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLL_L_X4Y147_SLICE_X5Y147_B5Q),
.O5(CLBLM_R_X7Y153_SLICE_X8Y153_CO5),
.O6(CLBLM_R_X7Y153_SLICE_X8Y153_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff4fff40004f0040)
  ) CLBLM_R_X7Y153_SLICE_X8Y153_BLUT (
.I0(CLBLM_R_X7Y155_SLICE_X8Y155_BO5),
.I1(CLBLM_R_X7Y153_SLICE_X8Y153_BQ),
.I2(CLBLM_R_X5Y155_SLICE_X7Y155_CO6),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y155_SLICE_X9Y155_AQ),
.I5(CLBLM_R_X3Y146_SLICE_X3Y146_CQ),
.O5(CLBLM_R_X7Y153_SLICE_X8Y153_BO5),
.O6(CLBLM_R_X7Y153_SLICE_X8Y153_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00ffffbfbf)
  ) CLBLM_R_X7Y153_SLICE_X8Y153_ALUT (
.I0(CLBLM_R_X5Y154_SLICE_X6Y154_BO6),
.I1(RIOB33_X105Y135_IOB_X1Y136_I),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(CLBLM_L_X10Y153_SLICE_X12Y153_DQ),
.I4(RIOB33_X105Y135_IOB_X1Y135_I),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X7Y153_SLICE_X8Y153_AO5),
.O6(CLBLM_R_X7Y153_SLICE_X8Y153_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y153_SLICE_X9Y153_A5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y153_SLICE_X9Y153_CO6),
.Q(CLBLM_R_X7Y153_SLICE_X9Y153_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y153_SLICE_X9Y153_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y153_SLICE_X9Y153_AO6),
.Q(CLBLM_R_X7Y153_SLICE_X9Y153_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y153_SLICE_X9Y153_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y153_SLICE_X9Y153_BO6),
.Q(CLBLM_R_X7Y153_SLICE_X9Y153_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y153_SLICE_X9Y153_D_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y153_SLICE_X9Y153_DO6),
.Q(CLBLM_R_X7Y153_SLICE_X9Y153_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'habbaabba01100110)
  ) CLBLM_R_X7Y153_SLICE_X9Y153_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLL_L_X4Y147_SLICE_X4Y147_CQ),
.I3(CLBLM_L_X8Y150_SLICE_X10Y150_DO6),
.I4(1'b1),
.I5(CLBLM_L_X8Y152_SLICE_X10Y152_AQ),
.O5(CLBLM_R_X7Y153_SLICE_X9Y153_DO5),
.O6(CLBLM_R_X7Y153_SLICE_X9Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0c000c50505050)
  ) CLBLM_R_X7Y153_SLICE_X9Y153_CLUT (
.I0(CLBLM_R_X3Y152_SLICE_X3Y152_CO6),
.I1(CLBLM_R_X7Y154_SLICE_X9Y154_AQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y153_SLICE_X8Y153_DQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y153_SLICE_X9Y153_CO5),
.O6(CLBLM_R_X7Y153_SLICE_X9Y153_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000cacacaca)
  ) CLBLM_R_X7Y153_SLICE_X9Y153_BLUT (
.I0(CLBLM_L_X8Y152_SLICE_X11Y152_AQ),
.I1(CLBLM_R_X7Y153_SLICE_X9Y153_BQ),
.I2(CLBLM_L_X8Y152_SLICE_X11Y152_BO6),
.I3(1'b1),
.I4(CLBLM_R_X5Y153_SLICE_X7Y153_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X7Y153_SLICE_X9Y153_BO5),
.O6(CLBLM_R_X7Y153_SLICE_X9Y153_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55ff55fa50ea40)
  ) CLBLM_R_X7Y153_SLICE_X9Y153_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y146_SLICE_X10Y146_BQ),
.I2(CLBLM_R_X7Y155_SLICE_X8Y155_BO5),
.I3(CLBLM_L_X8Y144_SLICE_X10Y144_BQ),
.I4(CLBLM_R_X5Y146_SLICE_X7Y146_BO6),
.I5(CLBLM_R_X7Y154_SLICE_X9Y154_CO6),
.O5(CLBLM_R_X7Y153_SLICE_X9Y153_AO5),
.O6(CLBLM_R_X7Y153_SLICE_X9Y153_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y154_SLICE_X8Y154_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y154_SLICE_X8Y154_AO6),
.Q(CLBLM_R_X7Y154_SLICE_X8Y154_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y154_SLICE_X8Y154_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y154_SLICE_X8Y154_BO6),
.Q(CLBLM_R_X7Y154_SLICE_X8Y154_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y154_SLICE_X8Y154_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y154_SLICE_X8Y154_CO6),
.Q(CLBLM_R_X7Y154_SLICE_X8Y154_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0050505055055051)
  ) CLBLM_R_X7Y154_SLICE_X8Y154_DLUT (
.I0(CLBLM_R_X5Y153_SLICE_X6Y153_CO6),
.I1(CLBLM_R_X7Y155_SLICE_X8Y155_A5Q),
.I2(CLBLL_L_X4Y147_SLICE_X5Y147_B5Q),
.I3(CLBLM_R_X7Y153_SLICE_X8Y153_CQ),
.I4(CLBLM_L_X10Y156_SLICE_X12Y156_CO6),
.I5(CLBLM_R_X7Y154_SLICE_X8Y154_BQ),
.O5(CLBLM_R_X7Y154_SLICE_X8Y154_DO5),
.O6(CLBLM_R_X7Y154_SLICE_X8Y154_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0e4e4a0a0e4e4)
  ) CLBLM_R_X7Y154_SLICE_X8Y154_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y154_SLICE_X8Y154_CQ),
.I2(CLBLM_R_X5Y152_SLICE_X6Y152_AQ),
.I3(1'b1),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y154_SLICE_X8Y154_CO5),
.O6(CLBLM_R_X7Y154_SLICE_X8Y154_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fcf0f6000c0006)
  ) CLBLM_R_X7Y154_SLICE_X8Y154_BLUT (
.I0(CLBLM_L_X10Y156_SLICE_X12Y156_CO6),
.I1(CLBLM_R_X7Y154_SLICE_X8Y154_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(CLBLM_L_X8Y154_SLICE_X10Y154_BO6),
.I5(CLBLM_R_X7Y150_SLICE_X8Y150_CQ),
.O5(CLBLM_R_X7Y154_SLICE_X8Y154_BO5),
.O6(CLBLM_R_X7Y154_SLICE_X8Y154_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd11fd31cc00ec20)
  ) CLBLM_R_X7Y154_SLICE_X8Y154_ALUT (
.I0(CLBLM_R_X5Y155_SLICE_X7Y155_CO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X7Y154_SLICE_X8Y154_AQ),
.I3(CLBLM_R_X7Y151_SLICE_X8Y151_A5Q),
.I4(CLBLM_R_X7Y155_SLICE_X8Y155_BO5),
.I5(CLBLM_R_X7Y153_SLICE_X8Y153_BQ),
.O5(CLBLM_R_X7Y154_SLICE_X8Y154_AO5),
.O6(CLBLM_R_X7Y154_SLICE_X8Y154_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y154_SLICE_X9Y154_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y154_SLICE_X9Y154_AO6),
.Q(CLBLM_R_X7Y154_SLICE_X9Y154_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y154_SLICE_X9Y154_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y154_SLICE_X9Y154_BO6),
.Q(CLBLM_R_X7Y154_SLICE_X9Y154_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha5a5b4b41eb41eb4)
  ) CLBLM_R_X7Y154_SLICE_X9Y154_DLUT (
.I0(CLBLM_R_X7Y153_SLICE_X9Y153_AQ),
.I1(CLBLM_R_X7Y155_SLICE_X8Y155_A5Q),
.I2(CLBLM_R_X7Y153_SLICE_X9Y153_CO5),
.I3(CLBLM_R_X7Y153_SLICE_X8Y153_CQ),
.I4(CLBLL_L_X4Y147_SLICE_X5Y147_B5Q),
.I5(CLBLM_R_X7Y154_SLICE_X8Y154_BQ),
.O5(CLBLM_R_X7Y154_SLICE_X9Y154_DO5),
.O6(CLBLM_R_X7Y154_SLICE_X9Y154_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5a5a4a4a5a5a4a48)
  ) CLBLM_R_X7Y154_SLICE_X9Y154_CLUT (
.I0(CLBLM_R_X7Y153_SLICE_X9Y153_AQ),
.I1(CLBLM_R_X7Y153_SLICE_X8Y153_CQ),
.I2(CLBLM_R_X5Y155_SLICE_X7Y155_BO5),
.I3(CLBLM_R_X7Y155_SLICE_X8Y155_A5Q),
.I4(CLBLL_L_X4Y147_SLICE_X5Y147_B5Q),
.I5(CLBLM_R_X7Y154_SLICE_X8Y154_BQ),
.O5(CLBLM_R_X7Y154_SLICE_X9Y154_CO5),
.O6(CLBLM_R_X7Y154_SLICE_X9Y154_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff0ffcc00f000cc)
  ) CLBLM_R_X7Y154_SLICE_X9Y154_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y155_SLICE_X9Y155_BO6),
.I2(CLBLM_R_X7Y151_SLICE_X9Y151_DO5),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y155_SLICE_X8Y155_BO5),
.I5(CLBLM_R_X11Y154_SLICE_X14Y154_AQ),
.O5(CLBLM_R_X7Y154_SLICE_X9Y154_BO5),
.O6(CLBLM_R_X7Y154_SLICE_X9Y154_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc00aacccc00aa)
  ) CLBLM_R_X7Y154_SLICE_X9Y154_ALUT (
.I0(CLBLM_L_X8Y154_SLICE_X10Y154_AQ),
.I1(CLBLM_L_X8Y152_SLICE_X11Y152_AQ),
.I2(1'b1),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y154_SLICE_X9Y154_AO5),
.O6(CLBLM_R_X7Y154_SLICE_X9Y154_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y155_SLICE_X8Y155_A5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y155_SLICE_X8Y155_AO5),
.Q(CLBLM_R_X7Y155_SLICE_X8Y155_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y155_SLICE_X8Y155_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y155_SLICE_X8Y155_AO6),
.Q(CLBLM_R_X7Y155_SLICE_X8Y155_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000551500005414)
  ) CLBLM_R_X7Y155_SLICE_X8Y155_DLUT (
.I0(RIOB33_X105Y121_IOB_X1Y121_I),
.I1(CLBLM_R_X7Y155_SLICE_X8Y155_AQ),
.I2(CLBLM_L_X8Y153_SLICE_X10Y153_AQ),
.I3(CLBLM_R_X5Y155_SLICE_X7Y155_CO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y155_SLICE_X8Y155_BO6),
.O5(CLBLM_R_X7Y155_SLICE_X8Y155_DO5),
.O6(CLBLM_R_X7Y155_SLICE_X8Y155_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000031ccff00)
  ) CLBLM_R_X7Y155_SLICE_X8Y155_CLUT (
.I0(CLBLM_R_X7Y154_SLICE_X8Y154_BQ),
.I1(CLBLM_R_X7Y155_SLICE_X8Y155_AQ),
.I2(CLBLM_L_X10Y156_SLICE_X12Y156_CO6),
.I3(CLBLM_R_X7Y155_SLICE_X8Y155_A5Q),
.I4(CLBLM_R_X5Y155_SLICE_X7Y155_BO5),
.I5(CLBLM_R_X5Y153_SLICE_X6Y153_CO6),
.O5(CLBLM_R_X7Y155_SLICE_X8Y155_CO5),
.O6(CLBLM_R_X7Y155_SLICE_X8Y155_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0002000000000003)
  ) CLBLM_R_X7Y155_SLICE_X8Y155_BLUT (
.I0(CLBLM_R_X5Y155_SLICE_X7Y155_BO5),
.I1(CLBLM_R_X7Y155_SLICE_X8Y155_A5Q),
.I2(CLBLM_R_X7Y153_SLICE_X8Y153_CQ),
.I3(CLBLL_L_X4Y147_SLICE_X5Y147_B5Q),
.I4(CLBLM_R_X7Y154_SLICE_X8Y154_BQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y155_SLICE_X8Y155_BO5),
.O6(CLBLM_R_X7Y155_SLICE_X8Y155_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfaaafaaaffffc0c0)
  ) CLBLM_R_X7Y155_SLICE_X8Y155_ALUT (
.I0(CLBLM_R_X7Y155_SLICE_X8Y155_DO6),
.I1(CLBLL_L_X4Y154_SLICE_X5Y154_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y150_SLICE_X12Y150_A5Q),
.I4(CLBLM_R_X7Y155_SLICE_X8Y155_CO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y155_SLICE_X8Y155_AO5),
.O6(CLBLM_R_X7Y155_SLICE_X8Y155_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y155_SLICE_X9Y155_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y155_SLICE_X9Y155_AO6),
.Q(CLBLM_R_X7Y155_SLICE_X9Y155_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y155_SLICE_X9Y155_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y155_SLICE_X9Y155_DO5),
.O6(CLBLM_R_X7Y155_SLICE_X9Y155_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfeff323200000000)
  ) CLBLM_R_X7Y155_SLICE_X9Y155_CLUT (
.I0(CLBLM_R_X7Y153_SLICE_X8Y153_CQ),
.I1(CLBLM_R_X7Y155_SLICE_X8Y155_A5Q),
.I2(CLBLL_L_X4Y147_SLICE_X5Y147_B5Q),
.I3(CLBLM_R_X7Y155_SLICE_X8Y155_AQ),
.I4(CLBLM_R_X7Y154_SLICE_X8Y154_BQ),
.I5(CLBLM_R_X5Y152_SLICE_X6Y152_BQ),
.O5(CLBLM_R_X7Y155_SLICE_X9Y155_CO5),
.O6(CLBLM_R_X7Y155_SLICE_X9Y155_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00ae0cff00ff0c)
  ) CLBLM_R_X7Y155_SLICE_X9Y155_BLUT (
.I0(CLBLM_R_X7Y154_SLICE_X9Y154_DO6),
.I1(CLBLL_L_X4Y147_SLICE_X5Y147_B5Q),
.I2(CLBLM_R_X7Y154_SLICE_X8Y154_BQ),
.I3(CLBLM_R_X7Y154_SLICE_X9Y154_BQ),
.I4(CLBLM_R_X7Y153_SLICE_X8Y153_CQ),
.I5(CLBLM_R_X7Y155_SLICE_X9Y155_CO6),
.O5(CLBLM_R_X7Y155_SLICE_X9Y155_BO5),
.O6(CLBLM_R_X7Y155_SLICE_X9Y155_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffff540000ff54)
  ) CLBLM_R_X7Y155_SLICE_X9Y155_ALUT (
.I0(CLBLM_R_X5Y155_SLICE_X7Y155_CO6),
.I1(CLBLM_L_X8Y153_SLICE_X10Y153_AQ),
.I2(CLBLM_R_X7Y155_SLICE_X9Y155_AQ),
.I3(CLBLM_R_X7Y155_SLICE_X8Y155_BO5),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X5Y152_SLICE_X6Y152_CQ),
.O5(CLBLM_R_X7Y155_SLICE_X9Y155_AO5),
.O6(CLBLM_R_X7Y155_SLICE_X9Y155_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y157_SLICE_X8Y157_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y157_SLICE_X14Y157_AO6),
.Q(CLBLM_R_X7Y157_SLICE_X8Y157_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y157_SLICE_X8Y157_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y157_SLICE_X8Y157_DO5),
.O6(CLBLM_R_X7Y157_SLICE_X8Y157_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y157_SLICE_X8Y157_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y157_SLICE_X8Y157_CO5),
.O6(CLBLM_R_X7Y157_SLICE_X8Y157_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y157_SLICE_X8Y157_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y157_SLICE_X8Y157_BO5),
.O6(CLBLM_R_X7Y157_SLICE_X8Y157_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y157_SLICE_X8Y157_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y157_SLICE_X8Y157_AO5),
.O6(CLBLM_R_X7Y157_SLICE_X8Y157_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y157_SLICE_X9Y157_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y157_SLICE_X9Y157_DO5),
.O6(CLBLM_R_X7Y157_SLICE_X9Y157_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y157_SLICE_X9Y157_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y157_SLICE_X9Y157_CO5),
.O6(CLBLM_R_X7Y157_SLICE_X9Y157_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y157_SLICE_X9Y157_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y157_SLICE_X9Y157_BO5),
.O6(CLBLM_R_X7Y157_SLICE_X9Y157_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y157_SLICE_X9Y157_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y157_SLICE_X9Y157_AO5),
.O6(CLBLM_R_X7Y157_SLICE_X9Y157_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y143_SLICE_X14Y143_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y143_SLICE_X14Y143_AO6),
.Q(CLBLM_R_X11Y143_SLICE_X14Y143_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y143_SLICE_X14Y143_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y143_SLICE_X14Y143_BO6),
.Q(CLBLM_R_X11Y143_SLICE_X14Y143_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y143_SLICE_X14Y143_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y143_SLICE_X14Y143_DO5),
.O6(CLBLM_R_X11Y143_SLICE_X14Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccc6fafaffff)
  ) CLBLM_R_X11Y143_SLICE_X14Y143_CLUT (
.I0(CLBLM_L_X12Y145_SLICE_X16Y145_AQ),
.I1(CLBLM_R_X7Y146_SLICE_X9Y146_CQ),
.I2(CLBLM_L_X12Y144_SLICE_X16Y144_BQ),
.I3(CLBLM_L_X12Y144_SLICE_X16Y144_CQ),
.I4(CLBLM_L_X12Y144_SLICE_X16Y144_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y143_SLICE_X14Y143_CO5),
.O6(CLBLM_R_X11Y143_SLICE_X14Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0f5a0e4a0f5a0e4)
  ) CLBLM_R_X11Y143_SLICE_X14Y143_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X11Y143_SLICE_X14Y143_BQ),
.I2(CLBLM_R_X11Y143_SLICE_X14Y143_AQ),
.I3(CLBLL_L_X4Y145_SLICE_X5Y145_DO6),
.I4(CLBLM_L_X10Y143_SLICE_X13Y143_BQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y143_SLICE_X14Y143_BO5),
.O6(CLBLM_R_X11Y143_SLICE_X14Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heeeaeeea44404440)
  ) CLBLM_R_X11Y143_SLICE_X14Y143_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y142_SLICE_X8Y142_DO6),
.I2(CLBLM_R_X11Y143_SLICE_X14Y143_AQ),
.I3(CLBLM_L_X8Y144_SLICE_X11Y144_AQ),
.I4(1'b1),
.I5(CLBLM_R_X11Y145_SLICE_X14Y145_BQ),
.O5(CLBLM_R_X11Y143_SLICE_X14Y143_AO5),
.O6(CLBLM_R_X11Y143_SLICE_X14Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y143_SLICE_X15Y143_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y143_SLICE_X15Y143_DO5),
.O6(CLBLM_R_X11Y143_SLICE_X15Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y143_SLICE_X15Y143_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y143_SLICE_X15Y143_CO5),
.O6(CLBLM_R_X11Y143_SLICE_X15Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y143_SLICE_X15Y143_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y143_SLICE_X15Y143_BO5),
.O6(CLBLM_R_X11Y143_SLICE_X15Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y143_SLICE_X15Y143_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y143_SLICE_X15Y143_AO5),
.O6(CLBLM_R_X11Y143_SLICE_X15Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y144_SLICE_X14Y144_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y144_SLICE_X14Y144_AO6),
.Q(CLBLM_R_X11Y144_SLICE_X14Y144_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y144_SLICE_X14Y144_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y144_SLICE_X14Y144_BO6),
.Q(CLBLM_R_X11Y144_SLICE_X14Y144_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffefefefe)
  ) CLBLM_R_X11Y144_SLICE_X14Y144_DLUT (
.I0(CLBLM_R_X11Y143_SLICE_X14Y143_BQ),
.I1(CLBLM_R_X7Y144_SLICE_X8Y144_DQ),
.I2(CLBLM_R_X11Y145_SLICE_X14Y145_BQ),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X12Y145_SLICE_X16Y145_BQ),
.O5(CLBLM_R_X11Y144_SLICE_X14Y144_DO5),
.O6(CLBLM_R_X11Y144_SLICE_X14Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00001e0000001eff)
  ) CLBLM_R_X11Y144_SLICE_X14Y144_CLUT (
.I0(CLBLM_L_X12Y144_SLICE_X16Y144_BQ),
.I1(CLBLM_R_X11Y144_SLICE_X15Y144_AO5),
.I2(CLBLM_R_X7Y144_SLICE_X8Y144_DQ),
.I3(CLBLM_R_X7Y142_SLICE_X8Y142_DO6),
.I4(CLBLM_R_X11Y144_SLICE_X14Y144_BQ),
.I5(CLBLM_R_X3Y145_SLICE_X3Y145_DQ),
.O5(CLBLM_R_X11Y144_SLICE_X14Y144_CO5),
.O6(CLBLM_R_X11Y144_SLICE_X14Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0f3f3c0f3)
  ) CLBLM_R_X11Y144_SLICE_X14Y144_BLUT (
.I0(1'b1),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X11Y144_SLICE_X14Y144_AQ),
.I3(RIOB33_X105Y141_IOB_X1Y142_I),
.I4(CLBLM_R_X5Y142_SLICE_X7Y142_AQ),
.I5(CLBLM_R_X11Y144_SLICE_X14Y144_CO6),
.O5(CLBLM_R_X11Y144_SLICE_X14Y144_BO5),
.O6(CLBLM_R_X11Y144_SLICE_X14Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffc000c0ffc000c0)
  ) CLBLM_R_X11Y144_SLICE_X14Y144_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X11Y144_SLICE_X14Y144_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X5Y145_SLICE_X6Y145_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y144_SLICE_X14Y144_AO5),
.O6(CLBLM_R_X11Y144_SLICE_X14Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6666676766666666)
  ) CLBLM_R_X11Y144_SLICE_X15Y144_DLUT (
.I0(CLBLM_R_X11Y145_SLICE_X15Y145_AQ),
.I1(CLBLM_L_X10Y144_SLICE_X13Y144_CQ),
.I2(CLBLM_R_X11Y144_SLICE_X14Y144_DO6),
.I3(1'b1),
.I4(CLBLM_R_X11Y145_SLICE_X15Y145_DO6),
.I5(CLBLM_R_X11Y144_SLICE_X15Y144_BO6),
.O5(CLBLM_R_X11Y144_SLICE_X15Y144_DO5),
.O6(CLBLM_R_X11Y144_SLICE_X15Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00002020ffffdfdf)
  ) CLBLM_R_X11Y144_SLICE_X15Y144_CLUT (
.I0(CLBLM_L_X12Y144_SLICE_X16Y144_AQ),
.I1(CLBLM_L_X12Y144_SLICE_X16Y144_BQ),
.I2(CLBLM_L_X12Y144_SLICE_X16Y144_CQ),
.I3(1'b1),
.I4(CLBLM_L_X12Y145_SLICE_X16Y145_AQ),
.I5(CLBLM_L_X10Y146_SLICE_X12Y146_BQ),
.O5(CLBLM_R_X11Y144_SLICE_X15Y144_CO5),
.O6(CLBLM_R_X11Y144_SLICE_X15Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000001)
  ) CLBLM_R_X11Y144_SLICE_X15Y144_BLUT (
.I0(CLBLM_L_X10Y145_SLICE_X13Y145_CQ),
.I1(CLBLM_L_X10Y146_SLICE_X12Y146_BQ),
.I2(CLBLM_L_X10Y143_SLICE_X13Y143_BQ),
.I3(CLBLM_R_X7Y142_SLICE_X8Y142_BQ),
.I4(CLBLM_R_X11Y146_SLICE_X15Y146_AQ),
.I5(CLBLM_R_X7Y142_SLICE_X8Y142_CQ),
.O5(CLBLM_R_X11Y144_SLICE_X15Y144_BO5),
.O6(CLBLM_R_X11Y144_SLICE_X15Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa9aaaaaffffff33)
  ) CLBLM_R_X11Y144_SLICE_X15Y144_ALUT (
.I0(CLBLM_L_X10Y145_SLICE_X13Y145_CQ),
.I1(CLBLM_L_X12Y144_SLICE_X16Y144_CQ),
.I2(CLBLM_L_X12Y144_SLICE_X16Y144_BQ),
.I3(CLBLM_L_X12Y144_SLICE_X16Y144_AQ),
.I4(CLBLM_L_X12Y145_SLICE_X16Y145_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y144_SLICE_X15Y144_AO5),
.O6(CLBLM_R_X11Y144_SLICE_X15Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y145_SLICE_X14Y145_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y145_SLICE_X14Y145_AO6),
.Q(CLBLM_R_X11Y145_SLICE_X14Y145_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y145_SLICE_X14Y145_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y145_SLICE_X14Y145_BO6),
.Q(CLBLM_R_X11Y145_SLICE_X14Y145_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h1010003323230033)
  ) CLBLM_R_X11Y145_SLICE_X14Y145_DLUT (
.I0(CLBLM_R_X11Y143_SLICE_X14Y143_CO5),
.I1(CLBLM_R_X11Y149_SLICE_X14Y149_CQ),
.I2(CLBLM_L_X12Y144_SLICE_X16Y144_CQ),
.I3(CLBLM_R_X11Y148_SLICE_X15Y148_A5Q),
.I4(CLBLM_R_X7Y142_SLICE_X8Y142_DO6),
.I5(CLBLM_L_X10Y146_SLICE_X12Y146_BQ),
.O5(CLBLM_R_X11Y145_SLICE_X14Y145_DO5),
.O6(CLBLM_R_X11Y145_SLICE_X14Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0132013200003333)
  ) CLBLM_R_X11Y145_SLICE_X14Y145_CLUT (
.I0(CLBLM_R_X11Y143_SLICE_X14Y143_CO5),
.I1(CLBLM_R_X11Y145_SLICE_X14Y145_AQ),
.I2(CLBLM_L_X12Y144_SLICE_X16Y144_CQ),
.I3(CLBLM_R_X7Y142_SLICE_X8Y142_CQ),
.I4(CLBLM_L_X10Y145_SLICE_X13Y145_A5Q),
.I5(CLBLM_R_X7Y142_SLICE_X8Y142_DO6),
.O5(CLBLM_R_X11Y145_SLICE_X14Y145_CO5),
.O6(CLBLM_R_X11Y145_SLICE_X14Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0e000eff0e000e)
  ) CLBLM_R_X11Y145_SLICE_X14Y145_BLUT (
.I0(CLBLM_R_X11Y143_SLICE_X14Y143_BQ),
.I1(CLBLM_R_X11Y145_SLICE_X14Y145_BQ),
.I2(CLBLL_L_X4Y145_SLICE_X5Y145_DO6),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X11Y149_SLICE_X14Y149_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y145_SLICE_X14Y145_BO5),
.O6(CLBLM_R_X11Y145_SLICE_X14Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00fa50ff55)
  ) CLBLM_R_X11Y145_SLICE_X14Y145_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(1'b1),
.I2(CLBLM_R_X5Y142_SLICE_X7Y142_AQ),
.I3(CLBLM_R_X11Y148_SLICE_X14Y148_AQ),
.I4(RIOB33_X105Y141_IOB_X1Y142_I),
.I5(CLBLM_R_X11Y145_SLICE_X14Y145_CO6),
.O5(CLBLM_R_X11Y145_SLICE_X14Y145_AO5),
.O6(CLBLM_R_X11Y145_SLICE_X14Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y145_SLICE_X15Y145_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y145_SLICE_X15Y145_AO6),
.Q(CLBLM_R_X11Y145_SLICE_X15Y145_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y145_SLICE_X15Y145_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y145_SLICE_X15Y145_BO6),
.Q(CLBLM_R_X11Y145_SLICE_X15Y145_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffeeffeeffeeffee)
  ) CLBLM_R_X11Y145_SLICE_X15Y145_DLUT (
.I0(CLBLM_R_X7Y146_SLICE_X9Y146_CQ),
.I1(CLBLM_L_X10Y148_SLICE_X12Y148_BQ),
.I2(1'b1),
.I3(CLBLM_R_X11Y145_SLICE_X15Y145_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y145_SLICE_X15Y145_DO5),
.O6(CLBLM_R_X11Y145_SLICE_X15Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000407300008cbf)
  ) CLBLM_R_X11Y145_SLICE_X15Y145_CLUT (
.I0(CLBLM_R_X11Y144_SLICE_X15Y144_AO5),
.I1(CLBLM_R_X7Y142_SLICE_X8Y142_DO6),
.I2(CLBLM_L_X12Y144_SLICE_X16Y144_BQ),
.I3(CLBLM_R_X15Y151_SLICE_X20Y151_AQ),
.I4(CLBLM_R_X11Y146_SLICE_X15Y146_BQ),
.I5(CLBLM_R_X7Y142_SLICE_X8Y142_BQ),
.O5(CLBLM_R_X11Y145_SLICE_X15Y145_CO5),
.O6(CLBLM_R_X11Y145_SLICE_X15Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0f5a0e4a0f5a0e4)
  ) CLBLM_R_X11Y145_SLICE_X15Y145_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X11Y145_SLICE_X15Y145_BQ),
.I2(CLBLM_L_X10Y154_SLICE_X12Y154_AQ),
.I3(CLBLL_L_X4Y145_SLICE_X5Y145_DO6),
.I4(CLBLM_L_X12Y145_SLICE_X16Y145_BQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y145_SLICE_X15Y145_BO5),
.O6(CLBLM_R_X11Y145_SLICE_X15Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haafeaafe00540054)
  ) CLBLM_R_X11Y145_SLICE_X15Y145_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X11Y145_SLICE_X15Y145_BQ),
.I2(CLBLM_R_X11Y145_SLICE_X15Y145_AQ),
.I3(CLBLL_L_X4Y145_SLICE_X5Y145_DO6),
.I4(1'b1),
.I5(CLBLM_L_X10Y147_SLICE_X12Y147_CQ),
.O5(CLBLM_R_X11Y145_SLICE_X15Y145_AO5),
.O6(CLBLM_R_X11Y145_SLICE_X15Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y146_SLICE_X14Y146_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y146_SLICE_X14Y146_AO6),
.Q(CLBLM_R_X11Y146_SLICE_X14Y146_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y146_SLICE_X14Y146_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y146_SLICE_X14Y146_BO6),
.Q(CLBLM_R_X11Y146_SLICE_X14Y146_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y146_SLICE_X14Y146_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y146_SLICE_X14Y146_CO6),
.Q(CLBLM_R_X11Y146_SLICE_X14Y146_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y146_SLICE_X14Y146_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y146_SLICE_X14Y146_DO6),
.Q(CLBLM_R_X11Y146_SLICE_X14Y146_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000aaaa3000)
  ) CLBLM_R_X11Y146_SLICE_X14Y146_DLUT (
.I0(CLBLM_R_X11Y146_SLICE_X14Y146_BQ),
.I1(CLBLM_L_X8Y147_SLICE_X11Y147_CO6),
.I2(CLBLM_L_X10Y147_SLICE_X13Y147_AQ),
.I3(CLBLM_R_X11Y146_SLICE_X15Y146_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X11Y146_SLICE_X14Y146_DO5),
.O6(CLBLM_R_X11Y146_SLICE_X14Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00aaccaac0)
  ) CLBLM_R_X11Y146_SLICE_X14Y146_CLUT (
.I0(CLBLM_R_X7Y146_SLICE_X9Y146_AQ),
.I1(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.I2(CLBLM_R_X11Y144_SLICE_X14Y144_BQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X11Y146_SLICE_X14Y146_CQ),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_R_X11Y146_SLICE_X14Y146_CO5),
.O6(CLBLM_R_X11Y146_SLICE_X14Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcffcccc30330000)
  ) CLBLM_R_X11Y146_SLICE_X14Y146_BLUT (
.I0(1'b1),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_R_X11Y146_SLICE_X14Y146_BQ),
.I5(CLBLM_L_X8Y146_SLICE_X10Y146_B5Q),
.O5(CLBLM_R_X11Y146_SLICE_X14Y146_BO5),
.O6(CLBLM_R_X11Y146_SLICE_X14Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaaccaaf0aac0)
  ) CLBLM_R_X11Y146_SLICE_X14Y146_ALUT (
.I0(CLBLM_R_X11Y146_SLICE_X14Y146_CQ),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_R_X11Y146_SLICE_X14Y146_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.I5(CLBLM_L_X8Y146_SLICE_X10Y146_B5Q),
.O5(CLBLM_R_X11Y146_SLICE_X14Y146_AO5),
.O6(CLBLM_R_X11Y146_SLICE_X14Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y146_SLICE_X15Y146_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y146_SLICE_X15Y146_AO6),
.Q(CLBLM_R_X11Y146_SLICE_X15Y146_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y146_SLICE_X15Y146_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y146_SLICE_X15Y146_BO6),
.Q(CLBLM_R_X11Y146_SLICE_X15Y146_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y146_SLICE_X15Y146_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y146_SLICE_X15Y146_CO6),
.Q(CLBLM_R_X11Y146_SLICE_X15Y146_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y146_SLICE_X15Y146_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y146_SLICE_X15Y146_DO6),
.Q(CLBLM_R_X11Y146_SLICE_X15Y146_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0cac0cac0cfc0cf)
  ) CLBLM_R_X11Y146_SLICE_X15Y146_DLUT (
.I0(CLBLM_R_X5Y142_SLICE_X7Y142_AQ),
.I1(CLBLM_L_X12Y148_SLICE_X16Y148_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y145_SLICE_X13Y145_DO6),
.I4(1'b1),
.I5(RIOB33_X105Y141_IOB_X1Y142_I),
.O5(CLBLM_R_X11Y146_SLICE_X15Y146_DO5),
.O6(CLBLM_R_X11Y146_SLICE_X15Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0f5a0a0a0e4a0)
  ) CLBLM_R_X11Y146_SLICE_X15Y146_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X11Y146_SLICE_X15Y146_CQ),
.I2(CLBLM_R_X11Y147_SLICE_X15Y147_DQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X11Y146_SLICE_X14Y146_DQ),
.I5(CLBLM_L_X8Y146_SLICE_X10Y146_CQ),
.O5(CLBLM_R_X11Y146_SLICE_X15Y146_CO5),
.O6(CLBLM_R_X11Y146_SLICE_X15Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc0000f0ff)
  ) CLBLM_R_X11Y146_SLICE_X15Y146_BLUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y146_SLICE_X5Y146_AQ),
.I2(CLBLM_R_X5Y142_SLICE_X7Y142_AQ),
.I3(RIOB33_X105Y141_IOB_X1Y142_I),
.I4(CLBLM_R_X11Y145_SLICE_X15Y145_CO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y146_SLICE_X15Y146_BO5),
.O6(CLBLM_R_X11Y146_SLICE_X15Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff33cc00fc30cc00)
  ) CLBLM_R_X11Y146_SLICE_X15Y146_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X11Y146_SLICE_X15Y146_AQ),
.I3(CLBLM_R_X11Y148_SLICE_X15Y148_AQ),
.I4(CLBLM_R_X7Y142_SLICE_X8Y142_DO6),
.I5(CLBLM_R_X7Y142_SLICE_X8Y142_CQ),
.O5(CLBLM_R_X11Y146_SLICE_X15Y146_AO5),
.O6(CLBLM_R_X11Y146_SLICE_X15Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y147_SLICE_X14Y147_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y147_SLICE_X14Y147_AO6),
.Q(CLBLM_R_X11Y147_SLICE_X14Y147_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y147_SLICE_X14Y147_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y147_SLICE_X14Y147_BO6),
.Q(CLBLM_R_X11Y147_SLICE_X14Y147_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6666999999996666)
  ) CLBLM_R_X11Y147_SLICE_X14Y147_DLUT (
.I0(CLBLM_R_X7Y145_SLICE_X9Y145_BQ),
.I1(CLBLM_R_X11Y147_SLICE_X14Y147_AQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_L_X12Y147_SLICE_X16Y147_AQ),
.I5(CLBLM_R_X7Y146_SLICE_X9Y146_BQ),
.O5(CLBLM_R_X11Y147_SLICE_X14Y147_DO5),
.O6(CLBLM_R_X11Y147_SLICE_X14Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000005000000050)
  ) CLBLM_R_X11Y147_SLICE_X14Y147_CLUT (
.I0(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.I1(1'b1),
.I2(CLBLM_R_X3Y147_SLICE_X2Y147_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_R_X11Y146_SLICE_X14Y146_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y147_SLICE_X14Y147_CO5),
.O6(CLBLM_R_X11Y147_SLICE_X14Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa03030c0c)
  ) CLBLM_R_X11Y147_SLICE_X14Y147_BLUT (
.I0(CLBLM_L_X12Y150_SLICE_X16Y150_BQ),
.I1(CLBLM_R_X11Y147_SLICE_X14Y147_BQ),
.I2(CLBLM_R_X11Y146_SLICE_X14Y146_AQ),
.I3(1'b1),
.I4(CLBLL_L_X4Y146_SLICE_X4Y146_DO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y147_SLICE_X14Y147_BO5),
.O6(CLBLM_R_X11Y147_SLICE_X14Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hb8b8b8b8b8b8bb88)
  ) CLBLM_R_X11Y147_SLICE_X14Y147_ALUT (
.I0(CLBLM_R_X7Y151_SLICE_X8Y151_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X11Y146_SLICE_X14Y146_CQ),
.I3(CLBLM_R_X11Y147_SLICE_X14Y147_AQ),
.I4(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_R_X11Y147_SLICE_X14Y147_AO5),
.O6(CLBLM_R_X11Y147_SLICE_X14Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y147_SLICE_X15Y147_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y147_SLICE_X15Y147_AO6),
.Q(CLBLM_R_X11Y147_SLICE_X15Y147_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y147_SLICE_X15Y147_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y147_SLICE_X15Y147_BO6),
.Q(CLBLM_R_X11Y147_SLICE_X15Y147_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y147_SLICE_X15Y147_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y147_SLICE_X15Y147_CO6),
.Q(CLBLM_R_X11Y147_SLICE_X15Y147_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y147_SLICE_X15Y147_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y147_SLICE_X15Y147_DO6),
.Q(CLBLM_R_X11Y147_SLICE_X15Y147_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffcffa800fc00a8)
  ) CLBLM_R_X11Y147_SLICE_X15Y147_DLUT (
.I0(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.I1(CLBLM_R_X5Y146_SLICE_X7Y146_DO6),
.I2(CLBLM_R_X11Y147_SLICE_X15Y147_DQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLM_L_X12Y152_SLICE_X17Y152_AQ),
.O5(CLBLM_R_X11Y147_SLICE_X15Y147_DO5),
.O6(CLBLM_R_X11Y147_SLICE_X15Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hee44fe54aa00aa00)
  ) CLBLM_R_X11Y147_SLICE_X15Y147_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X11Y147_SLICE_X15Y147_CQ),
.I2(CLBLM_R_X11Y146_SLICE_X14Y146_DQ),
.I3(CLBLM_L_X10Y143_SLICE_X13Y143_BQ),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X11Y147_SLICE_X15Y147_CO5),
.O6(CLBLM_R_X11Y147_SLICE_X15Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00fafac8c8)
  ) CLBLM_R_X11Y147_SLICE_X15Y147_BLUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_R_X11Y147_SLICE_X15Y147_BQ),
.I2(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.I3(CLBLM_R_X7Y145_SLICE_X8Y145_BQ),
.I4(CLBLM_L_X10Y147_SLICE_X13Y147_CO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y147_SLICE_X15Y147_BO5),
.O6(CLBLM_R_X11Y147_SLICE_X15Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffccf0cc55cc50)
  ) CLBLM_R_X11Y147_SLICE_X15Y147_ALUT (
.I0(CLBLM_R_X11Y148_SLICE_X15Y148_DO6),
.I1(CLBLM_R_X11Y147_SLICE_X15Y147_BQ),
.I2(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLM_L_X8Y147_SLICE_X11Y147_BO5),
.O5(CLBLM_R_X11Y147_SLICE_X15Y147_AO5),
.O6(CLBLM_R_X11Y147_SLICE_X15Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y148_SLICE_X14Y148_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y148_SLICE_X14Y148_AO6),
.Q(CLBLM_R_X11Y148_SLICE_X14Y148_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y148_SLICE_X14Y148_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y148_SLICE_X14Y148_BO6),
.Q(CLBLM_R_X11Y148_SLICE_X14Y148_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y148_SLICE_X14Y148_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y148_SLICE_X14Y148_CO6),
.Q(CLBLM_R_X11Y148_SLICE_X14Y148_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y148_SLICE_X14Y148_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y148_SLICE_X14Y148_DO6),
.Q(CLBLM_R_X11Y148_SLICE_X14Y148_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888dd88d888)
  ) CLBLM_R_X11Y148_SLICE_X14Y148_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y146_SLICE_X13Y146_AQ),
.I2(CLBLM_R_X11Y148_SLICE_X14Y148_DQ),
.I3(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.I4(CLBLM_R_X5Y148_SLICE_X7Y148_DO6),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_R_X11Y148_SLICE_X14Y148_DO5),
.O6(CLBLM_R_X11Y148_SLICE_X14Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hea40ea40ea40ea40)
  ) CLBLM_R_X11Y148_SLICE_X14Y148_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X11Y148_SLICE_X14Y148_CQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X11Y148_SLICE_X14Y148_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y148_SLICE_X14Y148_CO5),
.O6(CLBLM_R_X11Y148_SLICE_X14Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccfff0ccccaaa0)
  ) CLBLM_R_X11Y148_SLICE_X14Y148_BLUT (
.I0(CLBLM_R_X11Y148_SLICE_X14Y148_BQ),
.I1(CLBLM_R_X11Y147_SLICE_X14Y147_AQ),
.I2(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y148_SLICE_X11Y148_BO6),
.O5(CLBLM_R_X11Y148_SLICE_X14Y148_BO5),
.O6(CLBLM_R_X11Y148_SLICE_X14Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hddddddddd8d8d888)
  ) CLBLM_R_X11Y148_SLICE_X14Y148_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y146_SLICE_X12Y146_D5Q),
.I2(CLBLM_R_X11Y148_SLICE_X14Y148_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.I5(CLBLM_L_X10Y148_SLICE_X13Y148_DO6),
.O5(CLBLM_R_X11Y148_SLICE_X14Y148_AO5),
.O6(CLBLM_R_X11Y148_SLICE_X14Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y148_SLICE_X15Y148_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y150_SLICE_X16Y150_DO6),
.Q(CLBLM_R_X11Y148_SLICE_X15Y148_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y148_SLICE_X15Y148_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y148_SLICE_X15Y148_BO5),
.Q(CLBLM_R_X11Y148_SLICE_X15Y148_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y148_SLICE_X15Y148_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y148_SLICE_X15Y148_AO6),
.Q(CLBLM_R_X11Y148_SLICE_X15Y148_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y148_SLICE_X15Y148_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y148_SLICE_X15Y148_BO6),
.Q(CLBLM_R_X11Y148_SLICE_X15Y148_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y148_SLICE_X15Y148_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y148_SLICE_X15Y148_CO6),
.Q(CLBLM_R_X11Y148_SLICE_X15Y148_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h2121121212122121)
  ) CLBLM_R_X11Y148_SLICE_X15Y148_DLUT (
.I0(CLBLM_L_X10Y151_SLICE_X12Y151_AQ),
.I1(CLBLM_R_X11Y147_SLICE_X15Y147_AQ),
.I2(CLBLM_R_X11Y147_SLICE_X14Y147_DO6),
.I3(1'b1),
.I4(CLBLM_L_X12Y150_SLICE_X16Y150_AQ),
.I5(CLBLM_L_X12Y148_SLICE_X16Y148_CO6),
.O5(CLBLM_R_X11Y148_SLICE_X15Y148_DO5),
.O6(CLBLM_R_X11Y148_SLICE_X15Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffac80000fac8)
  ) CLBLM_R_X11Y148_SLICE_X15Y148_CLUT (
.I0(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.I1(CLBLM_R_X11Y148_SLICE_X15Y148_CQ),
.I2(RIOB33_X105Y117_IOB_X1Y118_I),
.I3(CLBLM_R_X7Y149_SLICE_X9Y149_CO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X11Y145_SLICE_X15Y145_BQ),
.O5(CLBLM_R_X11Y148_SLICE_X15Y148_CO5),
.O6(CLBLM_R_X11Y148_SLICE_X15Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafa0a0afc0cfc0c)
  ) CLBLM_R_X11Y148_SLICE_X15Y148_BLUT (
.I0(RIOB33_X105Y103_IOB_X1Y104_I),
.I1(CLBLM_L_X10Y146_SLICE_X12Y146_D5Q),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X11Y146_SLICE_X15Y146_BQ),
.I4(CLBLM_L_X12Y149_SLICE_X17Y149_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y148_SLICE_X15Y148_BO5),
.O6(CLBLM_R_X11Y148_SLICE_X15Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff3333fcec3020)
  ) CLBLM_R_X11Y148_SLICE_X15Y148_ALUT (
.I0(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X11Y148_SLICE_X15Y148_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_R_X11Y151_SLICE_X14Y151_AQ),
.I5(CLBLM_L_X10Y148_SLICE_X13Y148_DO6),
.O5(CLBLM_R_X11Y148_SLICE_X15Y148_AO5),
.O6(CLBLM_R_X11Y148_SLICE_X15Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y149_SLICE_X14Y149_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y149_SLICE_X14Y149_AO6),
.Q(CLBLM_R_X11Y149_SLICE_X14Y149_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y149_SLICE_X14Y149_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y149_SLICE_X14Y149_BO6),
.Q(CLBLM_R_X11Y149_SLICE_X14Y149_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y149_SLICE_X14Y149_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y149_SLICE_X14Y149_CO6),
.Q(CLBLM_R_X11Y149_SLICE_X14Y149_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffcfffc5faff5fa)
  ) CLBLM_R_X11Y149_SLICE_X14Y149_DLUT (
.I0(CLBLM_R_X11Y147_SLICE_X14Y147_AQ),
.I1(CLBLM_L_X12Y149_SLICE_X16Y149_AQ),
.I2(CLBLM_R_X11Y149_SLICE_X14Y149_BQ),
.I3(CLBLM_R_X11Y150_SLICE_X15Y150_AQ),
.I4(CLBLM_L_X12Y147_SLICE_X16Y147_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y149_SLICE_X14Y149_DO5),
.O6(CLBLM_R_X11Y149_SLICE_X14Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0fff05000f0005)
  ) CLBLM_R_X11Y149_SLICE_X14Y149_CLUT (
.I0(RIOB33_X105Y141_IOB_X1Y142_I),
.I1(1'b1),
.I2(CLBLM_R_X11Y145_SLICE_X14Y145_DO6),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X5Y142_SLICE_X7Y142_AQ),
.I5(CLBLM_R_X7Y151_SLICE_X9Y151_BQ),
.O5(CLBLM_R_X11Y149_SLICE_X14Y149_CO5),
.O6(CLBLM_R_X11Y149_SLICE_X14Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff880088fff000f0)
  ) CLBLM_R_X11Y149_SLICE_X14Y149_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X11Y149_SLICE_X14Y149_BQ),
.I2(CLBLM_R_X11Y149_SLICE_X14Y149_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y153_SLICE_X11Y153_BQ),
.I5(CLBLM_R_X11Y147_SLICE_X14Y147_CO6),
.O5(CLBLM_R_X11Y149_SLICE_X14Y149_BO5),
.O6(CLBLM_R_X11Y149_SLICE_X14Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccca0a0ccccff00)
  ) CLBLM_R_X11Y149_SLICE_X14Y149_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X5Y151_SLICE_X6Y151_BQ),
.I2(CLBLM_R_X11Y149_SLICE_X14Y149_AQ),
.I3(CLBLM_L_X10Y149_SLICE_X13Y149_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X11Y147_SLICE_X14Y147_CO6),
.O5(CLBLM_R_X11Y149_SLICE_X14Y149_AO5),
.O6(CLBLM_R_X11Y149_SLICE_X14Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffffaa)
  ) CLBLM_R_X11Y149_SLICE_X15Y149_DLUT (
.I0(CLBLM_R_X11Y149_SLICE_X14Y149_AQ),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_L_X12Y149_SLICE_X17Y149_BQ),
.I4(CLBLM_L_X10Y150_SLICE_X12Y150_AQ),
.I5(CLBLM_L_X12Y149_SLICE_X17Y149_CQ),
.O5(CLBLM_R_X11Y149_SLICE_X15Y149_DO5),
.O6(CLBLM_R_X11Y149_SLICE_X15Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0ff00ff50ff00ff0)
  ) CLBLM_R_X11Y149_SLICE_X15Y149_CLUT (
.I0(CLBLM_R_X11Y149_SLICE_X14Y149_DO6),
.I1(1'b1),
.I2(CLBLM_R_X11Y150_SLICE_X15Y150_BQ),
.I3(CLBLM_L_X10Y150_SLICE_X13Y150_BQ),
.I4(CLBLM_R_X11Y149_SLICE_X15Y149_DO6),
.I5(CLBLM_R_X11Y149_SLICE_X15Y149_BO6),
.O5(CLBLM_R_X11Y149_SLICE_X15Y149_CO5),
.O6(CLBLM_R_X11Y149_SLICE_X15Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000001)
  ) CLBLM_R_X11Y149_SLICE_X15Y149_BLUT (
.I0(CLBLM_L_X10Y151_SLICE_X12Y151_BQ),
.I1(CLBLM_L_X12Y149_SLICE_X17Y149_AQ),
.I2(CLBLM_L_X12Y148_SLICE_X16Y148_AQ),
.I3(CLBLM_L_X10Y149_SLICE_X13Y149_AQ),
.I4(CLBLM_L_X12Y148_SLICE_X16Y148_BQ),
.I5(CLBLM_L_X12Y150_SLICE_X16Y150_BQ),
.O5(CLBLM_R_X11Y149_SLICE_X15Y149_BO5),
.O6(CLBLM_R_X11Y149_SLICE_X15Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000100)
  ) CLBLM_R_X11Y149_SLICE_X15Y149_ALUT (
.I0(CLBLM_R_X11Y149_SLICE_X15Y149_DO6),
.I1(CLBLM_R_X11Y149_SLICE_X14Y149_BQ),
.I2(CLBLM_L_X12Y149_SLICE_X16Y149_AQ),
.I3(CLBLM_R_X11Y149_SLICE_X15Y149_BO6),
.I4(CLBLM_R_X11Y150_SLICE_X15Y150_AQ),
.I5(CLBLM_L_X10Y150_SLICE_X13Y150_BQ),
.O5(CLBLM_R_X11Y149_SLICE_X15Y149_AO5),
.O6(CLBLM_R_X11Y149_SLICE_X15Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000090900909)
  ) CLBLM_R_X11Y150_SLICE_X14Y150_DLUT (
.I0(CLBLM_L_X10Y151_SLICE_X12Y151_AQ),
.I1(CLBLM_L_X12Y148_SLICE_X16Y148_AQ),
.I2(CLBLM_L_X10Y149_SLICE_X13Y149_AQ),
.I3(1'b1),
.I4(CLBLM_L_X12Y150_SLICE_X16Y150_AQ),
.I5(CLBLM_R_X11Y149_SLICE_X14Y149_DO5),
.O5(CLBLM_R_X11Y150_SLICE_X14Y150_DO5),
.O6(CLBLM_R_X11Y150_SLICE_X14Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h009f0000009f0000)
  ) CLBLM_R_X11Y150_SLICE_X14Y150_CLUT (
.I0(CLBLM_L_X8Y147_SLICE_X11Y147_BO6),
.I1(CLBLM_R_X11Y149_SLICE_X15Y149_CO6),
.I2(CLBLM_R_X11Y151_SLICE_X14Y151_BO5),
.I3(CLBLM_L_X12Y149_SLICE_X16Y149_BO6),
.I4(CLBLM_R_X11Y150_SLICE_X14Y150_DO6),
.I5(1'b1),
.O5(CLBLM_R_X11Y150_SLICE_X14Y150_CO5),
.O6(CLBLM_R_X11Y150_SLICE_X14Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h55ff55ffd5ff75ff)
  ) CLBLM_R_X11Y150_SLICE_X14Y150_BLUT (
.I0(CLBLM_R_X11Y151_SLICE_X14Y151_BO5),
.I1(CLBLM_R_X11Y149_SLICE_X15Y149_CO6),
.I2(CLBLM_R_X11Y150_SLICE_X14Y150_DO6),
.I3(CLBLM_R_X11Y147_SLICE_X14Y147_CO6),
.I4(CLBLM_L_X8Y147_SLICE_X11Y147_BO6),
.I5(CLBLM_L_X12Y149_SLICE_X16Y149_BO6),
.O5(CLBLM_R_X11Y150_SLICE_X14Y150_BO5),
.O6(CLBLM_R_X11Y150_SLICE_X14Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000080000000)
  ) CLBLM_R_X11Y150_SLICE_X14Y150_ALUT (
.I0(CLBLM_R_X11Y147_SLICE_X14Y147_CO6),
.I1(CLBLM_L_X10Y151_SLICE_X13Y151_AQ),
.I2(CLBLM_L_X8Y151_SLICE_X11Y151_BQ),
.I3(CLBLM_R_X11Y151_SLICE_X15Y151_BQ),
.I4(CLBLM_L_X10Y151_SLICE_X13Y151_BQ),
.I5(CLBLM_R_X11Y150_SLICE_X14Y150_CO6),
.O5(CLBLM_R_X11Y150_SLICE_X14Y150_AO5),
.O6(CLBLM_R_X11Y150_SLICE_X14Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y150_SLICE_X15Y150_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y150_SLICE_X15Y150_AO6),
.Q(CLBLM_R_X11Y150_SLICE_X15Y150_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y150_SLICE_X15Y150_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y150_SLICE_X15Y150_BO6),
.Q(CLBLM_R_X11Y150_SLICE_X15Y150_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y150_SLICE_X15Y150_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y150_SLICE_X15Y150_CO6),
.Q(CLBLM_R_X11Y150_SLICE_X15Y150_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3afa3afa3a0a3a0a)
  ) CLBLM_R_X11Y150_SLICE_X15Y150_DLUT (
.I0(CLBLM_L_X8Y147_SLICE_X11Y147_BO6),
.I1(CLBLM_L_X10Y150_SLICE_X13Y150_BQ),
.I2(CLBLM_R_X11Y151_SLICE_X14Y151_BO5),
.I3(CLBLM_R_X11Y150_SLICE_X15Y150_BQ),
.I4(1'b1),
.I5(CLBLM_R_X11Y149_SLICE_X15Y149_AO6),
.O5(CLBLM_R_X11Y150_SLICE_X15Y150_DO5),
.O6(CLBLM_R_X11Y150_SLICE_X15Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff000000e0e0)
  ) CLBLM_R_X11Y150_SLICE_X15Y150_CLUT (
.I0(CLBLM_R_X11Y146_SLICE_X15Y146_BQ),
.I1(CLBLM_R_X11Y150_SLICE_X15Y150_CQ),
.I2(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.I3(CLBLM_R_X11Y150_SLICE_X15Y150_BQ),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y150_SLICE_X15Y150_CO5),
.O6(CLBLM_R_X11Y150_SLICE_X15Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3e2d1c0d1c0d1c0)
  ) CLBLM_R_X11Y150_SLICE_X15Y150_BLUT (
.I0(CLBLM_R_X11Y147_SLICE_X14Y147_CO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y147_SLICE_X13Y147_AQ),
.I3(CLBLM_L_X10Y150_SLICE_X13Y150_BQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X11Y150_SLICE_X15Y150_BQ),
.O5(CLBLM_R_X11Y150_SLICE_X15Y150_BO5),
.O6(CLBLM_R_X11Y150_SLICE_X15Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccf5a05500)
  ) CLBLM_R_X11Y150_SLICE_X15Y150_ALUT (
.I0(CLBLM_R_X11Y147_SLICE_X14Y147_CO6),
.I1(CLBLM_R_X11Y151_SLICE_X15Y151_AQ),
.I2(CLBLM_R_X11Y150_SLICE_X15Y150_AQ),
.I3(CLBLM_R_X11Y150_SLICE_X15Y150_DO6),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y150_SLICE_X15Y150_AO5),
.O6(CLBLM_R_X11Y150_SLICE_X15Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y151_SLICE_X14Y151_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y77_IOB_X0Y77_I),
.D(CLBLM_R_X11Y152_SLICE_X14Y152_CQ),
.Q(CLBLM_R_X11Y151_SLICE_X14Y151_AQ),
.R(CLBLM_R_X11Y151_SLICE_X15Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y151_SLICE_X14Y151_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y77_IOB_X0Y77_I),
.D(CLBLM_R_X11Y148_SLICE_X15Y148_BQ),
.Q(CLBLM_R_X11Y151_SLICE_X14Y151_BQ),
.R(CLBLM_R_X11Y151_SLICE_X15Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00f000ee00ee)
  ) CLBLM_R_X11Y151_SLICE_X14Y151_DLUT (
.I0(CLBLM_R_X11Y148_SLICE_X14Y148_AQ),
.I1(CLBLM_R_X11Y148_SLICE_X14Y148_DQ),
.I2(CLBLM_L_X10Y151_SLICE_X12Y151_DQ),
.I3(CLBLM_L_X8Y146_SLICE_X10Y146_BQ),
.I4(CLBLM_L_X8Y146_SLICE_X11Y146_BQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y151_SLICE_X14Y151_DO5),
.O6(CLBLM_R_X11Y151_SLICE_X14Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00700000007f0000)
  ) CLBLM_R_X11Y151_SLICE_X14Y151_CLUT (
.I0(CLBLM_L_X8Y151_SLICE_X11Y151_BQ),
.I1(CLBLM_L_X10Y151_SLICE_X13Y151_AQ),
.I2(CLBLM_L_X10Y151_SLICE_X13Y151_BQ),
.I3(CLBLM_R_X11Y147_SLICE_X14Y147_CO6),
.I4(CLBLM_R_X11Y151_SLICE_X15Y151_BQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y151_SLICE_X14Y151_CO5),
.O6(CLBLM_R_X11Y151_SLICE_X14Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0200000088000000)
  ) CLBLM_R_X11Y151_SLICE_X14Y151_BLUT (
.I0(CLBLM_L_X10Y151_SLICE_X13Y151_BQ),
.I1(CLBLM_L_X10Y151_SLICE_X13Y151_AQ),
.I2(CLBLM_R_X11Y147_SLICE_X14Y147_CO6),
.I3(CLBLM_R_X11Y151_SLICE_X15Y151_BQ),
.I4(CLBLM_L_X8Y151_SLICE_X11Y151_BQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y151_SLICE_X14Y151_BO5),
.O6(CLBLM_R_X11Y151_SLICE_X14Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccafccfa0000f0f0)
  ) CLBLM_R_X11Y151_SLICE_X14Y151_ALUT (
.I0(CLBLM_R_X11Y154_SLICE_X15Y154_CO6),
.I1(CLBLM_R_X11Y148_SLICE_X14Y148_CQ),
.I2(CLBLM_R_X7Y147_SLICE_X9Y147_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X11Y151_SLICE_X15Y151_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X11Y151_SLICE_X14Y151_AO5),
.O6(CLBLM_R_X11Y151_SLICE_X14Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y151_SLICE_X15Y151_A5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y151_SLICE_X14Y151_AO6),
.Q(CLBLM_R_X11Y151_SLICE_X15Y151_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y151_SLICE_X15Y151_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y151_SLICE_X15Y151_AO6),
.Q(CLBLM_R_X11Y151_SLICE_X15Y151_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y151_SLICE_X15Y151_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y151_SLICE_X15Y151_BO6),
.Q(CLBLM_R_X11Y151_SLICE_X15Y151_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y151_SLICE_X15Y151_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y151_SLICE_X15Y151_DO5),
.O6(CLBLM_R_X11Y151_SLICE_X15Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h2233223322332233)
  ) CLBLM_R_X11Y151_SLICE_X15Y151_CLUT (
.I0(CLBLM_R_X5Y142_SLICE_X7Y142_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(1'b1),
.I3(RIOB33_X105Y141_IOB_X1Y142_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y151_SLICE_X15Y151_CO5),
.O6(CLBLM_R_X11Y151_SLICE_X15Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf888faaaf888f222)
  ) CLBLM_R_X11Y151_SLICE_X15Y151_BLUT (
.I0(CLBLM_R_X5Y151_SLICE_X7Y151_DO6),
.I1(CLBLM_R_X11Y151_SLICE_X15Y151_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X11Y153_SLICE_X15Y153_BQ),
.I4(CLBLM_R_X11Y147_SLICE_X14Y147_CO6),
.I5(CLBLM_R_X11Y151_SLICE_X14Y151_BO5),
.O5(CLBLM_R_X11Y151_SLICE_X15Y151_BO5),
.O6(CLBLM_R_X11Y151_SLICE_X15Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa50ff55fa50fa50)
  ) CLBLM_R_X11Y151_SLICE_X15Y151_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(1'b1),
.I2(CLBLM_R_X11Y151_SLICE_X15Y151_AQ),
.I3(CLBLM_L_X10Y145_SLICE_X13Y145_A5Q),
.I4(CLBLM_R_X5Y142_SLICE_X7Y142_AQ),
.I5(RIOB33_X105Y141_IOB_X1Y142_I),
.O5(CLBLM_R_X11Y151_SLICE_X15Y151_AO5),
.O6(CLBLM_R_X11Y151_SLICE_X15Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y152_SLICE_X14Y152_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y152_SLICE_X14Y152_AO6),
.Q(CLBLM_R_X11Y152_SLICE_X14Y152_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y152_SLICE_X14Y152_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y152_SLICE_X14Y152_BO6),
.Q(CLBLM_R_X11Y152_SLICE_X14Y152_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y152_SLICE_X14Y152_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y152_SLICE_X14Y152_CO6),
.Q(CLBLM_R_X11Y152_SLICE_X14Y152_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y152_SLICE_X14Y152_D_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y152_SLICE_X14Y152_DO6),
.Q(CLBLM_R_X11Y152_SLICE_X14Y152_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hbabaffaa10105500)
  ) CLBLM_R_X11Y152_SLICE_X14Y152_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X11Y154_SLICE_X15Y154_CO6),
.I2(CLBLM_R_X11Y152_SLICE_X14Y152_DQ),
.I3(CLBLM_L_X10Y152_SLICE_X12Y152_BQ),
.I4(CLBLM_R_X11Y153_SLICE_X14Y153_BO5),
.I5(CLBLM_R_X11Y147_SLICE_X14Y147_BQ),
.O5(CLBLM_R_X11Y152_SLICE_X14Y152_DO5),
.O6(CLBLM_R_X11Y152_SLICE_X14Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaeefafa00445050)
  ) CLBLM_R_X11Y152_SLICE_X14Y152_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X11Y152_SLICE_X14Y152_CQ),
.I2(CLBLM_R_X11Y152_SLICE_X14Y152_BQ),
.I3(CLBLM_R_X11Y154_SLICE_X15Y154_CO6),
.I4(CLBLM_R_X11Y153_SLICE_X14Y153_BO5),
.I5(CLBLM_R_X7Y153_SLICE_X9Y153_DQ),
.O5(CLBLM_R_X11Y152_SLICE_X14Y152_CO5),
.O6(CLBLM_R_X11Y152_SLICE_X14Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc5cfc0cac5c5c0c0)
  ) CLBLM_R_X11Y152_SLICE_X14Y152_BLUT (
.I0(CLBLM_R_X11Y153_SLICE_X14Y153_BO5),
.I1(CLBLL_L_X2Y146_SLICE_X1Y146_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X11Y154_SLICE_X15Y154_CO6),
.I4(CLBLM_L_X10Y152_SLICE_X13Y152_BQ),
.I5(CLBLM_R_X11Y152_SLICE_X14Y152_BQ),
.O5(CLBLM_R_X11Y152_SLICE_X14Y152_BO5),
.O6(CLBLM_R_X11Y152_SLICE_X14Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff500050ffcc00cc)
  ) CLBLM_R_X11Y152_SLICE_X14Y152_ALUT (
.I0(CLBLM_R_X11Y154_SLICE_X15Y154_CO6),
.I1(CLBLM_R_X11Y152_SLICE_X14Y152_DQ),
.I2(CLBLM_R_X11Y152_SLICE_X14Y152_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y152_SLICE_X8Y152_DQ),
.I5(CLBLM_R_X11Y153_SLICE_X14Y153_BO5),
.O5(CLBLM_R_X11Y152_SLICE_X14Y152_AO5),
.O6(CLBLM_R_X11Y152_SLICE_X14Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y152_SLICE_X15Y152_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y152_SLICE_X15Y152_AO6),
.Q(CLBLM_R_X11Y152_SLICE_X15Y152_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y152_SLICE_X15Y152_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y152_SLICE_X15Y152_BO6),
.Q(CLBLM_R_X11Y152_SLICE_X15Y152_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y152_SLICE_X15Y152_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y152_SLICE_X15Y152_DO5),
.O6(CLBLM_R_X11Y152_SLICE_X15Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y152_SLICE_X15Y152_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y152_SLICE_X15Y152_CO5),
.O6(CLBLM_R_X11Y152_SLICE_X15Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaf0fcaaaaf3fc)
  ) CLBLM_R_X11Y152_SLICE_X15Y152_BLUT (
.I0(CLBLL_L_X4Y145_SLICE_X5Y145_AQ),
.I1(CLBLM_R_X11Y152_SLICE_X15Y152_BQ),
.I2(CLBLM_R_X11Y154_SLICE_X15Y154_CO6),
.I3(CLBLM_L_X12Y151_SLICE_X16Y151_DO5),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X11Y153_SLICE_X14Y153_CO6),
.O5(CLBLM_R_X11Y152_SLICE_X15Y152_BO5),
.O6(CLBLM_R_X11Y152_SLICE_X15Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc00facccc00af)
  ) CLBLM_R_X11Y152_SLICE_X15Y152_ALUT (
.I0(CLBLM_L_X10Y154_SLICE_X13Y154_CO5),
.I1(CLBLM_L_X8Y155_SLICE_X10Y155_BQ),
.I2(CLBLM_R_X11Y152_SLICE_X15Y152_AQ),
.I3(CLBLM_R_X11Y154_SLICE_X15Y154_CO5),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X12Y152_SLICE_X17Y152_DO6),
.O5(CLBLM_R_X11Y152_SLICE_X15Y152_AO5),
.O6(CLBLM_R_X11Y152_SLICE_X15Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y153_SLICE_X14Y153_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y77_IOB_X0Y77_I),
.D(CLBLM_R_X7Y155_SLICE_X8Y155_AQ),
.Q(CLBLM_R_X11Y153_SLICE_X14Y153_AQ),
.R(CLBLM_R_X11Y151_SLICE_X15Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y153_SLICE_X14Y153_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y77_IOB_X0Y77_I),
.D(CLBLM_R_X11Y154_SLICE_X15Y154_BQ),
.Q(CLBLM_R_X11Y153_SLICE_X14Y153_BQ),
.R(CLBLM_R_X11Y151_SLICE_X15Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y153_SLICE_X14Y153_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y77_IOB_X0Y77_I),
.D(CLBLM_R_X5Y150_SLICE_X7Y150_BQ),
.Q(CLBLM_R_X11Y153_SLICE_X14Y153_CQ),
.R(CLBLM_R_X11Y151_SLICE_X15Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafbffff00330033)
  ) CLBLM_R_X11Y153_SLICE_X14Y153_DLUT (
.I0(CLBLM_R_X11Y153_SLICE_X14Y153_AO6),
.I1(CLBLM_R_X11Y154_SLICE_X14Y154_CO6),
.I2(CLBLM_R_X11Y154_SLICE_X14Y154_DO6),
.I3(CLBLM_L_X10Y154_SLICE_X13Y154_AQ),
.I4(CLBLM_R_X7Y153_SLICE_X8Y153_DQ),
.I5(CLBLM_R_X11Y153_SLICE_X15Y153_BQ),
.O5(CLBLM_R_X11Y153_SLICE_X14Y153_DO5),
.O6(CLBLM_R_X11Y153_SLICE_X14Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0033003355575f5f)
  ) CLBLM_R_X11Y153_SLICE_X14Y153_CLUT (
.I0(CLBLM_L_X12Y151_SLICE_X16Y151_DO5),
.I1(CLBLM_R_X11Y154_SLICE_X15Y154_BQ),
.I2(CLBLM_R_X11Y154_SLICE_X14Y154_BO5),
.I3(CLBLM_R_X11Y154_SLICE_X14Y154_AQ),
.I4(CLBLM_R_X11Y152_SLICE_X15Y152_BQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y153_SLICE_X14Y153_CO5),
.O6(CLBLM_R_X11Y153_SLICE_X14Y153_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3133ffff44440000)
  ) CLBLM_R_X11Y153_SLICE_X14Y153_BLUT (
.I0(CLBLM_L_X10Y153_SLICE_X13Y153_BQ),
.I1(CLBLM_L_X10Y153_SLICE_X13Y153_CQ),
.I2(CLBLM_R_X11Y153_SLICE_X15Y153_CO5),
.I3(CLBLM_R_X11Y154_SLICE_X15Y154_AQ),
.I4(CLBLM_L_X12Y151_SLICE_X16Y151_DO5),
.I5(1'b1),
.O5(CLBLM_R_X11Y153_SLICE_X14Y153_BO5),
.O6(CLBLM_R_X11Y153_SLICE_X14Y153_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ab00ab01000000)
  ) CLBLM_R_X11Y153_SLICE_X14Y153_ALUT (
.I0(CLBLM_L_X10Y153_SLICE_X13Y153_BQ),
.I1(CLBLM_R_X11Y154_SLICE_X15Y154_BQ),
.I2(CLBLM_R_X11Y154_SLICE_X14Y154_AQ),
.I3(CLBLM_R_X11Y154_SLICE_X15Y154_AQ),
.I4(CLBLM_L_X12Y151_SLICE_X16Y151_DO5),
.I5(1'b1),
.O5(CLBLM_R_X11Y153_SLICE_X14Y153_AO5),
.O6(CLBLM_R_X11Y153_SLICE_X14Y153_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y153_SLICE_X15Y153_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y153_SLICE_X15Y153_AO6),
.Q(CLBLM_R_X11Y153_SLICE_X15Y153_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y153_SLICE_X15Y153_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y153_SLICE_X15Y153_BO6),
.Q(CLBLM_R_X11Y153_SLICE_X15Y153_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0ffff0ff03fffc)
  ) CLBLM_R_X11Y153_SLICE_X15Y153_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y153_SLICE_X12Y153_BQ),
.I2(CLBLM_L_X12Y153_SLICE_X16Y153_DO6),
.I3(CLBLM_L_X10Y154_SLICE_X13Y154_CO5),
.I4(CLBLM_R_X11Y153_SLICE_X15Y153_AQ),
.I5(CLBLM_R_X11Y153_SLICE_X14Y153_CO5),
.O5(CLBLM_R_X11Y153_SLICE_X15Y153_DO5),
.O6(CLBLM_R_X11Y153_SLICE_X15Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3202320232023202)
  ) CLBLM_R_X11Y153_SLICE_X15Y153_CLUT (
.I0(CLBLM_R_X13Y152_SLICE_X18Y152_AO6),
.I1(CLBLM_R_X11Y153_SLICE_X14Y153_CO5),
.I2(CLBLM_L_X12Y153_SLICE_X17Y153_AQ),
.I3(CLBLM_R_X13Y152_SLICE_X18Y152_BO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y153_SLICE_X15Y153_CO5),
.O6(CLBLM_R_X11Y153_SLICE_X15Y153_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00fcfcff000c0c)
  ) CLBLM_R_X11Y153_SLICE_X15Y153_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y153_SLICE_X14Y153_DO6),
.I2(CLBLM_R_X11Y154_SLICE_X15Y154_CO6),
.I3(CLBLM_L_X12Y153_SLICE_X17Y153_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLL_L_X4Y144_SLICE_X4Y144_CO6),
.O5(CLBLM_R_X11Y153_SLICE_X15Y153_BO5),
.O6(CLBLM_R_X11Y153_SLICE_X15Y153_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf2f20202f2f20202)
  ) CLBLM_R_X11Y153_SLICE_X15Y153_ALUT (
.I0(CLBLM_R_X11Y153_SLICE_X15Y153_DO6),
.I1(CLBLM_R_X11Y154_SLICE_X15Y154_CO5),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(CLBLM_R_X5Y143_SLICE_X7Y143_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y153_SLICE_X15Y153_AO5),
.O6(CLBLM_R_X11Y153_SLICE_X15Y153_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y154_SLICE_X14Y154_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y154_SLICE_X14Y154_AO6),
.Q(CLBLM_R_X11Y154_SLICE_X14Y154_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h33cca2ff55aaf7aa)
  ) CLBLM_R_X11Y154_SLICE_X14Y154_DLUT (
.I0(CLBLM_R_X11Y154_SLICE_X14Y154_CO5),
.I1(CLBLM_R_X11Y154_SLICE_X15Y154_AQ),
.I2(CLBLM_L_X10Y153_SLICE_X13Y153_CQ),
.I3(CLBLM_L_X10Y154_SLICE_X13Y154_DO6),
.I4(CLBLM_R_X11Y154_SLICE_X14Y154_AQ),
.I5(CLBLM_R_X11Y152_SLICE_X15Y152_BQ),
.O5(CLBLM_R_X11Y154_SLICE_X14Y154_DO5),
.O6(CLBLM_R_X11Y154_SLICE_X14Y154_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hefefefef00005f5f)
  ) CLBLM_R_X11Y154_SLICE_X14Y154_CLUT (
.I0(CLBLM_R_X11Y154_SLICE_X15Y154_AQ),
.I1(CLBLM_R_X11Y154_SLICE_X14Y154_AQ),
.I2(CLBLM_R_X11Y154_SLICE_X15Y154_BQ),
.I3(1'b1),
.I4(CLBLM_L_X10Y153_SLICE_X13Y153_BQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y154_SLICE_X14Y154_CO5),
.O6(CLBLM_R_X11Y154_SLICE_X14Y154_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0020000022220000)
  ) CLBLM_R_X11Y154_SLICE_X14Y154_BLUT (
.I0(CLBLM_L_X10Y153_SLICE_X13Y153_BQ),
.I1(CLBLM_L_X10Y153_SLICE_X13Y153_CQ),
.I2(CLBLM_R_X11Y153_SLICE_X15Y153_CO6),
.I3(CLBLM_L_X10Y154_SLICE_X13Y154_AQ),
.I4(CLBLM_R_X11Y154_SLICE_X15Y154_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y154_SLICE_X14Y154_BO5),
.O6(CLBLM_R_X11Y154_SLICE_X14Y154_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000aaaafc30)
  ) CLBLM_R_X11Y154_SLICE_X14Y154_ALUT (
.I0(CLBLM_R_X5Y152_SLICE_X7Y152_B5Q),
.I1(CLBLM_R_X11Y153_SLICE_X15Y153_CO6),
.I2(CLBLM_R_X11Y154_SLICE_X14Y154_AQ),
.I3(CLBLM_R_X11Y154_SLICE_X15Y154_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y121_IOB_X1Y121_I),
.O5(CLBLM_R_X11Y154_SLICE_X14Y154_AO5),
.O6(CLBLM_R_X11Y154_SLICE_X14Y154_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y154_SLICE_X15Y154_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y154_SLICE_X15Y154_AO6),
.Q(CLBLM_R_X11Y154_SLICE_X15Y154_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y154_SLICE_X15Y154_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y154_SLICE_X15Y154_BO6),
.Q(CLBLM_R_X11Y154_SLICE_X15Y154_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h77ffdd77575f5d57)
  ) CLBLM_R_X11Y154_SLICE_X15Y154_DLUT (
.I0(CLBLM_R_X11Y153_SLICE_X15Y153_CO5),
.I1(CLBLM_R_X11Y154_SLICE_X14Y154_AQ),
.I2(CLBLM_R_X11Y154_SLICE_X14Y154_BO5),
.I3(CLBLM_R_X11Y154_SLICE_X15Y154_BQ),
.I4(CLBLM_R_X11Y154_SLICE_X15Y154_AQ),
.I5(CLBLM_L_X10Y154_SLICE_X13Y154_AQ),
.O5(CLBLM_R_X11Y154_SLICE_X15Y154_DO5),
.O6(CLBLM_R_X11Y154_SLICE_X15Y154_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000355555554)
  ) CLBLM_R_X11Y154_SLICE_X15Y154_CLUT (
.I0(CLBLM_R_X11Y153_SLICE_X15Y153_CO5),
.I1(CLBLM_R_X11Y154_SLICE_X14Y154_AQ),
.I2(CLBLM_L_X10Y153_SLICE_X13Y153_BQ),
.I3(CLBLM_R_X11Y154_SLICE_X15Y154_BQ),
.I4(CLBLM_R_X11Y154_SLICE_X15Y154_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y154_SLICE_X15Y154_CO5),
.O6(CLBLM_R_X11Y154_SLICE_X15Y154_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0bbf000f099f000)
  ) CLBLM_R_X11Y154_SLICE_X15Y154_BLUT (
.I0(CLBLM_R_X11Y154_SLICE_X15Y154_DO6),
.I1(CLBLM_R_X11Y154_SLICE_X15Y154_BQ),
.I2(CLBLM_R_X11Y151_SLICE_X15Y151_BQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(CLBLM_R_X11Y154_SLICE_X15Y154_CO6),
.O5(CLBLM_R_X11Y154_SLICE_X15Y154_BO5),
.O6(CLBLM_R_X11Y154_SLICE_X15Y154_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00000faf60a06)
  ) CLBLM_R_X11Y154_SLICE_X15Y154_ALUT (
.I0(CLBLM_R_X11Y154_SLICE_X15Y154_AQ),
.I1(CLBLM_R_X11Y153_SLICE_X15Y153_CO5),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X12Y154_SLICE_X16Y154_BO6),
.I4(CLBLM_L_X10Y153_SLICE_X12Y153_AQ),
.I5(RIOB33_X105Y121_IOB_X1Y121_I),
.O5(CLBLM_R_X11Y154_SLICE_X15Y154_AO5),
.O6(CLBLM_R_X11Y154_SLICE_X15Y154_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y157_SLICE_X14Y157_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y157_SLICE_X14Y157_DO5),
.O6(CLBLM_R_X11Y157_SLICE_X14Y157_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y157_SLICE_X14Y157_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y157_SLICE_X14Y157_CO5),
.O6(CLBLM_R_X11Y157_SLICE_X14Y157_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y157_SLICE_X14Y157_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y157_SLICE_X14Y157_BO5),
.O6(CLBLM_R_X11Y157_SLICE_X14Y157_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc0cfc0cff00ffff)
  ) CLBLM_R_X11Y157_SLICE_X14Y157_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y145_SLICE_X6Y145_DO5),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X11Y153_SLICE_X14Y153_CQ),
.I4(RIOB33_X105Y143_IOB_X1Y143_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y157_SLICE_X14Y157_AO5),
.O6(CLBLM_R_X11Y157_SLICE_X14Y157_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y157_SLICE_X15Y157_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y157_SLICE_X15Y157_DO5),
.O6(CLBLM_R_X11Y157_SLICE_X15Y157_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y157_SLICE_X15Y157_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y157_SLICE_X15Y157_CO5),
.O6(CLBLM_R_X11Y157_SLICE_X15Y157_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y157_SLICE_X15Y157_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y157_SLICE_X15Y157_BO5),
.O6(CLBLM_R_X11Y157_SLICE_X15Y157_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y157_SLICE_X15Y157_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y157_SLICE_X15Y157_AO5),
.O6(CLBLM_R_X11Y157_SLICE_X15Y157_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y151_SLICE_X18Y151_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y151_SLICE_X18Y151_DO5),
.O6(CLBLM_R_X13Y151_SLICE_X18Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff7fffffff7fffff)
  ) CLBLM_R_X13Y151_SLICE_X18Y151_CLUT (
.I0(CLBLM_L_X12Y154_SLICE_X16Y154_AQ),
.I1(CLBLM_L_X12Y152_SLICE_X17Y152_BQ),
.I2(CLBLM_L_X12Y152_SLICE_X16Y152_AQ),
.I3(CLBLM_L_X12Y153_SLICE_X17Y153_CO6),
.I4(CLBLM_L_X12Y153_SLICE_X16Y153_AQ),
.I5(1'b1),
.O5(CLBLM_R_X13Y151_SLICE_X18Y151_CO5),
.O6(CLBLM_R_X13Y151_SLICE_X18Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hbfffffffffffffff)
  ) CLBLM_R_X13Y151_SLICE_X18Y151_BLUT (
.I0(CLBLM_L_X12Y154_SLICE_X16Y154_BO5),
.I1(CLBLM_L_X12Y152_SLICE_X16Y152_BQ),
.I2(CLBLM_R_X11Y153_SLICE_X15Y153_AQ),
.I3(CLBLM_L_X12Y153_SLICE_X16Y153_AQ),
.I4(CLBLM_L_X12Y154_SLICE_X16Y154_AQ),
.I5(CLBLM_R_X11Y152_SLICE_X15Y152_AQ),
.O5(CLBLM_R_X13Y151_SLICE_X18Y151_BO5),
.O6(CLBLM_R_X13Y151_SLICE_X18Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffd)
  ) CLBLM_R_X13Y151_SLICE_X18Y151_ALUT (
.I0(CLBLM_L_X12Y154_SLICE_X16Y154_BO5),
.I1(CLBLM_L_X12Y152_SLICE_X16Y152_BQ),
.I2(CLBLM_R_X11Y153_SLICE_X15Y153_AQ),
.I3(CLBLM_L_X12Y153_SLICE_X16Y153_AQ),
.I4(CLBLM_L_X12Y154_SLICE_X16Y154_AQ),
.I5(CLBLM_R_X11Y152_SLICE_X15Y152_AQ),
.O5(CLBLM_R_X13Y151_SLICE_X18Y151_AO5),
.O6(CLBLM_R_X13Y151_SLICE_X18Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y151_SLICE_X19Y151_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y151_SLICE_X19Y151_DO5),
.O6(CLBLM_R_X13Y151_SLICE_X19Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y151_SLICE_X19Y151_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y151_SLICE_X19Y151_CO5),
.O6(CLBLM_R_X13Y151_SLICE_X19Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y151_SLICE_X19Y151_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y151_SLICE_X19Y151_BO5),
.O6(CLBLM_R_X13Y151_SLICE_X19Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y151_SLICE_X19Y151_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y151_SLICE_X19Y151_AO5),
.O6(CLBLM_R_X13Y151_SLICE_X19Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y152_SLICE_X18Y152_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y152_SLICE_X18Y152_DO5),
.O6(CLBLM_R_X13Y152_SLICE_X18Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y152_SLICE_X18Y152_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y152_SLICE_X18Y152_CO5),
.O6(CLBLM_R_X13Y152_SLICE_X18Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000080000000)
  ) CLBLM_R_X13Y152_SLICE_X18Y152_BLUT (
.I0(CLBLM_L_X12Y153_SLICE_X16Y153_AQ),
.I1(CLBLM_L_X12Y152_SLICE_X17Y152_CQ),
.I2(CLBLM_L_X12Y154_SLICE_X16Y154_AQ),
.I3(CLBLM_L_X12Y152_SLICE_X16Y152_AQ),
.I4(CLBLM_L_X12Y152_SLICE_X17Y152_BQ),
.I5(CLBLM_L_X12Y153_SLICE_X17Y153_CO6),
.O5(CLBLM_R_X13Y152_SLICE_X18Y152_BO5),
.O6(CLBLM_R_X13Y152_SLICE_X18Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000001)
  ) CLBLM_R_X13Y152_SLICE_X18Y152_ALUT (
.I0(CLBLM_L_X12Y153_SLICE_X17Y153_DO6),
.I1(CLBLM_L_X12Y152_SLICE_X17Y152_CQ),
.I2(CLBLM_L_X12Y154_SLICE_X16Y154_AQ),
.I3(CLBLM_L_X12Y152_SLICE_X16Y152_AQ),
.I4(CLBLM_L_X12Y153_SLICE_X16Y153_AQ),
.I5(CLBLM_L_X12Y152_SLICE_X17Y152_BQ),
.O5(CLBLM_R_X13Y152_SLICE_X18Y152_AO5),
.O6(CLBLM_R_X13Y152_SLICE_X18Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y152_SLICE_X19Y152_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y152_SLICE_X19Y152_DO5),
.O6(CLBLM_R_X13Y152_SLICE_X19Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y152_SLICE_X19Y152_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y152_SLICE_X19Y152_CO5),
.O6(CLBLM_R_X13Y152_SLICE_X19Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y152_SLICE_X19Y152_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y152_SLICE_X19Y152_BO5),
.O6(CLBLM_R_X13Y152_SLICE_X19Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y152_SLICE_X19Y152_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y152_SLICE_X19Y152_AO5),
.O6(CLBLM_R_X13Y152_SLICE_X19Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X15Y151_SLICE_X20Y151_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X15Y153_SLICE_X20Y153_AO5),
.Q(CLBLM_R_X15Y151_SLICE_X20Y151_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y151_SLICE_X20Y151_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y151_SLICE_X20Y151_DO5),
.O6(CLBLM_R_X15Y151_SLICE_X20Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y151_SLICE_X20Y151_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y151_SLICE_X20Y151_CO5),
.O6(CLBLM_R_X15Y151_SLICE_X20Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y151_SLICE_X20Y151_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y151_SLICE_X20Y151_BO5),
.O6(CLBLM_R_X15Y151_SLICE_X20Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y151_SLICE_X20Y151_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y151_SLICE_X20Y151_AO5),
.O6(CLBLM_R_X15Y151_SLICE_X20Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y151_SLICE_X21Y151_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y151_SLICE_X21Y151_DO5),
.O6(CLBLM_R_X15Y151_SLICE_X21Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y151_SLICE_X21Y151_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y151_SLICE_X21Y151_CO5),
.O6(CLBLM_R_X15Y151_SLICE_X21Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y151_SLICE_X21Y151_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y151_SLICE_X21Y151_BO5),
.O6(CLBLM_R_X15Y151_SLICE_X21Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y151_SLICE_X21Y151_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y151_SLICE_X21Y151_AO5),
.O6(CLBLM_R_X15Y151_SLICE_X21Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y153_SLICE_X20Y153_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y153_SLICE_X20Y153_DO5),
.O6(CLBLM_R_X15Y153_SLICE_X20Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y153_SLICE_X20Y153_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y153_SLICE_X20Y153_CO5),
.O6(CLBLM_R_X15Y153_SLICE_X20Y153_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y153_SLICE_X20Y153_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y153_SLICE_X20Y153_BO5),
.O6(CLBLM_R_X15Y153_SLICE_X20Y153_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff00fffcfc3030)
  ) CLBLM_R_X15Y153_SLICE_X20Y153_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y150_SLICE_X12Y150_C5Q),
.I3(RIOB33_X105Y143_IOB_X1Y143_I),
.I4(CLBLM_R_X11Y153_SLICE_X14Y153_AQ),
.I5(1'b1),
.O5(CLBLM_R_X15Y153_SLICE_X20Y153_AO5),
.O6(CLBLM_R_X15Y153_SLICE_X20Y153_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y153_SLICE_X21Y153_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y153_SLICE_X21Y153_DO5),
.O6(CLBLM_R_X15Y153_SLICE_X21Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y153_SLICE_X21Y153_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y153_SLICE_X21Y153_CO5),
.O6(CLBLM_R_X15Y153_SLICE_X21Y153_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y153_SLICE_X21Y153_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y153_SLICE_X21Y153_BO5),
.O6(CLBLM_R_X15Y153_SLICE_X21Y153_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X15Y153_SLICE_X21Y153_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X15Y153_SLICE_X21Y153_AO5),
.O6(CLBLM_R_X15Y153_SLICE_X21Y153_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y141_SLICE_X162Y141_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y141_SLICE_X162Y141_DO5),
.O6(CLBLM_R_X103Y141_SLICE_X162Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y141_SLICE_X162Y141_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y141_SLICE_X162Y141_CO5),
.O6(CLBLM_R_X103Y141_SLICE_X162Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y141_SLICE_X162Y141_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y141_SLICE_X162Y141_BO5),
.O6(CLBLM_R_X103Y141_SLICE_X162Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y141_SLICE_X162Y141_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y141_SLICE_X162Y141_AO5),
.O6(CLBLM_R_X103Y141_SLICE_X162Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y141_SLICE_X163Y141_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y141_SLICE_X163Y141_DO5),
.O6(CLBLM_R_X103Y141_SLICE_X163Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y141_SLICE_X163Y141_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y141_SLICE_X163Y141_CO5),
.O6(CLBLM_R_X103Y141_SLICE_X163Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y141_SLICE_X163Y141_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y141_SLICE_X163Y141_BO5),
.O6(CLBLM_R_X103Y141_SLICE_X163Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha000a00088880000)
  ) CLBLM_R_X103Y141_SLICE_X163Y141_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(RIOB33_X105Y139_IOB_X1Y140_I),
.I2(RIOB33_X105Y139_IOB_X1Y139_I),
.I3(RIOB33_X105Y137_IOB_X1Y138_I),
.I4(RIOB33_X105Y141_IOB_X1Y141_I),
.I5(1'b1),
.O5(CLBLM_R_X103Y141_SLICE_X163Y141_AO5),
.O6(CLBLM_R_X103Y141_SLICE_X163Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y169_SLICE_X162Y169_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y169_SLICE_X162Y169_DO5),
.O6(CLBLM_R_X103Y169_SLICE_X162Y169_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y169_SLICE_X162Y169_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y169_SLICE_X162Y169_CO5),
.O6(CLBLM_R_X103Y169_SLICE_X162Y169_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y169_SLICE_X162Y169_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y169_SLICE_X162Y169_BO5),
.O6(CLBLM_R_X103Y169_SLICE_X162Y169_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y169_SLICE_X162Y169_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y169_SLICE_X162Y169_AO5),
.O6(CLBLM_R_X103Y169_SLICE_X162Y169_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y169_SLICE_X163Y169_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y169_SLICE_X163Y169_DO5),
.O6(CLBLM_R_X103Y169_SLICE_X163Y169_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y169_SLICE_X163Y169_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y169_SLICE_X163Y169_CO5),
.O6(CLBLM_R_X103Y169_SLICE_X163Y169_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y169_SLICE_X163Y169_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y169_SLICE_X163Y169_BO5),
.O6(CLBLM_R_X103Y169_SLICE_X163Y169_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcfcfcfcfcfcfcf)
  ) CLBLM_R_X103Y169_SLICE_X163Y169_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y151_SLICE_X14Y151_BQ),
.I2(RIOB33_X105Y143_IOB_X1Y143_I),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y169_SLICE_X163Y169_AO5),
.O6(CLBLM_R_X103Y169_SLICE_X163Y169_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y170_SLICE_X162Y170_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y170_SLICE_X162Y170_DO5),
.O6(CLBLM_R_X103Y170_SLICE_X162Y170_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y170_SLICE_X162Y170_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y170_SLICE_X162Y170_CO5),
.O6(CLBLM_R_X103Y170_SLICE_X162Y170_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y170_SLICE_X162Y170_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y170_SLICE_X162Y170_BO5),
.O6(CLBLM_R_X103Y170_SLICE_X162Y170_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y170_SLICE_X162Y170_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y170_SLICE_X162Y170_AO5),
.O6(CLBLM_R_X103Y170_SLICE_X162Y170_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y170_SLICE_X163Y170_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y170_SLICE_X163Y170_DO5),
.O6(CLBLM_R_X103Y170_SLICE_X163Y170_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y170_SLICE_X163Y170_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y170_SLICE_X163Y170_CO5),
.O6(CLBLM_R_X103Y170_SLICE_X163Y170_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y170_SLICE_X163Y170_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y170_SLICE_X163Y170_BO5),
.O6(CLBLM_R_X103Y170_SLICE_X163Y170_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ffffaaaaffff)
  ) CLBLM_R_X103Y170_SLICE_X163Y170_ALUT (
.I0(CLBLM_L_X12Y152_SLICE_X17Y152_AQ),
.I1(1'b1),
.I2(CLBLM_L_X10Y155_SLICE_X13Y155_AQ),
.I3(1'b1),
.I4(RIOB33_X105Y143_IOB_X1Y143_I),
.I5(1'b1),
.O5(CLBLM_R_X103Y170_SLICE_X163Y170_AO5),
.O6(CLBLM_R_X103Y170_SLICE_X163Y170_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y173_SLICE_X162Y173_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y173_SLICE_X162Y173_DO5),
.O6(CLBLM_R_X103Y173_SLICE_X162Y173_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y173_SLICE_X162Y173_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y173_SLICE_X162Y173_CO5),
.O6(CLBLM_R_X103Y173_SLICE_X162Y173_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y173_SLICE_X162Y173_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y173_SLICE_X162Y173_BO5),
.O6(CLBLM_R_X103Y173_SLICE_X162Y173_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y173_SLICE_X162Y173_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y173_SLICE_X162Y173_AO5),
.O6(CLBLM_R_X103Y173_SLICE_X162Y173_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y173_SLICE_X163Y173_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y173_SLICE_X163Y173_DO5),
.O6(CLBLM_R_X103Y173_SLICE_X163Y173_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y173_SLICE_X163Y173_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y173_SLICE_X163Y173_CO5),
.O6(CLBLM_R_X103Y173_SLICE_X163Y173_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y173_SLICE_X163Y173_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y173_SLICE_X163Y173_BO5),
.O6(CLBLM_R_X103Y173_SLICE_X163Y173_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccfffff0f0ffff)
  ) CLBLM_R_X103Y173_SLICE_X163Y173_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y149_SLICE_X12Y149_AQ),
.I2(CLBLM_R_X11Y151_SLICE_X15Y151_AQ),
.I3(1'b1),
.I4(RIOB33_X105Y143_IOB_X1Y143_I),
.I5(1'b1),
.O5(CLBLM_R_X103Y173_SLICE_X163Y173_AO5),
.O6(CLBLM_R_X103Y173_SLICE_X163Y173_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y176_SLICE_X162Y176_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y176_SLICE_X162Y176_DO5),
.O6(CLBLM_R_X103Y176_SLICE_X162Y176_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y176_SLICE_X162Y176_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y176_SLICE_X162Y176_CO5),
.O6(CLBLM_R_X103Y176_SLICE_X162Y176_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y176_SLICE_X162Y176_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y176_SLICE_X162Y176_BO5),
.O6(CLBLM_R_X103Y176_SLICE_X162Y176_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y176_SLICE_X162Y176_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y176_SLICE_X162Y176_AO5),
.O6(CLBLM_R_X103Y176_SLICE_X162Y176_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y176_SLICE_X163Y176_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y176_SLICE_X163Y176_DO5),
.O6(CLBLM_R_X103Y176_SLICE_X163Y176_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y176_SLICE_X163Y176_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y176_SLICE_X163Y176_CO5),
.O6(CLBLM_R_X103Y176_SLICE_X163Y176_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y176_SLICE_X163Y176_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y176_SLICE_X163Y176_BO5),
.O6(CLBLM_R_X103Y176_SLICE_X163Y176_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ffffff00ffff)
  ) CLBLM_R_X103Y176_SLICE_X163Y176_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_L_X12Y155_SLICE_X17Y155_AQ),
.I3(CLBLM_L_X12Y151_SLICE_X16Y151_AQ),
.I4(RIOB33_X105Y143_IOB_X1Y143_I),
.I5(1'b1),
.O5(CLBLM_R_X103Y176_SLICE_X163Y176_AO5),
.O6(CLBLM_R_X103Y176_SLICE_X163Y176_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y178_SLICE_X162Y178_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y178_SLICE_X162Y178_DO5),
.O6(CLBLM_R_X103Y178_SLICE_X162Y178_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y178_SLICE_X162Y178_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y178_SLICE_X162Y178_CO5),
.O6(CLBLM_R_X103Y178_SLICE_X162Y178_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y178_SLICE_X162Y178_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y178_SLICE_X162Y178_BO5),
.O6(CLBLM_R_X103Y178_SLICE_X162Y178_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y178_SLICE_X162Y178_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y178_SLICE_X162Y178_AO5),
.O6(CLBLM_R_X103Y178_SLICE_X162Y178_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y178_SLICE_X163Y178_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y178_SLICE_X163Y178_DO5),
.O6(CLBLM_R_X103Y178_SLICE_X163Y178_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y178_SLICE_X163Y178_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y178_SLICE_X163Y178_CO5),
.O6(CLBLM_R_X103Y178_SLICE_X163Y178_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y178_SLICE_X163Y178_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y178_SLICE_X163Y178_BO5),
.O6(CLBLM_R_X103Y178_SLICE_X163Y178_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ffffccccffff)
  ) CLBLM_R_X103Y178_SLICE_X163Y178_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y153_SLICE_X14Y153_BQ),
.I2(CLBLM_R_X11Y151_SLICE_X14Y151_AQ),
.I3(1'b1),
.I4(RIOB33_X105Y143_IOB_X1Y143_I),
.I5(1'b1),
.O5(CLBLM_R_X103Y178_SLICE_X163Y178_AO5),
.O6(CLBLM_R_X103Y178_SLICE_X163Y178_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFGCTRL" *)
  BUFGCTRL #(
    .INIT_OUT(0),
    .IS_CE0_INVERTED(0),
    .IS_CE1_INVERTED(1),
    .IS_IGNORE0_INVERTED(1),
    .IS_IGNORE1_INVERTED(0),
    .IS_S0_INVERTED(0),
    .IS_S1_INVERTED(1),
    .PRESELECT_I0("TRUE"),
    .PRESELECT_I1("FALSE")
  ) CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_BUFGCTRL (
.CE0(1'b1),
.CE1(1'b1),
.I0(LIOB33_X0Y77_IOB_X0Y78_I),
.I1(1'b1),
.IGNORE0(1'b1),
.IGNORE1(1'b1),
.O(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.S0(1'b1),
.S1(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFHCE" *)
  BUFHCE #(
    .CE_TYPE("SYNC"),
    .INIT_OUT(0),
    .IS_CE_INVERTED(0)
  ) CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_BUFHCE (
.CE(1'b1),
.I(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.O(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFHCE" *)
  BUFHCE #(
    .CE_TYPE("SYNC"),
    .INIT_OUT(0),
    .IS_CE_INVERTED(0)
  ) CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_BUFHCE (
.CE(1'b1),
.I(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.O(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y51_IOB_X0Y51_IBUF (
.I(LIOB33_X0Y51_IOB_X0Y51_IPAD),
.O(LIOB33_X0Y51_IOB_X0Y51_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y51_IOB_X0Y52_IBUF (
.I(LIOB33_X0Y51_IOB_X0Y52_IPAD),
.O(LIOB33_X0Y51_IOB_X0Y52_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y53_IOB_X0Y53_IBUF (
.I(LIOB33_X0Y53_IOB_X0Y53_IPAD),
.O(LIOB33_X0Y53_IOB_X0Y53_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y53_IOB_X0Y54_IBUF (
.I(LIOB33_X0Y53_IOB_X0Y54_IPAD),
.O(LIOB33_X0Y53_IOB_X0Y54_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y55_IOB_X0Y55_IBUF (
.I(LIOB33_X0Y55_IOB_X0Y55_IPAD),
.O(LIOB33_X0Y55_IOB_X0Y55_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y55_IOB_X0Y56_IBUF (
.I(LIOB33_X0Y55_IOB_X0Y56_IPAD),
.O(LIOB33_X0Y55_IOB_X0Y56_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y57_IOB_X0Y57_IBUF (
.I(LIOB33_X0Y57_IOB_X0Y57_IPAD),
.O(LIOB33_X0Y57_IOB_X0Y57_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y57_IOB_X0Y58_IBUF (
.I(LIOB33_X0Y57_IOB_X0Y58_IPAD),
.O(LIOB33_X0Y57_IOB_X0Y58_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y59_IOB_X0Y59_IBUF (
.I(LIOB33_X0Y59_IOB_X0Y59_IPAD),
.O(LIOB33_X0Y59_IOB_X0Y59_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y59_IOB_X0Y60_IBUF (
.I(LIOB33_X0Y59_IOB_X0Y60_IPAD),
.O(LIOB33_X0Y59_IOB_X0Y60_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y61_IOB_X0Y61_IBUF (
.I(LIOB33_X0Y61_IOB_X0Y61_IPAD),
.O(LIOB33_X0Y61_IOB_X0Y61_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y61_IOB_X0Y62_IBUF (
.I(LIOB33_X0Y61_IOB_X0Y62_IPAD),
.O(LIOB33_X0Y61_IOB_X0Y62_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y63_IOB_X0Y63_IBUF (
.I(LIOB33_X0Y63_IOB_X0Y63_IPAD),
.O(LIOB33_X0Y63_IOB_X0Y63_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y63_IOB_X0Y64_IBUF (
.I(LIOB33_X0Y63_IOB_X0Y64_IPAD),
.O(LIOB33_X0Y63_IOB_X0Y64_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y65_IOB_X0Y65_IBUF (
.I(LIOB33_X0Y65_IOB_X0Y65_IPAD),
.O(LIOB33_X0Y65_IOB_X0Y65_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y65_IOB_X0Y66_IBUF (
.I(LIOB33_X0Y65_IOB_X0Y66_IPAD),
.O(LIOB33_X0Y65_IOB_X0Y66_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y67_IOB_X0Y67_IBUF (
.I(LIOB33_X0Y67_IOB_X0Y67_IPAD),
.O(LIOB33_X0Y67_IOB_X0Y67_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y67_IOB_X0Y68_IBUF (
.I(LIOB33_X0Y67_IOB_X0Y68_IPAD),
.O(LIOB33_X0Y67_IOB_X0Y68_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y69_IOB_X0Y69_IBUF (
.I(LIOB33_X0Y69_IOB_X0Y69_IPAD),
.O(LIOB33_X0Y69_IOB_X0Y69_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y69_IOB_X0Y70_IBUF (
.I(LIOB33_X0Y69_IOB_X0Y70_IPAD),
.O(LIOB33_X0Y69_IOB_X0Y70_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y71_IOB_X0Y71_IBUF (
.I(LIOB33_X0Y71_IOB_X0Y71_IPAD),
.O(LIOB33_X0Y71_IOB_X0Y71_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y71_IOB_X0Y72_IBUF (
.I(LIOB33_X0Y71_IOB_X0Y72_IPAD),
.O(LIOB33_X0Y71_IOB_X0Y72_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y73_IOB_X0Y73_IBUF (
.I(LIOB33_X0Y73_IOB_X0Y73_IPAD),
.O(LIOB33_X0Y73_IOB_X0Y73_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y73_IOB_X0Y74_IBUF (
.I(LIOB33_X0Y73_IOB_X0Y74_IPAD),
.O(LIOB33_X0Y73_IOB_X0Y74_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y75_IOB_X0Y75_IBUF (
.I(LIOB33_X0Y75_IOB_X0Y75_IPAD),
.O(LIOB33_X0Y75_IOB_X0Y75_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y75_IOB_X0Y76_IBUF (
.I(LIOB33_X0Y75_IOB_X0Y76_IPAD),
.O(LIOB33_X0Y75_IOB_X0Y76_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y77_IOB_X0Y77_IBUF (
.I(LIOB33_X0Y77_IOB_X0Y77_IPAD),
.O(LIOB33_X0Y77_IOB_X0Y77_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y77_IOB_X0Y78_IBUF (
.I(LIOB33_X0Y77_IOB_X0Y78_IPAD),
.O(LIOB33_X0Y77_IOB_X0Y78_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y79_IOB_X0Y79_IBUF (
.I(LIOB33_X0Y79_IOB_X0Y79_IPAD),
.O(LIOB33_X0Y79_IOB_X0Y79_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y79_IOB_X0Y80_OBUF (
.I(CLBLL_L_X2Y138_SLICE_X0Y138_AO6),
.O(LIOB33_X0Y79_IOB_X0Y80_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y101_IOB_X0Y101_OBUF (
.I(CLBLL_L_X2Y138_SLICE_X0Y138_BO6),
.O(LIOB33_X0Y101_IOB_X0Y101_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y101_IOB_X0Y102_OBUF (
.I(CLBLL_L_X2Y138_SLICE_X0Y138_BO5),
.O(LIOB33_X0Y101_IOB_X0Y102_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y103_IOB_X0Y103_OBUF (
.I(CLBLL_L_X2Y141_SLICE_X0Y141_AO6),
.O(LIOB33_X0Y103_IOB_X0Y103_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y103_IOB_X0Y104_OBUF (
.I(CLBLL_L_X2Y141_SLICE_X0Y141_AO5),
.O(LIOB33_X0Y103_IOB_X0Y104_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y105_IOB_X0Y105_OBUF (
.I(CLBLL_L_X2Y138_SLICE_X0Y138_CO6),
.O(LIOB33_X0Y105_IOB_X0Y105_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y105_IOB_X0Y106_OBUF (
.I(CLBLL_L_X2Y138_SLICE_X0Y138_CO5),
.O(LIOB33_X0Y105_IOB_X0Y106_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y107_IOB_X0Y107_OBUF (
.I(CLBLL_L_X2Y120_SLICE_X0Y120_AO6),
.O(LIOB33_X0Y107_IOB_X0Y107_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y107_IOB_X0Y108_OBUF (
.I(CLBLM_R_X3Y152_SLICE_X2Y152_BO6),
.O(LIOB33_X0Y107_IOB_X0Y108_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y109_IOB_X0Y109_OBUF (
.I(CLBLL_L_X2Y134_SLICE_X0Y134_AO6),
.O(LIOB33_X0Y109_IOB_X0Y109_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y109_IOB_X0Y110_OBUF (
.I(CLBLL_L_X2Y134_SLICE_X0Y134_AO5),
.O(LIOB33_X0Y109_IOB_X0Y110_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y111_IOB_X0Y111_OBUF (
.I(1'b0),
.O(LIOB33_X0Y111_IOB_X0Y111_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y111_IOB_X0Y112_OBUF (
.I(CLBLM_R_X11Y148_SLICE_X15Y148_B5Q),
.O(LIOB33_X0Y111_IOB_X0Y112_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y113_IOB_X0Y113_OBUF (
.I(RIOB33_X105Y121_IOB_X1Y121_I),
.O(LIOB33_X0Y113_IOB_X0Y113_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y113_IOB_X0Y114_OBUF (
.I(CLBLM_R_X7Y143_SLICE_X8Y143_BQ),
.O(LIOB33_X0Y113_IOB_X0Y114_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y115_IOB_X0Y115_OBUF (
.I(CLBLM_R_X11Y148_SLICE_X15Y148_BQ),
.O(LIOB33_X0Y115_IOB_X0Y115_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y115_IOB_X0Y116_OBUF (
.I(CLBLM_L_X8Y142_SLICE_X10Y142_AQ),
.O(LIOB33_X0Y115_IOB_X0Y116_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y117_IOB_X0Y117_OBUF (
.I(CLBLM_R_X3Y144_SLICE_X2Y144_B5Q),
.O(LIOB33_X0Y117_IOB_X0Y117_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y117_IOB_X0Y118_OBUF (
.I(CLBLM_R_X3Y147_SLICE_X3Y147_CQ),
.O(LIOB33_X0Y117_IOB_X0Y118_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y119_IOB_X0Y119_OBUF (
.I(CLBLM_L_X10Y146_SLICE_X13Y146_BQ),
.O(LIOB33_X0Y119_IOB_X0Y119_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y119_IOB_X0Y120_OBUF (
.I(CLBLM_L_X10Y145_SLICE_X13Y145_AQ),
.O(LIOB33_X0Y119_IOB_X0Y120_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y121_IOB_X0Y121_OBUF (
.I(CLBLM_L_X8Y142_SLICE_X10Y142_A5Q),
.O(LIOB33_X0Y121_IOB_X0Y121_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y121_IOB_X0Y122_OBUF (
.I(CLBLM_R_X3Y144_SLICE_X2Y144_BQ),
.O(LIOB33_X0Y121_IOB_X0Y122_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y123_IOB_X0Y123_OBUF (
.I(CLBLM_R_X7Y143_SLICE_X8Y143_B5Q),
.O(LIOB33_X0Y123_IOB_X0Y123_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y123_IOB_X0Y124_OBUF (
.I(CLBLM_R_X3Y147_SLICE_X3Y147_C5Q),
.O(LIOB33_X0Y123_IOB_X0Y124_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y125_IOB_X0Y125_OBUF (
.I(CLBLM_L_X8Y145_SLICE_X11Y145_B5Q),
.O(LIOB33_X0Y125_IOB_X0Y125_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y125_IOB_X0Y126_OBUF (
.I(CLBLM_R_X3Y143_SLICE_X2Y143_BQ),
.O(LIOB33_X0Y125_IOB_X0Y126_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y127_IOB_X0Y127_OBUF (
.I(CLBLL_L_X4Y147_SLICE_X5Y147_CQ),
.O(LIOB33_X0Y127_IOB_X0Y127_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y127_IOB_X0Y128_OBUF (
.I(CLBLL_L_X2Y147_SLICE_X1Y147_AQ),
.O(LIOB33_X0Y127_IOB_X0Y128_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y129_IOB_X0Y129_OBUF (
.I(CLBLM_R_X3Y148_SLICE_X3Y148_AQ),
.O(LIOB33_X0Y129_IOB_X0Y129_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y129_IOB_X0Y130_OBUF (
.I(CLBLL_L_X52Y126_SLICE_X78Y126_AO6),
.O(LIOB33_X0Y129_IOB_X0Y130_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y131_IOB_X0Y131_OBUF (
.I(CLBLM_R_X7Y142_SLICE_X8Y142_AO5),
.O(LIOB33_X0Y131_IOB_X0Y131_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y131_IOB_X0Y132_OBUF (
.I(CLBLM_R_X5Y142_SLICE_X7Y142_AQ),
.O(LIOB33_X0Y131_IOB_X0Y132_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y133_IOB_X0Y133_OBUF (
.I(CLBLM_R_X3Y143_SLICE_X3Y143_A5Q),
.O(LIOB33_X0Y133_IOB_X0Y133_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y133_IOB_X0Y134_OBUF (
.I(CLBLM_R_X3Y143_SLICE_X2Y143_CQ),
.O(LIOB33_X0Y133_IOB_X0Y134_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y135_IOB_X0Y135_OBUF (
.I(CLBLM_R_X3Y142_SLICE_X2Y142_BQ),
.O(LIOB33_X0Y135_IOB_X0Y135_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y135_IOB_X0Y136_OBUF (
.I(CLBLL_L_X2Y145_SLICE_X1Y145_AQ),
.O(LIOB33_X0Y135_IOB_X0Y136_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y137_IOB_X0Y137_OBUF (
.I(CLBLM_R_X3Y142_SLICE_X2Y142_AQ),
.O(LIOB33_X0Y137_IOB_X0Y137_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y137_IOB_X0Y138_OBUF (
.I(CLBLM_R_X3Y143_SLICE_X3Y143_BQ),
.O(LIOB33_X0Y137_IOB_X0Y138_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y139_IOB_X0Y139_OBUF (
.I(CLBLM_R_X3Y143_SLICE_X3Y143_AQ),
.O(LIOB33_X0Y139_IOB_X0Y139_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y139_IOB_X0Y140_OBUF (
.I(CLBLM_R_X3Y142_SLICE_X2Y142_CQ),
.O(LIOB33_X0Y139_IOB_X0Y140_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y141_IOB_X0Y141_OBUF (
.I(CLBLM_R_X3Y143_SLICE_X2Y143_AQ),
.O(LIOB33_X0Y141_IOB_X0Y141_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y141_IOB_X0Y142_OBUF (
.I(LIOB33_X0Y53_IOB_X0Y54_I),
.O(LIOB33_X0Y141_IOB_X0Y142_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y143_IOB_X0Y143_OBUF (
.I(LIOB33_X0Y55_IOB_X0Y55_I),
.O(LIOB33_X0Y143_IOB_X0Y143_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y145_IOB_X0Y145_OBUF (
.I(LIOB33_X0Y57_IOB_X0Y58_I),
.O(LIOB33_X0Y145_IOB_X0Y145_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y145_IOB_X0Y146_OBUF (
.I(LIOB33_X0Y59_IOB_X0Y59_I),
.O(LIOB33_X0Y145_IOB_X0Y146_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y147_IOB_X0Y147_OBUF (
.I(LIOB33_X0Y71_IOB_X0Y71_I),
.O(LIOB33_X0Y147_IOB_X0Y147_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y147_IOB_X0Y148_OBUF (
.I(LIOB33_X0Y61_IOB_X0Y61_I),
.O(LIOB33_X0Y147_IOB_X0Y148_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y151_IOB_X0Y151_OBUF (
.I(LIOB33_X0Y65_IOB_X0Y65_I),
.O(LIOB33_X0Y151_IOB_X0Y151_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y151_IOB_X0Y152_OBUF (
.I(LIOB33_X0Y65_IOB_X0Y66_I),
.O(LIOB33_X0Y151_IOB_X0Y152_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y153_IOB_X0Y153_OBUF (
.I(LIOB33_X0Y67_IOB_X0Y67_I),
.O(LIOB33_X0Y153_IOB_X0Y153_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y153_IOB_X0Y154_OBUF (
.I(LIOB33_X0Y67_IOB_X0Y68_I),
.O(LIOB33_X0Y153_IOB_X0Y154_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y155_IOB_X0Y155_OBUF (
.I(LIOB33_X0Y69_IOB_X0Y70_I),
.O(LIOB33_X0Y155_IOB_X0Y155_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y155_IOB_X0Y156_OBUF (
.I(RIOB33_X105Y105_IOB_X1Y106_I),
.O(LIOB33_X0Y155_IOB_X0Y156_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y157_IOB_X0Y157_OBUF (
.I(RIOB33_X105Y115_IOB_X1Y115_I),
.O(LIOB33_X0Y157_IOB_X0Y157_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y157_IOB_X0Y158_OBUF (
.I(RIOB33_X105Y115_IOB_X1Y116_I),
.O(LIOB33_X0Y157_IOB_X0Y158_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y159_IOB_X0Y159_OBUF (
.I(RIOB33_X105Y117_IOB_X1Y117_I),
.O(LIOB33_X0Y159_IOB_X0Y159_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y159_IOB_X0Y160_OBUF (
.I(RIOB33_X105Y107_IOB_X1Y107_I),
.O(LIOB33_X0Y159_IOB_X0Y160_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y161_IOB_X0Y161_OBUF (
.I(RIOB33_X105Y107_IOB_X1Y108_I),
.O(LIOB33_X0Y161_IOB_X0Y161_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y161_IOB_X0Y162_OBUF (
.I(RIOB33_X105Y109_IOB_X1Y109_I),
.O(LIOB33_X0Y161_IOB_X0Y162_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y163_IOB_X0Y163_OBUF (
.I(RIOB33_X105Y109_IOB_X1Y110_I),
.O(LIOB33_X0Y163_IOB_X0Y163_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y163_IOB_X0Y164_OBUF (
.I(RIOB33_X105Y111_IOB_X1Y111_I),
.O(LIOB33_X0Y163_IOB_X0Y164_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y165_IOB_X0Y165_OBUF (
.I(RIOB33_X105Y111_IOB_X1Y112_I),
.O(LIOB33_X0Y165_IOB_X0Y165_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y165_IOB_X0Y166_OBUF (
.I(RIOB33_X105Y113_IOB_X1Y113_I),
.O(LIOB33_X0Y165_IOB_X0Y166_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y167_IOB_X0Y167_OBUF (
.I(RIOB33_X105Y113_IOB_X1Y114_I),
.O(LIOB33_X0Y167_IOB_X0Y167_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y167_IOB_X0Y168_OBUF (
.I(RIOB33_X105Y123_IOB_X1Y123_I),
.O(LIOB33_X0Y167_IOB_X0Y168_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y169_IOB_X0Y169_OBUF (
.I(RIOB33_X105Y121_IOB_X1Y122_I),
.O(LIOB33_X0Y169_IOB_X0Y169_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y169_IOB_X0Y170_OBUF (
.I(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.O(LIOB33_X0Y169_IOB_X0Y170_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y171_IOB_X0Y171_OBUF (
.I(LIOB33_SING_X0Y50_IOB_X0Y50_I),
.O(LIOB33_X0Y171_IOB_X0Y171_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y171_IOB_X0Y172_OBUF (
.I(CLBLM_R_X103Y141_SLICE_X163Y141_AO6),
.O(LIOB33_X0Y171_IOB_X0Y172_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y173_IOB_X0Y173_OBUF (
.I(CLBLM_R_X103Y141_SLICE_X163Y141_AO5),
.O(LIOB33_X0Y173_IOB_X0Y173_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y173_IOB_X0Y174_OBUF (
.I(CLBLM_L_X8Y159_SLICE_X10Y159_AO6),
.O(LIOB33_X0Y173_IOB_X0Y174_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y175_IOB_X0Y175_OBUF (
.I(RIOB33_X105Y127_IOB_X1Y127_I),
.O(LIOB33_X0Y175_IOB_X0Y175_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y175_IOB_X0Y176_OBUF (
.I(RIOB33_X105Y127_IOB_X1Y128_I),
.O(LIOB33_X0Y175_IOB_X0Y176_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y177_IOB_X0Y177_OBUF (
.I(RIOB33_X105Y129_IOB_X1Y129_I),
.O(LIOB33_X0Y177_IOB_X0Y177_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y177_IOB_X0Y178_OBUF (
.I(RIOB33_X105Y129_IOB_X1Y130_I),
.O(LIOB33_X0Y177_IOB_X0Y178_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y179_IOB_X0Y179_OBUF (
.I(RIOB33_X105Y131_IOB_X1Y131_I),
.O(LIOB33_X0Y179_IOB_X0Y179_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y179_IOB_X0Y180_OBUF (
.I(RIOB33_X105Y131_IOB_X1Y132_I),
.O(LIOB33_X0Y179_IOB_X0Y180_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y181_IOB_X0Y181_OBUF (
.I(RIOB33_X105Y133_IOB_X1Y133_I),
.O(LIOB33_X0Y181_IOB_X0Y181_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y181_IOB_X0Y182_OBUF (
.I(RIOB33_X105Y133_IOB_X1Y134_I),
.O(LIOB33_X0Y181_IOB_X0Y182_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y183_IOB_X0Y183_OBUF (
.I(RIOB33_X105Y135_IOB_X1Y135_I),
.O(LIOB33_X0Y183_IOB_X0Y183_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y183_IOB_X0Y184_OBUF (
.I(RIOB33_X105Y135_IOB_X1Y136_I),
.O(LIOB33_X0Y183_IOB_X0Y184_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y185_IOB_X0Y185_OBUF (
.I(RIOB33_X105Y137_IOB_X1Y137_I),
.O(LIOB33_X0Y185_IOB_X0Y185_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y185_IOB_X0Y186_OBUF (
.I(RIOB33_X105Y143_IOB_X1Y143_I),
.O(LIOB33_X0Y185_IOB_X0Y186_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y187_IOB_X0Y187_OBUF (
.I(RIOB33_X105Y143_IOB_X1Y144_I),
.O(LIOB33_X0Y187_IOB_X0Y187_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y187_IOB_X0Y188_OBUF (
.I(RIOB33_X105Y145_IOB_X1Y145_I),
.O(LIOB33_X0Y187_IOB_X0Y188_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y189_IOB_X0Y189_OBUF (
.I(RIOB33_X105Y145_IOB_X1Y146_I),
.O(LIOB33_X0Y189_IOB_X0Y189_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y189_IOB_X0Y190_OBUF (
.I(RIOB33_X105Y147_IOB_X1Y147_I),
.O(LIOB33_X0Y189_IOB_X0Y190_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y191_IOB_X0Y191_OBUF (
.I(RIOB33_X105Y147_IOB_X1Y148_I),
.O(LIOB33_X0Y191_IOB_X0Y191_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y191_IOB_X0Y192_OBUF (
.I(LIOB33_X0Y51_IOB_X0Y52_I),
.O(LIOB33_X0Y191_IOB_X0Y192_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y193_IOB_X0Y193_OBUF (
.I(LIOB33_X0Y55_IOB_X0Y56_I),
.O(LIOB33_X0Y193_IOB_X0Y193_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y193_IOB_X0Y194_OBUF (
.I(LIOB33_X0Y59_IOB_X0Y60_I),
.O(LIOB33_X0Y193_IOB_X0Y194_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y195_IOB_X0Y195_OBUF (
.I(LIOB33_X0Y63_IOB_X0Y64_I),
.O(LIOB33_X0Y195_IOB_X0Y195_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y195_IOB_X0Y196_OBUF (
.I(LIOB33_X0Y69_IOB_X0Y69_I),
.O(LIOB33_X0Y195_IOB_X0Y196_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y197_IOB_X0Y197_OBUF (
.I(LIOB33_X0Y71_IOB_X0Y72_I),
.O(LIOB33_X0Y197_IOB_X0Y197_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y197_IOB_X0Y198_OBUF (
.I(LIOB33_X0Y73_IOB_X0Y73_I),
.O(LIOB33_X0Y197_IOB_X0Y198_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_SING_X0Y50_IOB_X0Y50_IBUF (
.I(LIOB33_SING_X0Y50_IOB_X0Y50_IPAD),
.O(LIOB33_SING_X0Y50_IOB_X0Y50_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y100_IOB_X0Y100_OBUF (
.I(CLBLL_L_X2Y138_SLICE_X0Y138_AO5),
.O(LIOB33_SING_X0Y100_IOB_X0Y100_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y149_IOB_X0Y149_OBUF (
.I(LIOB33_X0Y61_IOB_X0Y62_I),
.O(LIOB33_SING_X0Y149_IOB_X0Y149_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y150_IOB_X0Y150_OBUF (
.I(LIOB33_X0Y63_IOB_X0Y63_I),
.O(LIOB33_SING_X0Y150_IOB_X0Y150_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y199_IOB_X0Y199_OBUF (
.I(LIOB33_X0Y73_IOB_X0Y74_I),
.O(LIOB33_SING_X0Y199_IOB_X0Y199_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y101_IOB_X1Y101_IBUF (
.I(RIOB33_X105Y101_IOB_X1Y101_IPAD),
.O(RIOB33_X105Y101_IOB_X1Y101_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y101_IOB_X1Y102_IBUF (
.I(RIOB33_X105Y101_IOB_X1Y102_IPAD),
.O(RIOB33_X105Y101_IOB_X1Y102_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y103_IOB_X1Y103_IBUF (
.I(RIOB33_X105Y103_IOB_X1Y103_IPAD),
.O(RIOB33_X105Y103_IOB_X1Y103_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y103_IOB_X1Y104_IBUF (
.I(RIOB33_X105Y103_IOB_X1Y104_IPAD),
.O(RIOB33_X105Y103_IOB_X1Y104_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y105_IOB_X1Y105_IBUF (
.I(RIOB33_X105Y105_IOB_X1Y105_IPAD),
.O(RIOB33_X105Y105_IOB_X1Y105_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y105_IOB_X1Y106_IBUF (
.I(RIOB33_X105Y105_IOB_X1Y106_IPAD),
.O(RIOB33_X105Y105_IOB_X1Y106_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y107_IOB_X1Y107_IBUF (
.I(RIOB33_X105Y107_IOB_X1Y107_IPAD),
.O(RIOB33_X105Y107_IOB_X1Y107_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y107_IOB_X1Y108_IBUF (
.I(RIOB33_X105Y107_IOB_X1Y108_IPAD),
.O(RIOB33_X105Y107_IOB_X1Y108_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y109_IOB_X1Y109_IBUF (
.I(RIOB33_X105Y109_IOB_X1Y109_IPAD),
.O(RIOB33_X105Y109_IOB_X1Y109_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y109_IOB_X1Y110_IBUF (
.I(RIOB33_X105Y109_IOB_X1Y110_IPAD),
.O(RIOB33_X105Y109_IOB_X1Y110_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y111_IOB_X1Y111_IBUF (
.I(RIOB33_X105Y111_IOB_X1Y111_IPAD),
.O(RIOB33_X105Y111_IOB_X1Y111_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y111_IOB_X1Y112_IBUF (
.I(RIOB33_X105Y111_IOB_X1Y112_IPAD),
.O(RIOB33_X105Y111_IOB_X1Y112_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y113_IOB_X1Y113_IBUF (
.I(RIOB33_X105Y113_IOB_X1Y113_IPAD),
.O(RIOB33_X105Y113_IOB_X1Y113_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y113_IOB_X1Y114_IBUF (
.I(RIOB33_X105Y113_IOB_X1Y114_IPAD),
.O(RIOB33_X105Y113_IOB_X1Y114_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y115_IOB_X1Y115_IBUF (
.I(RIOB33_X105Y115_IOB_X1Y115_IPAD),
.O(RIOB33_X105Y115_IOB_X1Y115_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y115_IOB_X1Y116_IBUF (
.I(RIOB33_X105Y115_IOB_X1Y116_IPAD),
.O(RIOB33_X105Y115_IOB_X1Y116_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y117_IOB_X1Y117_IBUF (
.I(RIOB33_X105Y117_IOB_X1Y117_IPAD),
.O(RIOB33_X105Y117_IOB_X1Y117_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y117_IOB_X1Y118_IBUF (
.I(RIOB33_X105Y117_IOB_X1Y118_IPAD),
.O(RIOB33_X105Y117_IOB_X1Y118_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y119_IOB_X1Y119_IBUF (
.I(RIOB33_X105Y119_IOB_X1Y119_IPAD),
.O(RIOB33_X105Y119_IOB_X1Y119_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y119_IOB_X1Y120_IBUF (
.I(RIOB33_X105Y119_IOB_X1Y120_IPAD),
.O(RIOB33_X105Y119_IOB_X1Y120_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y121_IOB_X1Y121_IBUF (
.I(RIOB33_X105Y121_IOB_X1Y121_IPAD),
.O(RIOB33_X105Y121_IOB_X1Y121_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y121_IOB_X1Y122_IBUF (
.I(RIOB33_X105Y121_IOB_X1Y122_IPAD),
.O(RIOB33_X105Y121_IOB_X1Y122_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y123_IOB_X1Y123_IBUF (
.I(RIOB33_X105Y123_IOB_X1Y123_IPAD),
.O(RIOB33_X105Y123_IOB_X1Y123_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y123_IOB_X1Y124_IBUF (
.I(RIOB33_X105Y123_IOB_X1Y124_IPAD),
.O(RIOB33_X105Y123_IOB_X1Y124_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y125_IOB_X1Y125_IBUF (
.I(RIOB33_X105Y125_IOB_X1Y125_IPAD),
.O(RIOB33_X105Y125_IOB_X1Y125_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y125_IOB_X1Y126_IBUF (
.I(RIOB33_X105Y125_IOB_X1Y126_IPAD),
.O(RIOB33_X105Y125_IOB_X1Y126_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y127_IOB_X1Y127_IBUF (
.I(RIOB33_X105Y127_IOB_X1Y127_IPAD),
.O(RIOB33_X105Y127_IOB_X1Y127_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y127_IOB_X1Y128_IBUF (
.I(RIOB33_X105Y127_IOB_X1Y128_IPAD),
.O(RIOB33_X105Y127_IOB_X1Y128_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y129_IOB_X1Y129_IBUF (
.I(RIOB33_X105Y129_IOB_X1Y129_IPAD),
.O(RIOB33_X105Y129_IOB_X1Y129_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y129_IOB_X1Y130_IBUF (
.I(RIOB33_X105Y129_IOB_X1Y130_IPAD),
.O(RIOB33_X105Y129_IOB_X1Y130_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y131_IOB_X1Y131_IBUF (
.I(RIOB33_X105Y131_IOB_X1Y131_IPAD),
.O(RIOB33_X105Y131_IOB_X1Y131_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y131_IOB_X1Y132_IBUF (
.I(RIOB33_X105Y131_IOB_X1Y132_IPAD),
.O(RIOB33_X105Y131_IOB_X1Y132_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y133_IOB_X1Y133_IBUF (
.I(RIOB33_X105Y133_IOB_X1Y133_IPAD),
.O(RIOB33_X105Y133_IOB_X1Y133_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y133_IOB_X1Y134_IBUF (
.I(RIOB33_X105Y133_IOB_X1Y134_IPAD),
.O(RIOB33_X105Y133_IOB_X1Y134_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y135_IOB_X1Y135_IBUF (
.I(RIOB33_X105Y135_IOB_X1Y135_IPAD),
.O(RIOB33_X105Y135_IOB_X1Y135_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y135_IOB_X1Y136_IBUF (
.I(RIOB33_X105Y135_IOB_X1Y136_IPAD),
.O(RIOB33_X105Y135_IOB_X1Y136_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y137_IOB_X1Y137_IBUF (
.I(RIOB33_X105Y137_IOB_X1Y137_IPAD),
.O(RIOB33_X105Y137_IOB_X1Y137_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y137_IOB_X1Y138_IBUF (
.I(RIOB33_X105Y137_IOB_X1Y138_IPAD),
.O(RIOB33_X105Y137_IOB_X1Y138_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y139_IOB_X1Y139_IBUF (
.I(RIOB33_X105Y139_IOB_X1Y139_IPAD),
.O(RIOB33_X105Y139_IOB_X1Y139_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y139_IOB_X1Y140_IBUF (
.I(RIOB33_X105Y139_IOB_X1Y140_IPAD),
.O(RIOB33_X105Y139_IOB_X1Y140_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y141_IOB_X1Y141_IBUF (
.I(RIOB33_X105Y141_IOB_X1Y141_IPAD),
.O(RIOB33_X105Y141_IOB_X1Y141_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y141_IOB_X1Y142_IBUF (
.I(RIOB33_X105Y141_IOB_X1Y142_IPAD),
.O(RIOB33_X105Y141_IOB_X1Y142_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y143_IOB_X1Y143_IBUF (
.I(RIOB33_X105Y143_IOB_X1Y143_IPAD),
.O(RIOB33_X105Y143_IOB_X1Y143_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y143_IOB_X1Y144_IBUF (
.I(RIOB33_X105Y143_IOB_X1Y144_IPAD),
.O(RIOB33_X105Y143_IOB_X1Y144_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y145_IOB_X1Y145_IBUF (
.I(RIOB33_X105Y145_IOB_X1Y145_IPAD),
.O(RIOB33_X105Y145_IOB_X1Y145_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y145_IOB_X1Y146_IBUF (
.I(RIOB33_X105Y145_IOB_X1Y146_IPAD),
.O(RIOB33_X105Y145_IOB_X1Y146_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y147_IOB_X1Y147_IBUF (
.I(RIOB33_X105Y147_IOB_X1Y147_IPAD),
.O(RIOB33_X105Y147_IOB_X1Y147_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y147_IOB_X1Y148_IBUF (
.I(RIOB33_X105Y147_IOB_X1Y148_IPAD),
.O(RIOB33_X105Y147_IOB_X1Y148_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y151_IOB_X1Y151_OBUF (
.I(LIOB33_X0Y75_IOB_X0Y76_I),
.O(RIOB33_X105Y151_IOB_X1Y151_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y151_IOB_X1Y152_OBUF (
.I(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.O(RIOB33_X105Y151_IOB_X1Y152_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y153_IOB_X1Y153_OBUF (
.I(RIOB33_X105Y101_IOB_X1Y101_I),
.O(RIOB33_X105Y153_IOB_X1Y153_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y153_IOB_X1Y154_OBUF (
.I(RIOB33_X105Y101_IOB_X1Y102_I),
.O(RIOB33_X105Y153_IOB_X1Y154_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y155_IOB_X1Y155_OBUF (
.I(RIOB33_X105Y103_IOB_X1Y103_I),
.O(RIOB33_X105Y155_IOB_X1Y155_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y155_IOB_X1Y156_OBUF (
.I(RIOB33_X105Y103_IOB_X1Y104_I),
.O(RIOB33_X105Y155_IOB_X1Y156_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y157_IOB_X1Y157_OBUF (
.I(RIOB33_X105Y125_IOB_X1Y126_I),
.O(RIOB33_X105Y157_IOB_X1Y157_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y157_IOB_X1Y158_OBUF (
.I(CLBLL_L_X36Y146_SLICE_X54Y146_AO6),
.O(RIOB33_X105Y157_IOB_X1Y158_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y159_IOB_X1Y159_OBUF (
.I(CLBLM_R_X11Y151_SLICE_X14Y151_DO6),
.O(RIOB33_X105Y159_IOB_X1Y159_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y159_IOB_X1Y160_OBUF (
.I(CLBLM_R_X11Y151_SLICE_X14Y151_DO5),
.O(RIOB33_X105Y159_IOB_X1Y160_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y161_IOB_X1Y161_OBUF (
.I(CLBLM_L_X10Y152_SLICE_X13Y152_CO6),
.O(RIOB33_X105Y161_IOB_X1Y161_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y161_IOB_X1Y162_OBUF (
.I(CLBLM_L_X10Y152_SLICE_X13Y152_CO5),
.O(RIOB33_X105Y161_IOB_X1Y162_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y163_IOB_X1Y163_OBUF (
.I(CLBLM_L_X10Y150_SLICE_X13Y150_DO6),
.O(RIOB33_X105Y163_IOB_X1Y163_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y163_IOB_X1Y164_OBUF (
.I(CLBLM_L_X10Y150_SLICE_X13Y150_DO5),
.O(RIOB33_X105Y163_IOB_X1Y164_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y165_IOB_X1Y165_OBUF (
.I(RIOB33_X105Y125_IOB_X1Y125_I),
.O(RIOB33_X105Y165_IOB_X1Y165_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y165_IOB_X1Y166_OBUF (
.I(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.O(RIOB33_X105Y165_IOB_X1Y166_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y167_IOB_X1Y167_OBUF (
.I(LIOB33_SING_X0Y50_IOB_X0Y50_I),
.O(RIOB33_X105Y167_IOB_X1Y167_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y167_IOB_X1Y168_OBUF (
.I(CLBLM_L_X8Y159_SLICE_X10Y159_AO6),
.O(RIOB33_X105Y167_IOB_X1Y168_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y169_IOB_X1Y169_OBUF (
.I(CLBLM_R_X103Y169_SLICE_X163Y169_AO6),
.O(RIOB33_X105Y169_IOB_X1Y169_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y169_IOB_X1Y170_OBUF (
.I(CLBLM_R_X103Y170_SLICE_X163Y170_AO6),
.O(RIOB33_X105Y169_IOB_X1Y170_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y171_IOB_X1Y171_OBUF (
.I(CLBLM_R_X11Y157_SLICE_X14Y157_AO5),
.O(RIOB33_X105Y171_IOB_X1Y171_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y171_IOB_X1Y172_OBUF (
.I(CLBLM_R_X103Y170_SLICE_X163Y170_AO5),
.O(RIOB33_X105Y171_IOB_X1Y172_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y173_IOB_X1Y173_OBUF (
.I(CLBLM_R_X103Y173_SLICE_X163Y173_AO6),
.O(RIOB33_X105Y173_IOB_X1Y173_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y173_IOB_X1Y174_OBUF (
.I(CLBLM_R_X103Y173_SLICE_X163Y173_AO5),
.O(RIOB33_X105Y173_IOB_X1Y174_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y175_IOB_X1Y175_OBUF (
.I(CLBLM_R_X15Y153_SLICE_X20Y153_AO6),
.O(RIOB33_X105Y175_IOB_X1Y175_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y175_IOB_X1Y176_OBUF (
.I(CLBLM_R_X103Y176_SLICE_X163Y176_AO6),
.O(RIOB33_X105Y175_IOB_X1Y176_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y177_IOB_X1Y177_OBUF (
.I(CLBLM_R_X103Y176_SLICE_X163Y176_AO5),
.O(RIOB33_X105Y177_IOB_X1Y177_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y177_IOB_X1Y178_OBUF (
.I(CLBLM_R_X103Y178_SLICE_X163Y178_AO6),
.O(RIOB33_X105Y177_IOB_X1Y178_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y179_IOB_X1Y179_OBUF (
.I(CLBLM_R_X103Y178_SLICE_X163Y178_AO5),
.O(RIOB33_X105Y179_IOB_X1Y179_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y179_IOB_X1Y180_OBUF (
.I(CLBLM_R_X11Y151_SLICE_X14Y151_DO6),
.O(RIOB33_X105Y179_IOB_X1Y180_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y181_IOB_X1Y181_OBUF (
.I(CLBLM_R_X11Y151_SLICE_X14Y151_DO5),
.O(RIOB33_X105Y181_IOB_X1Y181_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y181_IOB_X1Y182_OBUF (
.I(CLBLM_L_X10Y152_SLICE_X13Y152_CO6),
.O(RIOB33_X105Y181_IOB_X1Y182_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y183_IOB_X1Y183_OBUF (
.I(CLBLM_L_X10Y152_SLICE_X13Y152_CO5),
.O(RIOB33_X105Y183_IOB_X1Y183_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y183_IOB_X1Y184_OBUF (
.I(CLBLM_L_X10Y150_SLICE_X13Y150_DO6),
.O(RIOB33_X105Y183_IOB_X1Y184_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y185_IOB_X1Y185_OBUF (
.I(CLBLM_L_X10Y150_SLICE_X13Y150_DO5),
.O(RIOB33_X105Y185_IOB_X1Y185_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y185_IOB_X1Y186_OBUF (
.I(CLBLM_L_X12Y151_SLICE_X16Y151_AQ),
.O(RIOB33_X105Y185_IOB_X1Y186_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y187_IOB_X1Y187_OBUF (
.I(CLBLM_R_X11Y151_SLICE_X14Y151_BQ),
.O(RIOB33_X105Y187_IOB_X1Y187_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y187_IOB_X1Y188_OBUF (
.I(CLBLM_L_X10Y155_SLICE_X13Y155_AQ),
.O(RIOB33_X105Y187_IOB_X1Y188_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y189_IOB_X1Y189_OBUF (
.I(CLBLM_R_X11Y153_SLICE_X14Y153_CQ),
.O(RIOB33_X105Y189_IOB_X1Y189_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y189_IOB_X1Y190_OBUF (
.I(CLBLM_L_X12Y152_SLICE_X17Y152_AQ),
.O(RIOB33_X105Y189_IOB_X1Y190_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y191_IOB_X1Y191_OBUF (
.I(CLBLM_L_X10Y149_SLICE_X12Y149_AQ),
.O(RIOB33_X105Y191_IOB_X1Y191_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y191_IOB_X1Y192_OBUF (
.I(CLBLM_R_X11Y151_SLICE_X15Y151_AQ),
.O(RIOB33_X105Y191_IOB_X1Y192_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y193_IOB_X1Y193_OBUF (
.I(CLBLM_R_X11Y153_SLICE_X14Y153_AQ),
.O(RIOB33_X105Y193_IOB_X1Y193_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y193_IOB_X1Y194_OBUF (
.I(CLBLM_L_X12Y155_SLICE_X17Y155_AQ),
.O(RIOB33_X105Y193_IOB_X1Y194_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y195_IOB_X1Y195_OBUF (
.I(CLBLM_R_X11Y151_SLICE_X14Y151_AQ),
.O(RIOB33_X105Y195_IOB_X1Y195_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y195_IOB_X1Y196_OBUF (
.I(CLBLM_R_X11Y153_SLICE_X14Y153_BQ),
.O(RIOB33_X105Y195_IOB_X1Y196_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y197_IOB_X1Y197_OBUF (
.I(CLBLM_L_X16Y158_SLICE_X22Y158_AO6),
.O(RIOB33_X105Y197_IOB_X1Y197_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y197_IOB_X1Y198_OBUF (
.I(CLBLM_L_X16Y158_SLICE_X22Y158_AO6),
.O(RIOB33_X105Y197_IOB_X1Y198_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_SING_X105Y100_IOB_X1Y100_IBUF (
.I(RIOB33_SING_X105Y100_IOB_X1Y100_IPAD),
.O(RIOB33_SING_X105Y100_IOB_X1Y100_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_SING_X105Y149_IOB_X1Y149_IBUF (
.I(RIOB33_SING_X105Y149_IOB_X1Y149_IPAD),
.O(RIOB33_SING_X105Y149_IOB_X1Y149_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_SING_X105Y150_IOB_X1Y150_OBUF (
.I(LIOB33_X0Y75_IOB_X0Y75_I),
.O(RIOB33_SING_X105Y150_IOB_X1Y150_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_SING_X105Y199_IOB_X1Y199_OBUF (
.I(CLBLM_L_X12Y155_SLICE_X17Y155_AQ),
.O(RIOB33_SING_X105Y199_IOB_X1Y199_OPAD)
  );
  assign CLBLL_L_X2Y120_SLICE_X0Y120_A = CLBLL_L_X2Y120_SLICE_X0Y120_AO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_B = CLBLL_L_X2Y120_SLICE_X0Y120_BO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_C = CLBLL_L_X2Y120_SLICE_X0Y120_CO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_D = CLBLL_L_X2Y120_SLICE_X0Y120_DO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_A = CLBLL_L_X2Y120_SLICE_X1Y120_AO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_B = CLBLL_L_X2Y120_SLICE_X1Y120_BO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_C = CLBLL_L_X2Y120_SLICE_X1Y120_CO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_D = CLBLL_L_X2Y120_SLICE_X1Y120_DO6;
  assign CLBLL_L_X2Y134_SLICE_X0Y134_A = CLBLL_L_X2Y134_SLICE_X0Y134_AO6;
  assign CLBLL_L_X2Y134_SLICE_X0Y134_B = CLBLL_L_X2Y134_SLICE_X0Y134_BO6;
  assign CLBLL_L_X2Y134_SLICE_X0Y134_C = CLBLL_L_X2Y134_SLICE_X0Y134_CO6;
  assign CLBLL_L_X2Y134_SLICE_X0Y134_D = CLBLL_L_X2Y134_SLICE_X0Y134_DO6;
  assign CLBLL_L_X2Y134_SLICE_X0Y134_AMUX = CLBLL_L_X2Y134_SLICE_X0Y134_AO5;
  assign CLBLL_L_X2Y134_SLICE_X1Y134_A = CLBLL_L_X2Y134_SLICE_X1Y134_AO6;
  assign CLBLL_L_X2Y134_SLICE_X1Y134_B = CLBLL_L_X2Y134_SLICE_X1Y134_BO6;
  assign CLBLL_L_X2Y134_SLICE_X1Y134_C = CLBLL_L_X2Y134_SLICE_X1Y134_CO6;
  assign CLBLL_L_X2Y134_SLICE_X1Y134_D = CLBLL_L_X2Y134_SLICE_X1Y134_DO6;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_A = CLBLL_L_X2Y138_SLICE_X0Y138_AO6;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_B = CLBLL_L_X2Y138_SLICE_X0Y138_BO6;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_C = CLBLL_L_X2Y138_SLICE_X0Y138_CO6;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_D = CLBLL_L_X2Y138_SLICE_X0Y138_DO6;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_AMUX = CLBLL_L_X2Y138_SLICE_X0Y138_AO5;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_BMUX = CLBLL_L_X2Y138_SLICE_X0Y138_BO5;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_CMUX = CLBLL_L_X2Y138_SLICE_X0Y138_CO5;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_A = CLBLL_L_X2Y138_SLICE_X1Y138_AO6;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_B = CLBLL_L_X2Y138_SLICE_X1Y138_BO6;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_C = CLBLL_L_X2Y138_SLICE_X1Y138_CO6;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_D = CLBLL_L_X2Y138_SLICE_X1Y138_DO6;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_A = CLBLL_L_X2Y141_SLICE_X0Y141_AO6;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_B = CLBLL_L_X2Y141_SLICE_X0Y141_BO6;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_C = CLBLL_L_X2Y141_SLICE_X0Y141_CO6;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_D = CLBLL_L_X2Y141_SLICE_X0Y141_DO6;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_AMUX = CLBLL_L_X2Y141_SLICE_X0Y141_AO5;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_A = CLBLL_L_X2Y141_SLICE_X1Y141_AO6;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_B = CLBLL_L_X2Y141_SLICE_X1Y141_BO6;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_C = CLBLL_L_X2Y141_SLICE_X1Y141_CO6;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_D = CLBLL_L_X2Y141_SLICE_X1Y141_DO6;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_A = CLBLL_L_X2Y142_SLICE_X0Y142_AO6;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_B = CLBLL_L_X2Y142_SLICE_X0Y142_BO6;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_C = CLBLL_L_X2Y142_SLICE_X0Y142_CO6;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_D = CLBLL_L_X2Y142_SLICE_X0Y142_DO6;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_A = CLBLL_L_X2Y142_SLICE_X1Y142_AO6;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_B = CLBLL_L_X2Y142_SLICE_X1Y142_BO6;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_C = CLBLL_L_X2Y142_SLICE_X1Y142_CO6;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_D = CLBLL_L_X2Y142_SLICE_X1Y142_DO6;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_A = CLBLL_L_X2Y145_SLICE_X0Y145_AO6;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_B = CLBLL_L_X2Y145_SLICE_X0Y145_BO6;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_C = CLBLL_L_X2Y145_SLICE_X0Y145_CO6;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_D = CLBLL_L_X2Y145_SLICE_X0Y145_DO6;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_A = CLBLL_L_X2Y145_SLICE_X1Y145_AO6;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_B = CLBLL_L_X2Y145_SLICE_X1Y145_BO6;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_C = CLBLL_L_X2Y145_SLICE_X1Y145_CO6;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_D = CLBLL_L_X2Y145_SLICE_X1Y145_DO6;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_A = CLBLL_L_X2Y146_SLICE_X0Y146_AO6;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_B = CLBLL_L_X2Y146_SLICE_X0Y146_BO6;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_C = CLBLL_L_X2Y146_SLICE_X0Y146_CO6;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_D = CLBLL_L_X2Y146_SLICE_X0Y146_DO6;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_A = CLBLL_L_X2Y146_SLICE_X1Y146_AO6;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_B = CLBLL_L_X2Y146_SLICE_X1Y146_BO6;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_C = CLBLL_L_X2Y146_SLICE_X1Y146_CO6;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_D = CLBLL_L_X2Y146_SLICE_X1Y146_DO6;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_A = CLBLL_L_X2Y147_SLICE_X0Y147_AO6;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_B = CLBLL_L_X2Y147_SLICE_X0Y147_BO6;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_C = CLBLL_L_X2Y147_SLICE_X0Y147_CO6;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_D = CLBLL_L_X2Y147_SLICE_X0Y147_DO6;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_A = CLBLL_L_X2Y147_SLICE_X1Y147_AO6;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_B = CLBLL_L_X2Y147_SLICE_X1Y147_BO6;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_C = CLBLL_L_X2Y147_SLICE_X1Y147_CO6;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_D = CLBLL_L_X2Y147_SLICE_X1Y147_DO6;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_AMUX = CLBLL_L_X2Y147_SLICE_X1Y147_AO5;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_BMUX = CLBLL_L_X2Y147_SLICE_X1Y147_BO5;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_CMUX = CLBLL_L_X2Y147_SLICE_X1Y147_CO6;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_A = CLBLL_L_X2Y148_SLICE_X0Y148_AO6;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_B = CLBLL_L_X2Y148_SLICE_X0Y148_BO6;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_C = CLBLL_L_X2Y148_SLICE_X0Y148_CO6;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_D = CLBLL_L_X2Y148_SLICE_X0Y148_DO6;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_A = CLBLL_L_X2Y148_SLICE_X1Y148_AO6;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_B = CLBLL_L_X2Y148_SLICE_X1Y148_BO6;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_C = CLBLL_L_X2Y148_SLICE_X1Y148_CO6;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_D = CLBLL_L_X2Y148_SLICE_X1Y148_DO6;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_A = CLBLL_L_X2Y149_SLICE_X0Y149_AO6;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_B = CLBLL_L_X2Y149_SLICE_X0Y149_BO6;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_C = CLBLL_L_X2Y149_SLICE_X0Y149_CO6;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_D = CLBLL_L_X2Y149_SLICE_X0Y149_DO6;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_A = CLBLL_L_X2Y149_SLICE_X1Y149_AO6;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_B = CLBLL_L_X2Y149_SLICE_X1Y149_BO6;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_C = CLBLL_L_X2Y149_SLICE_X1Y149_CO6;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_D = CLBLL_L_X2Y149_SLICE_X1Y149_DO6;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_A = CLBLL_L_X2Y150_SLICE_X0Y150_AO6;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_B = CLBLL_L_X2Y150_SLICE_X0Y150_BO6;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_C = CLBLL_L_X2Y150_SLICE_X0Y150_CO6;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_D = CLBLL_L_X2Y150_SLICE_X0Y150_DO6;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_AMUX = CLBLL_L_X2Y150_SLICE_X0Y150_AO5;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_A = CLBLL_L_X2Y150_SLICE_X1Y150_AO6;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_B = CLBLL_L_X2Y150_SLICE_X1Y150_BO6;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_C = CLBLL_L_X2Y150_SLICE_X1Y150_CO6;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_D = CLBLL_L_X2Y150_SLICE_X1Y150_DO6;
  assign CLBLL_L_X2Y151_SLICE_X0Y151_A = CLBLL_L_X2Y151_SLICE_X0Y151_AO6;
  assign CLBLL_L_X2Y151_SLICE_X0Y151_B = CLBLL_L_X2Y151_SLICE_X0Y151_BO6;
  assign CLBLL_L_X2Y151_SLICE_X0Y151_C = CLBLL_L_X2Y151_SLICE_X0Y151_CO6;
  assign CLBLL_L_X2Y151_SLICE_X0Y151_D = CLBLL_L_X2Y151_SLICE_X0Y151_DO6;
  assign CLBLL_L_X2Y151_SLICE_X0Y151_AMUX = CLBLL_L_X2Y151_SLICE_X0Y151_AO5;
  assign CLBLL_L_X2Y151_SLICE_X0Y151_BMUX = CLBLL_L_X2Y151_SLICE_X0Y151_BO5;
  assign CLBLL_L_X2Y151_SLICE_X0Y151_CMUX = CLBLL_L_X2Y151_SLICE_X0Y151_CO5;
  assign CLBLL_L_X2Y151_SLICE_X0Y151_DMUX = CLBLL_L_X2Y151_SLICE_X0Y151_DO6;
  assign CLBLL_L_X2Y151_SLICE_X1Y151_A = CLBLL_L_X2Y151_SLICE_X1Y151_AO6;
  assign CLBLL_L_X2Y151_SLICE_X1Y151_B = CLBLL_L_X2Y151_SLICE_X1Y151_BO6;
  assign CLBLL_L_X2Y151_SLICE_X1Y151_C = CLBLL_L_X2Y151_SLICE_X1Y151_CO6;
  assign CLBLL_L_X2Y151_SLICE_X1Y151_D = CLBLL_L_X2Y151_SLICE_X1Y151_DO6;
  assign CLBLL_L_X2Y151_SLICE_X1Y151_AMUX = CLBLL_L_X2Y151_SLICE_X1Y151_AO5;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_A = CLBLL_L_X2Y152_SLICE_X0Y152_AO6;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_B = CLBLL_L_X2Y152_SLICE_X0Y152_BO6;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_C = CLBLL_L_X2Y152_SLICE_X0Y152_CO6;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_D = CLBLL_L_X2Y152_SLICE_X0Y152_DO6;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_A = CLBLL_L_X2Y152_SLICE_X1Y152_AO6;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_B = CLBLL_L_X2Y152_SLICE_X1Y152_BO6;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_C = CLBLL_L_X2Y152_SLICE_X1Y152_CO6;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_D = CLBLL_L_X2Y152_SLICE_X1Y152_DO6;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_AMUX = CLBLL_L_X2Y152_SLICE_X1Y152_AO5;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_BMUX = CLBLL_L_X2Y152_SLICE_X1Y152_BO5;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_A = CLBLL_L_X2Y153_SLICE_X0Y153_AO6;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_B = CLBLL_L_X2Y153_SLICE_X0Y153_BO6;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_C = CLBLL_L_X2Y153_SLICE_X0Y153_CO6;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_D = CLBLL_L_X2Y153_SLICE_X0Y153_DO6;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_A = CLBLL_L_X2Y153_SLICE_X1Y153_AO6;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_B = CLBLL_L_X2Y153_SLICE_X1Y153_BO6;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_C = CLBLL_L_X2Y153_SLICE_X1Y153_CO6;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_D = CLBLL_L_X2Y153_SLICE_X1Y153_DO6;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_AMUX = CLBLL_L_X2Y153_SLICE_X1Y153_AO6;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_CMUX = CLBLL_L_X2Y153_SLICE_X1Y153_CO6;
  assign CLBLL_L_X2Y154_SLICE_X0Y154_A = CLBLL_L_X2Y154_SLICE_X0Y154_AO6;
  assign CLBLL_L_X2Y154_SLICE_X0Y154_B = CLBLL_L_X2Y154_SLICE_X0Y154_BO6;
  assign CLBLL_L_X2Y154_SLICE_X0Y154_C = CLBLL_L_X2Y154_SLICE_X0Y154_CO6;
  assign CLBLL_L_X2Y154_SLICE_X0Y154_D = CLBLL_L_X2Y154_SLICE_X0Y154_DO6;
  assign CLBLL_L_X2Y154_SLICE_X1Y154_A = CLBLL_L_X2Y154_SLICE_X1Y154_AO6;
  assign CLBLL_L_X2Y154_SLICE_X1Y154_B = CLBLL_L_X2Y154_SLICE_X1Y154_BO6;
  assign CLBLL_L_X2Y154_SLICE_X1Y154_C = CLBLL_L_X2Y154_SLICE_X1Y154_CO6;
  assign CLBLL_L_X2Y154_SLICE_X1Y154_D = CLBLL_L_X2Y154_SLICE_X1Y154_DO6;
  assign CLBLL_L_X2Y154_SLICE_X1Y154_AMUX = CLBLL_L_X2Y154_SLICE_X1Y154_AO5;
  assign CLBLL_L_X2Y154_SLICE_X1Y154_BMUX = CLBLL_L_X2Y154_SLICE_X1Y154_BO5;
  assign CLBLL_L_X2Y154_SLICE_X1Y154_CMUX = CLBLL_L_X2Y154_SLICE_X1Y154_CO5;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_A = CLBLL_L_X2Y155_SLICE_X0Y155_AO6;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_B = CLBLL_L_X2Y155_SLICE_X0Y155_BO6;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_C = CLBLL_L_X2Y155_SLICE_X0Y155_CO6;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_D = CLBLL_L_X2Y155_SLICE_X0Y155_DO6;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_A = CLBLL_L_X2Y155_SLICE_X1Y155_AO6;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_B = CLBLL_L_X2Y155_SLICE_X1Y155_BO6;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_C = CLBLL_L_X2Y155_SLICE_X1Y155_CO6;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_D = CLBLL_L_X2Y155_SLICE_X1Y155_DO6;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_A = CLBLL_L_X4Y142_SLICE_X4Y142_AO6;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_B = CLBLL_L_X4Y142_SLICE_X4Y142_BO6;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_C = CLBLL_L_X4Y142_SLICE_X4Y142_CO6;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_D = CLBLL_L_X4Y142_SLICE_X4Y142_DO6;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_A = CLBLL_L_X4Y142_SLICE_X5Y142_AO6;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_B = CLBLL_L_X4Y142_SLICE_X5Y142_BO6;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_C = CLBLL_L_X4Y142_SLICE_X5Y142_CO6;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_D = CLBLL_L_X4Y142_SLICE_X5Y142_DO6;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_AMUX = CLBLL_L_X4Y142_SLICE_X5Y142_AO5;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_A = CLBLL_L_X4Y143_SLICE_X4Y143_AO6;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_B = CLBLL_L_X4Y143_SLICE_X4Y143_BO6;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_C = CLBLL_L_X4Y143_SLICE_X4Y143_CO6;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_D = CLBLL_L_X4Y143_SLICE_X4Y143_DO6;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_CMUX = CLBLL_L_X4Y143_SLICE_X4Y143_CO5;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_A = CLBLL_L_X4Y143_SLICE_X5Y143_AO6;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_B = CLBLL_L_X4Y143_SLICE_X5Y143_BO6;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_C = CLBLL_L_X4Y143_SLICE_X5Y143_CO6;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_D = CLBLL_L_X4Y143_SLICE_X5Y143_DO6;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_A = CLBLL_L_X4Y144_SLICE_X4Y144_AO6;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_B = CLBLL_L_X4Y144_SLICE_X4Y144_BO6;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_C = CLBLL_L_X4Y144_SLICE_X4Y144_CO6;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_D = CLBLL_L_X4Y144_SLICE_X4Y144_DO6;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_CMUX = CLBLL_L_X4Y144_SLICE_X4Y144_CO5;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_A = CLBLL_L_X4Y144_SLICE_X5Y144_AO6;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_B = CLBLL_L_X4Y144_SLICE_X5Y144_BO6;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_C = CLBLL_L_X4Y144_SLICE_X5Y144_CO6;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_D = CLBLL_L_X4Y144_SLICE_X5Y144_DO6;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_AMUX = CLBLL_L_X4Y144_SLICE_X5Y144_A5Q;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_CMUX = CLBLL_L_X4Y144_SLICE_X5Y144_CO5;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_A = CLBLL_L_X4Y145_SLICE_X4Y145_AO6;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_B = CLBLL_L_X4Y145_SLICE_X4Y145_BO6;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_C = CLBLL_L_X4Y145_SLICE_X4Y145_CO6;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_D = CLBLL_L_X4Y145_SLICE_X4Y145_DO6;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_AMUX = CLBLL_L_X4Y145_SLICE_X4Y145_A5Q;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_BMUX = CLBLL_L_X4Y145_SLICE_X4Y145_BO5;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_A = CLBLL_L_X4Y145_SLICE_X5Y145_AO6;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_B = CLBLL_L_X4Y145_SLICE_X5Y145_BO6;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_C = CLBLL_L_X4Y145_SLICE_X5Y145_CO6;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_D = CLBLL_L_X4Y145_SLICE_X5Y145_DO6;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_BMUX = CLBLL_L_X4Y145_SLICE_X5Y145_BO5;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_A = CLBLL_L_X4Y146_SLICE_X4Y146_AO6;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_B = CLBLL_L_X4Y146_SLICE_X4Y146_BO6;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_C = CLBLL_L_X4Y146_SLICE_X4Y146_CO6;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_D = CLBLL_L_X4Y146_SLICE_X4Y146_DO6;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_AMUX = CLBLL_L_X4Y146_SLICE_X4Y146_A5Q;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_CMUX = CLBLL_L_X4Y146_SLICE_X4Y146_CO5;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_A = CLBLL_L_X4Y146_SLICE_X5Y146_AO6;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_B = CLBLL_L_X4Y146_SLICE_X5Y146_BO6;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_C = CLBLL_L_X4Y146_SLICE_X5Y146_CO6;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_D = CLBLL_L_X4Y146_SLICE_X5Y146_DO6;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_AMUX = CLBLL_L_X4Y146_SLICE_X5Y146_A5Q;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_BMUX = CLBLL_L_X4Y146_SLICE_X5Y146_BO5;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_A = CLBLL_L_X4Y147_SLICE_X4Y147_AO6;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_B = CLBLL_L_X4Y147_SLICE_X4Y147_BO6;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_C = CLBLL_L_X4Y147_SLICE_X4Y147_CO6;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_D = CLBLL_L_X4Y147_SLICE_X4Y147_DO6;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_A = CLBLL_L_X4Y147_SLICE_X5Y147_AO6;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_B = CLBLL_L_X4Y147_SLICE_X5Y147_BO6;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_C = CLBLL_L_X4Y147_SLICE_X5Y147_CO6;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_D = CLBLL_L_X4Y147_SLICE_X5Y147_DO6;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_BMUX = CLBLL_L_X4Y147_SLICE_X5Y147_B5Q;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_A = CLBLL_L_X4Y148_SLICE_X4Y148_AO6;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_B = CLBLL_L_X4Y148_SLICE_X4Y148_BO6;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_C = CLBLL_L_X4Y148_SLICE_X4Y148_CO6;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_D = CLBLL_L_X4Y148_SLICE_X4Y148_DO6;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_CMUX = CLBLL_L_X4Y148_SLICE_X4Y148_C5Q;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_A = CLBLL_L_X4Y148_SLICE_X5Y148_AO6;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_B = CLBLL_L_X4Y148_SLICE_X5Y148_BO6;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_C = CLBLL_L_X4Y148_SLICE_X5Y148_CO6;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_D = CLBLL_L_X4Y148_SLICE_X5Y148_DO6;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_A = CLBLL_L_X4Y149_SLICE_X4Y149_AO6;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_B = CLBLL_L_X4Y149_SLICE_X4Y149_BO6;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_C = CLBLL_L_X4Y149_SLICE_X4Y149_CO6;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_D = CLBLL_L_X4Y149_SLICE_X4Y149_DO6;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_A = CLBLL_L_X4Y149_SLICE_X5Y149_AO6;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_B = CLBLL_L_X4Y149_SLICE_X5Y149_BO6;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_C = CLBLL_L_X4Y149_SLICE_X5Y149_CO6;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_D = CLBLL_L_X4Y149_SLICE_X5Y149_DO6;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_AMUX = CLBLL_L_X4Y149_SLICE_X5Y149_A5Q;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_BMUX = CLBLL_L_X4Y149_SLICE_X5Y149_BO5;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_A = CLBLL_L_X4Y150_SLICE_X4Y150_AO6;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_B = CLBLL_L_X4Y150_SLICE_X4Y150_BO6;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_C = CLBLL_L_X4Y150_SLICE_X4Y150_CO6;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_D = CLBLL_L_X4Y150_SLICE_X4Y150_DO6;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_BMUX = CLBLL_L_X4Y150_SLICE_X4Y150_B5Q;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_A = CLBLL_L_X4Y150_SLICE_X5Y150_AO6;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_B = CLBLL_L_X4Y150_SLICE_X5Y150_BO6;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_C = CLBLL_L_X4Y150_SLICE_X5Y150_CO6;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_D = CLBLL_L_X4Y150_SLICE_X5Y150_DO6;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_A = CLBLL_L_X4Y151_SLICE_X4Y151_AO6;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_B = CLBLL_L_X4Y151_SLICE_X4Y151_BO6;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_C = CLBLL_L_X4Y151_SLICE_X4Y151_CO6;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_D = CLBLL_L_X4Y151_SLICE_X4Y151_DO6;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_AMUX = CLBLL_L_X4Y151_SLICE_X4Y151_A5Q;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_A = CLBLL_L_X4Y151_SLICE_X5Y151_AO6;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_B = CLBLL_L_X4Y151_SLICE_X5Y151_BO6;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_C = CLBLL_L_X4Y151_SLICE_X5Y151_CO6;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_D = CLBLL_L_X4Y151_SLICE_X5Y151_DO6;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_BMUX = CLBLL_L_X4Y151_SLICE_X5Y151_B5Q;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_DMUX = CLBLL_L_X4Y151_SLICE_X5Y151_DO6;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_A = CLBLL_L_X4Y152_SLICE_X4Y152_AO6;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_B = CLBLL_L_X4Y152_SLICE_X4Y152_BO6;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_C = CLBLL_L_X4Y152_SLICE_X4Y152_CO6;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_D = CLBLL_L_X4Y152_SLICE_X4Y152_DO6;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_AMUX = CLBLL_L_X4Y152_SLICE_X4Y152_AO5;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_CMUX = CLBLL_L_X4Y152_SLICE_X4Y152_CO6;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_A = CLBLL_L_X4Y152_SLICE_X5Y152_AO6;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_B = CLBLL_L_X4Y152_SLICE_X5Y152_BO6;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_C = CLBLL_L_X4Y152_SLICE_X5Y152_CO6;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_D = CLBLL_L_X4Y152_SLICE_X5Y152_DO6;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_AMUX = CLBLL_L_X4Y152_SLICE_X5Y152_AO5;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_A = CLBLL_L_X4Y153_SLICE_X4Y153_AO6;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_B = CLBLL_L_X4Y153_SLICE_X4Y153_BO6;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_C = CLBLL_L_X4Y153_SLICE_X4Y153_CO6;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_D = CLBLL_L_X4Y153_SLICE_X4Y153_DO6;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_A = CLBLL_L_X4Y153_SLICE_X5Y153_AO6;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_B = CLBLL_L_X4Y153_SLICE_X5Y153_BO6;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_C = CLBLL_L_X4Y153_SLICE_X5Y153_CO6;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_D = CLBLL_L_X4Y153_SLICE_X5Y153_DO6;
  assign CLBLL_L_X4Y154_SLICE_X4Y154_A = CLBLL_L_X4Y154_SLICE_X4Y154_AO6;
  assign CLBLL_L_X4Y154_SLICE_X4Y154_B = CLBLL_L_X4Y154_SLICE_X4Y154_BO6;
  assign CLBLL_L_X4Y154_SLICE_X4Y154_C = CLBLL_L_X4Y154_SLICE_X4Y154_CO6;
  assign CLBLL_L_X4Y154_SLICE_X4Y154_D = CLBLL_L_X4Y154_SLICE_X4Y154_DO6;
  assign CLBLL_L_X4Y154_SLICE_X4Y154_AMUX = CLBLL_L_X4Y154_SLICE_X4Y154_AO6;
  assign CLBLL_L_X4Y154_SLICE_X5Y154_A = CLBLL_L_X4Y154_SLICE_X5Y154_AO6;
  assign CLBLL_L_X4Y154_SLICE_X5Y154_B = CLBLL_L_X4Y154_SLICE_X5Y154_BO6;
  assign CLBLL_L_X4Y154_SLICE_X5Y154_C = CLBLL_L_X4Y154_SLICE_X5Y154_CO6;
  assign CLBLL_L_X4Y154_SLICE_X5Y154_D = CLBLL_L_X4Y154_SLICE_X5Y154_DO6;
  assign CLBLL_L_X4Y154_SLICE_X5Y154_CMUX = CLBLL_L_X4Y154_SLICE_X5Y154_CO5;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_A = CLBLL_L_X4Y155_SLICE_X4Y155_AO6;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_B = CLBLL_L_X4Y155_SLICE_X4Y155_BO6;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_C = CLBLL_L_X4Y155_SLICE_X4Y155_CO6;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_D = CLBLL_L_X4Y155_SLICE_X4Y155_DO6;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_AMUX = CLBLL_L_X4Y155_SLICE_X4Y155_AO5;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_BMUX = CLBLL_L_X4Y155_SLICE_X4Y155_BO5;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_A = CLBLL_L_X4Y155_SLICE_X5Y155_AO6;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_B = CLBLL_L_X4Y155_SLICE_X5Y155_BO6;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_C = CLBLL_L_X4Y155_SLICE_X5Y155_CO6;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_D = CLBLL_L_X4Y155_SLICE_X5Y155_DO6;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_AMUX = CLBLL_L_X4Y155_SLICE_X5Y155_AO5;
  assign CLBLL_L_X36Y146_SLICE_X54Y146_A = CLBLL_L_X36Y146_SLICE_X54Y146_AO6;
  assign CLBLL_L_X36Y146_SLICE_X54Y146_B = CLBLL_L_X36Y146_SLICE_X54Y146_BO6;
  assign CLBLL_L_X36Y146_SLICE_X54Y146_C = CLBLL_L_X36Y146_SLICE_X54Y146_CO6;
  assign CLBLL_L_X36Y146_SLICE_X54Y146_D = CLBLL_L_X36Y146_SLICE_X54Y146_DO6;
  assign CLBLL_L_X36Y146_SLICE_X55Y146_A = CLBLL_L_X36Y146_SLICE_X55Y146_AO6;
  assign CLBLL_L_X36Y146_SLICE_X55Y146_B = CLBLL_L_X36Y146_SLICE_X55Y146_BO6;
  assign CLBLL_L_X36Y146_SLICE_X55Y146_C = CLBLL_L_X36Y146_SLICE_X55Y146_CO6;
  assign CLBLL_L_X36Y146_SLICE_X55Y146_D = CLBLL_L_X36Y146_SLICE_X55Y146_DO6;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_A = CLBLL_L_X52Y126_SLICE_X78Y126_AO6;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_B = CLBLL_L_X52Y126_SLICE_X78Y126_BO6;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_C = CLBLL_L_X52Y126_SLICE_X78Y126_CO6;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_D = CLBLL_L_X52Y126_SLICE_X78Y126_DO6;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_A = CLBLL_L_X52Y126_SLICE_X79Y126_AO6;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_B = CLBLL_L_X52Y126_SLICE_X79Y126_BO6;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_C = CLBLL_L_X52Y126_SLICE_X79Y126_CO6;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_D = CLBLL_L_X52Y126_SLICE_X79Y126_DO6;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_A = CLBLM_L_X8Y142_SLICE_X10Y142_AO6;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_B = CLBLM_L_X8Y142_SLICE_X10Y142_BO6;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_C = CLBLM_L_X8Y142_SLICE_X10Y142_CO6;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_D = CLBLM_L_X8Y142_SLICE_X10Y142_DO6;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_AMUX = CLBLM_L_X8Y142_SLICE_X10Y142_A5Q;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_A = CLBLM_L_X8Y142_SLICE_X11Y142_AO6;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_B = CLBLM_L_X8Y142_SLICE_X11Y142_BO6;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_C = CLBLM_L_X8Y142_SLICE_X11Y142_CO6;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_D = CLBLM_L_X8Y142_SLICE_X11Y142_DO6;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_A = CLBLM_L_X8Y143_SLICE_X10Y143_AO6;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_B = CLBLM_L_X8Y143_SLICE_X10Y143_BO6;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_C = CLBLM_L_X8Y143_SLICE_X10Y143_CO6;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_D = CLBLM_L_X8Y143_SLICE_X10Y143_DO6;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_A = CLBLM_L_X8Y143_SLICE_X11Y143_AO6;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_B = CLBLM_L_X8Y143_SLICE_X11Y143_BO6;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_C = CLBLM_L_X8Y143_SLICE_X11Y143_CO6;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_D = CLBLM_L_X8Y143_SLICE_X11Y143_DO6;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_BMUX = CLBLM_L_X8Y143_SLICE_X11Y143_BO6;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_A = CLBLM_L_X8Y144_SLICE_X10Y144_AO6;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_B = CLBLM_L_X8Y144_SLICE_X10Y144_BO6;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_C = CLBLM_L_X8Y144_SLICE_X10Y144_CO6;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_D = CLBLM_L_X8Y144_SLICE_X10Y144_DO6;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_A = CLBLM_L_X8Y144_SLICE_X11Y144_AO6;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_B = CLBLM_L_X8Y144_SLICE_X11Y144_BO6;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_C = CLBLM_L_X8Y144_SLICE_X11Y144_CO6;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_D = CLBLM_L_X8Y144_SLICE_X11Y144_DO6;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_A = CLBLM_L_X8Y145_SLICE_X10Y145_AO6;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_B = CLBLM_L_X8Y145_SLICE_X10Y145_BO6;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_C = CLBLM_L_X8Y145_SLICE_X10Y145_CO6;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_D = CLBLM_L_X8Y145_SLICE_X10Y145_DO6;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_AMUX = CLBLM_L_X8Y145_SLICE_X10Y145_A5Q;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_CMUX = CLBLM_L_X8Y145_SLICE_X10Y145_CO5;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_A = CLBLM_L_X8Y145_SLICE_X11Y145_AO6;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_B = CLBLM_L_X8Y145_SLICE_X11Y145_BO6;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_C = CLBLM_L_X8Y145_SLICE_X11Y145_CO6;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_D = CLBLM_L_X8Y145_SLICE_X11Y145_DO6;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_AMUX = CLBLM_L_X8Y145_SLICE_X11Y145_A5Q;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_BMUX = CLBLM_L_X8Y145_SLICE_X11Y145_B5Q;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_A = CLBLM_L_X8Y146_SLICE_X10Y146_AO6;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_B = CLBLM_L_X8Y146_SLICE_X10Y146_BO6;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_C = CLBLM_L_X8Y146_SLICE_X10Y146_CO6;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_D = CLBLM_L_X8Y146_SLICE_X10Y146_DO6;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_BMUX = CLBLM_L_X8Y146_SLICE_X10Y146_B5Q;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_A = CLBLM_L_X8Y146_SLICE_X11Y146_AO6;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_B = CLBLM_L_X8Y146_SLICE_X11Y146_BO6;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_C = CLBLM_L_X8Y146_SLICE_X11Y146_CO6;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_D = CLBLM_L_X8Y146_SLICE_X11Y146_DO6;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_A = CLBLM_L_X8Y147_SLICE_X10Y147_AO6;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_B = CLBLM_L_X8Y147_SLICE_X10Y147_BO6;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_C = CLBLM_L_X8Y147_SLICE_X10Y147_CO6;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_D = CLBLM_L_X8Y147_SLICE_X10Y147_DO6;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_A = CLBLM_L_X8Y147_SLICE_X11Y147_AO6;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_B = CLBLM_L_X8Y147_SLICE_X11Y147_BO6;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_C = CLBLM_L_X8Y147_SLICE_X11Y147_CO6;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_D = CLBLM_L_X8Y147_SLICE_X11Y147_DO6;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_AMUX = CLBLM_L_X8Y147_SLICE_X11Y147_AO5;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_BMUX = CLBLM_L_X8Y147_SLICE_X11Y147_BO5;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_CMUX = CLBLM_L_X8Y147_SLICE_X11Y147_CO6;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_A = CLBLM_L_X8Y148_SLICE_X10Y148_AO6;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_B = CLBLM_L_X8Y148_SLICE_X10Y148_BO6;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_C = CLBLM_L_X8Y148_SLICE_X10Y148_CO6;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_D = CLBLM_L_X8Y148_SLICE_X10Y148_DO6;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_AMUX = CLBLM_L_X8Y148_SLICE_X10Y148_A5Q;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_BMUX = CLBLM_L_X8Y148_SLICE_X10Y148_BO5;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_CMUX = CLBLM_L_X8Y148_SLICE_X10Y148_CO5;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_DMUX = CLBLM_L_X8Y148_SLICE_X10Y148_DO5;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_A = CLBLM_L_X8Y148_SLICE_X11Y148_AO6;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_B = CLBLM_L_X8Y148_SLICE_X11Y148_BO6;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_C = CLBLM_L_X8Y148_SLICE_X11Y148_CO6;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_D = CLBLM_L_X8Y148_SLICE_X11Y148_DO6;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_CMUX = CLBLM_L_X8Y148_SLICE_X11Y148_CO6;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_A = CLBLM_L_X8Y149_SLICE_X10Y149_AO6;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_B = CLBLM_L_X8Y149_SLICE_X10Y149_BO6;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_C = CLBLM_L_X8Y149_SLICE_X10Y149_CO6;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_D = CLBLM_L_X8Y149_SLICE_X10Y149_DO6;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_AMUX = CLBLM_L_X8Y149_SLICE_X10Y149_AO5;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_A = CLBLM_L_X8Y149_SLICE_X11Y149_AO6;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_B = CLBLM_L_X8Y149_SLICE_X11Y149_BO6;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_C = CLBLM_L_X8Y149_SLICE_X11Y149_CO6;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_D = CLBLM_L_X8Y149_SLICE_X11Y149_DO6;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_BMUX = CLBLM_L_X8Y149_SLICE_X11Y149_B5Q;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_A = CLBLM_L_X8Y150_SLICE_X10Y150_AO6;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_B = CLBLM_L_X8Y150_SLICE_X10Y150_BO6;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_C = CLBLM_L_X8Y150_SLICE_X10Y150_CO6;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_D = CLBLM_L_X8Y150_SLICE_X10Y150_DO6;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_A = CLBLM_L_X8Y150_SLICE_X11Y150_AO6;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_B = CLBLM_L_X8Y150_SLICE_X11Y150_BO6;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_C = CLBLM_L_X8Y150_SLICE_X11Y150_CO6;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_D = CLBLM_L_X8Y150_SLICE_X11Y150_DO6;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_A = CLBLM_L_X8Y151_SLICE_X10Y151_AO6;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_B = CLBLM_L_X8Y151_SLICE_X10Y151_BO6;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_C = CLBLM_L_X8Y151_SLICE_X10Y151_CO6;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_D = CLBLM_L_X8Y151_SLICE_X10Y151_DO6;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_BMUX = CLBLM_L_X8Y151_SLICE_X10Y151_B5Q;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_A = CLBLM_L_X8Y151_SLICE_X11Y151_AO6;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_B = CLBLM_L_X8Y151_SLICE_X11Y151_BO6;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_C = CLBLM_L_X8Y151_SLICE_X11Y151_CO6;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_D = CLBLM_L_X8Y151_SLICE_X11Y151_DO6;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_A = CLBLM_L_X8Y152_SLICE_X10Y152_AO6;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_B = CLBLM_L_X8Y152_SLICE_X10Y152_BO6;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_C = CLBLM_L_X8Y152_SLICE_X10Y152_CO6;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_D = CLBLM_L_X8Y152_SLICE_X10Y152_DO6;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_A = CLBLM_L_X8Y152_SLICE_X11Y152_AO6;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_B = CLBLM_L_X8Y152_SLICE_X11Y152_BO6;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_C = CLBLM_L_X8Y152_SLICE_X11Y152_CO6;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_D = CLBLM_L_X8Y152_SLICE_X11Y152_DO6;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_BMUX = CLBLM_L_X8Y152_SLICE_X11Y152_BO5;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_A = CLBLM_L_X8Y153_SLICE_X10Y153_AO6;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_B = CLBLM_L_X8Y153_SLICE_X10Y153_BO6;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_C = CLBLM_L_X8Y153_SLICE_X10Y153_CO6;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_D = CLBLM_L_X8Y153_SLICE_X10Y153_DO6;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_CMUX = CLBLM_L_X8Y153_SLICE_X10Y153_CO5;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_DMUX = CLBLM_L_X8Y153_SLICE_X10Y153_DO5;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_A = CLBLM_L_X8Y153_SLICE_X11Y153_AO6;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_B = CLBLM_L_X8Y153_SLICE_X11Y153_BO6;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_C = CLBLM_L_X8Y153_SLICE_X11Y153_CO6;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_D = CLBLM_L_X8Y153_SLICE_X11Y153_DO6;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_A = CLBLM_L_X8Y154_SLICE_X10Y154_AO6;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_B = CLBLM_L_X8Y154_SLICE_X10Y154_BO6;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_C = CLBLM_L_X8Y154_SLICE_X10Y154_CO6;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_D = CLBLM_L_X8Y154_SLICE_X10Y154_DO6;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_BMUX = CLBLM_L_X8Y154_SLICE_X10Y154_BO5;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_DMUX = CLBLM_L_X8Y154_SLICE_X10Y154_DO6;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_A = CLBLM_L_X8Y154_SLICE_X11Y154_AO6;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_B = CLBLM_L_X8Y154_SLICE_X11Y154_BO6;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_C = CLBLM_L_X8Y154_SLICE_X11Y154_CO6;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_D = CLBLM_L_X8Y154_SLICE_X11Y154_DO6;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_AMUX = CLBLM_L_X8Y154_SLICE_X11Y154_AO5;
  assign CLBLM_L_X8Y155_SLICE_X10Y155_A = CLBLM_L_X8Y155_SLICE_X10Y155_AO6;
  assign CLBLM_L_X8Y155_SLICE_X10Y155_B = CLBLM_L_X8Y155_SLICE_X10Y155_BO6;
  assign CLBLM_L_X8Y155_SLICE_X10Y155_C = CLBLM_L_X8Y155_SLICE_X10Y155_CO6;
  assign CLBLM_L_X8Y155_SLICE_X10Y155_D = CLBLM_L_X8Y155_SLICE_X10Y155_DO6;
  assign CLBLM_L_X8Y155_SLICE_X10Y155_CMUX = CLBLM_L_X8Y155_SLICE_X10Y155_CO6;
  assign CLBLM_L_X8Y155_SLICE_X11Y155_A = CLBLM_L_X8Y155_SLICE_X11Y155_AO6;
  assign CLBLM_L_X8Y155_SLICE_X11Y155_B = CLBLM_L_X8Y155_SLICE_X11Y155_BO6;
  assign CLBLM_L_X8Y155_SLICE_X11Y155_C = CLBLM_L_X8Y155_SLICE_X11Y155_CO6;
  assign CLBLM_L_X8Y155_SLICE_X11Y155_D = CLBLM_L_X8Y155_SLICE_X11Y155_DO6;
  assign CLBLM_L_X8Y159_SLICE_X10Y159_A = CLBLM_L_X8Y159_SLICE_X10Y159_AO6;
  assign CLBLM_L_X8Y159_SLICE_X10Y159_B = CLBLM_L_X8Y159_SLICE_X10Y159_BO6;
  assign CLBLM_L_X8Y159_SLICE_X10Y159_C = CLBLM_L_X8Y159_SLICE_X10Y159_CO6;
  assign CLBLM_L_X8Y159_SLICE_X10Y159_D = CLBLM_L_X8Y159_SLICE_X10Y159_DO6;
  assign CLBLM_L_X8Y159_SLICE_X11Y159_A = CLBLM_L_X8Y159_SLICE_X11Y159_AO6;
  assign CLBLM_L_X8Y159_SLICE_X11Y159_B = CLBLM_L_X8Y159_SLICE_X11Y159_BO6;
  assign CLBLM_L_X8Y159_SLICE_X11Y159_C = CLBLM_L_X8Y159_SLICE_X11Y159_CO6;
  assign CLBLM_L_X8Y159_SLICE_X11Y159_D = CLBLM_L_X8Y159_SLICE_X11Y159_DO6;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_A = CLBLM_L_X10Y141_SLICE_X12Y141_AO6;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_B = CLBLM_L_X10Y141_SLICE_X12Y141_BO6;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_C = CLBLM_L_X10Y141_SLICE_X12Y141_CO6;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_D = CLBLM_L_X10Y141_SLICE_X12Y141_DO6;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_AMUX = CLBLM_L_X10Y141_SLICE_X12Y141_AO5;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_BMUX = CLBLM_L_X10Y141_SLICE_X12Y141_BO5;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_A = CLBLM_L_X10Y141_SLICE_X13Y141_AO6;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_B = CLBLM_L_X10Y141_SLICE_X13Y141_BO6;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_C = CLBLM_L_X10Y141_SLICE_X13Y141_CO6;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_D = CLBLM_L_X10Y141_SLICE_X13Y141_DO6;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_A = CLBLM_L_X10Y142_SLICE_X12Y142_AO6;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_B = CLBLM_L_X10Y142_SLICE_X12Y142_BO6;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_C = CLBLM_L_X10Y142_SLICE_X12Y142_CO6;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_D = CLBLM_L_X10Y142_SLICE_X12Y142_DO6;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_A = CLBLM_L_X10Y142_SLICE_X13Y142_AO6;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_B = CLBLM_L_X10Y142_SLICE_X13Y142_BO6;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_C = CLBLM_L_X10Y142_SLICE_X13Y142_CO6;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_D = CLBLM_L_X10Y142_SLICE_X13Y142_DO6;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_BMUX = CLBLM_L_X10Y142_SLICE_X13Y142_BO5;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_CMUX = CLBLM_L_X10Y142_SLICE_X13Y142_CO6;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_DMUX = CLBLM_L_X10Y142_SLICE_X13Y142_DO6;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_A = CLBLM_L_X10Y143_SLICE_X12Y143_AO6;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_B = CLBLM_L_X10Y143_SLICE_X12Y143_BO6;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_C = CLBLM_L_X10Y143_SLICE_X12Y143_CO6;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_D = CLBLM_L_X10Y143_SLICE_X12Y143_DO6;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_A = CLBLM_L_X10Y143_SLICE_X13Y143_AO6;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_B = CLBLM_L_X10Y143_SLICE_X13Y143_BO6;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_C = CLBLM_L_X10Y143_SLICE_X13Y143_CO6;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_D = CLBLM_L_X10Y143_SLICE_X13Y143_DO6;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_CMUX = CLBLM_L_X10Y143_SLICE_X13Y143_CO5;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_DMUX = CLBLM_L_X10Y143_SLICE_X13Y143_DO6;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_A = CLBLM_L_X10Y144_SLICE_X12Y144_AO6;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_B = CLBLM_L_X10Y144_SLICE_X12Y144_BO6;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_C = CLBLM_L_X10Y144_SLICE_X12Y144_CO6;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_D = CLBLM_L_X10Y144_SLICE_X12Y144_DO6;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_A = CLBLM_L_X10Y144_SLICE_X13Y144_AO6;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_B = CLBLM_L_X10Y144_SLICE_X13Y144_BO6;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_C = CLBLM_L_X10Y144_SLICE_X13Y144_CO6;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_D = CLBLM_L_X10Y144_SLICE_X13Y144_DO6;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_A = CLBLM_L_X10Y145_SLICE_X12Y145_AO6;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_B = CLBLM_L_X10Y145_SLICE_X12Y145_BO6;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_C = CLBLM_L_X10Y145_SLICE_X12Y145_CO6;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_D = CLBLM_L_X10Y145_SLICE_X12Y145_DO6;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_CMUX = CLBLM_L_X10Y145_SLICE_X12Y145_C5Q;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_A = CLBLM_L_X10Y145_SLICE_X13Y145_AO6;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_B = CLBLM_L_X10Y145_SLICE_X13Y145_BO6;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_C = CLBLM_L_X10Y145_SLICE_X13Y145_CO6;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_D = CLBLM_L_X10Y145_SLICE_X13Y145_DO6;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_AMUX = CLBLM_L_X10Y145_SLICE_X13Y145_A5Q;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_A = CLBLM_L_X10Y146_SLICE_X12Y146_AO6;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_B = CLBLM_L_X10Y146_SLICE_X12Y146_BO6;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_C = CLBLM_L_X10Y146_SLICE_X12Y146_CO6;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_D = CLBLM_L_X10Y146_SLICE_X12Y146_DO6;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_AMUX = CLBLM_L_X10Y146_SLICE_X12Y146_A5Q;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_BMUX = CLBLM_L_X10Y146_SLICE_X12Y146_B5Q;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_CMUX = CLBLM_L_X10Y146_SLICE_X12Y146_C5Q;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_DMUX = CLBLM_L_X10Y146_SLICE_X12Y146_D5Q;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_A = CLBLM_L_X10Y146_SLICE_X13Y146_AO6;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_B = CLBLM_L_X10Y146_SLICE_X13Y146_BO6;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_C = CLBLM_L_X10Y146_SLICE_X13Y146_CO6;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_D = CLBLM_L_X10Y146_SLICE_X13Y146_DO6;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_AMUX = CLBLM_L_X10Y146_SLICE_X13Y146_A5Q;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_BMUX = CLBLM_L_X10Y146_SLICE_X13Y146_B5Q;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_A = CLBLM_L_X10Y147_SLICE_X12Y147_AO6;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_B = CLBLM_L_X10Y147_SLICE_X12Y147_BO6;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_C = CLBLM_L_X10Y147_SLICE_X12Y147_CO6;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_D = CLBLM_L_X10Y147_SLICE_X12Y147_DO6;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_AMUX = CLBLM_L_X10Y147_SLICE_X12Y147_A5Q;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_BMUX = CLBLM_L_X10Y147_SLICE_X12Y147_BO5;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_DMUX = CLBLM_L_X10Y147_SLICE_X12Y147_DO5;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_A = CLBLM_L_X10Y147_SLICE_X13Y147_AO6;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_B = CLBLM_L_X10Y147_SLICE_X13Y147_BO6;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_C = CLBLM_L_X10Y147_SLICE_X13Y147_CO6;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_D = CLBLM_L_X10Y147_SLICE_X13Y147_DO6;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_A = CLBLM_L_X10Y148_SLICE_X12Y148_AO6;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_B = CLBLM_L_X10Y148_SLICE_X12Y148_BO6;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_C = CLBLM_L_X10Y148_SLICE_X12Y148_CO6;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_D = CLBLM_L_X10Y148_SLICE_X12Y148_DO6;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_AMUX = CLBLM_L_X10Y148_SLICE_X12Y148_AO5;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_A = CLBLM_L_X10Y148_SLICE_X13Y148_AO6;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_B = CLBLM_L_X10Y148_SLICE_X13Y148_BO6;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_C = CLBLM_L_X10Y148_SLICE_X13Y148_CO6;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_D = CLBLM_L_X10Y148_SLICE_X13Y148_DO6;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_CMUX = CLBLM_L_X10Y148_SLICE_X13Y148_CO5;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_A = CLBLM_L_X10Y149_SLICE_X12Y149_AO6;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_B = CLBLM_L_X10Y149_SLICE_X12Y149_BO6;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_C = CLBLM_L_X10Y149_SLICE_X12Y149_CO6;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_D = CLBLM_L_X10Y149_SLICE_X12Y149_DO6;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_AMUX = CLBLM_L_X10Y149_SLICE_X12Y149_AO5;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_BMUX = CLBLM_L_X10Y149_SLICE_X12Y149_BO5;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_A = CLBLM_L_X10Y149_SLICE_X13Y149_AO6;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_B = CLBLM_L_X10Y149_SLICE_X13Y149_BO6;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_C = CLBLM_L_X10Y149_SLICE_X13Y149_CO6;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_D = CLBLM_L_X10Y149_SLICE_X13Y149_DO6;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_AMUX = CLBLM_L_X10Y149_SLICE_X13Y149_A5Q;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_CMUX = CLBLM_L_X10Y149_SLICE_X13Y149_CO5;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_A = CLBLM_L_X10Y150_SLICE_X12Y150_AO6;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_B = CLBLM_L_X10Y150_SLICE_X12Y150_BO6;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_C = CLBLM_L_X10Y150_SLICE_X12Y150_CO6;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_D = CLBLM_L_X10Y150_SLICE_X12Y150_DO6;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_AMUX = CLBLM_L_X10Y150_SLICE_X12Y150_A5Q;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_BMUX = CLBLM_L_X10Y150_SLICE_X12Y150_B5Q;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_CMUX = CLBLM_L_X10Y150_SLICE_X12Y150_C5Q;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_A = CLBLM_L_X10Y150_SLICE_X13Y150_AO6;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_B = CLBLM_L_X10Y150_SLICE_X13Y150_BO6;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_C = CLBLM_L_X10Y150_SLICE_X13Y150_CO6;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_D = CLBLM_L_X10Y150_SLICE_X13Y150_DO6;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_AMUX = CLBLM_L_X10Y150_SLICE_X13Y150_A5Q;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_DMUX = CLBLM_L_X10Y150_SLICE_X13Y150_DO5;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_A = CLBLM_L_X10Y151_SLICE_X12Y151_AO6;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_B = CLBLM_L_X10Y151_SLICE_X12Y151_BO6;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_C = CLBLM_L_X10Y151_SLICE_X12Y151_CO6;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_D = CLBLM_L_X10Y151_SLICE_X12Y151_DO6;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_A = CLBLM_L_X10Y151_SLICE_X13Y151_AO6;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_B = CLBLM_L_X10Y151_SLICE_X13Y151_BO6;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_C = CLBLM_L_X10Y151_SLICE_X13Y151_CO6;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_D = CLBLM_L_X10Y151_SLICE_X13Y151_DO6;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_A = CLBLM_L_X10Y152_SLICE_X12Y152_AO6;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_B = CLBLM_L_X10Y152_SLICE_X12Y152_BO6;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_C = CLBLM_L_X10Y152_SLICE_X12Y152_CO6;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_D = CLBLM_L_X10Y152_SLICE_X12Y152_DO6;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_CMUX = CLBLM_L_X10Y152_SLICE_X12Y152_CO5;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_DMUX = CLBLM_L_X10Y152_SLICE_X12Y152_D5Q;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_A = CLBLM_L_X10Y152_SLICE_X13Y152_AO6;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_B = CLBLM_L_X10Y152_SLICE_X13Y152_BO6;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_C = CLBLM_L_X10Y152_SLICE_X13Y152_CO6;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_D = CLBLM_L_X10Y152_SLICE_X13Y152_DO6;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_CMUX = CLBLM_L_X10Y152_SLICE_X13Y152_CO5;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_A = CLBLM_L_X10Y153_SLICE_X12Y153_AO6;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_B = CLBLM_L_X10Y153_SLICE_X12Y153_BO6;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_C = CLBLM_L_X10Y153_SLICE_X12Y153_CO6;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_D = CLBLM_L_X10Y153_SLICE_X12Y153_DO6;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_A = CLBLM_L_X10Y153_SLICE_X13Y153_AO6;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_B = CLBLM_L_X10Y153_SLICE_X13Y153_BO6;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_C = CLBLM_L_X10Y153_SLICE_X13Y153_CO6;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_D = CLBLM_L_X10Y153_SLICE_X13Y153_DO6;
  assign CLBLM_L_X10Y154_SLICE_X12Y154_A = CLBLM_L_X10Y154_SLICE_X12Y154_AO6;
  assign CLBLM_L_X10Y154_SLICE_X12Y154_B = CLBLM_L_X10Y154_SLICE_X12Y154_BO6;
  assign CLBLM_L_X10Y154_SLICE_X12Y154_C = CLBLM_L_X10Y154_SLICE_X12Y154_CO6;
  assign CLBLM_L_X10Y154_SLICE_X12Y154_D = CLBLM_L_X10Y154_SLICE_X12Y154_DO6;
  assign CLBLM_L_X10Y154_SLICE_X13Y154_A = CLBLM_L_X10Y154_SLICE_X13Y154_AO6;
  assign CLBLM_L_X10Y154_SLICE_X13Y154_B = CLBLM_L_X10Y154_SLICE_X13Y154_BO6;
  assign CLBLM_L_X10Y154_SLICE_X13Y154_C = CLBLM_L_X10Y154_SLICE_X13Y154_CO6;
  assign CLBLM_L_X10Y154_SLICE_X13Y154_D = CLBLM_L_X10Y154_SLICE_X13Y154_DO6;
  assign CLBLM_L_X10Y154_SLICE_X13Y154_CMUX = CLBLM_L_X10Y154_SLICE_X13Y154_CO5;
  assign CLBLM_L_X10Y155_SLICE_X12Y155_A = CLBLM_L_X10Y155_SLICE_X12Y155_AO6;
  assign CLBLM_L_X10Y155_SLICE_X12Y155_B = CLBLM_L_X10Y155_SLICE_X12Y155_BO6;
  assign CLBLM_L_X10Y155_SLICE_X12Y155_C = CLBLM_L_X10Y155_SLICE_X12Y155_CO6;
  assign CLBLM_L_X10Y155_SLICE_X12Y155_D = CLBLM_L_X10Y155_SLICE_X12Y155_DO6;
  assign CLBLM_L_X10Y155_SLICE_X13Y155_A = CLBLM_L_X10Y155_SLICE_X13Y155_AO6;
  assign CLBLM_L_X10Y155_SLICE_X13Y155_B = CLBLM_L_X10Y155_SLICE_X13Y155_BO6;
  assign CLBLM_L_X10Y155_SLICE_X13Y155_C = CLBLM_L_X10Y155_SLICE_X13Y155_CO6;
  assign CLBLM_L_X10Y155_SLICE_X13Y155_D = CLBLM_L_X10Y155_SLICE_X13Y155_DO6;
  assign CLBLM_L_X10Y156_SLICE_X12Y156_A = CLBLM_L_X10Y156_SLICE_X12Y156_AO6;
  assign CLBLM_L_X10Y156_SLICE_X12Y156_B = CLBLM_L_X10Y156_SLICE_X12Y156_BO6;
  assign CLBLM_L_X10Y156_SLICE_X12Y156_C = CLBLM_L_X10Y156_SLICE_X12Y156_CO6;
  assign CLBLM_L_X10Y156_SLICE_X12Y156_D = CLBLM_L_X10Y156_SLICE_X12Y156_DO6;
  assign CLBLM_L_X10Y156_SLICE_X12Y156_AMUX = CLBLM_L_X10Y156_SLICE_X12Y156_AO5;
  assign CLBLM_L_X10Y156_SLICE_X13Y156_A = CLBLM_L_X10Y156_SLICE_X13Y156_AO6;
  assign CLBLM_L_X10Y156_SLICE_X13Y156_B = CLBLM_L_X10Y156_SLICE_X13Y156_BO6;
  assign CLBLM_L_X10Y156_SLICE_X13Y156_C = CLBLM_L_X10Y156_SLICE_X13Y156_CO6;
  assign CLBLM_L_X10Y156_SLICE_X13Y156_D = CLBLM_L_X10Y156_SLICE_X13Y156_DO6;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_A = CLBLM_L_X12Y144_SLICE_X16Y144_AO6;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_B = CLBLM_L_X12Y144_SLICE_X16Y144_BO6;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_C = CLBLM_L_X12Y144_SLICE_X16Y144_CO6;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_D = CLBLM_L_X12Y144_SLICE_X16Y144_DO6;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_AMUX = CLBLM_L_X12Y144_SLICE_X16Y144_AO5;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_DMUX = CLBLM_L_X12Y144_SLICE_X16Y144_DO5;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_A = CLBLM_L_X12Y144_SLICE_X17Y144_AO6;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_B = CLBLM_L_X12Y144_SLICE_X17Y144_BO6;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_C = CLBLM_L_X12Y144_SLICE_X17Y144_CO6;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_D = CLBLM_L_X12Y144_SLICE_X17Y144_DO6;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_A = CLBLM_L_X12Y145_SLICE_X16Y145_AO6;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_B = CLBLM_L_X12Y145_SLICE_X16Y145_BO6;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_C = CLBLM_L_X12Y145_SLICE_X16Y145_CO6;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_D = CLBLM_L_X12Y145_SLICE_X16Y145_DO6;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_CMUX = CLBLM_L_X12Y145_SLICE_X16Y145_CO5;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_A = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_B = CLBLM_L_X12Y145_SLICE_X17Y145_BO6;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_C = CLBLM_L_X12Y145_SLICE_X17Y145_CO6;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_D = CLBLM_L_X12Y145_SLICE_X17Y145_DO6;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_A = CLBLM_L_X12Y146_SLICE_X16Y146_AO6;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_B = CLBLM_L_X12Y146_SLICE_X16Y146_BO6;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_C = CLBLM_L_X12Y146_SLICE_X16Y146_CO6;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_D = CLBLM_L_X12Y146_SLICE_X16Y146_DO6;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_A = CLBLM_L_X12Y146_SLICE_X17Y146_AO6;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_B = CLBLM_L_X12Y146_SLICE_X17Y146_BO6;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_C = CLBLM_L_X12Y146_SLICE_X17Y146_CO6;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_D = CLBLM_L_X12Y146_SLICE_X17Y146_DO6;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_A = CLBLM_L_X12Y147_SLICE_X16Y147_AO6;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_B = CLBLM_L_X12Y147_SLICE_X16Y147_BO6;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_C = CLBLM_L_X12Y147_SLICE_X16Y147_CO6;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_D = CLBLM_L_X12Y147_SLICE_X16Y147_DO6;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_A = CLBLM_L_X12Y147_SLICE_X17Y147_AO6;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_B = CLBLM_L_X12Y147_SLICE_X17Y147_BO6;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_C = CLBLM_L_X12Y147_SLICE_X17Y147_CO6;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_D = CLBLM_L_X12Y147_SLICE_X17Y147_DO6;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_A = CLBLM_L_X12Y148_SLICE_X16Y148_AO6;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_B = CLBLM_L_X12Y148_SLICE_X16Y148_BO6;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_C = CLBLM_L_X12Y148_SLICE_X16Y148_CO6;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_D = CLBLM_L_X12Y148_SLICE_X16Y148_DO6;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_A = CLBLM_L_X12Y148_SLICE_X17Y148_AO6;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_B = CLBLM_L_X12Y148_SLICE_X17Y148_BO6;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_C = CLBLM_L_X12Y148_SLICE_X17Y148_CO6;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_D = CLBLM_L_X12Y148_SLICE_X17Y148_DO6;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_A = CLBLM_L_X12Y149_SLICE_X16Y149_AO6;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_B = CLBLM_L_X12Y149_SLICE_X16Y149_BO6;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_C = CLBLM_L_X12Y149_SLICE_X16Y149_CO6;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_D = CLBLM_L_X12Y149_SLICE_X16Y149_DO6;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_A = CLBLM_L_X12Y149_SLICE_X17Y149_AO6;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_B = CLBLM_L_X12Y149_SLICE_X17Y149_BO6;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_C = CLBLM_L_X12Y149_SLICE_X17Y149_CO6;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_D = CLBLM_L_X12Y149_SLICE_X17Y149_DO6;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_A = CLBLM_L_X12Y150_SLICE_X16Y150_AO6;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_B = CLBLM_L_X12Y150_SLICE_X16Y150_BO6;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_C = CLBLM_L_X12Y150_SLICE_X16Y150_CO6;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_D = CLBLM_L_X12Y150_SLICE_X16Y150_DO6;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_DMUX = CLBLM_L_X12Y150_SLICE_X16Y150_DO5;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_A = CLBLM_L_X12Y150_SLICE_X17Y150_AO6;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_B = CLBLM_L_X12Y150_SLICE_X17Y150_BO6;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_C = CLBLM_L_X12Y150_SLICE_X17Y150_CO6;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_D = CLBLM_L_X12Y150_SLICE_X17Y150_DO6;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_A = CLBLM_L_X12Y151_SLICE_X16Y151_AO6;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_B = CLBLM_L_X12Y151_SLICE_X16Y151_BO6;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_C = CLBLM_L_X12Y151_SLICE_X16Y151_CO6;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_D = CLBLM_L_X12Y151_SLICE_X16Y151_DO6;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_DMUX = CLBLM_L_X12Y151_SLICE_X16Y151_DO5;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_A = CLBLM_L_X12Y151_SLICE_X17Y151_AO6;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_B = CLBLM_L_X12Y151_SLICE_X17Y151_BO6;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_C = CLBLM_L_X12Y151_SLICE_X17Y151_CO6;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_D = CLBLM_L_X12Y151_SLICE_X17Y151_DO6;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_A = CLBLM_L_X12Y152_SLICE_X16Y152_AO6;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_B = CLBLM_L_X12Y152_SLICE_X16Y152_BO6;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_C = CLBLM_L_X12Y152_SLICE_X16Y152_CO6;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_D = CLBLM_L_X12Y152_SLICE_X16Y152_DO6;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_A = CLBLM_L_X12Y152_SLICE_X17Y152_AO6;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_B = CLBLM_L_X12Y152_SLICE_X17Y152_BO6;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_C = CLBLM_L_X12Y152_SLICE_X17Y152_CO6;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_D = CLBLM_L_X12Y152_SLICE_X17Y152_DO6;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_A = CLBLM_L_X12Y153_SLICE_X16Y153_AO6;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_B = CLBLM_L_X12Y153_SLICE_X16Y153_BO6;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_C = CLBLM_L_X12Y153_SLICE_X16Y153_CO6;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_D = CLBLM_L_X12Y153_SLICE_X16Y153_DO6;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_A = CLBLM_L_X12Y153_SLICE_X17Y153_AO6;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_B = CLBLM_L_X12Y153_SLICE_X17Y153_BO6;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_C = CLBLM_L_X12Y153_SLICE_X17Y153_CO6;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_D = CLBLM_L_X12Y153_SLICE_X17Y153_DO6;
  assign CLBLM_L_X12Y154_SLICE_X16Y154_A = CLBLM_L_X12Y154_SLICE_X16Y154_AO6;
  assign CLBLM_L_X12Y154_SLICE_X16Y154_B = CLBLM_L_X12Y154_SLICE_X16Y154_BO6;
  assign CLBLM_L_X12Y154_SLICE_X16Y154_C = CLBLM_L_X12Y154_SLICE_X16Y154_CO6;
  assign CLBLM_L_X12Y154_SLICE_X16Y154_D = CLBLM_L_X12Y154_SLICE_X16Y154_DO6;
  assign CLBLM_L_X12Y154_SLICE_X16Y154_BMUX = CLBLM_L_X12Y154_SLICE_X16Y154_BO5;
  assign CLBLM_L_X12Y154_SLICE_X17Y154_A = CLBLM_L_X12Y154_SLICE_X17Y154_AO6;
  assign CLBLM_L_X12Y154_SLICE_X17Y154_B = CLBLM_L_X12Y154_SLICE_X17Y154_BO6;
  assign CLBLM_L_X12Y154_SLICE_X17Y154_C = CLBLM_L_X12Y154_SLICE_X17Y154_CO6;
  assign CLBLM_L_X12Y154_SLICE_X17Y154_D = CLBLM_L_X12Y154_SLICE_X17Y154_DO6;
  assign CLBLM_L_X12Y155_SLICE_X16Y155_A = CLBLM_L_X12Y155_SLICE_X16Y155_AO6;
  assign CLBLM_L_X12Y155_SLICE_X16Y155_B = CLBLM_L_X12Y155_SLICE_X16Y155_BO6;
  assign CLBLM_L_X12Y155_SLICE_X16Y155_C = CLBLM_L_X12Y155_SLICE_X16Y155_CO6;
  assign CLBLM_L_X12Y155_SLICE_X16Y155_D = CLBLM_L_X12Y155_SLICE_X16Y155_DO6;
  assign CLBLM_L_X12Y155_SLICE_X17Y155_A = CLBLM_L_X12Y155_SLICE_X17Y155_AO6;
  assign CLBLM_L_X12Y155_SLICE_X17Y155_B = CLBLM_L_X12Y155_SLICE_X17Y155_BO6;
  assign CLBLM_L_X12Y155_SLICE_X17Y155_C = CLBLM_L_X12Y155_SLICE_X17Y155_CO6;
  assign CLBLM_L_X12Y155_SLICE_X17Y155_D = CLBLM_L_X12Y155_SLICE_X17Y155_DO6;
  assign CLBLM_L_X16Y158_SLICE_X22Y158_A = CLBLM_L_X16Y158_SLICE_X22Y158_AO6;
  assign CLBLM_L_X16Y158_SLICE_X22Y158_B = CLBLM_L_X16Y158_SLICE_X22Y158_BO6;
  assign CLBLM_L_X16Y158_SLICE_X22Y158_C = CLBLM_L_X16Y158_SLICE_X22Y158_CO6;
  assign CLBLM_L_X16Y158_SLICE_X22Y158_D = CLBLM_L_X16Y158_SLICE_X22Y158_DO6;
  assign CLBLM_L_X16Y158_SLICE_X22Y158_AMUX = CLBLM_L_X16Y158_SLICE_X22Y158_AO5;
  assign CLBLM_L_X16Y158_SLICE_X23Y158_A = CLBLM_L_X16Y158_SLICE_X23Y158_AO6;
  assign CLBLM_L_X16Y158_SLICE_X23Y158_B = CLBLM_L_X16Y158_SLICE_X23Y158_BO6;
  assign CLBLM_L_X16Y158_SLICE_X23Y158_C = CLBLM_L_X16Y158_SLICE_X23Y158_CO6;
  assign CLBLM_L_X16Y158_SLICE_X23Y158_D = CLBLM_L_X16Y158_SLICE_X23Y158_DO6;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_A = CLBLM_R_X3Y141_SLICE_X2Y141_AO6;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_B = CLBLM_R_X3Y141_SLICE_X2Y141_BO6;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_C = CLBLM_R_X3Y141_SLICE_X2Y141_CO6;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_D = CLBLM_R_X3Y141_SLICE_X2Y141_DO6;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_A = CLBLM_R_X3Y141_SLICE_X3Y141_AO6;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_B = CLBLM_R_X3Y141_SLICE_X3Y141_BO6;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_C = CLBLM_R_X3Y141_SLICE_X3Y141_CO6;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_D = CLBLM_R_X3Y141_SLICE_X3Y141_DO6;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_A = CLBLM_R_X3Y142_SLICE_X2Y142_AO6;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_B = CLBLM_R_X3Y142_SLICE_X2Y142_BO6;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_C = CLBLM_R_X3Y142_SLICE_X2Y142_CO6;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_D = CLBLM_R_X3Y142_SLICE_X2Y142_DO6;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_DMUX = CLBLM_R_X3Y142_SLICE_X2Y142_DO5;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_A = CLBLM_R_X3Y142_SLICE_X3Y142_AO6;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_B = CLBLM_R_X3Y142_SLICE_X3Y142_BO6;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_C = CLBLM_R_X3Y142_SLICE_X3Y142_CO6;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_D = CLBLM_R_X3Y142_SLICE_X3Y142_DO6;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_A = CLBLM_R_X3Y143_SLICE_X2Y143_AO6;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_B = CLBLM_R_X3Y143_SLICE_X2Y143_BO6;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_C = CLBLM_R_X3Y143_SLICE_X2Y143_CO6;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_D = CLBLM_R_X3Y143_SLICE_X2Y143_DO6;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_A = CLBLM_R_X3Y143_SLICE_X3Y143_AO6;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_B = CLBLM_R_X3Y143_SLICE_X3Y143_BO6;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_C = CLBLM_R_X3Y143_SLICE_X3Y143_CO6;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_D = CLBLM_R_X3Y143_SLICE_X3Y143_DO6;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_AMUX = CLBLM_R_X3Y143_SLICE_X3Y143_A5Q;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_BMUX = CLBLM_R_X3Y143_SLICE_X3Y143_B5Q;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_CMUX = CLBLM_R_X3Y143_SLICE_X3Y143_CO5;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_DMUX = CLBLM_R_X3Y143_SLICE_X3Y143_DO5;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_A = CLBLM_R_X3Y144_SLICE_X2Y144_AO6;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_B = CLBLM_R_X3Y144_SLICE_X2Y144_BO6;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_C = CLBLM_R_X3Y144_SLICE_X2Y144_CO6;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_D = CLBLM_R_X3Y144_SLICE_X2Y144_DO6;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_AMUX = CLBLM_R_X3Y144_SLICE_X2Y144_A5Q;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_BMUX = CLBLM_R_X3Y144_SLICE_X2Y144_B5Q;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_A = CLBLM_R_X3Y144_SLICE_X3Y144_AO6;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_B = CLBLM_R_X3Y144_SLICE_X3Y144_BO6;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_C = CLBLM_R_X3Y144_SLICE_X3Y144_CO6;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_D = CLBLM_R_X3Y144_SLICE_X3Y144_DO6;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_BMUX = CLBLM_R_X3Y144_SLICE_X3Y144_BO5;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_A = CLBLM_R_X3Y145_SLICE_X2Y145_AO6;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_B = CLBLM_R_X3Y145_SLICE_X2Y145_BO6;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_C = CLBLM_R_X3Y145_SLICE_X2Y145_CO6;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_D = CLBLM_R_X3Y145_SLICE_X2Y145_DO6;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_AMUX = CLBLM_R_X3Y145_SLICE_X2Y145_A5Q;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_CMUX = CLBLM_R_X3Y145_SLICE_X2Y145_CO5;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_A = CLBLM_R_X3Y145_SLICE_X3Y145_AO6;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_B = CLBLM_R_X3Y145_SLICE_X3Y145_BO6;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_C = CLBLM_R_X3Y145_SLICE_X3Y145_CO6;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_D = CLBLM_R_X3Y145_SLICE_X3Y145_DO6;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_AMUX = CLBLM_R_X3Y145_SLICE_X3Y145_A5Q;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_DMUX = CLBLM_R_X3Y145_SLICE_X3Y145_D5Q;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_A = CLBLM_R_X3Y146_SLICE_X2Y146_AO6;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_B = CLBLM_R_X3Y146_SLICE_X2Y146_BO6;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_C = CLBLM_R_X3Y146_SLICE_X2Y146_CO6;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_D = CLBLM_R_X3Y146_SLICE_X2Y146_DO6;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_A = CLBLM_R_X3Y146_SLICE_X3Y146_AO6;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_B = CLBLM_R_X3Y146_SLICE_X3Y146_BO6;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_C = CLBLM_R_X3Y146_SLICE_X3Y146_CO6;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_D = CLBLM_R_X3Y146_SLICE_X3Y146_DO6;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_DMUX = CLBLM_R_X3Y146_SLICE_X3Y146_DO5;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_A = CLBLM_R_X3Y147_SLICE_X2Y147_AO6;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_B = CLBLM_R_X3Y147_SLICE_X2Y147_BO6;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_C = CLBLM_R_X3Y147_SLICE_X2Y147_CO6;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_D = CLBLM_R_X3Y147_SLICE_X2Y147_DO6;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_AMUX = CLBLM_R_X3Y147_SLICE_X2Y147_A5Q;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_BMUX = CLBLM_R_X3Y147_SLICE_X2Y147_BO5;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_A = CLBLM_R_X3Y147_SLICE_X3Y147_AO6;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_B = CLBLM_R_X3Y147_SLICE_X3Y147_BO6;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_C = CLBLM_R_X3Y147_SLICE_X3Y147_CO6;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_D = CLBLM_R_X3Y147_SLICE_X3Y147_DO6;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_CMUX = CLBLM_R_X3Y147_SLICE_X3Y147_C5Q;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_A = CLBLM_R_X3Y148_SLICE_X2Y148_AO6;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_B = CLBLM_R_X3Y148_SLICE_X2Y148_BO6;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_C = CLBLM_R_X3Y148_SLICE_X2Y148_CO6;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_D = CLBLM_R_X3Y148_SLICE_X2Y148_DO6;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_AMUX = CLBLM_R_X3Y148_SLICE_X2Y148_AO5;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_A = CLBLM_R_X3Y148_SLICE_X3Y148_AO6;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_B = CLBLM_R_X3Y148_SLICE_X3Y148_BO6;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_C = CLBLM_R_X3Y148_SLICE_X3Y148_CO6;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_D = CLBLM_R_X3Y148_SLICE_X3Y148_DO6;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_BMUX = CLBLM_R_X3Y148_SLICE_X3Y148_B5Q;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_DMUX = CLBLM_R_X3Y148_SLICE_X3Y148_DO6;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_A = CLBLM_R_X3Y149_SLICE_X2Y149_AO6;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_B = CLBLM_R_X3Y149_SLICE_X2Y149_BO6;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_C = CLBLM_R_X3Y149_SLICE_X2Y149_CO6;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_D = CLBLM_R_X3Y149_SLICE_X2Y149_DO6;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_A = CLBLM_R_X3Y149_SLICE_X3Y149_AO6;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_B = CLBLM_R_X3Y149_SLICE_X3Y149_BO6;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_C = CLBLM_R_X3Y149_SLICE_X3Y149_CO6;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_D = CLBLM_R_X3Y149_SLICE_X3Y149_DO6;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_BMUX = CLBLM_R_X3Y149_SLICE_X3Y149_B5Q;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_A = CLBLM_R_X3Y150_SLICE_X2Y150_AO6;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_B = CLBLM_R_X3Y150_SLICE_X2Y150_BO6;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_C = CLBLM_R_X3Y150_SLICE_X2Y150_CO6;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_D = CLBLM_R_X3Y150_SLICE_X2Y150_DO6;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_A = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_B = CLBLM_R_X3Y150_SLICE_X3Y150_BO6;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_C = CLBLM_R_X3Y150_SLICE_X3Y150_CO6;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_D = CLBLM_R_X3Y150_SLICE_X3Y150_DO6;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_AMUX = CLBLM_R_X3Y150_SLICE_X3Y150_A5Q;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_A = CLBLM_R_X3Y151_SLICE_X2Y151_AO6;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_B = CLBLM_R_X3Y151_SLICE_X2Y151_BO6;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_C = CLBLM_R_X3Y151_SLICE_X2Y151_CO6;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_D = CLBLM_R_X3Y151_SLICE_X2Y151_DO6;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_CMUX = CLBLM_R_X3Y151_SLICE_X2Y151_CO6;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_A = CLBLM_R_X3Y151_SLICE_X3Y151_AO6;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_B = CLBLM_R_X3Y151_SLICE_X3Y151_BO6;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_C = CLBLM_R_X3Y151_SLICE_X3Y151_CO6;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_D = CLBLM_R_X3Y151_SLICE_X3Y151_DO6;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_A = CLBLM_R_X3Y152_SLICE_X2Y152_AO6;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_B = CLBLM_R_X3Y152_SLICE_X2Y152_BO6;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_C = CLBLM_R_X3Y152_SLICE_X2Y152_CO6;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_D = CLBLM_R_X3Y152_SLICE_X2Y152_DO6;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_AMUX = CLBLM_R_X3Y152_SLICE_X2Y152_AO5;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_BMUX = CLBLM_R_X3Y152_SLICE_X2Y152_BO5;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_A = CLBLM_R_X3Y152_SLICE_X3Y152_AO6;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_B = CLBLM_R_X3Y152_SLICE_X3Y152_BO6;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_C = CLBLM_R_X3Y152_SLICE_X3Y152_CO6;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_D = CLBLM_R_X3Y152_SLICE_X3Y152_DO6;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_CMUX = CLBLM_R_X3Y152_SLICE_X3Y152_CO6;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_A = CLBLM_R_X3Y153_SLICE_X2Y153_AO6;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_B = CLBLM_R_X3Y153_SLICE_X2Y153_BO6;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_C = CLBLM_R_X3Y153_SLICE_X2Y153_CO6;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_D = CLBLM_R_X3Y153_SLICE_X2Y153_DO6;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_A = CLBLM_R_X3Y153_SLICE_X3Y153_AO6;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_B = CLBLM_R_X3Y153_SLICE_X3Y153_BO6;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_C = CLBLM_R_X3Y153_SLICE_X3Y153_CO6;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_D = CLBLM_R_X3Y153_SLICE_X3Y153_DO6;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_CMUX = CLBLM_R_X3Y153_SLICE_X3Y153_CO6;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_A = CLBLM_R_X3Y154_SLICE_X2Y154_AO6;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_B = CLBLM_R_X3Y154_SLICE_X2Y154_BO6;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_C = CLBLM_R_X3Y154_SLICE_X2Y154_CO6;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_D = CLBLM_R_X3Y154_SLICE_X2Y154_DO6;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_A = CLBLM_R_X3Y154_SLICE_X3Y154_AO6;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_B = CLBLM_R_X3Y154_SLICE_X3Y154_BO6;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_C = CLBLM_R_X3Y154_SLICE_X3Y154_CO6;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_D = CLBLM_R_X3Y154_SLICE_X3Y154_DO6;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_CMUX = CLBLM_R_X3Y154_SLICE_X3Y154_CO6;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_A = CLBLM_R_X3Y155_SLICE_X2Y155_AO6;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_B = CLBLM_R_X3Y155_SLICE_X2Y155_BO6;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_C = CLBLM_R_X3Y155_SLICE_X2Y155_CO6;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_D = CLBLM_R_X3Y155_SLICE_X2Y155_DO6;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_DMUX = CLBLM_R_X3Y155_SLICE_X2Y155_DO6;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_A = CLBLM_R_X3Y155_SLICE_X3Y155_AO6;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_B = CLBLM_R_X3Y155_SLICE_X3Y155_BO6;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_C = CLBLM_R_X3Y155_SLICE_X3Y155_CO6;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_D = CLBLM_R_X3Y155_SLICE_X3Y155_DO6;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_AMUX = CLBLM_R_X3Y155_SLICE_X3Y155_AO5;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_CMUX = CLBLM_R_X3Y155_SLICE_X3Y155_CO6;
  assign CLBLM_R_X3Y156_SLICE_X2Y156_A = CLBLM_R_X3Y156_SLICE_X2Y156_AO6;
  assign CLBLM_R_X3Y156_SLICE_X2Y156_B = CLBLM_R_X3Y156_SLICE_X2Y156_BO6;
  assign CLBLM_R_X3Y156_SLICE_X2Y156_C = CLBLM_R_X3Y156_SLICE_X2Y156_CO6;
  assign CLBLM_R_X3Y156_SLICE_X2Y156_D = CLBLM_R_X3Y156_SLICE_X2Y156_DO6;
  assign CLBLM_R_X3Y156_SLICE_X2Y156_AMUX = CLBLM_R_X3Y156_SLICE_X2Y156_AO5;
  assign CLBLM_R_X3Y156_SLICE_X3Y156_A = CLBLM_R_X3Y156_SLICE_X3Y156_AO6;
  assign CLBLM_R_X3Y156_SLICE_X3Y156_B = CLBLM_R_X3Y156_SLICE_X3Y156_BO6;
  assign CLBLM_R_X3Y156_SLICE_X3Y156_C = CLBLM_R_X3Y156_SLICE_X3Y156_CO6;
  assign CLBLM_R_X3Y156_SLICE_X3Y156_D = CLBLM_R_X3Y156_SLICE_X3Y156_DO6;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_A = CLBLM_R_X5Y142_SLICE_X6Y142_AO6;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_B = CLBLM_R_X5Y142_SLICE_X6Y142_BO6;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_C = CLBLM_R_X5Y142_SLICE_X6Y142_CO6;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_D = CLBLM_R_X5Y142_SLICE_X6Y142_DO6;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_A = CLBLM_R_X5Y142_SLICE_X7Y142_AO6;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_B = CLBLM_R_X5Y142_SLICE_X7Y142_BO6;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_C = CLBLM_R_X5Y142_SLICE_X7Y142_CO6;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_D = CLBLM_R_X5Y142_SLICE_X7Y142_DO6;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_A = CLBLM_R_X5Y143_SLICE_X6Y143_AO6;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_B = CLBLM_R_X5Y143_SLICE_X6Y143_BO6;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_C = CLBLM_R_X5Y143_SLICE_X6Y143_CO6;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_D = CLBLM_R_X5Y143_SLICE_X6Y143_DO6;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_A = CLBLM_R_X5Y143_SLICE_X7Y143_AO6;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_B = CLBLM_R_X5Y143_SLICE_X7Y143_BO6;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_C = CLBLM_R_X5Y143_SLICE_X7Y143_CO6;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_D = CLBLM_R_X5Y143_SLICE_X7Y143_DO6;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_BMUX = CLBLM_R_X5Y143_SLICE_X7Y143_BO5;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_A = CLBLM_R_X5Y144_SLICE_X6Y144_AO6;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_B = CLBLM_R_X5Y144_SLICE_X6Y144_BO6;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_C = CLBLM_R_X5Y144_SLICE_X6Y144_CO6;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_D = CLBLM_R_X5Y144_SLICE_X6Y144_DO6;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_BMUX = CLBLM_R_X5Y144_SLICE_X6Y144_BO5;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_A = CLBLM_R_X5Y144_SLICE_X7Y144_AO6;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_B = CLBLM_R_X5Y144_SLICE_X7Y144_BO6;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_C = CLBLM_R_X5Y144_SLICE_X7Y144_CO6;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_D = CLBLM_R_X5Y144_SLICE_X7Y144_DO6;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_BMUX = CLBLM_R_X5Y144_SLICE_X7Y144_B5Q;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_A = CLBLM_R_X5Y145_SLICE_X6Y145_AO6;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_B = CLBLM_R_X5Y145_SLICE_X6Y145_BO6;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_C = CLBLM_R_X5Y145_SLICE_X6Y145_CO6;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_D = CLBLM_R_X5Y145_SLICE_X6Y145_DO6;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_AMUX = CLBLM_R_X5Y145_SLICE_X6Y145_A5Q;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_BMUX = CLBLM_R_X5Y145_SLICE_X6Y145_BO5;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_DMUX = CLBLM_R_X5Y145_SLICE_X6Y145_DO5;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_A = CLBLM_R_X5Y145_SLICE_X7Y145_AO6;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_B = CLBLM_R_X5Y145_SLICE_X7Y145_BO6;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_C = CLBLM_R_X5Y145_SLICE_X7Y145_CO6;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_D = CLBLM_R_X5Y145_SLICE_X7Y145_DO6;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_DMUX = CLBLM_R_X5Y145_SLICE_X7Y145_DO5;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_A = CLBLM_R_X5Y146_SLICE_X6Y146_AO6;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_B = CLBLM_R_X5Y146_SLICE_X6Y146_BO6;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_C = CLBLM_R_X5Y146_SLICE_X6Y146_CO6;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_D = CLBLM_R_X5Y146_SLICE_X6Y146_DO6;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_AMUX = CLBLM_R_X5Y146_SLICE_X6Y146_A5Q;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_BMUX = CLBLM_R_X5Y146_SLICE_X6Y146_BO5;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_A = CLBLM_R_X5Y146_SLICE_X7Y146_AO6;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_B = CLBLM_R_X5Y146_SLICE_X7Y146_BO6;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_C = CLBLM_R_X5Y146_SLICE_X7Y146_CO6;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_D = CLBLM_R_X5Y146_SLICE_X7Y146_DO6;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_AMUX = CLBLM_R_X5Y146_SLICE_X7Y146_AO5;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_CMUX = CLBLM_R_X5Y146_SLICE_X7Y146_CO6;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_DMUX = CLBLM_R_X5Y146_SLICE_X7Y146_DO6;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_A = CLBLM_R_X5Y147_SLICE_X6Y147_AO6;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_B = CLBLM_R_X5Y147_SLICE_X6Y147_BO6;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_C = CLBLM_R_X5Y147_SLICE_X6Y147_CO6;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_D = CLBLM_R_X5Y147_SLICE_X6Y147_DO6;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_A = CLBLM_R_X5Y147_SLICE_X7Y147_AO6;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_B = CLBLM_R_X5Y147_SLICE_X7Y147_BO6;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_C = CLBLM_R_X5Y147_SLICE_X7Y147_CO6;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_D = CLBLM_R_X5Y147_SLICE_X7Y147_DO6;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_DMUX = CLBLM_R_X5Y147_SLICE_X7Y147_D5Q;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_A = CLBLM_R_X5Y148_SLICE_X6Y148_AO6;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_B = CLBLM_R_X5Y148_SLICE_X6Y148_BO6;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_C = CLBLM_R_X5Y148_SLICE_X6Y148_CO6;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_D = CLBLM_R_X5Y148_SLICE_X6Y148_DO6;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_A = CLBLM_R_X5Y148_SLICE_X7Y148_AO6;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_B = CLBLM_R_X5Y148_SLICE_X7Y148_BO6;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_C = CLBLM_R_X5Y148_SLICE_X7Y148_CO6;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_D = CLBLM_R_X5Y148_SLICE_X7Y148_DO6;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_CMUX = CLBLM_R_X5Y148_SLICE_X7Y148_C5Q;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_A = CLBLM_R_X5Y149_SLICE_X6Y149_AO6;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_B = CLBLM_R_X5Y149_SLICE_X6Y149_BO6;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_C = CLBLM_R_X5Y149_SLICE_X6Y149_CO6;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_D = CLBLM_R_X5Y149_SLICE_X6Y149_DO6;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_CMUX = CLBLM_R_X5Y149_SLICE_X6Y149_CO5;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_A = CLBLM_R_X5Y149_SLICE_X7Y149_AO6;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_B = CLBLM_R_X5Y149_SLICE_X7Y149_BO6;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_C = CLBLM_R_X5Y149_SLICE_X7Y149_CO6;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_D = CLBLM_R_X5Y149_SLICE_X7Y149_DO6;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_A = CLBLM_R_X5Y150_SLICE_X6Y150_AO6;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_B = CLBLM_R_X5Y150_SLICE_X6Y150_BO6;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_C = CLBLM_R_X5Y150_SLICE_X6Y150_CO6;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_D = CLBLM_R_X5Y150_SLICE_X6Y150_DO6;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_AMUX = CLBLM_R_X5Y150_SLICE_X6Y150_A5Q;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_A = CLBLM_R_X5Y150_SLICE_X7Y150_AO6;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_B = CLBLM_R_X5Y150_SLICE_X7Y150_BO6;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_C = CLBLM_R_X5Y150_SLICE_X7Y150_CO6;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_D = CLBLM_R_X5Y150_SLICE_X7Y150_DO6;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_DMUX = CLBLM_R_X5Y150_SLICE_X7Y150_DO6;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_A = CLBLM_R_X5Y151_SLICE_X6Y151_AO6;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_B = CLBLM_R_X5Y151_SLICE_X6Y151_BO6;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_C = CLBLM_R_X5Y151_SLICE_X6Y151_CO6;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_D = CLBLM_R_X5Y151_SLICE_X6Y151_DO6;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_A = CLBLM_R_X5Y151_SLICE_X7Y151_AO6;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_B = CLBLM_R_X5Y151_SLICE_X7Y151_BO6;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_C = CLBLM_R_X5Y151_SLICE_X7Y151_CO6;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_D = CLBLM_R_X5Y151_SLICE_X7Y151_DO6;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_DMUX = CLBLM_R_X5Y151_SLICE_X7Y151_DO5;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_A = CLBLM_R_X5Y152_SLICE_X6Y152_AO6;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_B = CLBLM_R_X5Y152_SLICE_X6Y152_BO6;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_C = CLBLM_R_X5Y152_SLICE_X6Y152_CO6;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_D = CLBLM_R_X5Y152_SLICE_X6Y152_DO6;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_AMUX = CLBLM_R_X5Y152_SLICE_X6Y152_A5Q;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_A = CLBLM_R_X5Y152_SLICE_X7Y152_AO6;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_B = CLBLM_R_X5Y152_SLICE_X7Y152_BO6;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_C = CLBLM_R_X5Y152_SLICE_X7Y152_CO6;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_D = CLBLM_R_X5Y152_SLICE_X7Y152_DO6;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_BMUX = CLBLM_R_X5Y152_SLICE_X7Y152_B5Q;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_DMUX = CLBLM_R_X5Y152_SLICE_X7Y152_DO5;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_A = CLBLM_R_X5Y153_SLICE_X6Y153_AO6;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_B = CLBLM_R_X5Y153_SLICE_X6Y153_BO6;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_C = CLBLM_R_X5Y153_SLICE_X6Y153_CO6;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_D = CLBLM_R_X5Y153_SLICE_X6Y153_DO6;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_AMUX = CLBLM_R_X5Y153_SLICE_X6Y153_A5Q;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_CMUX = CLBLM_R_X5Y153_SLICE_X6Y153_CO5;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_A = CLBLM_R_X5Y153_SLICE_X7Y153_AO6;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_B = CLBLM_R_X5Y153_SLICE_X7Y153_BO6;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_C = CLBLM_R_X5Y153_SLICE_X7Y153_CO6;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_D = CLBLM_R_X5Y153_SLICE_X7Y153_DO6;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_A = CLBLM_R_X5Y154_SLICE_X6Y154_AO6;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_B = CLBLM_R_X5Y154_SLICE_X6Y154_BO6;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_C = CLBLM_R_X5Y154_SLICE_X6Y154_CO6;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_D = CLBLM_R_X5Y154_SLICE_X6Y154_DO6;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_A = CLBLM_R_X5Y154_SLICE_X7Y154_AO6;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_B = CLBLM_R_X5Y154_SLICE_X7Y154_BO6;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_C = CLBLM_R_X5Y154_SLICE_X7Y154_CO6;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_D = CLBLM_R_X5Y154_SLICE_X7Y154_DO6;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_AMUX = CLBLM_R_X5Y154_SLICE_X7Y154_AO5;
  assign CLBLM_R_X5Y155_SLICE_X6Y155_A = CLBLM_R_X5Y155_SLICE_X6Y155_AO6;
  assign CLBLM_R_X5Y155_SLICE_X6Y155_B = CLBLM_R_X5Y155_SLICE_X6Y155_BO6;
  assign CLBLM_R_X5Y155_SLICE_X6Y155_C = CLBLM_R_X5Y155_SLICE_X6Y155_CO6;
  assign CLBLM_R_X5Y155_SLICE_X6Y155_D = CLBLM_R_X5Y155_SLICE_X6Y155_DO6;
  assign CLBLM_R_X5Y155_SLICE_X7Y155_A = CLBLM_R_X5Y155_SLICE_X7Y155_AO6;
  assign CLBLM_R_X5Y155_SLICE_X7Y155_B = CLBLM_R_X5Y155_SLICE_X7Y155_BO6;
  assign CLBLM_R_X5Y155_SLICE_X7Y155_C = CLBLM_R_X5Y155_SLICE_X7Y155_CO6;
  assign CLBLM_R_X5Y155_SLICE_X7Y155_D = CLBLM_R_X5Y155_SLICE_X7Y155_DO6;
  assign CLBLM_R_X5Y155_SLICE_X7Y155_BMUX = CLBLM_R_X5Y155_SLICE_X7Y155_BO5;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_A = CLBLM_R_X7Y142_SLICE_X8Y142_AO6;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_B = CLBLM_R_X7Y142_SLICE_X8Y142_BO6;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_C = CLBLM_R_X7Y142_SLICE_X8Y142_CO6;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_D = CLBLM_R_X7Y142_SLICE_X8Y142_DO6;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_AMUX = CLBLM_R_X7Y142_SLICE_X8Y142_AO5;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_DMUX = CLBLM_R_X7Y142_SLICE_X8Y142_DO6;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_A = CLBLM_R_X7Y142_SLICE_X9Y142_AO6;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_B = CLBLM_R_X7Y142_SLICE_X9Y142_BO6;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_C = CLBLM_R_X7Y142_SLICE_X9Y142_CO6;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_D = CLBLM_R_X7Y142_SLICE_X9Y142_DO6;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_A = CLBLM_R_X7Y143_SLICE_X8Y143_AO6;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_B = CLBLM_R_X7Y143_SLICE_X8Y143_BO6;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_C = CLBLM_R_X7Y143_SLICE_X8Y143_CO6;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_D = CLBLM_R_X7Y143_SLICE_X8Y143_DO6;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_BMUX = CLBLM_R_X7Y143_SLICE_X8Y143_B5Q;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_A = CLBLM_R_X7Y143_SLICE_X9Y143_AO6;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_B = CLBLM_R_X7Y143_SLICE_X9Y143_BO6;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_C = CLBLM_R_X7Y143_SLICE_X9Y143_CO6;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_D = CLBLM_R_X7Y143_SLICE_X9Y143_DO6;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_A = CLBLM_R_X7Y144_SLICE_X8Y144_AO6;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_B = CLBLM_R_X7Y144_SLICE_X8Y144_BO6;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_C = CLBLM_R_X7Y144_SLICE_X8Y144_CO6;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_D = CLBLM_R_X7Y144_SLICE_X8Y144_DO6;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_A = CLBLM_R_X7Y144_SLICE_X9Y144_AO6;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_B = CLBLM_R_X7Y144_SLICE_X9Y144_BO6;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_C = CLBLM_R_X7Y144_SLICE_X9Y144_CO6;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_D = CLBLM_R_X7Y144_SLICE_X9Y144_DO6;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_AMUX = CLBLM_R_X7Y144_SLICE_X9Y144_A5Q;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_DMUX = CLBLM_R_X7Y144_SLICE_X9Y144_DO5;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_A = CLBLM_R_X7Y145_SLICE_X8Y145_AO6;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_B = CLBLM_R_X7Y145_SLICE_X8Y145_BO6;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_C = CLBLM_R_X7Y145_SLICE_X8Y145_CO6;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_D = CLBLM_R_X7Y145_SLICE_X8Y145_DO6;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_CMUX = CLBLM_R_X7Y145_SLICE_X8Y145_C5Q;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_DMUX = CLBLM_R_X7Y145_SLICE_X8Y145_DO6;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_A = CLBLM_R_X7Y145_SLICE_X9Y145_AO6;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_B = CLBLM_R_X7Y145_SLICE_X9Y145_BO6;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_C = CLBLM_R_X7Y145_SLICE_X9Y145_CO6;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_D = CLBLM_R_X7Y145_SLICE_X9Y145_DO6;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_CMUX = CLBLM_R_X7Y145_SLICE_X9Y145_C5Q;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_A = CLBLM_R_X7Y146_SLICE_X8Y146_AO6;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_B = CLBLM_R_X7Y146_SLICE_X8Y146_BO6;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_C = CLBLM_R_X7Y146_SLICE_X8Y146_CO6;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_D = CLBLM_R_X7Y146_SLICE_X8Y146_DO6;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_BMUX = CLBLM_R_X7Y146_SLICE_X8Y146_BO5;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_CMUX = CLBLM_R_X7Y146_SLICE_X8Y146_C5Q;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_A = CLBLM_R_X7Y146_SLICE_X9Y146_AO6;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_B = CLBLM_R_X7Y146_SLICE_X9Y146_BO6;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_C = CLBLM_R_X7Y146_SLICE_X9Y146_CO6;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_D = CLBLM_R_X7Y146_SLICE_X9Y146_DO6;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_A = CLBLM_R_X7Y147_SLICE_X8Y147_AO6;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_B = CLBLM_R_X7Y147_SLICE_X8Y147_BO6;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_C = CLBLM_R_X7Y147_SLICE_X8Y147_CO6;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_D = CLBLM_R_X7Y147_SLICE_X8Y147_DO6;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_BMUX = CLBLM_R_X7Y147_SLICE_X8Y147_B5Q;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_CMUX = CLBLM_R_X7Y147_SLICE_X8Y147_C5Q;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_A = CLBLM_R_X7Y147_SLICE_X9Y147_AO6;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_B = CLBLM_R_X7Y147_SLICE_X9Y147_BO6;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_C = CLBLM_R_X7Y147_SLICE_X9Y147_CO6;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_D = CLBLM_R_X7Y147_SLICE_X9Y147_DO6;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_CMUX = CLBLM_R_X7Y147_SLICE_X9Y147_CO5;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_A = CLBLM_R_X7Y148_SLICE_X8Y148_AO6;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_B = CLBLM_R_X7Y148_SLICE_X8Y148_BO6;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_C = CLBLM_R_X7Y148_SLICE_X8Y148_CO6;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_D = CLBLM_R_X7Y148_SLICE_X8Y148_DO6;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_BMUX = CLBLM_R_X7Y148_SLICE_X8Y148_BO5;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_DMUX = CLBLM_R_X7Y148_SLICE_X8Y148_D5Q;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_A = CLBLM_R_X7Y148_SLICE_X9Y148_AO6;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_B = CLBLM_R_X7Y148_SLICE_X9Y148_BO6;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_C = CLBLM_R_X7Y148_SLICE_X9Y148_CO6;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_D = CLBLM_R_X7Y148_SLICE_X9Y148_DO6;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_A = CLBLM_R_X7Y149_SLICE_X8Y149_AO6;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_B = CLBLM_R_X7Y149_SLICE_X8Y149_BO6;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_C = CLBLM_R_X7Y149_SLICE_X8Y149_CO6;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_D = CLBLM_R_X7Y149_SLICE_X8Y149_DO6;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_A = CLBLM_R_X7Y149_SLICE_X9Y149_AO6;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_B = CLBLM_R_X7Y149_SLICE_X9Y149_BO6;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_C = CLBLM_R_X7Y149_SLICE_X9Y149_CO6;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_D = CLBLM_R_X7Y149_SLICE_X9Y149_DO6;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_A = CLBLM_R_X7Y150_SLICE_X8Y150_AO6;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_B = CLBLM_R_X7Y150_SLICE_X8Y150_BO6;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_C = CLBLM_R_X7Y150_SLICE_X8Y150_CO6;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_D = CLBLM_R_X7Y150_SLICE_X8Y150_DO6;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_A = CLBLM_R_X7Y150_SLICE_X9Y150_AO6;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_B = CLBLM_R_X7Y150_SLICE_X9Y150_BO6;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_C = CLBLM_R_X7Y150_SLICE_X9Y150_CO6;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_D = CLBLM_R_X7Y150_SLICE_X9Y150_DO6;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_AMUX = CLBLM_R_X7Y150_SLICE_X9Y150_A5Q;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_BMUX = CLBLM_R_X7Y150_SLICE_X9Y150_BO5;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_CMUX = CLBLM_R_X7Y150_SLICE_X9Y150_CO5;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_A = CLBLM_R_X7Y151_SLICE_X8Y151_AO6;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_B = CLBLM_R_X7Y151_SLICE_X8Y151_BO6;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_C = CLBLM_R_X7Y151_SLICE_X8Y151_CO6;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_D = CLBLM_R_X7Y151_SLICE_X8Y151_DO6;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_AMUX = CLBLM_R_X7Y151_SLICE_X8Y151_A5Q;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_CMUX = CLBLM_R_X7Y151_SLICE_X8Y151_CO5;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_DMUX = CLBLM_R_X7Y151_SLICE_X8Y151_DO5;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_A = CLBLM_R_X7Y151_SLICE_X9Y151_AO6;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_B = CLBLM_R_X7Y151_SLICE_X9Y151_BO6;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_C = CLBLM_R_X7Y151_SLICE_X9Y151_CO6;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_D = CLBLM_R_X7Y151_SLICE_X9Y151_DO6;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_DMUX = CLBLM_R_X7Y151_SLICE_X9Y151_DO5;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_A = CLBLM_R_X7Y152_SLICE_X8Y152_AO6;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_B = CLBLM_R_X7Y152_SLICE_X8Y152_BO6;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_C = CLBLM_R_X7Y152_SLICE_X8Y152_CO6;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_D = CLBLM_R_X7Y152_SLICE_X8Y152_DO6;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_A = CLBLM_R_X7Y152_SLICE_X9Y152_AO6;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_B = CLBLM_R_X7Y152_SLICE_X9Y152_BO6;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_C = CLBLM_R_X7Y152_SLICE_X9Y152_CO6;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_D = CLBLM_R_X7Y152_SLICE_X9Y152_DO6;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_A = CLBLM_R_X7Y153_SLICE_X8Y153_AO6;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_B = CLBLM_R_X7Y153_SLICE_X8Y153_BO6;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_C = CLBLM_R_X7Y153_SLICE_X8Y153_CO6;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_D = CLBLM_R_X7Y153_SLICE_X8Y153_DO6;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_A = CLBLM_R_X7Y153_SLICE_X9Y153_AO6;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_B = CLBLM_R_X7Y153_SLICE_X9Y153_BO6;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_C = CLBLM_R_X7Y153_SLICE_X9Y153_CO6;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_D = CLBLM_R_X7Y153_SLICE_X9Y153_DO6;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_AMUX = CLBLM_R_X7Y153_SLICE_X9Y153_A5Q;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_CMUX = CLBLM_R_X7Y153_SLICE_X9Y153_CO5;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_A = CLBLM_R_X7Y154_SLICE_X8Y154_AO6;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_B = CLBLM_R_X7Y154_SLICE_X8Y154_BO6;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_C = CLBLM_R_X7Y154_SLICE_X8Y154_CO6;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_D = CLBLM_R_X7Y154_SLICE_X8Y154_DO6;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_A = CLBLM_R_X7Y154_SLICE_X9Y154_AO6;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_B = CLBLM_R_X7Y154_SLICE_X9Y154_BO6;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_C = CLBLM_R_X7Y154_SLICE_X9Y154_CO6;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_D = CLBLM_R_X7Y154_SLICE_X9Y154_DO6;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_A = CLBLM_R_X7Y155_SLICE_X8Y155_AO6;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_B = CLBLM_R_X7Y155_SLICE_X8Y155_BO6;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_C = CLBLM_R_X7Y155_SLICE_X8Y155_CO6;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_D = CLBLM_R_X7Y155_SLICE_X8Y155_DO6;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_AMUX = CLBLM_R_X7Y155_SLICE_X8Y155_A5Q;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_BMUX = CLBLM_R_X7Y155_SLICE_X8Y155_BO5;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_CMUX = CLBLM_R_X7Y155_SLICE_X8Y155_CO6;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_A = CLBLM_R_X7Y155_SLICE_X9Y155_AO6;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_B = CLBLM_R_X7Y155_SLICE_X9Y155_BO6;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_C = CLBLM_R_X7Y155_SLICE_X9Y155_CO6;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_D = CLBLM_R_X7Y155_SLICE_X9Y155_DO6;
  assign CLBLM_R_X7Y157_SLICE_X8Y157_A = CLBLM_R_X7Y157_SLICE_X8Y157_AO6;
  assign CLBLM_R_X7Y157_SLICE_X8Y157_B = CLBLM_R_X7Y157_SLICE_X8Y157_BO6;
  assign CLBLM_R_X7Y157_SLICE_X8Y157_C = CLBLM_R_X7Y157_SLICE_X8Y157_CO6;
  assign CLBLM_R_X7Y157_SLICE_X8Y157_D = CLBLM_R_X7Y157_SLICE_X8Y157_DO6;
  assign CLBLM_R_X7Y157_SLICE_X9Y157_A = CLBLM_R_X7Y157_SLICE_X9Y157_AO6;
  assign CLBLM_R_X7Y157_SLICE_X9Y157_B = CLBLM_R_X7Y157_SLICE_X9Y157_BO6;
  assign CLBLM_R_X7Y157_SLICE_X9Y157_C = CLBLM_R_X7Y157_SLICE_X9Y157_CO6;
  assign CLBLM_R_X7Y157_SLICE_X9Y157_D = CLBLM_R_X7Y157_SLICE_X9Y157_DO6;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_A = CLBLM_R_X11Y143_SLICE_X14Y143_AO6;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_B = CLBLM_R_X11Y143_SLICE_X14Y143_BO6;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_C = CLBLM_R_X11Y143_SLICE_X14Y143_CO6;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_D = CLBLM_R_X11Y143_SLICE_X14Y143_DO6;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_CMUX = CLBLM_R_X11Y143_SLICE_X14Y143_CO5;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_A = CLBLM_R_X11Y143_SLICE_X15Y143_AO6;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_B = CLBLM_R_X11Y143_SLICE_X15Y143_BO6;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_C = CLBLM_R_X11Y143_SLICE_X15Y143_CO6;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_D = CLBLM_R_X11Y143_SLICE_X15Y143_DO6;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_A = CLBLM_R_X11Y144_SLICE_X14Y144_AO6;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_B = CLBLM_R_X11Y144_SLICE_X14Y144_BO6;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_C = CLBLM_R_X11Y144_SLICE_X14Y144_CO6;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_D = CLBLM_R_X11Y144_SLICE_X14Y144_DO6;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_A = CLBLM_R_X11Y144_SLICE_X15Y144_AO6;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_B = CLBLM_R_X11Y144_SLICE_X15Y144_BO6;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_C = CLBLM_R_X11Y144_SLICE_X15Y144_CO6;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_D = CLBLM_R_X11Y144_SLICE_X15Y144_DO6;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_AMUX = CLBLM_R_X11Y144_SLICE_X15Y144_AO5;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_A = CLBLM_R_X11Y145_SLICE_X14Y145_AO6;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_B = CLBLM_R_X11Y145_SLICE_X14Y145_BO6;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_C = CLBLM_R_X11Y145_SLICE_X14Y145_CO6;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_D = CLBLM_R_X11Y145_SLICE_X14Y145_DO6;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_A = CLBLM_R_X11Y145_SLICE_X15Y145_AO6;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_B = CLBLM_R_X11Y145_SLICE_X15Y145_BO6;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_C = CLBLM_R_X11Y145_SLICE_X15Y145_CO6;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_D = CLBLM_R_X11Y145_SLICE_X15Y145_DO6;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_A = CLBLM_R_X11Y146_SLICE_X14Y146_AO6;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_B = CLBLM_R_X11Y146_SLICE_X14Y146_BO6;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_C = CLBLM_R_X11Y146_SLICE_X14Y146_CO6;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_D = CLBLM_R_X11Y146_SLICE_X14Y146_DO6;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_A = CLBLM_R_X11Y146_SLICE_X15Y146_AO6;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_B = CLBLM_R_X11Y146_SLICE_X15Y146_BO6;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_C = CLBLM_R_X11Y146_SLICE_X15Y146_CO6;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_D = CLBLM_R_X11Y146_SLICE_X15Y146_DO6;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_A = CLBLM_R_X11Y147_SLICE_X14Y147_AO6;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_B = CLBLM_R_X11Y147_SLICE_X14Y147_BO6;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_C = CLBLM_R_X11Y147_SLICE_X14Y147_CO6;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_D = CLBLM_R_X11Y147_SLICE_X14Y147_DO6;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_A = CLBLM_R_X11Y147_SLICE_X15Y147_AO6;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_B = CLBLM_R_X11Y147_SLICE_X15Y147_BO6;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_C = CLBLM_R_X11Y147_SLICE_X15Y147_CO6;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_D = CLBLM_R_X11Y147_SLICE_X15Y147_DO6;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_A = CLBLM_R_X11Y148_SLICE_X14Y148_AO6;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_B = CLBLM_R_X11Y148_SLICE_X14Y148_BO6;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_C = CLBLM_R_X11Y148_SLICE_X14Y148_CO6;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_D = CLBLM_R_X11Y148_SLICE_X14Y148_DO6;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_A = CLBLM_R_X11Y148_SLICE_X15Y148_AO6;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_B = CLBLM_R_X11Y148_SLICE_X15Y148_BO6;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_C = CLBLM_R_X11Y148_SLICE_X15Y148_CO6;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_D = CLBLM_R_X11Y148_SLICE_X15Y148_DO6;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_AMUX = CLBLM_R_X11Y148_SLICE_X15Y148_A5Q;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_BMUX = CLBLM_R_X11Y148_SLICE_X15Y148_B5Q;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_A = CLBLM_R_X11Y149_SLICE_X14Y149_AO6;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_B = CLBLM_R_X11Y149_SLICE_X14Y149_BO6;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_C = CLBLM_R_X11Y149_SLICE_X14Y149_CO6;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_D = CLBLM_R_X11Y149_SLICE_X14Y149_DO6;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_DMUX = CLBLM_R_X11Y149_SLICE_X14Y149_DO5;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_A = CLBLM_R_X11Y149_SLICE_X15Y149_AO6;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_B = CLBLM_R_X11Y149_SLICE_X15Y149_BO6;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_C = CLBLM_R_X11Y149_SLICE_X15Y149_CO6;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_D = CLBLM_R_X11Y149_SLICE_X15Y149_DO6;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_A = CLBLM_R_X11Y150_SLICE_X14Y150_AO6;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_B = CLBLM_R_X11Y150_SLICE_X14Y150_BO6;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_C = CLBLM_R_X11Y150_SLICE_X14Y150_CO6;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_D = CLBLM_R_X11Y150_SLICE_X14Y150_DO6;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_A = CLBLM_R_X11Y150_SLICE_X15Y150_AO6;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_B = CLBLM_R_X11Y150_SLICE_X15Y150_BO6;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_C = CLBLM_R_X11Y150_SLICE_X15Y150_CO6;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_D = CLBLM_R_X11Y150_SLICE_X15Y150_DO6;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_DMUX = CLBLM_R_X11Y150_SLICE_X15Y150_DO6;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_A = CLBLM_R_X11Y151_SLICE_X14Y151_AO6;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_B = CLBLM_R_X11Y151_SLICE_X14Y151_BO6;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_C = CLBLM_R_X11Y151_SLICE_X14Y151_CO6;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_D = CLBLM_R_X11Y151_SLICE_X14Y151_DO6;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_AMUX = CLBLM_R_X11Y151_SLICE_X14Y151_AO5;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_BMUX = CLBLM_R_X11Y151_SLICE_X14Y151_BO5;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_CMUX = CLBLM_R_X11Y151_SLICE_X14Y151_CO5;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_DMUX = CLBLM_R_X11Y151_SLICE_X14Y151_DO5;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_A = CLBLM_R_X11Y151_SLICE_X15Y151_AO6;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_B = CLBLM_R_X11Y151_SLICE_X15Y151_BO6;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_C = CLBLM_R_X11Y151_SLICE_X15Y151_CO6;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_D = CLBLM_R_X11Y151_SLICE_X15Y151_DO6;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_AMUX = CLBLM_R_X11Y151_SLICE_X15Y151_A5Q;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_CMUX = CLBLM_R_X11Y151_SLICE_X15Y151_CO6;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_A = CLBLM_R_X11Y152_SLICE_X14Y152_AO6;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_B = CLBLM_R_X11Y152_SLICE_X14Y152_BO6;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_C = CLBLM_R_X11Y152_SLICE_X14Y152_CO6;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_D = CLBLM_R_X11Y152_SLICE_X14Y152_DO6;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_A = CLBLM_R_X11Y152_SLICE_X15Y152_AO6;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_B = CLBLM_R_X11Y152_SLICE_X15Y152_BO6;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_C = CLBLM_R_X11Y152_SLICE_X15Y152_CO6;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_D = CLBLM_R_X11Y152_SLICE_X15Y152_DO6;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_A = CLBLM_R_X11Y153_SLICE_X14Y153_AO6;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_B = CLBLM_R_X11Y153_SLICE_X14Y153_BO6;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_C = CLBLM_R_X11Y153_SLICE_X14Y153_CO6;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_D = CLBLM_R_X11Y153_SLICE_X14Y153_DO6;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_AMUX = CLBLM_R_X11Y153_SLICE_X14Y153_AO5;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_BMUX = CLBLM_R_X11Y153_SLICE_X14Y153_BO5;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_CMUX = CLBLM_R_X11Y153_SLICE_X14Y153_CO5;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_DMUX = CLBLM_R_X11Y153_SLICE_X14Y153_DO6;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_A = CLBLM_R_X11Y153_SLICE_X15Y153_AO6;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_B = CLBLM_R_X11Y153_SLICE_X15Y153_BO6;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_C = CLBLM_R_X11Y153_SLICE_X15Y153_CO6;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_D = CLBLM_R_X11Y153_SLICE_X15Y153_DO6;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_CMUX = CLBLM_R_X11Y153_SLICE_X15Y153_CO5;
  assign CLBLM_R_X11Y154_SLICE_X14Y154_A = CLBLM_R_X11Y154_SLICE_X14Y154_AO6;
  assign CLBLM_R_X11Y154_SLICE_X14Y154_B = CLBLM_R_X11Y154_SLICE_X14Y154_BO6;
  assign CLBLM_R_X11Y154_SLICE_X14Y154_C = CLBLM_R_X11Y154_SLICE_X14Y154_CO6;
  assign CLBLM_R_X11Y154_SLICE_X14Y154_D = CLBLM_R_X11Y154_SLICE_X14Y154_DO6;
  assign CLBLM_R_X11Y154_SLICE_X14Y154_BMUX = CLBLM_R_X11Y154_SLICE_X14Y154_BO5;
  assign CLBLM_R_X11Y154_SLICE_X14Y154_CMUX = CLBLM_R_X11Y154_SLICE_X14Y154_CO5;
  assign CLBLM_R_X11Y154_SLICE_X15Y154_A = CLBLM_R_X11Y154_SLICE_X15Y154_AO6;
  assign CLBLM_R_X11Y154_SLICE_X15Y154_B = CLBLM_R_X11Y154_SLICE_X15Y154_BO6;
  assign CLBLM_R_X11Y154_SLICE_X15Y154_C = CLBLM_R_X11Y154_SLICE_X15Y154_CO6;
  assign CLBLM_R_X11Y154_SLICE_X15Y154_D = CLBLM_R_X11Y154_SLICE_X15Y154_DO6;
  assign CLBLM_R_X11Y154_SLICE_X15Y154_CMUX = CLBLM_R_X11Y154_SLICE_X15Y154_CO5;
  assign CLBLM_R_X11Y157_SLICE_X14Y157_A = CLBLM_R_X11Y157_SLICE_X14Y157_AO6;
  assign CLBLM_R_X11Y157_SLICE_X14Y157_B = CLBLM_R_X11Y157_SLICE_X14Y157_BO6;
  assign CLBLM_R_X11Y157_SLICE_X14Y157_C = CLBLM_R_X11Y157_SLICE_X14Y157_CO6;
  assign CLBLM_R_X11Y157_SLICE_X14Y157_D = CLBLM_R_X11Y157_SLICE_X14Y157_DO6;
  assign CLBLM_R_X11Y157_SLICE_X14Y157_AMUX = CLBLM_R_X11Y157_SLICE_X14Y157_AO5;
  assign CLBLM_R_X11Y157_SLICE_X15Y157_A = CLBLM_R_X11Y157_SLICE_X15Y157_AO6;
  assign CLBLM_R_X11Y157_SLICE_X15Y157_B = CLBLM_R_X11Y157_SLICE_X15Y157_BO6;
  assign CLBLM_R_X11Y157_SLICE_X15Y157_C = CLBLM_R_X11Y157_SLICE_X15Y157_CO6;
  assign CLBLM_R_X11Y157_SLICE_X15Y157_D = CLBLM_R_X11Y157_SLICE_X15Y157_DO6;
  assign CLBLM_R_X13Y151_SLICE_X18Y151_A = CLBLM_R_X13Y151_SLICE_X18Y151_AO6;
  assign CLBLM_R_X13Y151_SLICE_X18Y151_B = CLBLM_R_X13Y151_SLICE_X18Y151_BO6;
  assign CLBLM_R_X13Y151_SLICE_X18Y151_C = CLBLM_R_X13Y151_SLICE_X18Y151_CO6;
  assign CLBLM_R_X13Y151_SLICE_X18Y151_D = CLBLM_R_X13Y151_SLICE_X18Y151_DO6;
  assign CLBLM_R_X13Y151_SLICE_X19Y151_A = CLBLM_R_X13Y151_SLICE_X19Y151_AO6;
  assign CLBLM_R_X13Y151_SLICE_X19Y151_B = CLBLM_R_X13Y151_SLICE_X19Y151_BO6;
  assign CLBLM_R_X13Y151_SLICE_X19Y151_C = CLBLM_R_X13Y151_SLICE_X19Y151_CO6;
  assign CLBLM_R_X13Y151_SLICE_X19Y151_D = CLBLM_R_X13Y151_SLICE_X19Y151_DO6;
  assign CLBLM_R_X13Y152_SLICE_X18Y152_A = CLBLM_R_X13Y152_SLICE_X18Y152_AO6;
  assign CLBLM_R_X13Y152_SLICE_X18Y152_B = CLBLM_R_X13Y152_SLICE_X18Y152_BO6;
  assign CLBLM_R_X13Y152_SLICE_X18Y152_C = CLBLM_R_X13Y152_SLICE_X18Y152_CO6;
  assign CLBLM_R_X13Y152_SLICE_X18Y152_D = CLBLM_R_X13Y152_SLICE_X18Y152_DO6;
  assign CLBLM_R_X13Y152_SLICE_X19Y152_A = CLBLM_R_X13Y152_SLICE_X19Y152_AO6;
  assign CLBLM_R_X13Y152_SLICE_X19Y152_B = CLBLM_R_X13Y152_SLICE_X19Y152_BO6;
  assign CLBLM_R_X13Y152_SLICE_X19Y152_C = CLBLM_R_X13Y152_SLICE_X19Y152_CO6;
  assign CLBLM_R_X13Y152_SLICE_X19Y152_D = CLBLM_R_X13Y152_SLICE_X19Y152_DO6;
  assign CLBLM_R_X15Y151_SLICE_X20Y151_A = CLBLM_R_X15Y151_SLICE_X20Y151_AO6;
  assign CLBLM_R_X15Y151_SLICE_X20Y151_B = CLBLM_R_X15Y151_SLICE_X20Y151_BO6;
  assign CLBLM_R_X15Y151_SLICE_X20Y151_C = CLBLM_R_X15Y151_SLICE_X20Y151_CO6;
  assign CLBLM_R_X15Y151_SLICE_X20Y151_D = CLBLM_R_X15Y151_SLICE_X20Y151_DO6;
  assign CLBLM_R_X15Y151_SLICE_X21Y151_A = CLBLM_R_X15Y151_SLICE_X21Y151_AO6;
  assign CLBLM_R_X15Y151_SLICE_X21Y151_B = CLBLM_R_X15Y151_SLICE_X21Y151_BO6;
  assign CLBLM_R_X15Y151_SLICE_X21Y151_C = CLBLM_R_X15Y151_SLICE_X21Y151_CO6;
  assign CLBLM_R_X15Y151_SLICE_X21Y151_D = CLBLM_R_X15Y151_SLICE_X21Y151_DO6;
  assign CLBLM_R_X15Y153_SLICE_X20Y153_A = CLBLM_R_X15Y153_SLICE_X20Y153_AO6;
  assign CLBLM_R_X15Y153_SLICE_X20Y153_B = CLBLM_R_X15Y153_SLICE_X20Y153_BO6;
  assign CLBLM_R_X15Y153_SLICE_X20Y153_C = CLBLM_R_X15Y153_SLICE_X20Y153_CO6;
  assign CLBLM_R_X15Y153_SLICE_X20Y153_D = CLBLM_R_X15Y153_SLICE_X20Y153_DO6;
  assign CLBLM_R_X15Y153_SLICE_X20Y153_AMUX = CLBLM_R_X15Y153_SLICE_X20Y153_AO5;
  assign CLBLM_R_X15Y153_SLICE_X21Y153_A = CLBLM_R_X15Y153_SLICE_X21Y153_AO6;
  assign CLBLM_R_X15Y153_SLICE_X21Y153_B = CLBLM_R_X15Y153_SLICE_X21Y153_BO6;
  assign CLBLM_R_X15Y153_SLICE_X21Y153_C = CLBLM_R_X15Y153_SLICE_X21Y153_CO6;
  assign CLBLM_R_X15Y153_SLICE_X21Y153_D = CLBLM_R_X15Y153_SLICE_X21Y153_DO6;
  assign CLBLM_R_X103Y141_SLICE_X162Y141_A = CLBLM_R_X103Y141_SLICE_X162Y141_AO6;
  assign CLBLM_R_X103Y141_SLICE_X162Y141_B = CLBLM_R_X103Y141_SLICE_X162Y141_BO6;
  assign CLBLM_R_X103Y141_SLICE_X162Y141_C = CLBLM_R_X103Y141_SLICE_X162Y141_CO6;
  assign CLBLM_R_X103Y141_SLICE_X162Y141_D = CLBLM_R_X103Y141_SLICE_X162Y141_DO6;
  assign CLBLM_R_X103Y141_SLICE_X163Y141_A = CLBLM_R_X103Y141_SLICE_X163Y141_AO6;
  assign CLBLM_R_X103Y141_SLICE_X163Y141_B = CLBLM_R_X103Y141_SLICE_X163Y141_BO6;
  assign CLBLM_R_X103Y141_SLICE_X163Y141_C = CLBLM_R_X103Y141_SLICE_X163Y141_CO6;
  assign CLBLM_R_X103Y141_SLICE_X163Y141_D = CLBLM_R_X103Y141_SLICE_X163Y141_DO6;
  assign CLBLM_R_X103Y141_SLICE_X163Y141_AMUX = CLBLM_R_X103Y141_SLICE_X163Y141_AO5;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_A = CLBLM_R_X103Y169_SLICE_X162Y169_AO6;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_B = CLBLM_R_X103Y169_SLICE_X162Y169_BO6;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_C = CLBLM_R_X103Y169_SLICE_X162Y169_CO6;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_D = CLBLM_R_X103Y169_SLICE_X162Y169_DO6;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_A = CLBLM_R_X103Y169_SLICE_X163Y169_AO6;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_B = CLBLM_R_X103Y169_SLICE_X163Y169_BO6;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_C = CLBLM_R_X103Y169_SLICE_X163Y169_CO6;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_D = CLBLM_R_X103Y169_SLICE_X163Y169_DO6;
  assign CLBLM_R_X103Y170_SLICE_X162Y170_A = CLBLM_R_X103Y170_SLICE_X162Y170_AO6;
  assign CLBLM_R_X103Y170_SLICE_X162Y170_B = CLBLM_R_X103Y170_SLICE_X162Y170_BO6;
  assign CLBLM_R_X103Y170_SLICE_X162Y170_C = CLBLM_R_X103Y170_SLICE_X162Y170_CO6;
  assign CLBLM_R_X103Y170_SLICE_X162Y170_D = CLBLM_R_X103Y170_SLICE_X162Y170_DO6;
  assign CLBLM_R_X103Y170_SLICE_X163Y170_A = CLBLM_R_X103Y170_SLICE_X163Y170_AO6;
  assign CLBLM_R_X103Y170_SLICE_X163Y170_B = CLBLM_R_X103Y170_SLICE_X163Y170_BO6;
  assign CLBLM_R_X103Y170_SLICE_X163Y170_C = CLBLM_R_X103Y170_SLICE_X163Y170_CO6;
  assign CLBLM_R_X103Y170_SLICE_X163Y170_D = CLBLM_R_X103Y170_SLICE_X163Y170_DO6;
  assign CLBLM_R_X103Y170_SLICE_X163Y170_AMUX = CLBLM_R_X103Y170_SLICE_X163Y170_AO5;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_A = CLBLM_R_X103Y173_SLICE_X162Y173_AO6;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_B = CLBLM_R_X103Y173_SLICE_X162Y173_BO6;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_C = CLBLM_R_X103Y173_SLICE_X162Y173_CO6;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_D = CLBLM_R_X103Y173_SLICE_X162Y173_DO6;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_A = CLBLM_R_X103Y173_SLICE_X163Y173_AO6;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_B = CLBLM_R_X103Y173_SLICE_X163Y173_BO6;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_C = CLBLM_R_X103Y173_SLICE_X163Y173_CO6;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_D = CLBLM_R_X103Y173_SLICE_X163Y173_DO6;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_AMUX = CLBLM_R_X103Y173_SLICE_X163Y173_AO5;
  assign CLBLM_R_X103Y176_SLICE_X162Y176_A = CLBLM_R_X103Y176_SLICE_X162Y176_AO6;
  assign CLBLM_R_X103Y176_SLICE_X162Y176_B = CLBLM_R_X103Y176_SLICE_X162Y176_BO6;
  assign CLBLM_R_X103Y176_SLICE_X162Y176_C = CLBLM_R_X103Y176_SLICE_X162Y176_CO6;
  assign CLBLM_R_X103Y176_SLICE_X162Y176_D = CLBLM_R_X103Y176_SLICE_X162Y176_DO6;
  assign CLBLM_R_X103Y176_SLICE_X163Y176_A = CLBLM_R_X103Y176_SLICE_X163Y176_AO6;
  assign CLBLM_R_X103Y176_SLICE_X163Y176_B = CLBLM_R_X103Y176_SLICE_X163Y176_BO6;
  assign CLBLM_R_X103Y176_SLICE_X163Y176_C = CLBLM_R_X103Y176_SLICE_X163Y176_CO6;
  assign CLBLM_R_X103Y176_SLICE_X163Y176_D = CLBLM_R_X103Y176_SLICE_X163Y176_DO6;
  assign CLBLM_R_X103Y176_SLICE_X163Y176_AMUX = CLBLM_R_X103Y176_SLICE_X163Y176_AO5;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_A = CLBLM_R_X103Y178_SLICE_X162Y178_AO6;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_B = CLBLM_R_X103Y178_SLICE_X162Y178_BO6;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_C = CLBLM_R_X103Y178_SLICE_X162Y178_CO6;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_D = CLBLM_R_X103Y178_SLICE_X162Y178_DO6;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_A = CLBLM_R_X103Y178_SLICE_X163Y178_AO6;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_B = CLBLM_R_X103Y178_SLICE_X163Y178_BO6;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_C = CLBLM_R_X103Y178_SLICE_X163Y178_CO6;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_D = CLBLM_R_X103Y178_SLICE_X163Y178_DO6;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_AMUX = CLBLM_R_X103Y178_SLICE_X163Y178_AO5;
  assign LIOI3_X0Y51_ILOGIC_X0Y52_O = LIOB33_X0Y51_IOB_X0Y52_I;
  assign LIOI3_X0Y51_ILOGIC_X0Y51_O = LIOB33_X0Y51_IOB_X0Y51_I;
  assign LIOI3_X0Y53_ILOGIC_X0Y54_O = LIOB33_X0Y53_IOB_X0Y54_I;
  assign LIOI3_X0Y53_ILOGIC_X0Y53_O = LIOB33_X0Y53_IOB_X0Y53_I;
  assign LIOI3_X0Y55_ILOGIC_X0Y56_O = LIOB33_X0Y55_IOB_X0Y56_I;
  assign LIOI3_X0Y55_ILOGIC_X0Y55_O = LIOB33_X0Y55_IOB_X0Y55_I;
  assign LIOI3_X0Y59_ILOGIC_X0Y60_O = LIOB33_X0Y59_IOB_X0Y60_I;
  assign LIOI3_X0Y59_ILOGIC_X0Y59_O = LIOB33_X0Y59_IOB_X0Y59_I;
  assign LIOI3_X0Y61_ILOGIC_X0Y62_O = LIOB33_X0Y61_IOB_X0Y62_I;
  assign LIOI3_X0Y61_ILOGIC_X0Y61_O = LIOB33_X0Y61_IOB_X0Y61_I;
  assign LIOI3_X0Y65_ILOGIC_X0Y66_O = LIOB33_X0Y65_IOB_X0Y66_I;
  assign LIOI3_X0Y65_ILOGIC_X0Y65_O = LIOB33_X0Y65_IOB_X0Y65_I;
  assign LIOI3_X0Y67_ILOGIC_X0Y68_O = LIOB33_X0Y67_IOB_X0Y68_I;
  assign LIOI3_X0Y67_ILOGIC_X0Y67_O = LIOB33_X0Y67_IOB_X0Y67_I;
  assign LIOI3_X0Y71_ILOGIC_X0Y72_O = LIOB33_X0Y71_IOB_X0Y72_I;
  assign LIOI3_X0Y71_ILOGIC_X0Y71_O = LIOB33_X0Y71_IOB_X0Y71_I;
  assign LIOI3_X0Y73_ILOGIC_X0Y74_O = LIOB33_X0Y73_IOB_X0Y74_I;
  assign LIOI3_X0Y73_ILOGIC_X0Y73_O = LIOB33_X0Y73_IOB_X0Y73_I;
  assign LIOI3_X0Y75_ILOGIC_X0Y76_O = LIOB33_X0Y75_IOB_X0Y76_I;
  assign LIOI3_X0Y75_ILOGIC_X0Y75_O = LIOB33_X0Y75_IOB_X0Y75_I;
  assign LIOI3_X0Y77_ILOGIC_X0Y78_O = LIOB33_X0Y77_IOB_X0Y78_I;
  assign LIOI3_X0Y77_ILOGIC_X0Y77_O = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOI3_X0Y79_ILOGIC_X0Y79_O = LIOB33_X0Y79_IOB_X0Y79_I;
  assign LIOI3_X0Y79_OLOGIC_X0Y80_OQ = CLBLL_L_X2Y138_SLICE_X0Y138_AO6;
  assign LIOI3_X0Y79_OLOGIC_X0Y80_TQ = 1'b1;
  assign LIOI3_X0Y101_OLOGIC_X0Y102_OQ = CLBLL_L_X2Y138_SLICE_X0Y138_BO5;
  assign LIOI3_X0Y101_OLOGIC_X0Y102_TQ = 1'b1;
  assign LIOI3_X0Y101_OLOGIC_X0Y101_OQ = CLBLL_L_X2Y138_SLICE_X0Y138_BO6;
  assign LIOI3_X0Y101_OLOGIC_X0Y101_TQ = 1'b1;
  assign LIOI3_X0Y103_OLOGIC_X0Y104_OQ = CLBLL_L_X2Y141_SLICE_X0Y141_AO5;
  assign LIOI3_X0Y103_OLOGIC_X0Y104_TQ = 1'b1;
  assign LIOI3_X0Y103_OLOGIC_X0Y103_OQ = CLBLL_L_X2Y141_SLICE_X0Y141_AO6;
  assign LIOI3_X0Y103_OLOGIC_X0Y103_TQ = 1'b1;
  assign LIOI3_X0Y105_OLOGIC_X0Y106_OQ = CLBLL_L_X2Y138_SLICE_X0Y138_CO5;
  assign LIOI3_X0Y105_OLOGIC_X0Y106_TQ = 1'b1;
  assign LIOI3_X0Y105_OLOGIC_X0Y105_OQ = CLBLL_L_X2Y138_SLICE_X0Y138_CO6;
  assign LIOI3_X0Y105_OLOGIC_X0Y105_TQ = 1'b1;
  assign LIOI3_X0Y109_OLOGIC_X0Y110_OQ = CLBLL_L_X2Y134_SLICE_X0Y134_AO5;
  assign LIOI3_X0Y109_OLOGIC_X0Y110_TQ = 1'b1;
  assign LIOI3_X0Y109_OLOGIC_X0Y109_OQ = CLBLL_L_X2Y134_SLICE_X0Y134_AO6;
  assign LIOI3_X0Y109_OLOGIC_X0Y109_TQ = 1'b1;
  assign LIOI3_X0Y111_OLOGIC_X0Y112_OQ = CLBLM_R_X11Y148_SLICE_X15Y148_B5Q;
  assign LIOI3_X0Y111_OLOGIC_X0Y112_TQ = 1'b1;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_OQ = 1'b0;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_TQ = 1'b1;
  assign LIOI3_X0Y115_OLOGIC_X0Y116_OQ = CLBLM_L_X8Y142_SLICE_X10Y142_AQ;
  assign LIOI3_X0Y115_OLOGIC_X0Y116_TQ = 1'b1;
  assign LIOI3_X0Y115_OLOGIC_X0Y115_OQ = CLBLM_R_X11Y148_SLICE_X15Y148_BQ;
  assign LIOI3_X0Y115_OLOGIC_X0Y115_TQ = 1'b1;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_OQ = CLBLM_R_X3Y147_SLICE_X3Y147_CQ;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_TQ = 1'b1;
  assign LIOI3_X0Y117_OLOGIC_X0Y117_OQ = CLBLM_R_X3Y144_SLICE_X2Y144_B5Q;
  assign LIOI3_X0Y117_OLOGIC_X0Y117_TQ = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_OQ = CLBLM_R_X3Y144_SLICE_X2Y144_BQ;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_TQ = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_OQ = CLBLM_L_X8Y142_SLICE_X10Y142_A5Q;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_TQ = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_OQ = CLBLM_R_X3Y147_SLICE_X3Y147_C5Q;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_TQ = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_OQ = CLBLM_R_X7Y143_SLICE_X8Y143_B5Q;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_TQ = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_OQ = CLBLM_R_X3Y143_SLICE_X2Y143_BQ;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_TQ = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_OQ = CLBLM_L_X8Y145_SLICE_X11Y145_B5Q;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_TQ = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_OQ = CLBLL_L_X2Y147_SLICE_X1Y147_AQ;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_TQ = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_OQ = CLBLL_L_X4Y147_SLICE_X5Y147_CQ;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_TQ = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_OQ = CLBLL_L_X52Y126_SLICE_X78Y126_AO6;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_TQ = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_OQ = CLBLM_R_X3Y148_SLICE_X3Y148_AQ;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_TQ = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_OQ = CLBLM_R_X3Y143_SLICE_X2Y143_CQ;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_TQ = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_OQ = CLBLM_R_X3Y143_SLICE_X3Y143_A5Q;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_TQ = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_OQ = CLBLL_L_X2Y145_SLICE_X1Y145_AQ;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_TQ = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_OQ = CLBLM_R_X3Y142_SLICE_X2Y142_BQ;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_TQ = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_OQ = CLBLM_R_X3Y142_SLICE_X2Y142_CQ;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_TQ = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_OQ = CLBLM_R_X3Y143_SLICE_X3Y143_AQ;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_TQ = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_OQ = LIOB33_X0Y53_IOB_X0Y54_I;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_TQ = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_OQ = CLBLM_R_X3Y143_SLICE_X2Y143_AQ;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_TQ = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_OQ = LIOB33_X0Y59_IOB_X0Y59_I;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_TQ = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_OQ = LIOB33_X0Y57_IOB_X0Y58_I;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_TQ = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_OQ = LIOB33_X0Y61_IOB_X0Y61_I;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_TQ = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_OQ = LIOB33_X0Y71_IOB_X0Y71_I;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_TQ = 1'b1;
  assign LIOI3_X0Y151_OLOGIC_X0Y152_OQ = LIOB33_X0Y65_IOB_X0Y66_I;
  assign LIOI3_X0Y151_OLOGIC_X0Y152_TQ = 1'b1;
  assign LIOI3_X0Y151_OLOGIC_X0Y151_OQ = LIOB33_X0Y65_IOB_X0Y65_I;
  assign LIOI3_X0Y151_OLOGIC_X0Y151_TQ = 1'b1;
  assign LIOI3_X0Y153_OLOGIC_X0Y154_OQ = LIOB33_X0Y67_IOB_X0Y68_I;
  assign LIOI3_X0Y153_OLOGIC_X0Y154_TQ = 1'b1;
  assign LIOI3_X0Y153_OLOGIC_X0Y153_OQ = LIOB33_X0Y67_IOB_X0Y67_I;
  assign LIOI3_X0Y153_OLOGIC_X0Y153_TQ = 1'b1;
  assign LIOI3_X0Y155_OLOGIC_X0Y156_OQ = RIOB33_X105Y105_IOB_X1Y106_I;
  assign LIOI3_X0Y155_OLOGIC_X0Y156_TQ = 1'b1;
  assign LIOI3_X0Y155_OLOGIC_X0Y155_OQ = LIOB33_X0Y69_IOB_X0Y70_I;
  assign LIOI3_X0Y155_OLOGIC_X0Y155_TQ = 1'b1;
  assign LIOI3_X0Y159_OLOGIC_X0Y160_OQ = RIOB33_X105Y107_IOB_X1Y107_I;
  assign LIOI3_X0Y159_OLOGIC_X0Y160_TQ = 1'b1;
  assign LIOI3_X0Y159_OLOGIC_X0Y159_OQ = RIOB33_X105Y117_IOB_X1Y117_I;
  assign LIOI3_X0Y159_OLOGIC_X0Y159_TQ = 1'b1;
  assign LIOI3_X0Y161_OLOGIC_X0Y162_OQ = RIOB33_X105Y109_IOB_X1Y109_I;
  assign LIOI3_X0Y161_OLOGIC_X0Y162_TQ = 1'b1;
  assign LIOI3_X0Y161_OLOGIC_X0Y161_OQ = RIOB33_X105Y107_IOB_X1Y108_I;
  assign LIOI3_X0Y161_OLOGIC_X0Y161_TQ = 1'b1;
  assign LIOI3_X0Y165_OLOGIC_X0Y166_OQ = RIOB33_X105Y113_IOB_X1Y113_I;
  assign LIOI3_X0Y165_OLOGIC_X0Y166_TQ = 1'b1;
  assign LIOI3_X0Y165_OLOGIC_X0Y165_OQ = RIOB33_X105Y111_IOB_X1Y112_I;
  assign LIOI3_X0Y165_OLOGIC_X0Y165_TQ = 1'b1;
  assign LIOI3_X0Y167_OLOGIC_X0Y168_OQ = RIOB33_X105Y123_IOB_X1Y123_I;
  assign LIOI3_X0Y167_OLOGIC_X0Y168_TQ = 1'b1;
  assign LIOI3_X0Y167_OLOGIC_X0Y167_OQ = RIOB33_X105Y113_IOB_X1Y114_I;
  assign LIOI3_X0Y167_OLOGIC_X0Y167_TQ = 1'b1;
  assign LIOI3_X0Y171_OLOGIC_X0Y172_OQ = CLBLM_R_X103Y141_SLICE_X163Y141_AO6;
  assign LIOI3_X0Y171_OLOGIC_X0Y172_TQ = 1'b1;
  assign LIOI3_X0Y171_OLOGIC_X0Y171_OQ = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign LIOI3_X0Y171_OLOGIC_X0Y171_TQ = 1'b1;
  assign LIOI3_X0Y173_OLOGIC_X0Y174_OQ = CLBLM_L_X8Y159_SLICE_X10Y159_AO6;
  assign LIOI3_X0Y173_OLOGIC_X0Y174_TQ = 1'b1;
  assign LIOI3_X0Y173_OLOGIC_X0Y173_OQ = CLBLM_R_X103Y141_SLICE_X163Y141_AO5;
  assign LIOI3_X0Y173_OLOGIC_X0Y173_TQ = 1'b1;
  assign LIOI3_X0Y175_OLOGIC_X0Y176_OQ = RIOB33_X105Y127_IOB_X1Y128_I;
  assign LIOI3_X0Y175_OLOGIC_X0Y176_TQ = 1'b1;
  assign LIOI3_X0Y175_OLOGIC_X0Y175_OQ = RIOB33_X105Y127_IOB_X1Y127_I;
  assign LIOI3_X0Y175_OLOGIC_X0Y175_TQ = 1'b1;
  assign LIOI3_X0Y177_OLOGIC_X0Y178_OQ = RIOB33_X105Y129_IOB_X1Y130_I;
  assign LIOI3_X0Y177_OLOGIC_X0Y178_TQ = 1'b1;
  assign LIOI3_X0Y177_OLOGIC_X0Y177_OQ = RIOB33_X105Y129_IOB_X1Y129_I;
  assign LIOI3_X0Y177_OLOGIC_X0Y177_TQ = 1'b1;
  assign LIOI3_X0Y179_OLOGIC_X0Y180_OQ = RIOB33_X105Y131_IOB_X1Y132_I;
  assign LIOI3_X0Y179_OLOGIC_X0Y180_TQ = 1'b1;
  assign LIOI3_X0Y179_OLOGIC_X0Y179_OQ = RIOB33_X105Y131_IOB_X1Y131_I;
  assign LIOI3_X0Y179_OLOGIC_X0Y179_TQ = 1'b1;
  assign LIOI3_X0Y183_OLOGIC_X0Y184_OQ = RIOB33_X105Y135_IOB_X1Y136_I;
  assign LIOI3_X0Y183_OLOGIC_X0Y184_TQ = 1'b1;
  assign LIOI3_X0Y183_OLOGIC_X0Y183_OQ = RIOB33_X105Y135_IOB_X1Y135_I;
  assign LIOI3_X0Y183_OLOGIC_X0Y183_TQ = 1'b1;
  assign LIOI3_X0Y185_OLOGIC_X0Y186_OQ = RIOB33_X105Y143_IOB_X1Y143_I;
  assign LIOI3_X0Y185_OLOGIC_X0Y186_TQ = 1'b1;
  assign LIOI3_X0Y185_OLOGIC_X0Y185_OQ = RIOB33_X105Y137_IOB_X1Y137_I;
  assign LIOI3_X0Y185_OLOGIC_X0Y185_TQ = 1'b1;
  assign LIOI3_X0Y189_OLOGIC_X0Y190_OQ = RIOB33_X105Y147_IOB_X1Y147_I;
  assign LIOI3_X0Y189_OLOGIC_X0Y190_TQ = 1'b1;
  assign LIOI3_X0Y189_OLOGIC_X0Y189_OQ = RIOB33_X105Y145_IOB_X1Y146_I;
  assign LIOI3_X0Y189_OLOGIC_X0Y189_TQ = 1'b1;
  assign LIOI3_X0Y191_OLOGIC_X0Y192_OQ = LIOB33_X0Y51_IOB_X0Y52_I;
  assign LIOI3_X0Y191_OLOGIC_X0Y192_TQ = 1'b1;
  assign LIOI3_X0Y191_OLOGIC_X0Y191_OQ = RIOB33_X105Y147_IOB_X1Y148_I;
  assign LIOI3_X0Y191_OLOGIC_X0Y191_TQ = 1'b1;
  assign LIOI3_X0Y195_OLOGIC_X0Y196_OQ = LIOB33_X0Y69_IOB_X0Y69_I;
  assign LIOI3_X0Y195_OLOGIC_X0Y196_TQ = 1'b1;
  assign LIOI3_X0Y195_OLOGIC_X0Y195_OQ = LIOB33_X0Y63_IOB_X0Y64_I;
  assign LIOI3_X0Y195_OLOGIC_X0Y195_TQ = 1'b1;
  assign LIOI3_X0Y197_OLOGIC_X0Y198_OQ = LIOB33_X0Y73_IOB_X0Y73_I;
  assign LIOI3_X0Y197_OLOGIC_X0Y198_TQ = 1'b1;
  assign LIOI3_X0Y197_OLOGIC_X0Y197_OQ = LIOB33_X0Y71_IOB_X0Y72_I;
  assign LIOI3_X0Y197_OLOGIC_X0Y197_TQ = 1'b1;
  assign LIOI3_SING_X0Y50_ILOGIC_X0Y50_O = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign LIOI3_SING_X0Y100_OLOGIC_X0Y100_OQ = CLBLL_L_X2Y138_SLICE_X0Y138_AO5;
  assign LIOI3_SING_X0Y100_OLOGIC_X0Y100_TQ = 1'b1;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_OQ = LIOB33_X0Y61_IOB_X0Y62_I;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_TQ = 1'b1;
  assign LIOI3_SING_X0Y150_OLOGIC_X0Y150_OQ = LIOB33_X0Y63_IOB_X0Y63_I;
  assign LIOI3_SING_X0Y150_OLOGIC_X0Y150_TQ = 1'b1;
  assign LIOI3_SING_X0Y199_OLOGIC_X0Y199_OQ = LIOB33_X0Y73_IOB_X0Y74_I;
  assign LIOI3_SING_X0Y199_OLOGIC_X0Y199_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y58_O = LIOB33_X0Y57_IOB_X0Y58_I;
  assign LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y57_O = LIOB33_X0Y57_IOB_X0Y57_I;
  assign LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y70_O = LIOB33_X0Y69_IOB_X0Y70_I;
  assign LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y69_O = LIOB33_X0Y69_IOB_X0Y69_I;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_OQ = CLBLM_R_X3Y152_SLICE_X2Y152_BO6;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_OQ = CLBLL_L_X2Y120_SLICE_X0Y120_AO6;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_OQ = CLBLM_L_X10Y145_SLICE_X13Y145_AQ;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_OQ = CLBLM_L_X10Y146_SLICE_X13Y146_BQ;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_OQ = CLBLM_R_X5Y142_SLICE_X7Y142_AQ;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_OQ = CLBLM_R_X7Y142_SLICE_X8Y142_AO5;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_OQ = LIOB33_X0Y57_IOB_X0Y57_I;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_OQ = LIOB33_X0Y55_IOB_X0Y55_I;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_OQ = RIOB33_X105Y115_IOB_X1Y116_I;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_OQ = RIOB33_X105Y115_IOB_X1Y115_I;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_OQ = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_OQ = RIOB33_X105Y121_IOB_X1Y122_I;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_OQ = RIOB33_X105Y133_IOB_X1Y134_I;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_OQ = RIOB33_X105Y133_IOB_X1Y133_I;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_OQ = LIOB33_X0Y59_IOB_X0Y60_I;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_OQ = LIOB33_X0Y55_IOB_X0Y56_I;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y64_O = LIOB33_X0Y63_IOB_X0Y64_I;
  assign LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y63_O = LIOB33_X0Y63_IOB_X0Y63_I;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_OQ = CLBLM_R_X7Y143_SLICE_X8Y143_BQ;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_OQ = RIOB33_X105Y121_IOB_X1Y121_I;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_OQ = CLBLM_R_X3Y143_SLICE_X3Y143_BQ;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_OQ = CLBLM_R_X3Y142_SLICE_X2Y142_AQ;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_OQ = RIOB33_X105Y111_IOB_X1Y111_I;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_OQ = RIOB33_X105Y109_IOB_X1Y110_I;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_OQ = RIOB33_X105Y145_IOB_X1Y145_I;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_OQ = RIOB33_X105Y143_IOB_X1Y144_I;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_TQ = 1'b1;
  assign RIOI3_X105Y101_ILOGIC_X1Y102_O = RIOB33_X105Y101_IOB_X1Y102_I;
  assign RIOI3_X105Y101_ILOGIC_X1Y101_O = RIOB33_X105Y101_IOB_X1Y101_I;
  assign RIOI3_X105Y103_ILOGIC_X1Y104_O = RIOB33_X105Y103_IOB_X1Y104_I;
  assign RIOI3_X105Y103_ILOGIC_X1Y103_O = RIOB33_X105Y103_IOB_X1Y103_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y106_O = RIOB33_X105Y105_IOB_X1Y106_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y105_O = RIOB33_X105Y105_IOB_X1Y105_I;
  assign RIOI3_X105Y109_ILOGIC_X1Y110_O = RIOB33_X105Y109_IOB_X1Y110_I;
  assign RIOI3_X105Y109_ILOGIC_X1Y109_O = RIOB33_X105Y109_IOB_X1Y109_I;
  assign RIOI3_X105Y111_ILOGIC_X1Y112_O = RIOB33_X105Y111_IOB_X1Y112_I;
  assign RIOI3_X105Y111_ILOGIC_X1Y111_O = RIOB33_X105Y111_IOB_X1Y111_I;
  assign RIOI3_X105Y115_ILOGIC_X1Y116_O = RIOB33_X105Y115_IOB_X1Y116_I;
  assign RIOI3_X105Y115_ILOGIC_X1Y115_O = RIOB33_X105Y115_IOB_X1Y115_I;
  assign RIOI3_X105Y117_ILOGIC_X1Y118_O = RIOB33_X105Y117_IOB_X1Y118_I;
  assign RIOI3_X105Y117_ILOGIC_X1Y117_O = RIOB33_X105Y117_IOB_X1Y117_I;
  assign RIOI3_X105Y121_ILOGIC_X1Y122_O = RIOB33_X105Y121_IOB_X1Y122_I;
  assign RIOI3_X105Y121_ILOGIC_X1Y121_O = RIOB33_X105Y121_IOB_X1Y121_I;
  assign RIOI3_X105Y123_ILOGIC_X1Y124_O = RIOB33_X105Y123_IOB_X1Y124_I;
  assign RIOI3_X105Y123_ILOGIC_X1Y123_O = RIOB33_X105Y123_IOB_X1Y123_I;
  assign RIOI3_X105Y125_ILOGIC_X1Y126_O = RIOB33_X105Y125_IOB_X1Y126_I;
  assign RIOI3_X105Y125_ILOGIC_X1Y125_O = RIOB33_X105Y125_IOB_X1Y125_I;
  assign RIOI3_X105Y127_ILOGIC_X1Y128_O = RIOB33_X105Y127_IOB_X1Y128_I;
  assign RIOI3_X105Y127_ILOGIC_X1Y127_O = RIOB33_X105Y127_IOB_X1Y127_I;
  assign RIOI3_X105Y129_ILOGIC_X1Y130_O = RIOB33_X105Y129_IOB_X1Y130_I;
  assign RIOI3_X105Y129_ILOGIC_X1Y129_O = RIOB33_X105Y129_IOB_X1Y129_I;
  assign RIOI3_X105Y133_ILOGIC_X1Y134_O = RIOB33_X105Y133_IOB_X1Y134_I;
  assign RIOI3_X105Y133_ILOGIC_X1Y133_O = RIOB33_X105Y133_IOB_X1Y133_I;
  assign RIOI3_X105Y135_ILOGIC_X1Y136_O = RIOB33_X105Y135_IOB_X1Y136_I;
  assign RIOI3_X105Y135_ILOGIC_X1Y135_O = RIOB33_X105Y135_IOB_X1Y135_I;
  assign RIOI3_X105Y139_ILOGIC_X1Y140_O = RIOB33_X105Y139_IOB_X1Y140_I;
  assign RIOI3_X105Y139_ILOGIC_X1Y139_O = RIOB33_X105Y139_IOB_X1Y139_I;
  assign RIOI3_X105Y141_ILOGIC_X1Y142_O = RIOB33_X105Y141_IOB_X1Y142_I;
  assign RIOI3_X105Y141_ILOGIC_X1Y141_O = RIOB33_X105Y141_IOB_X1Y141_I;
  assign RIOI3_X105Y145_ILOGIC_X1Y146_O = RIOB33_X105Y145_IOB_X1Y146_I;
  assign RIOI3_X105Y145_ILOGIC_X1Y145_O = RIOB33_X105Y145_IOB_X1Y145_I;
  assign RIOI3_X105Y147_ILOGIC_X1Y148_O = RIOB33_X105Y147_IOB_X1Y148_I;
  assign RIOI3_X105Y147_ILOGIC_X1Y147_O = RIOB33_X105Y147_IOB_X1Y147_I;
  assign RIOI3_X105Y151_OLOGIC_X1Y152_OQ = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign RIOI3_X105Y151_OLOGIC_X1Y152_TQ = 1'b1;
  assign RIOI3_X105Y151_OLOGIC_X1Y151_OQ = LIOB33_X0Y75_IOB_X0Y76_I;
  assign RIOI3_X105Y151_OLOGIC_X1Y151_TQ = 1'b1;
  assign RIOI3_X105Y153_OLOGIC_X1Y154_OQ = RIOB33_X105Y101_IOB_X1Y102_I;
  assign RIOI3_X105Y153_OLOGIC_X1Y154_TQ = 1'b1;
  assign RIOI3_X105Y153_OLOGIC_X1Y153_OQ = RIOB33_X105Y101_IOB_X1Y101_I;
  assign RIOI3_X105Y153_OLOGIC_X1Y153_TQ = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y156_OQ = RIOB33_X105Y103_IOB_X1Y104_I;
  assign RIOI3_X105Y155_OLOGIC_X1Y156_TQ = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y155_OQ = RIOB33_X105Y103_IOB_X1Y103_I;
  assign RIOI3_X105Y155_OLOGIC_X1Y155_TQ = 1'b1;
  assign RIOI3_X105Y159_OLOGIC_X1Y160_OQ = CLBLM_R_X11Y151_SLICE_X14Y151_DO5;
  assign RIOI3_X105Y159_OLOGIC_X1Y160_TQ = 1'b1;
  assign RIOI3_X105Y159_OLOGIC_X1Y159_OQ = CLBLM_R_X11Y151_SLICE_X14Y151_DO6;
  assign RIOI3_X105Y159_OLOGIC_X1Y159_TQ = 1'b1;
  assign RIOI3_X105Y161_OLOGIC_X1Y162_OQ = CLBLM_L_X10Y152_SLICE_X13Y152_CO5;
  assign RIOI3_X105Y161_OLOGIC_X1Y162_TQ = 1'b1;
  assign RIOI3_X105Y161_OLOGIC_X1Y161_OQ = CLBLM_L_X10Y152_SLICE_X13Y152_CO6;
  assign RIOI3_X105Y161_OLOGIC_X1Y161_TQ = 1'b1;
  assign RIOI3_X105Y165_OLOGIC_X1Y166_OQ = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign RIOI3_X105Y165_OLOGIC_X1Y166_TQ = 1'b1;
  assign RIOI3_X105Y165_OLOGIC_X1Y165_OQ = RIOB33_X105Y125_IOB_X1Y125_I;
  assign RIOI3_X105Y165_OLOGIC_X1Y165_TQ = 1'b1;
  assign RIOI3_X105Y167_OLOGIC_X1Y168_OQ = CLBLM_L_X8Y159_SLICE_X10Y159_AO6;
  assign RIOI3_X105Y167_OLOGIC_X1Y168_TQ = 1'b1;
  assign RIOI3_X105Y167_OLOGIC_X1Y167_OQ = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign RIOI3_X105Y167_OLOGIC_X1Y167_TQ = 1'b1;
  assign RIOI3_X105Y171_OLOGIC_X1Y172_OQ = CLBLM_R_X103Y170_SLICE_X163Y170_AO5;
  assign RIOI3_X105Y171_OLOGIC_X1Y172_TQ = 1'b1;
  assign RIOI3_X105Y171_OLOGIC_X1Y171_OQ = CLBLM_R_X11Y157_SLICE_X14Y157_AO5;
  assign RIOI3_X105Y171_OLOGIC_X1Y171_TQ = 1'b1;
  assign RIOI3_X105Y173_OLOGIC_X1Y174_OQ = CLBLM_R_X103Y173_SLICE_X163Y173_AO5;
  assign RIOI3_X105Y173_OLOGIC_X1Y174_TQ = 1'b1;
  assign RIOI3_X105Y173_OLOGIC_X1Y173_OQ = CLBLM_R_X103Y173_SLICE_X163Y173_AO6;
  assign RIOI3_X105Y173_OLOGIC_X1Y173_TQ = 1'b1;
  assign RIOI3_X105Y175_OLOGIC_X1Y176_OQ = CLBLM_R_X103Y176_SLICE_X163Y176_AO6;
  assign RIOI3_X105Y175_OLOGIC_X1Y176_TQ = 1'b1;
  assign RIOI3_X105Y175_OLOGIC_X1Y175_OQ = CLBLM_R_X15Y153_SLICE_X20Y153_AO6;
  assign RIOI3_X105Y175_OLOGIC_X1Y175_TQ = 1'b1;
  assign RIOI3_X105Y177_OLOGIC_X1Y178_OQ = CLBLM_R_X103Y178_SLICE_X163Y178_AO6;
  assign RIOI3_X105Y177_OLOGIC_X1Y178_TQ = 1'b1;
  assign RIOI3_X105Y177_OLOGIC_X1Y177_OQ = CLBLM_R_X103Y176_SLICE_X163Y176_AO5;
  assign RIOI3_X105Y177_OLOGIC_X1Y177_TQ = 1'b1;
  assign RIOI3_X105Y179_OLOGIC_X1Y180_OQ = CLBLM_R_X11Y151_SLICE_X14Y151_DO6;
  assign RIOI3_X105Y179_OLOGIC_X1Y180_TQ = 1'b1;
  assign RIOI3_X105Y179_OLOGIC_X1Y179_OQ = CLBLM_R_X103Y178_SLICE_X163Y178_AO5;
  assign RIOI3_X105Y179_OLOGIC_X1Y179_TQ = 1'b1;
  assign RIOI3_X105Y183_OLOGIC_X1Y184_OQ = CLBLM_L_X10Y150_SLICE_X13Y150_DO6;
  assign RIOI3_X105Y183_OLOGIC_X1Y184_TQ = 1'b1;
  assign RIOI3_X105Y183_OLOGIC_X1Y183_OQ = CLBLM_L_X10Y152_SLICE_X13Y152_CO5;
  assign RIOI3_X105Y183_OLOGIC_X1Y183_TQ = 1'b1;
  assign RIOI3_X105Y185_OLOGIC_X1Y186_OQ = CLBLM_L_X12Y151_SLICE_X16Y151_AQ;
  assign RIOI3_X105Y185_OLOGIC_X1Y186_TQ = 1'b1;
  assign RIOI3_X105Y185_OLOGIC_X1Y185_OQ = CLBLM_L_X10Y150_SLICE_X13Y150_DO5;
  assign RIOI3_X105Y185_OLOGIC_X1Y185_TQ = 1'b1;
  assign RIOI3_X105Y189_OLOGIC_X1Y190_OQ = CLBLM_L_X12Y152_SLICE_X17Y152_AQ;
  assign RIOI3_X105Y189_OLOGIC_X1Y190_TQ = 1'b1;
  assign RIOI3_X105Y189_OLOGIC_X1Y189_OQ = CLBLM_R_X11Y153_SLICE_X14Y153_CQ;
  assign RIOI3_X105Y189_OLOGIC_X1Y189_TQ = 1'b1;
  assign RIOI3_X105Y191_OLOGIC_X1Y192_OQ = CLBLM_R_X11Y151_SLICE_X15Y151_AQ;
  assign RIOI3_X105Y191_OLOGIC_X1Y192_TQ = 1'b1;
  assign RIOI3_X105Y191_OLOGIC_X1Y191_OQ = CLBLM_L_X10Y149_SLICE_X12Y149_AQ;
  assign RIOI3_X105Y191_OLOGIC_X1Y191_TQ = 1'b1;
  assign RIOI3_X105Y195_OLOGIC_X1Y196_OQ = CLBLM_R_X11Y153_SLICE_X14Y153_BQ;
  assign RIOI3_X105Y195_OLOGIC_X1Y196_TQ = 1'b1;
  assign RIOI3_X105Y195_OLOGIC_X1Y195_OQ = CLBLM_R_X11Y151_SLICE_X14Y151_AQ;
  assign RIOI3_X105Y195_OLOGIC_X1Y195_TQ = 1'b1;
  assign RIOI3_X105Y197_OLOGIC_X1Y198_OQ = CLBLM_L_X16Y158_SLICE_X22Y158_AO6;
  assign RIOI3_X105Y197_OLOGIC_X1Y198_TQ = 1'b1;
  assign RIOI3_X105Y197_OLOGIC_X1Y197_OQ = CLBLM_L_X16Y158_SLICE_X22Y158_AO6;
  assign RIOI3_X105Y197_OLOGIC_X1Y197_TQ = 1'b1;
  assign RIOI3_SING_X105Y100_ILOGIC_X1Y100_O = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign RIOI3_SING_X105Y149_ILOGIC_X1Y149_O = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign RIOI3_SING_X105Y150_OLOGIC_X1Y150_OQ = LIOB33_X0Y75_IOB_X0Y75_I;
  assign RIOI3_SING_X105Y150_OLOGIC_X1Y150_TQ = 1'b1;
  assign RIOI3_SING_X105Y199_OLOGIC_X1Y199_OQ = CLBLM_L_X12Y155_SLICE_X17Y155_AQ;
  assign RIOI3_SING_X105Y199_OLOGIC_X1Y199_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_O = RIOB33_X105Y107_IOB_X1Y108_I;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_O = RIOB33_X105Y107_IOB_X1Y107_I;
  assign RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_O = RIOB33_X105Y119_IOB_X1Y119_I;
  assign RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y132_O = RIOB33_X105Y131_IOB_X1Y132_I;
  assign RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y131_O = RIOB33_X105Y131_IOB_X1Y131_I;
  assign RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y144_O = RIOB33_X105Y143_IOB_X1Y144_I;
  assign RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y143_O = RIOB33_X105Y143_IOB_X1Y143_I;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_OQ = CLBLL_L_X36Y146_SLICE_X54Y146_AO6;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_OQ = RIOB33_X105Y125_IOB_X1Y126_I;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_OQ = CLBLM_R_X103Y170_SLICE_X163Y170_AO6;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_OQ = CLBLM_R_X103Y169_SLICE_X163Y169_AO6;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_OQ = CLBLM_L_X10Y152_SLICE_X13Y152_CO6;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_OQ = CLBLM_R_X11Y151_SLICE_X14Y151_DO5;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_OQ = CLBLM_L_X12Y155_SLICE_X17Y155_AQ;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_OQ = CLBLM_R_X11Y153_SLICE_X14Y153_AQ;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y114_O = RIOB33_X105Y113_IOB_X1Y114_I;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_O = RIOB33_X105Y113_IOB_X1Y113_I;
  assign RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y138_O = RIOB33_X105Y137_IOB_X1Y138_I;
  assign RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y137_O = RIOB33_X105Y137_IOB_X1Y137_I;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_OQ = CLBLM_L_X10Y150_SLICE_X13Y150_DO5;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_OQ = CLBLM_L_X10Y150_SLICE_X13Y150_DO6;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_OQ = CLBLM_L_X10Y155_SLICE_X13Y155_AQ;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_OQ = CLBLM_R_X11Y151_SLICE_X14Y151_BQ;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_TQ = 1'b1;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_B1 = CLBLL_L_X4Y145_SLICE_X5Y145_DO6;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_B2 = CLBLM_L_X8Y145_SLICE_X10Y145_BQ;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_B4 = CLBLM_L_X8Y144_SLICE_X10Y144_DO6;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_B5 = 1'b1;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_B6 = CLBLM_R_X7Y153_SLICE_X9Y153_BQ;
  assign CLBLM_L_X10Y155_SLICE_X12Y155_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X10Y155_SLICE_X12Y155_D1 = CLBLM_L_X8Y155_SLICE_X10Y155_CO6;
  assign CLBLM_L_X10Y155_SLICE_X12Y155_D2 = CLBLM_L_X8Y153_SLICE_X11Y153_BQ;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_C1 = CLBLM_L_X10Y144_SLICE_X13Y144_AQ;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_C2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_C3 = CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_C4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_C5 = CLBLM_R_X5Y144_SLICE_X7Y144_AQ;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_C6 = 1'b1;
  assign CLBLM_L_X10Y155_SLICE_X12Y155_D3 = CLBLM_L_X8Y155_SLICE_X11Y155_DO6;
  assign CLBLM_L_X10Y155_SLICE_X12Y155_D4 = CLBLM_L_X8Y155_SLICE_X11Y155_CO6;
  assign CLBLM_L_X10Y155_SLICE_X12Y155_D5 = CLBLM_L_X10Y154_SLICE_X12Y154_AQ;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y155_SLICE_X12Y155_D6 = CLBLM_L_X8Y154_SLICE_X11Y154_DO6;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_D1 = CLBLM_L_X10Y144_SLICE_X13Y144_AQ;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_D2 = CLBLM_L_X8Y148_SLICE_X10Y148_CO6;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_D3 = CLBLL_L_X4Y154_SLICE_X4Y154_CO6;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_D4 = CLBLM_L_X8Y145_SLICE_X10Y145_CO6;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_D5 = CLBLM_R_X5Y144_SLICE_X7Y144_AQ;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_D6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_A1 = CLBLM_R_X11Y149_SLICE_X15Y149_DO6;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_A2 = CLBLM_R_X11Y149_SLICE_X14Y149_BQ;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_A3 = CLBLM_L_X12Y149_SLICE_X16Y149_AQ;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_A4 = CLBLM_R_X11Y149_SLICE_X15Y149_BO6;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_A5 = CLBLM_R_X11Y150_SLICE_X15Y150_AQ;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_A6 = CLBLM_L_X10Y150_SLICE_X13Y150_BQ;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_B1 = CLBLM_L_X10Y151_SLICE_X12Y151_BQ;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_B2 = CLBLM_L_X12Y149_SLICE_X17Y149_AQ;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_B3 = CLBLM_L_X12Y148_SLICE_X16Y148_AQ;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_B4 = CLBLM_L_X10Y149_SLICE_X13Y149_AQ;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_B5 = CLBLM_L_X12Y148_SLICE_X16Y148_BQ;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_B6 = CLBLM_L_X12Y150_SLICE_X16Y150_BQ;
  assign LIOI3_X0Y155_OLOGIC_X0Y156_D1 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_C1 = CLBLM_R_X11Y149_SLICE_X14Y149_DO6;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_C2 = 1'b1;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_C3 = CLBLM_R_X11Y150_SLICE_X15Y150_BQ;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_C4 = CLBLM_L_X10Y150_SLICE_X13Y150_BQ;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_C5 = CLBLM_R_X11Y149_SLICE_X15Y149_DO6;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_A1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_A2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_A3 = CLBLL_L_X2Y152_SLICE_X1Y152_AO6;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_A4 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_A5 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_A6 = 1'b1;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_C6 = CLBLM_R_X11Y149_SLICE_X15Y149_BO6;
  assign LIOI3_X0Y155_OLOGIC_X0Y156_T1 = 1'b1;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_B1 = CLBLL_L_X2Y151_SLICE_X1Y151_AO6;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_B2 = CLBLM_R_X5Y147_SLICE_X7Y147_BQ;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_B3 = CLBLL_L_X2Y151_SLICE_X0Y151_CO5;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_B4 = CLBLL_L_X2Y155_SLICE_X1Y155_DO6;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_B5 = CLBLL_L_X2Y152_SLICE_X1Y152_AO6;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_B6 = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_D1 = CLBLM_R_X11Y149_SLICE_X14Y149_AQ;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_D2 = 1'b1;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_D3 = 1'b1;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_C1 = CLBLL_L_X2Y151_SLICE_X0Y151_CO5;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_C2 = CLBLL_L_X4Y149_SLICE_X5Y149_CQ;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_C3 = 1'b1;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_C4 = CLBLL_L_X4Y153_SLICE_X5Y153_AQ;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_C5 = CLBLL_L_X2Y154_SLICE_X1Y154_BO5;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_C6 = CLBLL_L_X2Y155_SLICE_X1Y155_DO6;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_A1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_A2 = CLBLM_R_X5Y151_SLICE_X6Y151_BQ;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_A3 = CLBLM_R_X11Y149_SLICE_X14Y149_AQ;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_A4 = CLBLM_L_X10Y149_SLICE_X13Y149_AQ;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_A6 = CLBLM_R_X11Y147_SLICE_X14Y147_CO6;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_D1 = 1'b1;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_D2 = CLBLL_L_X4Y152_SLICE_X5Y152_AO5;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_D3 = CLBLM_L_X10Y152_SLICE_X12Y152_D5Q;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_D4 = 1'b1;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_D5 = CLBLM_R_X3Y146_SLICE_X3Y146_AQ;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_D6 = CLBLL_L_X2Y152_SLICE_X1Y152_BO6;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_B3 = CLBLM_R_X11Y149_SLICE_X14Y149_AQ;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_B5 = CLBLM_L_X8Y153_SLICE_X11Y153_BQ;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_B6 = CLBLM_R_X11Y147_SLICE_X14Y147_CO6;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_C1 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_C2 = 1'b1;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_C3 = CLBLM_R_X11Y145_SLICE_X14Y145_DO6;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_C5 = CLBLM_R_X5Y142_SLICE_X7Y142_AQ;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_C6 = CLBLM_R_X7Y151_SLICE_X9Y151_BQ;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_D1 = CLBLM_R_X11Y147_SLICE_X14Y147_AQ;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_D2 = CLBLM_L_X12Y149_SLICE_X16Y149_AQ;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_D3 = CLBLM_R_X11Y149_SLICE_X14Y149_BQ;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_D4 = CLBLM_R_X11Y150_SLICE_X15Y150_AQ;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_D5 = CLBLM_L_X12Y147_SLICE_X16Y147_AQ;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_D6 = 1'b1;
  assign RIOB33_SING_X105Y150_IOB_X1Y150_O = LIOB33_X0Y75_IOB_X0Y75_I;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_D1 = CLBLM_L_X10Y152_SLICE_X13Y152_CO6;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_A1 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_A2 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_A3 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_A4 = CLBLL_L_X2Y155_SLICE_X1Y155_DO6;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_A5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_A6 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_A4 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_A5 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_A1 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_A2 = CLBLM_R_X3Y154_SLICE_X2Y154_BO6;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_A3 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_A4 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_A5 = CLBLL_L_X2Y153_SLICE_X1Y153_DO6;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_A6 = 1'b1;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_B1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_B2 = CLBLL_L_X2Y155_SLICE_X1Y155_DO6;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_B3 = CLBLL_L_X2Y152_SLICE_X1Y152_AO6;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_C1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_C2 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_C3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_B1 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_C5 = CLBLL_L_X2Y155_SLICE_X1Y155_DO6;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_C6 = CLBLL_L_X4Y147_SLICE_X5Y147_AQ;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_B2 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_B3 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_B4 = CLBLL_L_X2Y151_SLICE_X1Y151_BO6;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_B5 = CLBLM_R_X3Y151_SLICE_X3Y151_AO6;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_B6 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_C1 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_C2 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_C3 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_C4 = CLBLM_R_X3Y152_SLICE_X3Y152_CO6;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_C5 = CLBLM_R_X3Y153_SLICE_X2Y153_DO6;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_C6 = 1'b1;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_D1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_D2 = CLBLM_L_X8Y150_SLICE_X11Y150_BQ;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_D3 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_D4 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_D5 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_D1 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_D2 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_D3 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_D4 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_D5 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_D6 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_B3 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_B4 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_B5 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_B6 = 1'b1;
  assign CLBLM_L_X10Y156_SLICE_X13Y156_A1 = 1'b1;
  assign CLBLM_L_X10Y156_SLICE_X13Y156_A2 = 1'b1;
  assign CLBLM_L_X10Y156_SLICE_X13Y156_A3 = 1'b1;
  assign CLBLM_L_X10Y156_SLICE_X13Y156_A4 = 1'b1;
  assign CLBLM_L_X10Y156_SLICE_X13Y156_A5 = 1'b1;
  assign CLBLM_L_X10Y156_SLICE_X13Y156_A6 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_A1 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_A2 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_A3 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_A4 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_A5 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_A6 = 1'b1;
  assign CLBLM_L_X10Y156_SLICE_X13Y156_B1 = 1'b1;
  assign CLBLM_L_X10Y156_SLICE_X13Y156_B2 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_B1 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_B2 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_B3 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_B4 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_B5 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_B6 = 1'b1;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_A1 = CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_A2 = CLBLM_L_X8Y145_SLICE_X11Y145_DQ;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_A3 = CLBLM_L_X8Y146_SLICE_X11Y146_AQ;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_C1 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_C2 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_C3 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_C4 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_C5 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_C6 = 1'b1;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_A5 = 1'b1;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_A6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_B1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_B2 = CLBLM_L_X8Y146_SLICE_X11Y146_BQ;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_B3 = CLBLM_L_X8Y146_SLICE_X11Y146_AQ;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_B4 = CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_D1 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_D2 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_D3 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_D4 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_D5 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_D6 = 1'b1;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_C1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_C2 = CLBLM_L_X8Y145_SLICE_X11Y145_DQ;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_C3 = CLBLM_R_X5Y149_SLICE_X6Y149_CO6;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_C4 = CLBLM_L_X10Y147_SLICE_X13Y147_AQ;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_C5 = CLBLM_L_X8Y146_SLICE_X11Y146_DO6;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_C6 = CLBLM_R_X3Y153_SLICE_X2Y153_DO6;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_D1 = CLBLL_L_X4Y150_SLICE_X4Y150_AQ;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_D2 = CLBLL_L_X4Y149_SLICE_X4Y149_DQ;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_D3 = 1'b1;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_D4 = CLBLM_L_X8Y146_SLICE_X11Y146_AQ;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_D5 = CLBLM_R_X11Y146_SLICE_X14Y146_BQ;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_D6 = 1'b1;
  assign CLBLM_L_X10Y156_SLICE_X12Y156_B1 = CLBLM_L_X10Y156_SLICE_X12Y156_DO6;
  assign CLBLM_L_X10Y156_SLICE_X12Y156_B2 = CLBLM_L_X10Y155_SLICE_X12Y155_AQ;
  assign CLBLM_L_X10Y156_SLICE_X12Y156_B3 = CLBLM_L_X8Y154_SLICE_X11Y154_DO6;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_A1 = CLBLM_L_X8Y147_SLICE_X11Y147_AO5;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_A2 = CLBLM_L_X8Y152_SLICE_X10Y152_DQ;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_A5 = 1'b1;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_A6 = CLBLM_R_X7Y146_SLICE_X8Y146_DQ;
  assign CLBLM_L_X10Y156_SLICE_X12Y156_C1 = CLBLM_L_X10Y156_SLICE_X12Y156_AO6;
  assign CLBLM_L_X10Y156_SLICE_X12Y156_C2 = CLBLM_L_X10Y155_SLICE_X13Y155_CQ;
  assign CLBLM_L_X10Y156_SLICE_X12Y156_C3 = CLBLM_L_X8Y154_SLICE_X11Y154_DO6;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_B1 = CLBLM_R_X7Y146_SLICE_X8Y146_CQ;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_B2 = CLBLM_R_X3Y148_SLICE_X2Y148_CQ;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_B4 = RIOB33_X105Y119_IOB_X1Y119_I;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_B5 = CLBLM_L_X8Y146_SLICE_X10Y146_BQ;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_B6 = 1'b1;
  assign CLBLM_L_X10Y156_SLICE_X12Y156_D1 = CLBLM_L_X8Y155_SLICE_X11Y155_CO6;
  assign CLBLM_L_X10Y156_SLICE_X12Y156_D2 = CLBLM_L_X10Y154_SLICE_X12Y154_DQ;
  assign CLBLM_L_X10Y156_SLICE_X12Y156_D3 = CLBLM_L_X8Y153_SLICE_X11Y153_BQ;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_C1 = CLBLM_L_X8Y147_SLICE_X11Y147_CO6;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_C2 = CLBLM_L_X10Y147_SLICE_X13Y147_AQ;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_C5 = 1'b1;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_C6 = CLBLM_L_X8Y142_SLICE_X10Y142_A5Q;
  assign CLBLM_L_X10Y156_SLICE_X12Y156_D4 = CLBLM_L_X10Y155_SLICE_X13Y155_CQ;
  assign CLBLM_L_X10Y156_SLICE_X12Y156_D5 = CLBLM_L_X8Y155_SLICE_X10Y155_AQ;
  assign CLBLM_L_X10Y156_SLICE_X12Y156_D6 = CLBLM_L_X10Y155_SLICE_X13Y155_BQ;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_D1 = CLBLM_L_X8Y148_SLICE_X10Y148_CO5;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_D2 = CLBLL_L_X2Y153_SLICE_X1Y153_DO6;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_D3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_D4 = CLBLM_R_X5Y144_SLICE_X7Y144_AQ;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_D5 = 1'b1;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_D6 = CLBLM_L_X10Y144_SLICE_X13Y144_AQ;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_A1 = CLBLM_R_X11Y147_SLICE_X14Y147_CO6;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_A2 = CLBLM_R_X11Y151_SLICE_X15Y151_AQ;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_A3 = CLBLM_R_X11Y150_SLICE_X15Y150_AQ;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_A4 = CLBLM_R_X11Y150_SLICE_X15Y150_DO6;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_B1 = CLBLM_R_X11Y147_SLICE_X14Y147_CO6;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_B3 = CLBLM_L_X10Y147_SLICE_X13Y147_AQ;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_B4 = CLBLM_L_X10Y150_SLICE_X13Y150_BQ;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_B6 = CLBLM_R_X11Y150_SLICE_X15Y150_BQ;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_A1 = CLBLL_L_X4Y148_SLICE_X4Y148_DQ;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_A2 = CLBLM_R_X5Y153_SLICE_X6Y153_BQ;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_A3 = CLBLL_L_X2Y151_SLICE_X0Y151_CO5;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_A4 = CLBLL_L_X2Y152_SLICE_X1Y152_AO6;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_A5 = CLBLL_L_X2Y154_SLICE_X1Y154_BO5;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_A6 = CLBLL_L_X2Y155_SLICE_X1Y155_DO6;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_C1 = CLBLM_R_X11Y146_SLICE_X15Y146_BQ;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_C2 = CLBLM_R_X11Y150_SLICE_X15Y150_CQ;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_C3 = CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_B1 = CLBLM_R_X3Y155_SLICE_X3Y155_DO6;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_B2 = CLBLL_L_X4Y149_SLICE_X4Y149_BQ;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_B3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_B4 = CLBLL_L_X2Y155_SLICE_X1Y155_DO6;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_B5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_B6 = CLBLM_L_X8Y152_SLICE_X10Y152_AQ;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_D1 = CLBLM_L_X8Y147_SLICE_X11Y147_BO6;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_C1 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_C2 = CLBLL_L_X2Y152_SLICE_X1Y152_AO5;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_C3 = CLBLM_R_X5Y153_SLICE_X7Y153_BQ;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_C4 = CLBLL_L_X4Y155_SLICE_X4Y155_BO6;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_C5 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_C6 = CLBLL_L_X4Y150_SLICE_X4Y150_BQ;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_D3 = CLBLM_R_X11Y151_SLICE_X14Y151_BO5;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_D4 = CLBLM_R_X11Y150_SLICE_X15Y150_BQ;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_A1 = CLBLM_R_X11Y147_SLICE_X14Y147_CO6;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_A2 = CLBLM_L_X10Y151_SLICE_X13Y151_AQ;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_A3 = CLBLM_L_X8Y151_SLICE_X11Y151_BQ;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_A4 = CLBLM_R_X11Y151_SLICE_X15Y151_BQ;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_A5 = CLBLM_L_X10Y151_SLICE_X13Y151_BQ;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_A6 = CLBLM_R_X11Y150_SLICE_X14Y150_CO6;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_D1 = CLBLL_L_X4Y155_SLICE_X5Y155_AO6;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_D2 = CLBLM_R_X5Y153_SLICE_X6Y153_BQ;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_D3 = CLBLL_L_X4Y154_SLICE_X5Y154_AQ;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_D4 = CLBLL_L_X4Y152_SLICE_X4Y152_AO6;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_D5 = CLBLL_L_X4Y148_SLICE_X4Y148_DQ;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_D6 = CLBLM_R_X3Y152_SLICE_X2Y152_AO5;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_B1 = CLBLM_R_X11Y151_SLICE_X14Y151_BO5;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_B2 = CLBLM_R_X11Y149_SLICE_X15Y149_CO6;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_B3 = CLBLM_R_X11Y150_SLICE_X14Y150_DO6;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_B4 = CLBLM_R_X11Y147_SLICE_X14Y147_CO6;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_B5 = CLBLM_L_X8Y147_SLICE_X11Y147_BO6;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_B6 = CLBLM_L_X12Y149_SLICE_X16Y149_BO6;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_C1 = CLBLM_L_X8Y147_SLICE_X11Y147_BO6;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_C2 = CLBLM_R_X11Y149_SLICE_X15Y149_CO6;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_C3 = CLBLM_R_X11Y151_SLICE_X14Y151_BO5;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_C1 = CLBLM_L_X12Y153_SLICE_X16Y153_DO6;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_C4 = CLBLM_L_X12Y149_SLICE_X16Y149_BO6;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_C5 = CLBLM_R_X11Y150_SLICE_X14Y150_DO6;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_C6 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_C2 = CLBLM_R_X11Y153_SLICE_X14Y153_CO5;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_D1 = CLBLM_L_X10Y151_SLICE_X12Y151_AQ;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_D2 = CLBLM_L_X12Y148_SLICE_X16Y148_AQ;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_D3 = CLBLM_L_X10Y149_SLICE_X13Y149_AQ;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_D4 = 1'b1;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_A1 = CLBLL_L_X4Y153_SLICE_X5Y153_AQ;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_A2 = CLBLM_R_X5Y153_SLICE_X6Y153_AQ;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_A3 = CLBLM_R_X5Y151_SLICE_X6Y151_BQ;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_A5 = CLBLM_R_X5Y152_SLICE_X7Y152_DO5;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_A6 = 1'b1;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_D5 = CLBLM_L_X12Y150_SLICE_X16Y150_AQ;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_D6 = CLBLM_R_X11Y149_SLICE_X14Y149_DO5;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_B1 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_B2 = CLBLM_R_X5Y153_SLICE_X7Y153_AQ;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_B3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_B4 = CLBLL_L_X2Y155_SLICE_X1Y155_DO6;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_B5 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_B6 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_C1 = CLBLL_L_X4Y152_SLICE_X5Y152_AO6;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_C2 = CLBLM_R_X5Y153_SLICE_X6Y153_AQ;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_C3 = CLBLL_L_X2Y154_SLICE_X1Y154_AO5;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_C4 = CLBLM_R_X7Y151_SLICE_X9Y151_AQ;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_C5 = CLBLL_L_X4Y152_SLICE_X5Y152_DO6;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_C6 = CLBLL_L_X4Y153_SLICE_X5Y153_BO6;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_D1 = CLBLL_L_X4Y152_SLICE_X5Y152_AO6;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_D2 = CLBLM_L_X8Y152_SLICE_X10Y152_AQ;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_D3 = CLBLL_L_X4Y146_SLICE_X5Y146_AQ;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_D4 = CLBLL_L_X4Y149_SLICE_X4Y149_BQ;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_D5 = CLBLM_R_X5Y154_SLICE_X7Y154_AO6;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_D6 = CLBLL_L_X2Y152_SLICE_X1Y152_BO6;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_C4 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_C5 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_C6 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_D3 = CLBLM_L_X12Y153_SLICE_X17Y153_DO6;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_D4 = CLBLM_L_X12Y153_SLICE_X16Y153_AQ;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_A1 = CLBLM_L_X10Y151_SLICE_X12Y151_BQ;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_A3 = CLBLM_R_X5Y148_SLICE_X6Y148_BQ;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_A4 = CLBLM_R_X7Y144_SLICE_X8Y144_BQ;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_A5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_A6 = 1'b1;
  assign LIOB33_X0Y153_IOB_X0Y154_O = LIOB33_X0Y67_IOB_X0Y68_I;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_B1 = CLBLM_R_X5Y149_SLICE_X6Y149_CO6;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_B2 = CLBLM_R_X7Y145_SLICE_X9Y145_BQ;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_B3 = CLBLL_L_X2Y153_SLICE_X1Y153_DO6;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_B4 = 1'b1;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_B5 = CLBLM_L_X8Y151_SLICE_X10Y151_AQ;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_B6 = 1'b1;
  assign LIOB33_X0Y153_IOB_X0Y153_O = LIOB33_X0Y67_IOB_X0Y67_I;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_C1 = CLBLM_R_X7Y146_SLICE_X9Y146_DO6;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_C2 = CLBLM_R_X7Y147_SLICE_X9Y147_DO6;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_C3 = CLBLM_L_X10Y146_SLICE_X12Y146_DQ;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_C4 = CLBLM_L_X10Y149_SLICE_X13Y149_DQ;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_C5 = CLBLM_L_X8Y147_SLICE_X11Y147_DO6;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_C6 = CLBLM_L_X10Y150_SLICE_X12Y150_BQ;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_D1 = CLBLM_L_X10Y146_SLICE_X13Y146_AQ;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_D2 = CLBLM_L_X10Y147_SLICE_X13Y147_BQ;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_D3 = CLBLM_R_X7Y147_SLICE_X8Y147_CQ;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_D4 = CLBLL_L_X4Y148_SLICE_X4Y148_CQ;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_D5 = CLBLM_L_X8Y145_SLICE_X10Y145_AQ;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_D6 = CLBLM_R_X5Y148_SLICE_X6Y148_BQ;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_A1 = CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_A2 = CLBLL_L_X4Y144_SLICE_X5Y144_A5Q;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_A3 = CLBLM_L_X8Y147_SLICE_X10Y147_AQ;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_A5 = CLBLM_R_X7Y149_SLICE_X9Y149_DO6;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_A6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_B1 = CLBLM_L_X8Y152_SLICE_X11Y152_BO6;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_B2 = CLBLM_L_X8Y147_SLICE_X10Y147_BQ;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_B3 = CLBLM_L_X8Y145_SLICE_X10Y145_AQ;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_B4 = CLBLM_R_X7Y145_SLICE_X8Y145_CQ;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_B5 = 1'b1;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_C1 = CLBLM_L_X10Y152_SLICE_X12Y152_AQ;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_C1 = CLBLM_L_X8Y148_SLICE_X11Y148_CO6;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_C2 = CLBLM_L_X8Y147_SLICE_X10Y147_CQ;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_C3 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_C4 = CLBLM_L_X12Y150_SLICE_X16Y150_CQ;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_C5 = CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_D1 = CLBLM_L_X8Y150_SLICE_X10Y150_BQ;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_D2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_D3 = CLBLM_L_X8Y147_SLICE_X10Y147_DQ;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_D4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_D5 = 1'b1;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_D6 = 1'b1;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_A2 = 1'b1;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_A3 = CLBLM_R_X11Y151_SLICE_X15Y151_AQ;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_A4 = CLBLM_L_X10Y145_SLICE_X13Y145_A5Q;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_A5 = CLBLM_R_X5Y142_SLICE_X7Y142_AQ;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_A6 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_AX = CLBLM_R_X11Y151_SLICE_X14Y151_AO6;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_B1 = CLBLM_R_X5Y151_SLICE_X7Y151_DO6;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_B2 = CLBLM_R_X11Y151_SLICE_X15Y151_BQ;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_B4 = CLBLM_R_X11Y153_SLICE_X15Y153_BQ;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_B5 = CLBLM_R_X11Y147_SLICE_X14Y147_CO6;
  assign CLBLL_L_X4Y154_SLICE_X4Y154_A1 = CLBLL_L_X2Y155_SLICE_X1Y155_DO6;
  assign CLBLL_L_X4Y154_SLICE_X4Y154_A2 = CLBLL_L_X4Y155_SLICE_X4Y155_BO6;
  assign CLBLL_L_X4Y154_SLICE_X4Y154_A3 = CLBLL_L_X2Y151_SLICE_X1Y151_AO6;
  assign CLBLL_L_X4Y154_SLICE_X4Y154_A4 = CLBLL_L_X2Y152_SLICE_X1Y152_AO6;
  assign CLBLL_L_X4Y154_SLICE_X4Y154_A5 = CLBLL_L_X4Y150_SLICE_X5Y150_AQ;
  assign CLBLL_L_X4Y154_SLICE_X4Y154_A6 = CLBLM_R_X3Y148_SLICE_X3Y148_B5Q;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_C3 = CLBLM_R_X11Y154_SLICE_X15Y154_CO6;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_B6 = CLBLM_R_X11Y151_SLICE_X14Y151_BO5;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_D4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X4Y154_SLICE_X4Y154_B1 = 1'b1;
  assign CLBLL_L_X4Y154_SLICE_X4Y154_B2 = CLBLL_L_X4Y152_SLICE_X4Y152_BO6;
  assign CLBLL_L_X4Y154_SLICE_X4Y154_B3 = CLBLL_L_X4Y153_SLICE_X4Y153_AO6;
  assign CLBLL_L_X4Y154_SLICE_X4Y154_B4 = CLBLM_R_X3Y152_SLICE_X2Y152_AO5;
  assign CLBLL_L_X4Y154_SLICE_X4Y154_B5 = CLBLL_L_X4Y154_SLICE_X5Y154_AQ;
  assign CLBLL_L_X4Y154_SLICE_X4Y154_B6 = CLBLL_L_X4Y154_SLICE_X4Y154_AO6;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_C5 = CLBLM_L_X12Y151_SLICE_X16Y151_DO6;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_C4 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_C6 = 1'b1;
  assign CLBLL_L_X4Y154_SLICE_X4Y154_C1 = CLBLL_L_X2Y150_SLICE_X1Y150_CO6;
  assign CLBLL_L_X4Y154_SLICE_X4Y154_C2 = CLBLM_R_X5Y154_SLICE_X7Y154_DO6;
  assign CLBLL_L_X4Y154_SLICE_X4Y154_C3 = CLBLL_L_X4Y153_SLICE_X4Y153_DO6;
  assign CLBLL_L_X4Y154_SLICE_X4Y154_C4 = 1'b1;
  assign CLBLL_L_X4Y154_SLICE_X4Y154_C5 = CLBLL_L_X4Y154_SLICE_X4Y154_DO6;
  assign CLBLL_L_X4Y154_SLICE_X4Y154_C6 = CLBLM_R_X3Y155_SLICE_X2Y155_DO6;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_D1 = 1'b1;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_D2 = 1'b1;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_D3 = 1'b1;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_D4 = 1'b1;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_D5 = 1'b1;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_D6 = 1'b1;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_A1 = CLBLM_R_X11Y154_SLICE_X15Y154_CO6;
  assign CLBLL_L_X4Y154_SLICE_X4Y154_D1 = CLBLL_L_X4Y150_SLICE_X5Y150_AQ;
  assign CLBLL_L_X4Y154_SLICE_X4Y154_D2 = CLBLL_L_X4Y155_SLICE_X5Y155_AO5;
  assign CLBLL_L_X4Y154_SLICE_X4Y154_D3 = CLBLL_L_X2Y152_SLICE_X1Y152_BO5;
  assign CLBLL_L_X4Y154_SLICE_X4Y154_D4 = CLBLL_L_X4Y152_SLICE_X4Y152_BO6;
  assign CLBLL_L_X4Y154_SLICE_X4Y154_D5 = 1'b1;
  assign CLBLL_L_X4Y154_SLICE_X4Y154_D6 = CLBLM_R_X3Y148_SLICE_X3Y148_B5Q;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_A2 = CLBLM_R_X11Y148_SLICE_X14Y148_CQ;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_A3 = CLBLM_R_X7Y147_SLICE_X9Y147_AQ;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_A5 = CLBLM_R_X11Y151_SLICE_X15Y151_A5Q;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_A6 = 1'b1;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_AX = CLBLM_R_X11Y152_SLICE_X14Y152_CQ;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_B1 = CLBLM_L_X10Y151_SLICE_X13Y151_BQ;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_B2 = CLBLM_L_X10Y151_SLICE_X13Y151_AQ;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_B3 = CLBLM_R_X11Y147_SLICE_X14Y147_CO6;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_B4 = CLBLM_R_X11Y151_SLICE_X15Y151_BQ;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_B5 = CLBLM_L_X8Y151_SLICE_X11Y151_BQ;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_B6 = 1'b1;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_BX = CLBLM_R_X11Y148_SLICE_X15Y148_BQ;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_C1 = CLBLM_L_X8Y151_SLICE_X11Y151_BQ;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_C2 = CLBLM_L_X10Y151_SLICE_X13Y151_AQ;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_C3 = CLBLM_L_X10Y151_SLICE_X13Y151_BQ;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_C4 = CLBLM_R_X11Y147_SLICE_X14Y147_CO6;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_C5 = CLBLM_R_X11Y151_SLICE_X15Y151_BQ;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_C6 = 1'b1;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_CE = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLL_L_X4Y154_SLICE_X5Y154_A1 = 1'b1;
  assign CLBLL_L_X4Y154_SLICE_X5Y154_A2 = CLBLL_L_X4Y153_SLICE_X5Y153_AQ;
  assign CLBLL_L_X4Y154_SLICE_X5Y154_A3 = CLBLL_L_X4Y154_SLICE_X5Y154_AQ;
  assign CLBLL_L_X4Y154_SLICE_X5Y154_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y154_SLICE_X5Y154_A5 = CLBLM_R_X5Y150_SLICE_X7Y150_BQ;
  assign CLBLL_L_X4Y154_SLICE_X5Y154_A6 = CLBLM_R_X5Y152_SLICE_X7Y152_DO5;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_D1 = CLBLM_R_X11Y148_SLICE_X14Y148_AQ;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_D2 = CLBLM_R_X11Y148_SLICE_X14Y148_DQ;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_D3 = CLBLM_L_X10Y151_SLICE_X12Y151_DQ;
  assign CLBLL_L_X4Y154_SLICE_X5Y154_B1 = CLBLL_L_X4Y154_SLICE_X5Y154_BQ;
  assign CLBLL_L_X4Y154_SLICE_X5Y154_B2 = CLBLM_R_X3Y144_SLICE_X2Y144_CO6;
  assign CLBLL_L_X4Y154_SLICE_X5Y154_B3 = 1'b1;
  assign CLBLL_L_X4Y154_SLICE_X5Y154_B4 = CLBLL_L_X4Y147_SLICE_X5Y147_AQ;
  assign CLBLL_L_X4Y154_SLICE_X5Y154_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y154_SLICE_X5Y154_B6 = CLBLM_R_X7Y145_SLICE_X8Y145_C5Q;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_D3 = CLBLM_R_X7Y147_SLICE_X9Y147_AQ;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_A6 = CLBLM_R_X5Y154_SLICE_X6Y154_BO6;
  assign CLBLL_L_X4Y154_SLICE_X5Y154_C1 = 1'b1;
  assign CLBLL_L_X4Y154_SLICE_X5Y154_C2 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y154_SLICE_X5Y154_C3 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X4Y154_SLICE_X5Y154_C4 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X4Y154_SLICE_X5Y154_C5 = CLBLL_L_X2Y155_SLICE_X1Y155_DO6;
  assign CLBLL_L_X4Y154_SLICE_X5Y154_C6 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_D4 = CLBLM_L_X12Y150_SLICE_X16Y150_CQ;
  assign CLBLL_L_X4Y154_SLICE_X5Y154_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLL_L_X4Y154_SLICE_X5Y154_D1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y154_SLICE_X5Y154_D2 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X4Y154_SLICE_X5Y154_D3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y154_SLICE_X5Y154_D4 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X4Y154_SLICE_X5Y154_D5 = CLBLL_L_X4Y146_SLICE_X5Y146_AQ;
  assign CLBLL_L_X4Y154_SLICE_X5Y154_D6 = CLBLL_L_X2Y152_SLICE_X1Y152_AO6;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_B1 = CLBLM_L_X8Y153_SLICE_X11Y153_DQ;
  assign LIOI3_X0Y159_OLOGIC_X0Y160_D1 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign LIOI3_X0Y159_OLOGIC_X0Y160_T1 = 1'b1;
  assign LIOI3_X0Y159_OLOGIC_X0Y159_D1 = RIOB33_X105Y117_IOB_X1Y117_I;
  assign LIOI3_X0Y159_OLOGIC_X0Y159_T1 = 1'b1;
  assign LIOB33_X0Y155_IOB_X0Y156_O = RIOB33_X105Y105_IOB_X1Y106_I;
  assign LIOB33_X0Y155_IOB_X0Y155_O = LIOB33_X0Y69_IOB_X0Y70_I;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_C1 = CLBLM_R_X11Y154_SLICE_X15Y154_AQ;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_A1 = CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_A2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_A3 = CLBLM_L_X8Y148_SLICE_X11Y148_AQ;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_A4 = CLBLL_L_X4Y148_SLICE_X4Y148_BQ;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_A6 = CLBLM_R_X5Y148_SLICE_X7Y148_DO6;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_B1 = CLBLM_R_X7Y143_SLICE_X8Y143_AQ;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_B2 = CLBLM_L_X8Y149_SLICE_X10Y149_AO6;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_B3 = CLBLM_R_X7Y145_SLICE_X8Y145_BQ;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_B4 = CLBLM_R_X7Y152_SLICE_X9Y152_CQ;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_B5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_B6 = CLBLM_L_X8Y145_SLICE_X11Y145_A5Q;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_C4 = CLBLM_L_X10Y153_SLICE_X13Y153_CQ;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_D1 = CLBLM_L_X12Y155_SLICE_X17Y155_AQ;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_C1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_C2 = CLBLM_L_X8Y147_SLICE_X10Y147_DQ;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_C3 = CLBLL_L_X4Y143_SLICE_X4Y143_BQ;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_C4 = CLBLM_R_X5Y145_SLICE_X6Y145_CQ;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_C5 = CLBLM_R_X7Y147_SLICE_X8Y147_CQ;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_C6 = CLBLM_L_X8Y148_SLICE_X11Y148_DO6;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_T1 = 1'b1;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_D1 = CLBLM_R_X7Y145_SLICE_X8Y145_BQ;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_D2 = 1'b1;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_D3 = 1'b1;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_D4 = CLBLM_R_X7Y143_SLICE_X8Y143_AQ;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_D5 = 1'b1;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_D6 = 1'b1;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_B4 = CLBLM_R_X5Y152_SLICE_X7Y152_DO5;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_D1 = CLBLM_R_X11Y153_SLICE_X14Y153_AQ;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_A1 = CLBLM_L_X8Y148_SLICE_X10Y148_AQ;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_A3 = CLBLM_L_X10Y155_SLICE_X13Y155_AQ;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_A5 = CLBLM_R_X5Y147_SLICE_X7Y147_AQ;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_A6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_T1 = 1'b1;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_B1 = CLBLM_R_X7Y149_SLICE_X8Y149_CQ;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_B2 = CLBLM_R_X7Y146_SLICE_X9Y146_BQ;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_B4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_B5 = CLBLM_L_X8Y147_SLICE_X10Y147_AQ;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_B6 = 1'b1;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_BX = CLBLM_L_X8Y153_SLICE_X10Y153_CO6;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_C1 = CLBLM_L_X10Y146_SLICE_X12Y146_DQ;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_C2 = CLBLM_R_X11Y148_SLICE_X14Y148_BQ;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_C3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_C4 = CLBLM_L_X8Y152_SLICE_X10Y152_CQ;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_C5 = CLBLM_R_X7Y147_SLICE_X8Y147_CQ;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_C6 = 1'b1;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_D1 = CLBLM_R_X7Y145_SLICE_X8Y145_BQ;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_D2 = CLBLM_R_X7Y143_SLICE_X8Y143_AQ;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_D3 = CLBLM_L_X8Y148_SLICE_X10Y148_AQ;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_D4 = CLBLM_R_X5Y145_SLICE_X6Y145_CQ;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_D5 = CLBLL_L_X4Y143_SLICE_X4Y143_BQ;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_D6 = 1'b1;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_D3 = CLBLM_R_X11Y154_SLICE_X15Y154_BQ;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_D4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_D5 = CLBLM_L_X10Y153_SLICE_X13Y153_BQ;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_D6 = CLBLM_R_X7Y148_SLICE_X9Y148_BQ;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_A1 = CLBLM_L_X10Y154_SLICE_X13Y154_CO5;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_A2 = CLBLM_L_X8Y155_SLICE_X10Y155_BQ;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_A3 = CLBLM_R_X11Y152_SLICE_X15Y152_AQ;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_A4 = CLBLM_R_X11Y154_SLICE_X15Y154_CO5;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_A6 = CLBLM_L_X12Y152_SLICE_X17Y152_DO6;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_A1 = CLBLL_L_X4Y151_SLICE_X5Y151_B5Q;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_A2 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_A3 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_A4 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_A5 = 1'b1;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_A6 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_B3 = CLBLM_R_X11Y154_SLICE_X15Y154_CO6;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_B4 = CLBLM_L_X12Y151_SLICE_X16Y151_DO5;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_B1 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_B2 = CLBLL_L_X2Y152_SLICE_X1Y152_AO6;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_B3 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_B4 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_B5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_B6 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_A1 = CLBLL_L_X2Y151_SLICE_X1Y151_BO6;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_A2 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_A3 = CLBLM_R_X3Y152_SLICE_X3Y152_CO6;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_C1 = CLBLL_L_X4Y154_SLICE_X5Y154_BQ;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_C2 = LIOB33_X0Y67_IOB_X0Y68_I;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_C3 = CLBLL_L_X2Y154_SLICE_X1Y154_BO5;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_C4 = CLBLL_L_X2Y152_SLICE_X1Y152_AO5;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_C5 = CLBLL_L_X4Y155_SLICE_X4Y155_AO6;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_C6 = CLBLL_L_X4Y155_SLICE_X4Y155_BO6;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_B1 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_B2 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_B3 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_B4 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_B5 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_B6 = 1'b1;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_D1 = CLBLL_L_X4Y154_SLICE_X5Y154_BQ;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_D2 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_D3 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_D4 = CLBLL_L_X2Y152_SLICE_X1Y152_AO5;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_D5 = CLBLL_L_X4Y151_SLICE_X5Y151_B5Q;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_D6 = CLBLL_L_X4Y155_SLICE_X4Y155_BO6;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_C3 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_C4 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_C6 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_D1 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_D2 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_D3 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_D4 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_D5 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_D6 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_B1 = CLBLM_R_X11Y153_SLICE_X14Y153_BO5;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_B2 = CLBLL_L_X2Y146_SLICE_X1Y146_CQ;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_A1 = CLBLM_R_X7Y144_SLICE_X8Y144_DQ;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_A2 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_A3 = CLBLM_R_X5Y142_SLICE_X7Y142_AQ;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_A5 = CLBLM_R_X7Y147_SLICE_X8Y147_B5Q;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_A6 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_C2 = CLBLM_R_X11Y152_SLICE_X14Y152_CQ;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_C3 = CLBLM_R_X11Y152_SLICE_X14Y152_BQ;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_B1 = CLBLM_R_X7Y144_SLICE_X8Y144_DQ;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_A1 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_A2 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_A3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_A4 = CLBLL_L_X2Y155_SLICE_X1Y155_DO6;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_A5 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_A6 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_B2 = CLBLM_L_X8Y142_SLICE_X10Y142_AQ;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_B4 = CLBLM_R_X7Y142_SLICE_X8Y142_DO6;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_A1 = CLBLL_L_X4Y154_SLICE_X4Y154_CO6;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_A2 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_A3 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_A4 = CLBLM_R_X3Y150_SLICE_X2Y150_BO6;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_A5 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_A6 = 1'b1;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_B1 = 1'b1;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_B2 = 1'b1;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_B3 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_B1 = CLBLL_L_X4Y154_SLICE_X4Y154_CO6;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_B2 = CLBLL_L_X2Y151_SLICE_X1Y151_BO6;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_B3 = LIOB33_X0Y51_IOB_X0Y51_I;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_B4 = CLBLM_R_X3Y148_SLICE_X3Y148_BQ;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_B6 = CLBLM_R_X3Y141_SLICE_X2Y141_BO6;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_C1 = 1'b1;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_C2 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_C1 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_C2 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_C3 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_C4 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_C5 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_C6 = 1'b1;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_D1 = 1'b1;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_D2 = 1'b1;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_D3 = 1'b1;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_D6 = 1'b1;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_D4 = 1'b1;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_D5 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_D1 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_D2 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_D3 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_D4 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_D5 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X0Y141_D6 = 1'b1;
  assign LIOB33_X0Y157_IOB_X0Y158_O = RIOB33_X105Y115_IOB_X1Y116_I;
  assign LIOB33_X0Y157_IOB_X0Y157_O = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_B2 = CLBLM_R_X11Y149_SLICE_X14Y149_BQ;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_A1 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_A2 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_A3 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_A4 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_A5 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_A6 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_B1 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_B2 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_B3 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_B4 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_B5 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_B6 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_C1 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_C2 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_C3 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_C4 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_C5 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_C6 = 1'b1;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_A1 = 1'b1;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_A2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_A3 = CLBLM_L_X8Y149_SLICE_X11Y149_AQ;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_A4 = CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_A5 = CLBLM_L_X12Y149_SLICE_X17Y149_CQ;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_D1 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_D2 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_D3 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_D4 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_D5 = 1'b1;
  assign CLBLL_L_X2Y141_SLICE_X1Y141_D6 = 1'b1;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_B1 = CLBLM_R_X3Y151_SLICE_X3Y151_AO6;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_B3 = CLBLM_L_X10Y150_SLICE_X12Y150_DQ;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_B4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_B5 = CLBLM_L_X8Y149_SLICE_X11Y149_BQ;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_B6 = 1'b1;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_C1 = CLBLM_L_X8Y146_SLICE_X11Y146_CO6;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_C2 = CLBLM_L_X8Y149_SLICE_X11Y149_CQ;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_C4 = CLBLM_R_X7Y149_SLICE_X8Y149_BQ;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_C5 = CLBLM_L_X10Y149_SLICE_X12Y149_AO5;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_C6 = CLBLM_L_X8Y149_SLICE_X11Y149_DO6;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_D5 = CLBLM_L_X8Y151_SLICE_X11Y151_CQ;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_D6 = 1'b1;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_D1 = CLBLM_L_X8Y149_SLICE_X11Y149_BQ;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_D2 = CLBLM_L_X8Y149_SLICE_X11Y149_AQ;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_D3 = CLBLM_L_X8Y149_SLICE_X10Y149_DO6;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_D4 = CLBLM_L_X8Y149_SLICE_X10Y149_AO6;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_D5 = CLBLM_L_X8Y151_SLICE_X11Y151_DQ;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_D6 = CLBLM_L_X8Y148_SLICE_X11Y148_DO6;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_A1 = CLBLL_L_X4Y143_SLICE_X4Y143_BQ;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_A2 = 1'b1;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_A3 = CLBLM_R_X5Y145_SLICE_X6Y145_CQ;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_A4 = 1'b1;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_A5 = 1'b1;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_A6 = 1'b1;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_D4 = CLBLM_R_X5Y144_SLICE_X6Y144_DO6;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_B1 = CLBLM_L_X8Y145_SLICE_X11Y145_A5Q;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_B2 = CLBLM_L_X8Y151_SLICE_X10Y151_BQ;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_B3 = CLBLM_L_X8Y148_SLICE_X10Y148_AQ;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_B4 = CLBLM_R_X7Y152_SLICE_X9Y152_BQ;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_B5 = CLBLM_R_X7Y148_SLICE_X9Y148_AQ;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_B6 = CLBLM_R_X11Y148_SLICE_X14Y148_CQ;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_D1 = 1'b1;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_C1 = CLBLM_R_X3Y149_SLICE_X3Y149_BQ;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_C2 = CLBLM_L_X8Y149_SLICE_X10Y149_AO6;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_C3 = CLBLM_R_X7Y143_SLICE_X8Y143_AQ;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_C4 = CLBLM_R_X7Y145_SLICE_X8Y145_BQ;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_C5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_C6 = CLBLM_R_X5Y148_SLICE_X6Y148_BQ;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_D1 = CLBLM_R_X3Y149_SLICE_X3Y149_BQ;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_D2 = CLBLM_R_X7Y154_SLICE_X8Y154_CQ;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_D3 = CLBLM_L_X8Y151_SLICE_X11Y151_DQ;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_D4 = CLBLM_L_X8Y144_SLICE_X11Y144_CO6;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_D5 = CLBLM_R_X5Y149_SLICE_X7Y149_CQ;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_D6 = CLBLM_L_X8Y149_SLICE_X10Y149_BO6;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_D2 = 1'b1;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_C4 = CLBLL_L_X2Y155_SLICE_X1Y155_DO6;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_C5 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_D3 = 1'b1;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_C6 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_A1 = CLBLM_R_X11Y153_SLICE_X15Y153_DO6;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_A2 = CLBLM_R_X11Y154_SLICE_X15Y154_CO5;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_A4 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_A5 = CLBLM_R_X5Y143_SLICE_X7Y143_AQ;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_A6 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_B1 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_B2 = CLBLM_R_X11Y153_SLICE_X14Y153_DO6;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_B3 = CLBLM_R_X11Y154_SLICE_X15Y154_CO6;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_B4 = CLBLM_L_X12Y153_SLICE_X17Y153_AQ;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_B6 = CLBLL_L_X4Y144_SLICE_X4Y144_CO6;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_D4 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_A1 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_A2 = CLBLM_R_X7Y143_SLICE_X9Y143_BQ;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_A3 = CLBLM_R_X7Y143_SLICE_X9Y143_AQ;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_A5 = CLBLM_R_X7Y144_SLICE_X9Y144_AQ;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_A6 = CLBLM_R_X5Y143_SLICE_X7Y143_CO6;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_C1 = CLBLM_R_X13Y152_SLICE_X18Y152_AO6;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_C2 = CLBLM_R_X11Y153_SLICE_X14Y153_CO5;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_C3 = CLBLM_L_X12Y153_SLICE_X17Y153_AQ;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_B1 = CLBLM_R_X3Y149_SLICE_X3Y149_B5Q;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_B2 = CLBLM_R_X7Y143_SLICE_X9Y143_BQ;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_B3 = CLBLM_R_X5Y143_SLICE_X7Y143_CO6;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_B4 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_B6 = CLBLM_L_X8Y143_SLICE_X10Y143_BQ;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_D1 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_C2 = CLBLM_R_X7Y143_SLICE_X9Y143_CQ;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_C3 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_C4 = CLBLM_R_X5Y143_SLICE_X7Y143_CO6;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_C5 = CLBLM_R_X7Y143_SLICE_X9Y143_AQ;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_B3 = CLBLM_R_X11Y146_SLICE_X15Y146_AQ;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_C6 = CLBLM_R_X7Y143_SLICE_X8Y143_BQ;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_D5 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_A1 = CLBLM_L_X10Y153_SLICE_X13Y153_BQ;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_A2 = CLBLM_R_X11Y154_SLICE_X15Y154_BQ;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_A3 = CLBLM_R_X11Y154_SLICE_X14Y154_AQ;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_A4 = CLBLM_R_X11Y154_SLICE_X15Y154_AQ;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_D2 = CLBLM_R_X11Y147_SLICE_X15Y147_CQ;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_B5 = CLBLM_L_X10Y143_SLICE_X13Y143_AQ;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_D1 = CLBLM_L_X8Y143_SLICE_X11Y143_AQ;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_D2 = CLBLM_R_X5Y143_SLICE_X7Y143_AQ;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_D3 = CLBLM_R_X7Y143_SLICE_X9Y143_BQ;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_D4 = CLBLM_R_X7Y143_SLICE_X9Y143_AQ;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_B6 = CLBLM_L_X10Y141_SLICE_X12Y141_AO5;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_D5 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_D6 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_AX = CLBLM_R_X7Y155_SLICE_X8Y155_AQ;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_B1 = CLBLM_L_X10Y153_SLICE_X13Y153_BQ;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_B2 = CLBLM_L_X10Y153_SLICE_X13Y153_CQ;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_B3 = CLBLM_R_X11Y153_SLICE_X15Y153_CO5;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_D5 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_A1 = CLBLM_L_X8Y147_SLICE_X10Y147_DQ;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_A2 = CLBLM_R_X5Y148_SLICE_X7Y148_CQ;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_A3 = CLBLM_R_X7Y143_SLICE_X8Y143_AQ;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_D6 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_A5 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_D6 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_C1 = CLBLM_L_X12Y151_SLICE_X16Y151_DO5;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_B1 = CLBLL_L_X4Y148_SLICE_X4Y148_AQ;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_B2 = CLBLM_R_X7Y144_SLICE_X9Y144_BQ;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_B3 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_B4 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_B6 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_A1 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_A2 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_A3 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_A4 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_A5 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_A6 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_C1 = CLBLM_R_X5Y142_SLICE_X7Y142_AQ;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_B1 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_B2 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_B3 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_B4 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_B5 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_B6 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_C3 = CLBLM_R_X7Y145_SLICE_X8Y145_CQ;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_C4 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_C1 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_C2 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_C3 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_C4 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_C5 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_C6 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_D1 = CLBLM_R_X7Y142_SLICE_X8Y142_DO6;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_D2 = CLBLM_R_X7Y143_SLICE_X8Y143_CQ;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_D3 = CLBLM_L_X12Y144_SLICE_X16Y144_CQ;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_D4 = CLBLM_L_X8Y145_SLICE_X11Y145_BQ;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_D5 = CLBLM_R_X7Y146_SLICE_X9Y146_CQ;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_D6 = CLBLM_L_X10Y142_SLICE_X13Y142_BO6;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_D1 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_D2 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_D3 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_D4 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_D5 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X0Y142_D6 = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_T1 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_A1 = CLBLM_R_X3Y143_SLICE_X3Y143_A5Q;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_A2 = CLBLM_R_X3Y143_SLICE_X2Y143_CQ;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_A3 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_A4 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_A5 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_A6 = CLBLM_R_X3Y142_SLICE_X2Y142_BQ;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_A3 = CLBLL_L_X4Y144_SLICE_X5Y144_BQ;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_B1 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_B2 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_B3 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_B4 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_B5 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_B6 = 1'b1;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_A4 = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y155_D1 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_C1 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_C2 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_C3 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_C4 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_C5 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_C6 = 1'b1;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_A6 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_A1 = CLBLM_L_X12Y151_SLICE_X16Y151_CQ;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_D1 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_D2 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_D3 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_D4 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_D5 = 1'b1;
  assign CLBLL_L_X2Y142_SLICE_X1Y142_D6 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_A2 = CLBLM_L_X10Y147_SLICE_X12Y147_CQ;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_A3 = CLBLM_L_X8Y150_SLICE_X11Y150_AQ;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_A5 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_A6 = CLBLM_L_X8Y152_SLICE_X11Y152_BO6;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_B1 = CLBLM_R_X7Y148_SLICE_X8Y148_CQ;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_B6 = CLBLM_L_X8Y152_SLICE_X11Y152_BO6;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_B2 = CLBLM_L_X8Y150_SLICE_X11Y150_BQ;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_B3 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_B5 = CLBLM_L_X10Y149_SLICE_X13Y149_AQ;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_C1 = CLBLM_R_X7Y148_SLICE_X9Y148_CQ;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_C2 = CLBLM_L_X8Y152_SLICE_X10Y152_DQ;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_C3 = CLBLM_L_X8Y152_SLICE_X11Y152_BO5;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_C4 = CLBLM_L_X10Y150_SLICE_X12Y150_CQ;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_C5 = CLBLM_L_X8Y150_SLICE_X11Y150_DO6;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_C6 = CLBLM_R_X7Y149_SLICE_X8Y149_BQ;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_D1 = CLBLM_L_X8Y152_SLICE_X11Y152_AQ;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_D2 = CLBLM_L_X10Y147_SLICE_X12Y147_CQ;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_D3 = CLBLM_L_X10Y150_SLICE_X12Y150_DQ;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_D4 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_D5 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_D6 = CLBLM_R_X7Y150_SLICE_X8Y150_CQ;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_B5 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_A1 = CLBLM_L_X8Y149_SLICE_X10Y149_CO6;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_A3 = CLBLM_L_X8Y150_SLICE_X10Y150_AQ;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_A4 = CLBLM_L_X10Y153_SLICE_X13Y153_AQ;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_A5 = CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_A6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_C4 = CLBLM_R_X5Y153_SLICE_X6Y153_A5Q;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_C5 = CLBLM_L_X10Y154_SLICE_X12Y154_BQ;
  assign LIOI3_X0Y161_OLOGIC_X0Y162_D1 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_B1 = CLBLM_L_X8Y149_SLICE_X10Y149_CO6;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_B3 = CLBLM_L_X10Y145_SLICE_X12Y145_BQ;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_B4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_B5 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_B6 = CLBLM_R_X7Y151_SLICE_X9Y151_CQ;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_C6 = 1'b1;
  assign LIOI3_X0Y161_OLOGIC_X0Y162_T1 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_C1 = CLBLM_L_X8Y152_SLICE_X11Y152_AQ;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_C2 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_C3 = CLBLM_L_X8Y148_SLICE_X10Y148_BO5;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_C5 = CLBLM_R_X7Y144_SLICE_X8Y144_AQ;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOI3_X0Y101_OLOGIC_X0Y102_D1 = CLBLL_L_X2Y138_SLICE_X0Y138_BO5;
  assign LIOI3_X0Y161_OLOGIC_X0Y161_D1 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign LIOI3_X0Y101_OLOGIC_X0Y102_T1 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_A1 = CLBLM_R_X11Y154_SLICE_X15Y154_CO6;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_D1 = CLBLM_L_X8Y149_SLICE_X10Y149_AO5;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_D2 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_D3 = CLBLM_R_X7Y154_SLICE_X8Y154_CQ;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_D4 = CLBLM_R_X7Y149_SLICE_X8Y149_CQ;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_D5 = CLBLM_R_X7Y145_SLICE_X8Y145_BQ;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_D6 = CLBLM_R_X7Y143_SLICE_X8Y143_AQ;
  assign LIOI3_X0Y161_OLOGIC_X0Y161_T1 = 1'b1;
  assign LIOI3_X0Y101_OLOGIC_X0Y101_D1 = CLBLL_L_X2Y138_SLICE_X0Y138_BO6;
  assign LIOI3_X0Y101_OLOGIC_X0Y101_T1 = 1'b1;
  assign CLBLM_R_X11Y154_SLICE_X15Y154_A1 = CLBLM_R_X11Y154_SLICE_X15Y154_AQ;
  assign CLBLM_R_X11Y154_SLICE_X15Y154_A2 = CLBLM_R_X11Y153_SLICE_X15Y153_CO5;
  assign CLBLM_R_X11Y154_SLICE_X15Y154_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y154_SLICE_X15Y154_A4 = CLBLM_L_X12Y154_SLICE_X16Y154_BO6;
  assign CLBLM_R_X11Y154_SLICE_X15Y154_A5 = CLBLM_L_X10Y153_SLICE_X12Y153_AQ;
  assign CLBLM_R_X11Y154_SLICE_X15Y154_A6 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X11Y154_SLICE_X15Y154_B1 = CLBLM_R_X11Y154_SLICE_X15Y154_DO6;
  assign CLBLM_R_X11Y154_SLICE_X15Y154_B2 = CLBLM_R_X11Y154_SLICE_X15Y154_BQ;
  assign CLBLM_R_X11Y154_SLICE_X15Y154_B3 = CLBLM_R_X11Y151_SLICE_X15Y151_BQ;
  assign CLBLM_R_X11Y154_SLICE_X15Y154_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y154_SLICE_X15Y154_B5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X11Y154_SLICE_X15Y154_B6 = CLBLM_R_X11Y154_SLICE_X15Y154_CO6;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_A1 = CLBLM_R_X7Y144_SLICE_X9Y144_AQ;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_A3 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_A4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_A5 = CLBLM_R_X3Y150_SLICE_X3Y150_AQ;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_A6 = CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  assign CLBLM_R_X11Y154_SLICE_X15Y154_C3 = CLBLM_L_X10Y153_SLICE_X13Y153_BQ;
  assign CLBLM_R_X11Y154_SLICE_X15Y154_C4 = CLBLM_R_X11Y154_SLICE_X15Y154_BQ;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_AX = CLBLM_L_X8Y148_SLICE_X10Y148_BO6;
  assign CLBLM_R_X11Y154_SLICE_X15Y154_C5 = CLBLM_R_X11Y154_SLICE_X15Y154_AQ;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_B1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_B2 = CLBLM_R_X7Y144_SLICE_X9Y144_BQ;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_B3 = CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_B4 = CLBLM_L_X8Y150_SLICE_X10Y150_AQ;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_B5 = CLBLM_L_X10Y144_SLICE_X12Y144_AQ;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y154_SLICE_X15Y154_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X11Y154_SLICE_X15Y154_D1 = CLBLM_R_X11Y153_SLICE_X15Y153_CO5;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_C1 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_C2 = CLBLM_R_X7Y144_SLICE_X9Y144_CQ;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_C3 = CLBLM_R_X5Y144_SLICE_X7Y144_B5Q;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_C5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_C6 = 1'b1;
  assign CLBLM_R_X11Y154_SLICE_X15Y154_D3 = CLBLM_R_X11Y154_SLICE_X14Y154_BO5;
  assign CLBLM_R_X11Y154_SLICE_X15Y154_D4 = CLBLM_R_X11Y154_SLICE_X15Y154_BQ;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y154_SLICE_X14Y154_A1 = CLBLM_R_X5Y152_SLICE_X7Y152_B5Q;
  assign CLBLM_R_X11Y154_SLICE_X14Y154_A2 = CLBLM_R_X11Y153_SLICE_X15Y153_CO6;
  assign CLBLM_R_X11Y154_SLICE_X14Y154_A3 = CLBLM_R_X11Y154_SLICE_X14Y154_AQ;
  assign CLBLM_R_X11Y154_SLICE_X14Y154_A4 = CLBLM_R_X11Y154_SLICE_X15Y154_BQ;
  assign CLBLM_R_X11Y154_SLICE_X14Y154_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_D1 = CLBLL_L_X2Y146_SLICE_X1Y146_AQ;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_D2 = CLBLM_L_X8Y144_SLICE_X11Y144_BO6;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_D3 = CLBLL_L_X4Y143_SLICE_X4Y143_CO6;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_D4 = CLBLM_L_X10Y144_SLICE_X12Y144_DO6;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_D5 = CLBLM_R_X7Y142_SLICE_X8Y142_DO6;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_D6 = 1'b1;
  assign CLBLM_R_X11Y154_SLICE_X14Y154_A6 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X11Y154_SLICE_X14Y154_B1 = CLBLM_L_X10Y153_SLICE_X13Y153_BQ;
  assign CLBLM_R_X11Y154_SLICE_X14Y154_B2 = CLBLM_L_X10Y153_SLICE_X13Y153_CQ;
  assign CLBLM_R_X11Y154_SLICE_X14Y154_B3 = CLBLM_R_X11Y153_SLICE_X15Y153_CO6;
  assign CLBLM_R_X11Y154_SLICE_X14Y154_B4 = CLBLM_L_X10Y154_SLICE_X13Y154_AQ;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_A1 = CLBLM_R_X5Y144_SLICE_X7Y144_DO6;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_A2 = CLBLM_R_X3Y144_SLICE_X2Y144_BQ;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_A3 = CLBLM_R_X7Y144_SLICE_X8Y144_AQ;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_A5 = CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_A6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_C5 = CLBLM_R_X7Y155_SLICE_X8Y155_A5Q;
  assign CLBLM_R_X11Y154_SLICE_X14Y154_C1 = CLBLM_R_X11Y154_SLICE_X15Y154_AQ;
  assign CLBLM_R_X11Y154_SLICE_X14Y154_C2 = CLBLM_R_X11Y154_SLICE_X14Y154_AQ;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_B1 = CLBLM_R_X5Y144_SLICE_X7Y144_DO6;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_B2 = CLBLM_R_X7Y144_SLICE_X8Y144_BQ;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_B3 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_B5 = CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_B6 = CLBLL_L_X4Y148_SLICE_X4Y148_CQ;
  assign CLBLM_R_X11Y154_SLICE_X14Y154_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X11Y154_SLICE_X14Y154_D1 = CLBLM_R_X11Y154_SLICE_X14Y154_CO5;
  assign CLBLM_R_X11Y154_SLICE_X14Y154_D2 = CLBLM_R_X11Y154_SLICE_X15Y154_AQ;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_C1 = CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_C2 = CLBLM_R_X7Y144_SLICE_X8Y144_CQ;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_C3 = CLBLM_R_X3Y145_SLICE_X3Y145_A5Q;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_C5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_C6 = CLBLM_L_X10Y144_SLICE_X13Y144_BQ;
  assign CLBLM_R_X11Y154_SLICE_X14Y154_D3 = CLBLM_L_X10Y153_SLICE_X13Y153_CQ;
  assign CLBLM_R_X11Y154_SLICE_X14Y154_D4 = CLBLM_L_X10Y154_SLICE_X13Y154_DO6;
  assign CLBLM_R_X11Y154_SLICE_X14Y154_D5 = CLBLM_R_X11Y154_SLICE_X14Y154_AQ;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y154_SLICE_X14Y154_D6 = CLBLM_R_X11Y152_SLICE_X15Y152_BQ;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_D1 = CLBLM_R_X11Y144_SLICE_X15Y144_DO6;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_D2 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_D3 = CLBLM_R_X7Y144_SLICE_X8Y144_DQ;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_D4 = CLBLM_R_X7Y142_SLICE_X8Y142_DO6;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_D5 = CLBLM_R_X3Y145_SLICE_X2Y145_A5Q;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_D6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_B1 = CLBLL_L_X4Y154_SLICE_X4Y154_CO6;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_B2 = CLBLM_R_X3Y153_SLICE_X2Y153_DO6;
  assign RIOI3_X105Y145_ILOGIC_X1Y146_D = RIOB33_X105Y145_IOB_X1Y146_I;
  assign RIOI3_X105Y145_ILOGIC_X1Y145_D = RIOB33_X105Y145_IOB_X1Y145_I;
  assign LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y64_D = LIOB33_X0Y63_IOB_X0Y64_I;
  assign LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y63_D = LIOB33_X0Y63_IOB_X0Y63_I;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_A1 = 1'b1;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_A2 = CLBLM_R_X5Y145_SLICE_X6Y145_CQ;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_A3 = CLBLM_L_X10Y150_SLICE_X12Y150_DQ;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_A4 = CLBLM_L_X8Y151_SLICE_X11Y151_AQ;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_A6 = CLBLM_L_X8Y152_SLICE_X11Y152_BO6;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_C6 = CLBLM_R_X5Y152_SLICE_X7Y152_DO5;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_B1 = CLBLM_R_X5Y152_SLICE_X7Y152_BQ;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_B2 = CLBLM_L_X8Y151_SLICE_X11Y151_BQ;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_B4 = CLBLM_R_X11Y151_SLICE_X14Y151_CO6;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_B6 = CLBLM_R_X7Y153_SLICE_X9Y153_A5Q;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_C4 = CLBLM_R_X5Y152_SLICE_X7Y152_B5Q;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_C1 = CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_C2 = CLBLM_L_X8Y151_SLICE_X11Y151_CQ;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_C3 = CLBLM_L_X10Y151_SLICE_X13Y151_DQ;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_C4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_C5 = CLBLM_L_X8Y148_SLICE_X11Y148_AQ;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_C5 = CLBLL_L_X4Y144_SLICE_X5Y144_DO6;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_C6 = CLBLM_R_X5Y143_SLICE_X7Y143_BO6;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_D1 = 1'b1;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_D2 = CLBLM_L_X12Y152_SLICE_X16Y152_AQ;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_D3 = CLBLM_L_X8Y151_SLICE_X11Y151_DQ;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_D4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_D5 = 1'b1;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_D6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_A1 = CLBLM_L_X8Y151_SLICE_X10Y151_B5Q;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_A2 = CLBLM_L_X10Y151_SLICE_X12Y151_CQ;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_A3 = CLBLM_L_X8Y151_SLICE_X10Y151_AQ;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_A5 = CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_A6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X103Y176_SLICE_X162Y176_D2 = 1'b1;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_B2 = CLBLM_L_X10Y150_SLICE_X12Y150_AQ;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_B4 = CLBLL_L_X4Y148_SLICE_X5Y148_CQ;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_B5 = CLBLM_L_X8Y151_SLICE_X10Y151_BQ;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_B6 = 1'b1;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_C1 = CLBLM_R_X11Y150_SLICE_X14Y150_BO6;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_C2 = CLBLM_L_X8Y151_SLICE_X10Y151_CQ;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_C4 = CLBLM_L_X8Y148_SLICE_X10Y148_A5Q;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_C5 = CLBLM_R_X11Y147_SLICE_X14Y147_BQ;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_C6 = CLBLM_R_X7Y152_SLICE_X9Y152_BQ;
  assign LIOI3_X0Y179_OLOGIC_X0Y180_T1 = 1'b1;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_D1 = CLBLM_L_X10Y144_SLICE_X13Y144_CQ;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_D2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_D3 = CLBLM_L_X8Y151_SLICE_X10Y151_DQ;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_D4 = CLBLM_R_X11Y150_SLICE_X14Y150_BO6;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_D5 = CLBLM_R_X5Y145_SLICE_X7Y145_AQ;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_D6 = CLBLM_L_X8Y148_SLICE_X10Y148_A5Q;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_A1 = CLBLM_R_X7Y148_SLICE_X9Y148_CQ;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_A2 = CLBLM_L_X8Y152_SLICE_X11Y152_BO6;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_A3 = CLBLM_R_X7Y145_SLICE_X9Y145_AQ;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_A5 = 1'b1;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_A6 = CLBLM_L_X8Y145_SLICE_X11Y145_BQ;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_B1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_B2 = CLBLM_R_X7Y145_SLICE_X9Y145_BQ;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_B3 = CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_B4 = CLBLM_R_X7Y144_SLICE_X9Y144_BQ;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_B6 = CLBLM_R_X3Y144_SLICE_X2Y144_AQ;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_C2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_C3 = CLBLM_R_X7Y147_SLICE_X8Y147_DQ;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_C4 = CLBLM_L_X12Y149_SLICE_X16Y149_AQ;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_C5 = CLBLM_L_X8Y145_SLICE_X10Y145_A5Q;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_C6 = 1'b1;
  assign LIOB33_X0Y163_IOB_X0Y163_O = RIOB33_X105Y109_IOB_X1Y110_I;
  assign LIOB33_X0Y163_IOB_X0Y164_O = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_D1 = CLBLM_R_X7Y153_SLICE_X9Y153_CO5;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_D2 = CLBLL_L_X2Y151_SLICE_X1Y151_BO6;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_D3 = CLBLL_L_X4Y154_SLICE_X4Y154_CO6;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_D4 = 1'b1;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_D5 = CLBLM_R_X5Y149_SLICE_X6Y149_CO6;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_D6 = CLBLM_R_X5Y145_SLICE_X6Y145_DO6;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_A1 = CLBLM_R_X5Y145_SLICE_X7Y145_DO6;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_A2 = CLBLM_L_X12Y145_SLICE_X16Y145_BQ;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_A3 = CLBLM_R_X7Y145_SLICE_X8Y145_AQ;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_A4 = CLBLM_R_X11Y146_SLICE_X14Y146_AQ;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_A5 = 1'b1;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_B1 = CLBLM_R_X7Y145_SLICE_X8Y145_BQ;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_B2 = CLBLM_R_X5Y148_SLICE_X7Y148_CQ;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_B4 = CLBLM_R_X7Y147_SLICE_X8Y147_BQ;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_C1 = CLBLM_L_X10Y154_SLICE_X13Y154_CO5;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_B5 = 1'b1;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_C1 = CLBLM_R_X3Y145_SLICE_X2Y145_A5Q;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_C2 = CLBLM_R_X5Y147_SLICE_X6Y147_CQ;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_C3 = CLBLM_R_X7Y148_SLICE_X9Y148_CQ;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_C6 = 1'b1;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_D1 = CLBLM_R_X7Y143_SLICE_X8Y143_AQ;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_D2 = CLBLM_R_X11Y148_SLICE_X14Y148_CQ;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_D3 = CLBLL_L_X4Y143_SLICE_X4Y143_BQ;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_D4 = CLBLM_R_X5Y145_SLICE_X6Y145_CQ;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_D5 = CLBLM_R_X7Y145_SLICE_X8Y145_BQ;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_D6 = CLBLL_L_X4Y145_SLICE_X4Y145_BQ;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_C5 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_A1 = CLBLM_L_X8Y153_SLICE_X10Y153_BQ;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_A3 = 1'b1;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_A4 = CLBLM_R_X7Y149_SLICE_X8Y149_BQ;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_A5 = CLBLM_L_X10Y149_SLICE_X13Y149_CO5;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_A6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_B1 = 1'b1;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_B2 = CLBLM_R_X11Y147_SLICE_X15Y147_CQ;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_B3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_B4 = CLBLM_R_X11Y146_SLICE_X14Y146_DQ;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_B6 = 1'b1;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_C1 = 1'b1;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_C2 = 1'b1;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_C3 = 1'b1;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_C4 = 1'b1;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_C5 = 1'b1;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_C6 = 1'b1;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_D1 = 1'b1;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_D2 = 1'b1;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_D3 = 1'b1;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_D4 = 1'b1;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_D5 = 1'b1;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_D6 = 1'b1;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_A1 = CLBLM_L_X10Y153_SLICE_X13Y153_DQ;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_A2 = CLBLM_L_X8Y152_SLICE_X11Y152_BO6;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_A3 = CLBLM_L_X8Y152_SLICE_X10Y152_AQ;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_A5 = 1'b1;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_A6 = CLBLM_L_X8Y152_SLICE_X10Y152_DQ;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_A4 = CLBLM_R_X7Y152_SLICE_X9Y152_CQ;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_A5 = CLBLM_L_X12Y151_SLICE_X17Y151_AO6;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_B1 = 1'b1;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_B2 = CLBLM_L_X8Y152_SLICE_X10Y152_BQ;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_B3 = CLBLM_L_X12Y149_SLICE_X17Y149_BQ;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_B5 = CLBLM_L_X8Y152_SLICE_X11Y152_BO6;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_B6 = CLBLM_L_X10Y150_SLICE_X12Y150_CQ;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_A6 = CLBLM_R_X11Y154_SLICE_X15Y154_CO5;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_C1 = CLBLM_L_X8Y154_SLICE_X10Y154_AQ;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_C2 = CLBLM_L_X8Y152_SLICE_X10Y152_CQ;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_C3 = CLBLM_L_X8Y150_SLICE_X10Y150_DO6;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_C4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_C5 = CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_D2 = CLBLM_L_X10Y152_SLICE_X12Y152_CO5;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_D3 = CLBLM_R_X7Y152_SLICE_X9Y152_AQ;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_D4 = CLBLM_L_X8Y150_SLICE_X10Y150_CQ;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_D5 = 1'b1;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_D6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_B1 = CLBLM_L_X12Y152_SLICE_X16Y152_DO6;
  assign LIOB33_X0Y165_IOB_X0Y166_O = RIOB33_X105Y113_IOB_X1Y113_I;
  assign LIOB33_X0Y165_IOB_X0Y165_O = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_C1 = CLBLM_L_X12Y153_SLICE_X16Y153_DO6;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_A1 = CLBLM_R_X5Y148_SLICE_X6Y148_AQ;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_A2 = CLBLM_R_X7Y143_SLICE_X9Y143_AQ;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_A3 = CLBLM_L_X8Y148_SLICE_X10Y148_CO5;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_A6 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_B1 = CLBLL_L_X4Y146_SLICE_X4Y146_BQ;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_B2 = CLBLM_R_X7Y146_SLICE_X9Y146_BQ;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_B3 = CLBLM_R_X7Y147_SLICE_X9Y147_AQ;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_B4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_B5 = CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_C1 = CLBLM_R_X5Y148_SLICE_X7Y148_AQ;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_C2 = CLBLM_R_X7Y146_SLICE_X9Y146_CQ;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_C3 = CLBLM_L_X10Y148_SLICE_X12Y148_BQ;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_C4 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_C5 = CLBLL_L_X4Y145_SLICE_X5Y145_DO6;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOI3_X0Y165_OLOGIC_X0Y166_D1 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y165_OLOGIC_X0Y166_T1 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_D1 = CLBLM_R_X7Y145_SLICE_X9Y145_C5Q;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_D2 = CLBLM_R_X7Y152_SLICE_X9Y152_CQ;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_D3 = CLBLM_R_X7Y147_SLICE_X8Y147_DQ;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_D4 = CLBLM_R_X7Y149_SLICE_X8Y149_CQ;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_D5 = CLBLM_R_X7Y146_SLICE_X8Y146_DQ;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_D6 = CLBLL_L_X4Y146_SLICE_X5Y146_A5Q;
  assign LIOI3_X0Y103_OLOGIC_X0Y104_D1 = CLBLL_L_X2Y141_SLICE_X0Y141_AO5;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_D1 = LIOB33_X0Y59_IOB_X0Y59_I;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign LIOI3_X0Y165_OLOGIC_X0Y165_D1 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_A1 = RIOB33_X105Y119_IOB_X1Y119_I;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_A1 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_A2 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_A3 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_A4 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_A5 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_A6 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_A3 = CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_A4 = CLBLM_R_X7Y146_SLICE_X8Y146_CQ;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_A5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_B1 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_B2 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_B3 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_B4 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_B5 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_B6 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_B1 = CLBLM_R_X11Y146_SLICE_X15Y146_DQ;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_C1 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_C2 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_C3 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_C4 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_C5 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_C6 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_C1 = CLBLM_R_X7Y146_SLICE_X8Y146_C5Q;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_C2 = RIOB33_X105Y119_IOB_X1Y119_I;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_C3 = CLBLM_L_X10Y146_SLICE_X13Y146_B5Q;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_C5 = CLBLM_R_X5Y146_SLICE_X6Y146_DQ;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_C6 = 1'b1;
  assign CLBLM_L_X10Y154_SLICE_X12Y154_A5 = CLBLM_L_X8Y147_SLICE_X10Y147_AQ;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_D1 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_D2 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_D3 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_D4 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_D5 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_D6 = 1'b1;
  assign CLBLM_L_X10Y154_SLICE_X12Y154_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_D1 = CLBLM_L_X8Y145_SLICE_X11Y145_AQ;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_D4 = CLBLM_L_X12Y152_SLICE_X16Y152_BQ;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_D2 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_D3 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_D4 = CLBLM_R_X7Y152_SLICE_X9Y152_CQ;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_D5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_D6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_A2 = CLBLM_R_X5Y152_SLICE_X6Y152_BQ;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_A3 = CLBLL_L_X2Y145_SLICE_X1Y145_AQ;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_A4 = CLBLM_R_X3Y145_SLICE_X3Y145_D5Q;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_A5 = CLBLL_L_X2Y142_SLICE_X1Y142_AO6;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_A6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y154_SLICE_X12Y154_B3 = CLBLM_L_X10Y154_SLICE_X12Y154_AQ;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_B2 = CLBLL_L_X2Y145_SLICE_X1Y145_BQ;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_B3 = CLBLM_R_X3Y144_SLICE_X2Y144_CO6;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_B4 = CLBLM_R_X5Y146_SLICE_X6Y146_CQ;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_B5 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_B6 = CLBLL_L_X4Y145_SLICE_X4Y145_A5Q;
  assign CLBLM_R_X103Y176_SLICE_X163Y176_D3 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X163Y176_D4 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_C1 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_C2 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_C3 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_C4 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_C5 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_C6 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X163Y176_D5 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X103Y176_SLICE_X163Y176_D6 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_D1 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_D2 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_D3 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_D4 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_D5 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_D6 = 1'b1;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_A1 = CLBLM_R_X3Y147_SLICE_X2Y147_AQ;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_A3 = 1'b1;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_A4 = CLBLM_L_X8Y154_SLICE_X11Y154_BO6;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_A5 = CLBLM_L_X8Y153_SLICE_X10Y153_DO6;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_A6 = CLBLM_L_X8Y153_SLICE_X10Y153_CO5;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_B1 = CLBLM_L_X8Y154_SLICE_X10Y154_DO6;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_B3 = CLBLM_L_X8Y153_SLICE_X10Y153_CO5;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_B4 = CLBLM_L_X8Y153_SLICE_X10Y153_DO6;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_B5 = CLBLM_R_X5Y145_SLICE_X7Y145_AQ;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_B6 = 1'b1;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_C1 = CLBLM_L_X8Y153_SLICE_X10Y153_DO6;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_C2 = CLBLM_L_X8Y153_SLICE_X11Y153_CQ;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_C3 = CLBLM_L_X8Y154_SLICE_X11Y154_CO6;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_C4 = CLBLM_R_X7Y154_SLICE_X8Y154_CQ;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_C5 = CLBLM_L_X8Y153_SLICE_X10Y153_CO5;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_D1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_D2 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_D3 = CLBLM_R_X7Y153_SLICE_X9Y153_AQ;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_D4 = CLBLM_L_X8Y153_SLICE_X11Y153_DQ;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_D5 = CLBLM_R_X11Y146_SLICE_X14Y146_DQ;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_D6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_A2 = CLBLM_L_X8Y153_SLICE_X10Y153_BQ;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_A3 = CLBLM_L_X8Y153_SLICE_X10Y153_AQ;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_A4 = CLBLM_R_X5Y155_SLICE_X7Y155_CO6;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_A5 = CLBLM_R_X7Y155_SLICE_X8Y155_BO5;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_A6 = CLBLM_L_X10Y146_SLICE_X13Y146_BQ;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_B1 = CLBLM_R_X5Y153_SLICE_X7Y153_BQ;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_B2 = CLBLM_L_X8Y153_SLICE_X10Y153_BQ;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_B3 = CLBLM_L_X10Y153_SLICE_X13Y153_AQ;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_B4 = CLBLM_R_X5Y155_SLICE_X7Y155_CO6;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_B5 = CLBLM_R_X7Y155_SLICE_X8Y155_BO5;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_C1 = CLBLM_L_X8Y153_SLICE_X11Y153_AQ;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_C2 = CLBLM_L_X8Y154_SLICE_X10Y154_BO5;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_C3 = CLBLM_L_X10Y156_SLICE_X12Y156_CO6;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_C5 = CLBLM_L_X10Y150_SLICE_X12Y150_B5Q;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_C6 = 1'b1;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_D1 = CLBLM_R_X7Y155_SLICE_X8Y155_A5Q;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_D2 = CLBLL_L_X4Y147_SLICE_X5Y147_B5Q;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_D3 = CLBLM_R_X7Y153_SLICE_X8Y153_CQ;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_D4 = CLBLM_L_X10Y156_SLICE_X12Y156_CO6;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_D5 = CLBLM_R_X7Y154_SLICE_X8Y154_BQ;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_D6 = 1'b1;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_C4 = CLBLM_R_X11Y150_SLICE_X15Y150_BQ;
  assign RIOI3_X105Y147_ILOGIC_X1Y148_D = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_C5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X103Y176_SLICE_X162Y176_B5 = 1'b1;
  assign RIOI3_X105Y147_ILOGIC_X1Y147_D = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X103Y176_SLICE_X162Y176_B6 = 1'b1;
  assign LIOB33_X0Y167_IOB_X0Y168_O = RIOB33_X105Y123_IOB_X1Y123_I;
  assign LIOB33_X0Y167_IOB_X0Y167_O = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLM_R_X11Y157_SLICE_X15Y157_A1 = 1'b1;
  assign CLBLM_R_X11Y157_SLICE_X15Y157_A2 = 1'b1;
  assign CLBLM_R_X11Y157_SLICE_X15Y157_A3 = 1'b1;
  assign CLBLM_R_X11Y157_SLICE_X15Y157_A4 = 1'b1;
  assign CLBLM_R_X11Y157_SLICE_X15Y157_A5 = 1'b1;
  assign CLBLM_R_X11Y157_SLICE_X15Y157_A6 = 1'b1;
  assign CLBLM_R_X11Y157_SLICE_X15Y157_B1 = 1'b1;
  assign CLBLM_R_X11Y157_SLICE_X15Y157_B2 = 1'b1;
  assign CLBLM_R_X11Y157_SLICE_X15Y157_B3 = 1'b1;
  assign CLBLM_R_X11Y157_SLICE_X15Y157_B4 = 1'b1;
  assign CLBLM_R_X11Y157_SLICE_X15Y157_B5 = 1'b1;
  assign CLBLM_R_X11Y157_SLICE_X15Y157_B6 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X162Y176_C3 = 1'b1;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_A1 = 1'b1;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_A3 = CLBLM_L_X8Y146_SLICE_X10Y146_AQ;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_A4 = CLBLM_R_X7Y147_SLICE_X8Y147_BQ;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_A5 = CLBLM_R_X11Y153_SLICE_X14Y153_AO6;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_A6 = 1'b1;
  assign CLBLM_R_X11Y157_SLICE_X15Y157_C1 = 1'b1;
  assign CLBLM_R_X11Y157_SLICE_X15Y157_C2 = 1'b1;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_D2 = CLBLM_L_X10Y150_SLICE_X13Y150_BQ;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_B1 = 1'b1;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_B3 = CLBLM_L_X10Y151_SLICE_X12Y151_AQ;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_B4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_B5 = CLBLM_R_X7Y145_SLICE_X9Y145_C5Q;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_B6 = 1'b1;
  assign CLBLM_R_X11Y157_SLICE_X15Y157_D1 = 1'b1;
  assign CLBLM_R_X11Y157_SLICE_X15Y157_D2 = 1'b1;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_C1 = CLBLM_R_X7Y145_SLICE_X9Y145_C5Q;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_C2 = CLBLL_L_X4Y147_SLICE_X4Y147_AQ;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_C3 = CLBLM_R_X7Y149_SLICE_X8Y149_CQ;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_C4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_C5 = CLBLM_L_X8Y150_SLICE_X10Y150_AQ;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_C6 = 1'b1;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_D5 = 1'b1;
  assign CLBLM_R_X11Y157_SLICE_X15Y157_D4 = 1'b1;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_D6 = CLBLM_R_X11Y149_SLICE_X15Y149_AO6;
  assign CLBLM_R_X11Y157_SLICE_X14Y157_A1 = 1'b1;
  assign CLBLM_R_X11Y157_SLICE_X14Y157_A2 = CLBLM_R_X5Y145_SLICE_X6Y145_DO5;
  assign CLBLM_R_X11Y157_SLICE_X14Y157_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y157_SLICE_X14Y157_A4 = CLBLM_R_X11Y153_SLICE_X14Y153_CQ;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_D1 = CLBLM_R_X5Y148_SLICE_X7Y148_C5Q;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_D2 = CLBLM_L_X10Y146_SLICE_X13Y146_B5Q;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_D3 = CLBLM_R_X7Y147_SLICE_X9Y147_BQ;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_D4 = CLBLM_R_X5Y148_SLICE_X7Y148_BQ;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_D5 = CLBLM_L_X10Y146_SLICE_X13Y146_DO6;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_D6 = 1'b1;
  assign CLBLM_R_X11Y157_SLICE_X14Y157_A5 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_R_X11Y157_SLICE_X14Y157_A6 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_A1 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_A2 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_A3 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_A4 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_A5 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_A6 = 1'b1;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_A1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_A2 = CLBLM_L_X8Y150_SLICE_X10Y150_CQ;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_A3 = CLBLM_R_X7Y147_SLICE_X8Y147_AQ;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_B1 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_B2 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_B3 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_B4 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_B5 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_B6 = 1'b1;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_A5 = CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_A6 = CLBLM_R_X11Y146_SLICE_X14Y146_AQ;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_C1 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_C2 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_C3 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_C4 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_C5 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_C6 = 1'b1;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_B5 = CLBLM_R_X5Y147_SLICE_X7Y147_DQ;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_B6 = 1'b1;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_C2 = CLBLM_R_X7Y147_SLICE_X9Y147_BQ;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_C4 = CLBLM_R_X7Y153_SLICE_X8Y153_CQ;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_D1 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_D2 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_D3 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_D4 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_D5 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_D6 = 1'b1;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_D1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_D2 = CLBLM_R_X5Y152_SLICE_X7Y152_CQ;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_D3 = 1'b1;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_D4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_D5 = 1'b1;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_D6 = CLBLM_L_X10Y146_SLICE_X13Y146_B5Q;
  assign CLBLM_R_X103Y176_SLICE_X162Y176_D5 = 1'b1;
  assign RIOI3_X105Y123_ILOGIC_X1Y123_D = RIOB33_X105Y123_IOB_X1Y123_I;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_C1 = CLBLM_R_X7Y150_SLICE_X9Y150_AQ;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_C2 = CLBLM_L_X10Y150_SLICE_X12Y150_BQ;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_A1 = CLBLL_L_X4Y144_SLICE_X4Y144_DO6;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_A2 = CLBLL_L_X2Y146_SLICE_X1Y146_BQ;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_A3 = CLBLL_L_X2Y146_SLICE_X1Y146_AQ;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_A4 = CLBLM_R_X3Y144_SLICE_X3Y144_BO6;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_A5 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_C4 = 1'b1;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_C5 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_B1 = CLBLL_L_X4Y146_SLICE_X4Y146_BQ;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_B2 = CLBLL_L_X2Y146_SLICE_X1Y146_BQ;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_B3 = CLBLM_R_X3Y144_SLICE_X2Y144_DO6;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_B4 = CLBLL_L_X2Y147_SLICE_X1Y147_BO6;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_B5 = CLBLM_R_X3Y144_SLICE_X3Y144_BO6;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_C6 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_C1 = CLBLM_R_X3Y144_SLICE_X3Y144_BO6;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_C2 = CLBLL_L_X2Y146_SLICE_X1Y146_CQ;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_C3 = CLBLL_L_X4Y144_SLICE_X4Y144_DO6;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_C4 = CLBLL_L_X4Y146_SLICE_X5Y146_CQ;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_C5 = CLBLL_L_X2Y146_SLICE_X1Y146_AQ;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_D1 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_D2 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_D3 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_D4 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_D5 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_D6 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_C6 = 1'b1;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_A1 = CLBLM_R_X7Y155_SLICE_X8Y155_AQ;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_A2 = CLBLM_R_X7Y153_SLICE_X8Y153_CQ;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_A3 = CLBLL_L_X4Y147_SLICE_X5Y147_B5Q;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_A4 = CLBLM_R_X7Y155_SLICE_X8Y155_A5Q;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_A5 = CLBLM_R_X7Y154_SLICE_X8Y154_BQ;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_A6 = 1'b1;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_D1 = CLBLM_L_X8Y150_SLICE_X10Y150_BQ;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_B1 = CLBLM_L_X8Y154_SLICE_X11Y154_DO6;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_B2 = CLBLM_R_X7Y153_SLICE_X8Y153_BQ;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_B3 = CLBLM_L_X8Y153_SLICE_X11Y153_AQ;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_B4 = CLBLM_L_X8Y155_SLICE_X10Y155_BQ;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_B5 = CLBLM_L_X8Y154_SLICE_X11Y154_AO6;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_B6 = CLBLM_L_X8Y155_SLICE_X10Y155_CO6;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_D2 = CLBLM_R_X5Y152_SLICE_X6Y152_CQ;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_D3 = CLBLM_L_X8Y154_SLICE_X10Y154_AQ;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_C1 = CLBLM_L_X8Y154_SLICE_X11Y154_AO6;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_C2 = CLBLM_R_X7Y154_SLICE_X8Y154_AQ;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_C3 = CLBLM_L_X8Y155_SLICE_X10Y155_CO6;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_C4 = CLBLM_L_X8Y153_SLICE_X11Y153_AQ;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_C5 = CLBLM_L_X8Y154_SLICE_X11Y154_DO6;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_C6 = CLBLM_L_X8Y155_SLICE_X10Y155_BQ;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_D4 = CLBLM_R_X7Y154_SLICE_X9Y154_AQ;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_D5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_D6 = CLBLM_R_X7Y151_SLICE_X8Y151_DO5;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_D1 = CLBLM_R_X7Y153_SLICE_X8Y153_CQ;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_D2 = CLBLL_L_X4Y147_SLICE_X5Y147_B5Q;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_D3 = CLBLM_R_X5Y155_SLICE_X7Y155_BO5;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_D4 = CLBLM_L_X8Y154_SLICE_X11Y154_AO5;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_D5 = CLBLM_R_X7Y153_SLICE_X9Y153_AQ;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_D6 = 1'b1;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_A1 = CLBLM_L_X10Y154_SLICE_X12Y154_CQ;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_A2 = 1'b1;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_A3 = CLBLM_R_X5Y150_SLICE_X7Y150_BQ;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_A5 = 1'b1;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_A6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_B1 = CLBLM_R_X7Y155_SLICE_X8Y155_AQ;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_B2 = CLBLM_R_X7Y153_SLICE_X8Y153_CQ;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_B3 = CLBLM_R_X7Y155_SLICE_X8Y155_A5Q;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_B4 = CLBLL_L_X4Y147_SLICE_X5Y147_B5Q;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_B5 = CLBLM_R_X7Y154_SLICE_X8Y154_BQ;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_B6 = 1'b1;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_C1 = CLBLM_L_X8Y153_SLICE_X11Y153_AQ;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_C2 = CLBLM_L_X8Y153_SLICE_X11Y153_CQ;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_C3 = CLBLM_R_X7Y154_SLICE_X8Y154_BQ;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_C4 = CLBLL_L_X4Y147_SLICE_X5Y147_B5Q;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_C5 = CLBLM_R_X7Y153_SLICE_X8Y153_CQ;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_C6 = CLBLM_L_X8Y155_SLICE_X10Y155_BQ;
  assign LIOB33_X0Y169_IOB_X0Y170_O = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X103Y141_SLICE_X163Y141_A1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X103Y141_SLICE_X163Y141_A2 = RIOB33_X105Y139_IOB_X1Y140_I;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X103Y141_SLICE_X163Y141_A3 = RIOB33_X105Y139_IOB_X1Y139_I;
  assign CLBLM_R_X103Y141_SLICE_X163Y141_A4 = RIOB33_X105Y137_IOB_X1Y138_I;
  assign CLBLM_R_X103Y141_SLICE_X163Y141_A5 = RIOB33_X105Y141_IOB_X1Y141_I;
  assign CLBLM_R_X103Y141_SLICE_X163Y141_A6 = 1'b1;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_A3 = CLBLM_R_X7Y152_SLICE_X8Y152_AQ;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_D1 = CLBLM_L_X8Y153_SLICE_X11Y153_BQ;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_D2 = CLBLM_L_X10Y154_SLICE_X12Y154_CQ;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_D3 = CLBLM_L_X8Y154_SLICE_X11Y154_DO6;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_D4 = CLBLM_L_X8Y154_SLICE_X10Y154_CO6;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_D5 = CLBLM_L_X8Y155_SLICE_X10Y155_CO6;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_D6 = 1'b1;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_A4 = CLBLM_R_X5Y151_SLICE_X6Y151_AQ;
  assign CLBLM_R_X103Y141_SLICE_X163Y141_B1 = 1'b1;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X103Y141_SLICE_X163Y141_B2 = 1'b1;
  assign CLBLM_R_X103Y141_SLICE_X163Y141_B3 = 1'b1;
  assign CLBLM_R_X103Y141_SLICE_X163Y141_B4 = 1'b1;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_A6 = CLBLM_R_X7Y149_SLICE_X8Y149_BQ;
  assign CLBLM_R_X103Y141_SLICE_X163Y141_B6 = 1'b1;
  assign CLBLM_R_X103Y141_SLICE_X163Y141_C1 = 1'b1;
  assign CLBLM_R_X103Y141_SLICE_X163Y141_C2 = 1'b1;
  assign CLBLM_R_X103Y141_SLICE_X163Y141_C3 = 1'b1;
  assign CLBLM_R_X103Y141_SLICE_X163Y141_C4 = 1'b1;
  assign CLBLM_R_X103Y141_SLICE_X163Y141_C5 = 1'b1;
  assign CLBLM_R_X103Y141_SLICE_X163Y141_C6 = 1'b1;
  assign CLBLM_R_X103Y141_SLICE_X163Y141_D1 = 1'b1;
  assign CLBLM_R_X103Y141_SLICE_X163Y141_D2 = 1'b1;
  assign CLBLM_R_X103Y141_SLICE_X163Y141_D3 = 1'b1;
  assign CLBLM_R_X103Y141_SLICE_X163Y141_D4 = 1'b1;
  assign CLBLM_R_X103Y141_SLICE_X163Y141_D5 = 1'b1;
  assign CLBLM_R_X103Y141_SLICE_X163Y141_D6 = 1'b1;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_B6 = CLBLM_L_X8Y146_SLICE_X10Y146_DO6;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_C4 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X103Y141_SLICE_X162Y141_A1 = 1'b1;
  assign CLBLM_R_X103Y141_SLICE_X162Y141_A2 = 1'b1;
  assign CLBLM_R_X103Y141_SLICE_X162Y141_A3 = 1'b1;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_C5 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_B1 = CLBLM_L_X8Y154_SLICE_X10Y154_AQ;
  assign CLBLM_R_X103Y141_SLICE_X162Y141_A4 = 1'b1;
  assign CLBLM_R_X103Y141_SLICE_X162Y141_A5 = 1'b1;
  assign CLBLM_R_X103Y141_SLICE_X162Y141_A6 = 1'b1;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_C6 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_B2 = CLBLM_L_X10Y151_SLICE_X13Y151_DQ;
  assign CLBLM_R_X103Y141_SLICE_X162Y141_B1 = 1'b1;
  assign CLBLM_R_X103Y141_SLICE_X162Y141_B2 = 1'b1;
  assign CLBLM_R_X103Y141_SLICE_X162Y141_B3 = 1'b1;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X103Y141_SLICE_X162Y141_B4 = 1'b1;
  assign CLBLL_L_X36Y146_SLICE_X54Y146_A1 = CLBLM_R_X7Y146_SLICE_X8Y146_CQ;
  assign CLBLL_L_X36Y146_SLICE_X54Y146_A2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X36Y146_SLICE_X54Y146_A3 = 1'b1;
  assign CLBLL_L_X36Y146_SLICE_X54Y146_A4 = 1'b1;
  assign CLBLL_L_X36Y146_SLICE_X54Y146_A5 = RIOB33_X105Y119_IOB_X1Y119_I;
  assign CLBLL_L_X36Y146_SLICE_X54Y146_A6 = 1'b1;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_A2 = 1'b1;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_A3 = CLBLM_R_X7Y148_SLICE_X9Y148_AQ;
  assign CLBLL_L_X36Y146_SLICE_X54Y146_B1 = 1'b1;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_B4 = CLBLM_R_X5Y152_SLICE_X7Y152_AQ;
  assign CLBLL_L_X36Y146_SLICE_X54Y146_B2 = 1'b1;
  assign CLBLL_L_X36Y146_SLICE_X54Y146_B3 = 1'b1;
  assign CLBLL_L_X36Y146_SLICE_X54Y146_B4 = 1'b1;
  assign CLBLL_L_X36Y146_SLICE_X54Y146_B5 = 1'b1;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_B5 = CLBLL_L_X4Y154_SLICE_X5Y154_CO5;
  assign CLBLL_L_X36Y146_SLICE_X54Y146_B6 = 1'b1;
  assign CLBLL_L_X36Y146_SLICE_X54Y146_C1 = 1'b1;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_B6 = CLBLM_R_X5Y150_SLICE_X6Y150_BQ;
  assign CLBLL_L_X36Y146_SLICE_X54Y146_C2 = 1'b1;
  assign CLBLL_L_X36Y146_SLICE_X54Y146_C3 = 1'b1;
  assign CLBLL_L_X36Y146_SLICE_X54Y146_C4 = 1'b1;
  assign CLBLL_L_X36Y146_SLICE_X54Y146_C5 = 1'b1;
  assign CLBLL_L_X36Y146_SLICE_X54Y146_C6 = 1'b1;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_C3 = CLBLM_R_X7Y148_SLICE_X9Y148_BQ;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_C4 = CLBLM_R_X5Y146_SLICE_X6Y146_CQ;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_C5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_C6 = 1'b1;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_C2 = CLBLM_L_X10Y148_SLICE_X12Y148_AO5;
  assign CLBLL_L_X36Y146_SLICE_X54Y146_D1 = 1'b1;
  assign CLBLL_L_X36Y146_SLICE_X54Y146_D2 = 1'b1;
  assign CLBLL_L_X36Y146_SLICE_X54Y146_D3 = 1'b1;
  assign CLBLL_L_X36Y146_SLICE_X54Y146_D4 = 1'b1;
  assign CLBLL_L_X36Y146_SLICE_X54Y146_D5 = 1'b1;
  assign CLBLL_L_X36Y146_SLICE_X54Y146_D6 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_A1 = CLBLM_R_X3Y147_SLICE_X2Y147_BO5;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_A2 = CLBLL_L_X2Y153_SLICE_X1Y153_DO6;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_A3 = CLBLL_L_X2Y147_SLICE_X1Y147_CO6;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_A4 = CLBLL_L_X4Y154_SLICE_X4Y154_CO6;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_A5 = CLBLL_L_X4Y150_SLICE_X4Y150_B5Q;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_A6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_D3 = CLBLM_R_X7Y148_SLICE_X9Y148_DQ;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_D4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_A1 = CLBLM_R_X5Y154_SLICE_X6Y154_BO6;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_B1 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_B2 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_B3 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_B4 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_B5 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_B6 = 1'b1;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_C4 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_D5 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_C1 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_C2 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_C3 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_C4 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_C5 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_C6 = 1'b1;
  assign CLBLL_L_X36Y146_SLICE_X55Y146_A1 = 1'b1;
  assign CLBLL_L_X36Y146_SLICE_X55Y146_A2 = 1'b1;
  assign CLBLL_L_X36Y146_SLICE_X55Y146_A3 = 1'b1;
  assign CLBLL_L_X36Y146_SLICE_X55Y146_A4 = 1'b1;
  assign CLBLL_L_X36Y146_SLICE_X55Y146_A5 = 1'b1;
  assign CLBLL_L_X36Y146_SLICE_X55Y146_A6 = 1'b1;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_D6 = CLBLM_R_X5Y154_SLICE_X7Y154_BO6;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_D1 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_D2 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_D3 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_D4 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_D5 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_D6 = 1'b1;
  assign CLBLL_L_X36Y146_SLICE_X55Y146_B1 = 1'b1;
  assign CLBLL_L_X36Y146_SLICE_X55Y146_B2 = 1'b1;
  assign CLBLL_L_X36Y146_SLICE_X55Y146_B3 = 1'b1;
  assign CLBLL_L_X36Y146_SLICE_X55Y146_B4 = 1'b1;
  assign CLBLL_L_X36Y146_SLICE_X55Y146_B5 = 1'b1;
  assign CLBLL_L_X36Y146_SLICE_X55Y146_B6 = 1'b1;
  assign CLBLL_L_X36Y146_SLICE_X55Y146_C1 = 1'b1;
  assign CLBLL_L_X36Y146_SLICE_X55Y146_C2 = 1'b1;
  assign CLBLL_L_X36Y146_SLICE_X55Y146_C3 = 1'b1;
  assign CLBLL_L_X36Y146_SLICE_X55Y146_C4 = 1'b1;
  assign CLBLL_L_X36Y146_SLICE_X55Y146_C5 = 1'b1;
  assign CLBLL_L_X36Y146_SLICE_X55Y146_C6 = 1'b1;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_D2 = CLBLM_L_X10Y154_SLICE_X12Y154_DQ;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_D3 = CLBLL_L_X2Y146_SLICE_X1Y146_AQ;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_D4 = 1'b1;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_D6 = 1'b1;
  assign CLBLL_L_X36Y146_SLICE_X55Y146_D1 = 1'b1;
  assign CLBLL_L_X36Y146_SLICE_X55Y146_D2 = 1'b1;
  assign CLBLL_L_X36Y146_SLICE_X55Y146_D3 = 1'b1;
  assign CLBLL_L_X36Y146_SLICE_X55Y146_D4 = 1'b1;
  assign CLBLL_L_X36Y146_SLICE_X55Y146_D5 = 1'b1;
  assign CLBLL_L_X36Y146_SLICE_X55Y146_D6 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_A1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_A2 = CLBLM_R_X5Y144_SLICE_X7Y144_BQ;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_A3 = CLBLL_L_X4Y150_SLICE_X4Y150_B5Q;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_A4 = CLBLM_R_X5Y152_SLICE_X7Y152_BQ;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_A5 = CLBLM_R_X3Y148_SLICE_X3Y148_AQ;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_A6 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_AX = CLBLL_L_X2Y147_SLICE_X1Y147_BO5;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_B1 = CLBLL_L_X2Y146_SLICE_X1Y146_AQ;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_B3 = CLBLM_R_X3Y144_SLICE_X3Y144_AQ;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_B4 = CLBLL_L_X2Y146_SLICE_X1Y146_BQ;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_B5 = CLBLL_L_X2Y146_SLICE_X1Y146_CQ;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_B6 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_C1 = CLBLM_R_X3Y143_SLICE_X2Y143_BQ;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_C2 = CLBLM_R_X3Y154_SLICE_X2Y154_BO6;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_C3 = CLBLM_R_X11Y147_SLICE_X15Y147_AQ;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_C4 = CLBLL_L_X2Y147_SLICE_X1Y147_AO5;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_C5 = CLBLM_R_X3Y152_SLICE_X3Y152_CO6;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_C6 = CLBLM_R_X3Y153_SLICE_X2Y153_DO6;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_D3 = CLBLM_R_X7Y152_SLICE_X8Y152_DQ;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_D4 = CLBLM_L_X10Y150_SLICE_X13Y150_CQ;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y167_OLOGIC_X0Y168_D1 = RIOB33_X105Y123_IOB_X1Y123_I;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_D5 = 1'b1;
  assign LIOB33_X0Y179_IOB_X0Y180_O = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_D6 = CLBLL_L_X2Y155_SLICE_X1Y155_DO6;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_D1 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_D2 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_D3 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_D4 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_D5 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_D6 = 1'b1;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_D6 = CLBLM_R_X5Y152_SLICE_X7Y152_DO5;
  assign LIOB33_X0Y179_IOB_X0Y179_O = RIOB33_X105Y131_IOB_X1Y131_I;
  assign LIOI3_X0Y105_OLOGIC_X0Y106_D1 = CLBLL_L_X2Y138_SLICE_X0Y138_CO5;
  assign LIOI3_X0Y167_OLOGIC_X0Y168_T1 = 1'b1;
  assign LIOI3_X0Y167_OLOGIC_X0Y167_D1 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign LIOI3_X0Y105_OLOGIC_X0Y106_T1 = 1'b1;
  assign RIOI3_X105Y151_OLOGIC_X1Y152_D1 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_L_X8Y155_SLICE_X11Y155_A1 = CLBLM_L_X8Y155_SLICE_X11Y155_DO6;
  assign CLBLM_L_X8Y155_SLICE_X11Y155_A2 = CLBLM_L_X10Y154_SLICE_X12Y154_DQ;
  assign CLBLM_L_X8Y155_SLICE_X11Y155_A3 = CLBLM_L_X8Y155_SLICE_X10Y155_CO6;
  assign CLBLM_L_X8Y155_SLICE_X11Y155_A4 = CLBLM_L_X8Y155_SLICE_X11Y155_BO6;
  assign CLBLM_L_X8Y155_SLICE_X11Y155_A5 = CLBLM_L_X10Y154_SLICE_X12Y154_BQ;
  assign CLBLM_L_X8Y155_SLICE_X11Y155_A6 = CLBLM_L_X8Y154_SLICE_X11Y154_DO6;
  assign LIOI3_X0Y167_OLOGIC_X0Y167_T1 = 1'b1;
  assign LIOI3_X0Y105_OLOGIC_X0Y105_D1 = CLBLL_L_X2Y138_SLICE_X0Y138_CO6;
  assign CLBLM_L_X8Y155_SLICE_X11Y155_B1 = CLBLM_L_X8Y155_SLICE_X10Y155_BQ;
  assign CLBLM_L_X8Y155_SLICE_X11Y155_B2 = CLBLM_L_X8Y154_SLICE_X11Y154_AO6;
  assign CLBLM_L_X8Y155_SLICE_X11Y155_B3 = CLBLM_L_X8Y153_SLICE_X11Y153_AQ;
  assign CLBLM_L_X8Y155_SLICE_X11Y155_B4 = CLBLM_L_X10Y154_SLICE_X12Y154_DQ;
  assign CLBLM_L_X8Y155_SLICE_X11Y155_B5 = CLBLM_L_X8Y153_SLICE_X11Y153_BQ;
  assign CLBLM_L_X8Y155_SLICE_X11Y155_B6 = CLBLM_L_X8Y153_SLICE_X11Y153_CQ;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_B5 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_B6 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_L_X8Y155_SLICE_X11Y155_C1 = CLBLM_L_X8Y153_SLICE_X11Y153_CQ;
  assign CLBLM_L_X8Y155_SLICE_X11Y155_C2 = CLBLM_R_X7Y154_SLICE_X8Y154_BQ;
  assign CLBLM_L_X8Y155_SLICE_X11Y155_C3 = CLBLM_R_X7Y153_SLICE_X8Y153_CQ;
  assign CLBLM_L_X8Y155_SLICE_X11Y155_C4 = CLBLM_L_X8Y153_SLICE_X11Y153_AQ;
  assign CLBLM_L_X8Y155_SLICE_X11Y155_C5 = CLBLM_L_X8Y155_SLICE_X10Y155_BQ;
  assign CLBLM_L_X8Y155_SLICE_X11Y155_C6 = CLBLL_L_X4Y147_SLICE_X5Y147_B5Q;
  assign LIOI3_X0Y105_OLOGIC_X0Y105_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_T1 = 1'b1;
  assign RIOI3_X105Y151_OLOGIC_X1Y151_D1 = LIOB33_X0Y75_IOB_X0Y76_I;
  assign RIOI3_X105Y151_OLOGIC_X1Y151_T1 = 1'b1;
  assign CLBLM_L_X8Y155_SLICE_X11Y155_D1 = CLBLM_L_X8Y153_SLICE_X11Y153_CQ;
  assign CLBLM_L_X8Y155_SLICE_X11Y155_D2 = CLBLM_L_X8Y155_SLICE_X10Y155_BQ;
  assign CLBLM_L_X8Y155_SLICE_X11Y155_D3 = CLBLM_L_X8Y153_SLICE_X11Y153_BQ;
  assign CLBLM_L_X8Y155_SLICE_X11Y155_D4 = 1'b1;
  assign CLBLM_L_X8Y155_SLICE_X11Y155_D5 = CLBLM_L_X8Y153_SLICE_X11Y153_AQ;
  assign CLBLM_L_X8Y155_SLICE_X11Y155_D6 = CLBLM_L_X8Y154_SLICE_X11Y154_AO6;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_D1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign LIOB33_X0Y171_IOB_X0Y172_O = CLBLM_R_X103Y141_SLICE_X163Y141_AO6;
  assign LIOB33_X0Y171_IOB_X0Y171_O = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign CLBLM_L_X8Y155_SLICE_X10Y155_A1 = CLBLM_R_X5Y152_SLICE_X7Y152_BQ;
  assign CLBLM_L_X8Y155_SLICE_X10Y155_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y155_SLICE_X10Y155_A3 = CLBLM_L_X8Y155_SLICE_X11Y155_AO6;
  assign CLBLM_L_X8Y155_SLICE_X10Y155_A4 = CLBLM_L_X8Y155_SLICE_X10Y155_AQ;
  assign CLBLM_L_X8Y155_SLICE_X10Y155_A5 = CLBLM_L_X8Y153_SLICE_X10Y153_CO5;
  assign CLBLM_L_X8Y155_SLICE_X10Y155_A6 = CLBLM_L_X8Y153_SLICE_X10Y153_DO6;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_T1 = 1'b1;
  assign CLBLM_L_X8Y155_SLICE_X10Y155_B1 = CLBLM_L_X8Y155_SLICE_X10Y155_DO6;
  assign CLBLM_L_X8Y155_SLICE_X10Y155_B2 = CLBLM_L_X8Y151_SLICE_X10Y151_DQ;
  assign CLBLM_L_X8Y155_SLICE_X10Y155_B3 = CLBLM_L_X8Y153_SLICE_X10Y153_CO5;
  assign CLBLM_L_X8Y155_SLICE_X10Y155_B4 = 1'b1;
  assign CLBLM_L_X8Y155_SLICE_X10Y155_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y155_SLICE_X10Y155_B6 = CLBLM_L_X8Y153_SLICE_X10Y153_DO6;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_C4 = 1'b1;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_C5 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_A4 = 1'b1;
  assign CLBLM_L_X8Y155_SLICE_X10Y155_C1 = CLBLL_L_X4Y147_SLICE_X5Y147_B5Q;
  assign CLBLM_L_X8Y155_SLICE_X10Y155_C2 = CLBLM_R_X5Y155_SLICE_X7Y155_BO5;
  assign CLBLM_L_X8Y155_SLICE_X10Y155_C3 = CLBLM_R_X7Y153_SLICE_X8Y153_CQ;
  assign CLBLM_L_X8Y155_SLICE_X10Y155_C4 = CLBLM_R_X7Y154_SLICE_X8Y154_BQ;
  assign CLBLM_L_X8Y155_SLICE_X10Y155_C5 = CLBLM_R_X7Y155_SLICE_X8Y155_A5Q;
  assign CLBLM_L_X8Y155_SLICE_X10Y155_C6 = CLBLM_R_X7Y155_SLICE_X8Y155_AQ;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_C6 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_A5 = 1'b1;
  assign CLBLM_L_X8Y155_SLICE_X10Y155_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_A6 = 1'b1;
  assign CLBLM_L_X8Y155_SLICE_X10Y155_D1 = CLBLM_L_X8Y155_SLICE_X10Y155_CO6;
  assign CLBLM_L_X8Y155_SLICE_X10Y155_D2 = 1'b1;
  assign CLBLM_L_X8Y155_SLICE_X10Y155_D3 = CLBLM_L_X8Y155_SLICE_X10Y155_BQ;
  assign CLBLM_L_X8Y155_SLICE_X10Y155_D4 = CLBLM_L_X8Y154_SLICE_X11Y154_DO6;
  assign CLBLM_L_X8Y155_SLICE_X10Y155_D5 = CLBLM_R_X7Y155_SLICE_X9Y155_AQ;
  assign CLBLM_L_X8Y155_SLICE_X10Y155_D6 = 1'b1;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_D3 = CLBLM_L_X10Y146_SLICE_X12Y146_DQ;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_D4 = CLBLM_R_X5Y149_SLICE_X7Y149_CQ;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_A1 = CLBLM_R_X3Y143_SLICE_X3Y143_B5Q;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_A2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_A3 = CLBLM_R_X7Y150_SLICE_X9Y150_DO6;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_A4 = CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_A6 = CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_D5 = CLBLM_R_X7Y145_SLICE_X8Y145_BQ;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_C1 = 1'b1;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_B1 = CLBLM_L_X8Y149_SLICE_X10Y149_AO5;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_B2 = CLBLL_L_X4Y146_SLICE_X5Y146_A5Q;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_B3 = CLBLM_R_X7Y143_SLICE_X8Y143_AQ;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_C2 = 1'b1;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_B4 = CLBLM_R_X7Y145_SLICE_X8Y145_BQ;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_B5 = CLBLM_R_X7Y152_SLICE_X9Y152_BQ;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_B6 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_C1 = 1'b1;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_C2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_C3 = CLBLM_R_X5Y144_SLICE_X7Y144_AQ;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_C4 = CLBLL_L_X2Y151_SLICE_X1Y151_BO6;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_C5 = CLBLL_L_X4Y146_SLICE_X4Y146_CO5;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_C6 = CLBLM_L_X10Y144_SLICE_X13Y144_AQ;
  assign CLBLM_R_X103Y176_SLICE_X162Y176_C4 = 1'b1;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_C5 = 1'b1;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_D6 = CLBLM_R_X7Y143_SLICE_X8Y143_AQ;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_A1 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_A2 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_A3 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_A4 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_A5 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_A6 = 1'b1;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_D1 = CLBLM_R_X7Y153_SLICE_X9Y153_CO5;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_D2 = CLBLM_L_X10Y149_SLICE_X12Y149_AO5;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_D3 = CLBLM_R_X5Y144_SLICE_X7Y144_AQ;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_B1 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_B2 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_B3 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_B4 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_B5 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_B6 = 1'b1;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_A2 = CLBLM_L_X10Y149_SLICE_X13Y149_BQ;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_A3 = CLBLM_R_X7Y149_SLICE_X8Y149_DQ;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_C1 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_C2 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_C3 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_C4 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_C5 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_C6 = 1'b1;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_A5 = 1'b1;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_A6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_B1 = CLBLM_R_X7Y148_SLICE_X8Y148_BO5;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_B2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_B3 = 1'b1;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_B4 = CLBLL_L_X4Y149_SLICE_X4Y149_DQ;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_D1 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_D2 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_D3 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_D4 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_D5 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_D6 = 1'b1;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_C2 = 1'b1;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_C3 = CLBLM_R_X3Y149_SLICE_X2Y149_AQ;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_C5 = CLBLM_L_X10Y148_SLICE_X13Y148_BQ;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_C6 = 1'b1;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_D1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_D2 = CLBLM_R_X7Y150_SLICE_X8Y150_DO6;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_D3 = 1'b1;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_D4 = CLBLM_L_X8Y146_SLICE_X11Y146_CO6;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_D6 = CLBLM_R_X5Y148_SLICE_X7Y148_BQ;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_B6 = CLBLM_R_X7Y152_SLICE_X8Y152_BQ;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_A4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_A5 = CLBLM_R_X11Y146_SLICE_X14Y146_AQ;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_A2 = CLBLM_L_X12Y153_SLICE_X16Y153_AQ;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_A3 = CLBLL_L_X2Y148_SLICE_X1Y148_AQ;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_A4 = CLBLM_R_X3Y144_SLICE_X2Y144_CO6;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_A5 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_A6 = CLBLM_R_X3Y144_SLICE_X2Y144_AQ;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_A6 = CLBLM_R_X3Y143_SLICE_X3Y143_A5Q;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_B2 = CLBLM_R_X3Y148_SLICE_X3Y148_AQ;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_B3 = CLBLM_R_X5Y152_SLICE_X7Y152_BQ;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_B4 = CLBLM_R_X5Y144_SLICE_X7Y144_BQ;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_B6 = CLBLL_L_X4Y150_SLICE_X4Y150_B5Q;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_C1 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_C2 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_C3 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_C4 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_C5 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_C6 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_D1 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_D2 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_D3 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_D4 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_D5 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_D6 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_C1 = CLBLM_R_X7Y143_SLICE_X8Y143_B5Q;
  assign LIOB33_X0Y173_IOB_X0Y173_O = CLBLM_R_X103Y141_SLICE_X163Y141_AO5;
  assign LIOB33_X0Y173_IOB_X0Y174_O = CLBLM_L_X8Y159_SLICE_X10Y159_AO6;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_C2 = CLBLM_R_X5Y144_SLICE_X7Y144_CQ;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_C5 = CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_C6 = CLBLM_R_X5Y146_SLICE_X7Y146_DO6;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_B5 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_B6 = CLBLM_R_X7Y142_SLICE_X8Y142_BQ;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_C1 = CLBLM_R_X3Y148_SLICE_X3Y148_AQ;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_C2 = CLBLM_R_X7Y142_SLICE_X8Y142_CQ;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_C4 = CLBLM_R_X7Y142_SLICE_X8Y142_BQ;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_C5 = CLBLM_R_X7Y142_SLICE_X8Y142_DO6;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_C6 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_A1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_A2 = CLBLM_L_X8Y150_SLICE_X11Y150_CO6;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_A3 = CLBLM_R_X7Y150_SLICE_X9Y150_AQ;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_A4 = CLBLM_L_X8Y143_SLICE_X10Y143_BQ;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_A6 = CLBLM_R_X7Y150_SLICE_X9Y150_CO6;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_C4 = 1'b1;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_AX = CLBLM_R_X7Y150_SLICE_X9Y150_BO6;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_B1 = CLBLM_L_X8Y150_SLICE_X10Y150_CQ;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_B2 = CLBLM_R_X7Y145_SLICE_X8Y145_CQ;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_B4 = CLBLM_R_X11Y153_SLICE_X14Y153_BQ;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_B6 = 1'b1;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_C1 = CLBLM_R_X7Y148_SLICE_X8Y148_CQ;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_C2 = CLBLM_R_X5Y146_SLICE_X6Y146_CQ;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_C3 = CLBLM_L_X8Y146_SLICE_X10Y146_AQ;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_C4 = CLBLM_R_X7Y150_SLICE_X9Y150_A5Q;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_C5 = CLBLM_R_X7Y150_SLICE_X9Y150_BO5;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_D1 = CLBLM_R_X3Y152_SLICE_X3Y152_CO6;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_C6 = 1'b1;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_A1 = CLBLL_L_X2Y152_SLICE_X1Y152_AO5;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_A2 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_A3 = CLBLL_L_X2Y148_SLICE_X1Y148_AQ;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_A4 = CLBLL_L_X2Y150_SLICE_X0Y150_AO5;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_A5 = LIOB33_X0Y55_IOB_X0Y55_I;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_A6 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_D2 = CLBLM_R_X5Y145_SLICE_X6Y145_DO6;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_D3 = CLBLM_R_X5Y143_SLICE_X7Y143_BO6;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_B1 = CLBLL_L_X2Y152_SLICE_X1Y152_AO5;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_B2 = CLBLM_R_X3Y143_SLICE_X2Y143_DQ;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_B3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_B4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_B5 = LIOB33_X0Y57_IOB_X0Y57_I;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_B6 = CLBLL_L_X2Y150_SLICE_X0Y150_AO5;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_D4 = CLBLL_L_X2Y151_SLICE_X1Y151_BO6;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_D5 = CLBLM_R_X5Y144_SLICE_X6Y144_DO6;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_C1 = CLBLL_L_X2Y152_SLICE_X1Y152_AO5;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_C2 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_C3 = LIOB33_X0Y63_IOB_X0Y63_I;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_C4 = CLBLM_R_X5Y149_SLICE_X6Y149_CO5;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_C5 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_C6 = LIOB33_X0Y57_IOB_X0Y58_I;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_D6 = 1'b1;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_A1 = CLBLM_L_X8Y151_SLICE_X11Y151_DQ;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_A3 = CLBLM_R_X7Y150_SLICE_X8Y150_AQ;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_A4 = CLBLL_L_X4Y151_SLICE_X4Y151_AQ;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_A5 = CLBLM_L_X8Y149_SLICE_X11Y149_AQ;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_A6 = CLBLM_R_X7Y145_SLICE_X8Y145_AQ;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_D1 = 1'b1;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_D2 = 1'b1;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_D3 = 1'b1;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_D4 = 1'b1;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_D5 = 1'b1;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_D6 = 1'b1;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_B5 = 1'b1;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_C2 = CLBLM_R_X7Y150_SLICE_X8Y150_CQ;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_C3 = CLBLM_R_X7Y148_SLICE_X8Y148_DQ;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_C4 = CLBLM_R_X7Y148_SLICE_X9Y148_CQ;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_C5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_C6 = CLBLM_R_X7Y150_SLICE_X9Y150_CO5;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign LIOB33_X0Y109_IOB_X0Y110_O = CLBLL_L_X2Y134_SLICE_X0Y134_AO5;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_C3 = CLBLM_R_X11Y154_SLICE_X14Y154_AQ;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_D1 = CLBLM_L_X8Y154_SLICE_X10Y154_AQ;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_D2 = CLBLM_R_X7Y153_SLICE_X9Y153_A5Q;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_D3 = 1'b1;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_D4 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_B6 = 1'b1;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_D5 = CLBLM_R_X7Y149_SLICE_X8Y149_DQ;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_D6 = CLBLM_R_X5Y150_SLICE_X7Y150_BQ;
  assign CLBLM_R_X103Y176_SLICE_X162Y176_D3 = 1'b1;
  assign LIOB33_X0Y109_IOB_X0Y109_O = CLBLL_L_X2Y134_SLICE_X0Y134_AO6;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_A1 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_A2 = CLBLL_L_X4Y155_SLICE_X4Y155_BO6;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_A3 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_A4 = CLBLM_R_X5Y150_SLICE_X6Y150_AQ;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_A5 = CLBLM_R_X3Y144_SLICE_X3Y144_AQ;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_A6 = CLBLL_L_X2Y152_SLICE_X1Y152_AO5;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_B1 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_B2 = CLBLM_R_X3Y148_SLICE_X3Y148_CQ;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_B3 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_B4 = CLBLM_R_X3Y145_SLICE_X3Y145_AQ;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_B5 = CLBLL_L_X2Y151_SLICE_X0Y151_CO5;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_B6 = CLBLL_L_X2Y152_SLICE_X1Y152_AO5;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X103Y176_SLICE_X162Y176_D4 = 1'b1;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_C1 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_C2 = CLBLL_L_X4Y155_SLICE_X4Y155_BO6;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_C3 = CLBLL_L_X2Y151_SLICE_X1Y151_AO5;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_C4 = CLBLL_L_X4Y146_SLICE_X5Y146_CQ;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_C5 = CLBLL_L_X2Y152_SLICE_X1Y152_AO5;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_C6 = CLBLL_L_X2Y146_SLICE_X1Y146_BQ;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_C3 = CLBLM_R_X3Y144_SLICE_X2Y144_AQ;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_D1 = CLBLL_L_X2Y145_SLICE_X1Y145_BQ;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_D2 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_D3 = CLBLL_L_X2Y152_SLICE_X1Y152_AO5;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_D4 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_D5 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_D6 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_C4 = CLBLM_R_X7Y145_SLICE_X8Y145_C5Q;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_C5 = CLBLM_R_X3Y144_SLICE_X2Y144_A5Q;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_C6 = CLBLM_R_X3Y143_SLICE_X3Y143_B5Q;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_D1 = CLBLM_R_X11Y154_SLICE_X14Y154_AQ;
  assign LIOB33_X0Y175_IOB_X0Y176_O = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_D2 = CLBLM_R_X11Y154_SLICE_X15Y154_AQ;
  assign LIOB33_X0Y175_IOB_X0Y175_O = RIOB33_X105Y127_IOB_X1Y127_I;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_D4 = CLBLM_R_X11Y152_SLICE_X15Y152_AQ;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_D5 = CLBLM_R_X11Y153_SLICE_X15Y153_AQ;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_A1 = CLBLM_R_X7Y154_SLICE_X9Y154_AQ;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_D5 = CLBLM_L_X8Y146_SLICE_X10Y146_DO6;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_C2 = CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_D6 = CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  assign LIOI3_X0Y171_OLOGIC_X0Y172_D1 = CLBLM_R_X103Y141_SLICE_X163Y141_AO6;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_C3 = CLBLM_R_X11Y144_SLICE_X14Y144_BQ;
  assign RIOI3_SING_X105Y100_ILOGIC_X1Y100_D = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_L_X10Y155_SLICE_X13Y155_C3 = CLBLM_R_X11Y148_SLICE_X15Y148_CQ;
  assign LIOI3_X0Y171_OLOGIC_X0Y172_T1 = 1'b1;
  assign LIOI3_X0Y109_OLOGIC_X0Y110_D1 = CLBLL_L_X2Y134_SLICE_X0Y134_AO5;
  assign LIOI3_X0Y171_OLOGIC_X0Y171_D1 = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign LIOI3_X0Y109_OLOGIC_X0Y110_T1 = 1'b1;
  assign RIOI3_X105Y153_OLOGIC_X1Y154_D1 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign LIOI3_X0Y171_OLOGIC_X0Y171_T1 = 1'b1;
  assign CLBLM_L_X10Y155_SLICE_X13Y155_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign LIOI3_X0Y109_OLOGIC_X0Y109_D1 = CLBLL_L_X2Y134_SLICE_X0Y134_AO6;
  assign RIOI3_X105Y153_OLOGIC_X1Y154_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_D1 = CLBLM_R_X3Y143_SLICE_X3Y143_BQ;
  assign LIOI3_X0Y109_OLOGIC_X0Y109_T1 = 1'b1;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_C5 = CLBLM_R_X11Y146_SLICE_X14Y146_CQ;
  assign RIOI3_X105Y153_OLOGIC_X1Y153_D1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_T1 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_A1 = CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_A2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_A3 = CLBLM_R_X7Y151_SLICE_X9Y151_AQ;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_A4 = CLBLL_L_X4Y151_SLICE_X4Y151_AQ;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_A5 = CLBLM_R_X7Y153_SLICE_X9Y153_CO5;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_D1 = CLBLM_R_X3Y142_SLICE_X2Y142_AQ;
  assign CLBLM_L_X10Y155_SLICE_X13Y155_D1 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_B1 = CLBLM_L_X10Y152_SLICE_X13Y152_BQ;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_B2 = CLBLM_R_X7Y151_SLICE_X9Y151_BQ;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_B4 = CLBLL_L_X4Y151_SLICE_X4Y151_AQ;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_B5 = CLBLM_L_X8Y149_SLICE_X11Y149_AQ;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_B6 = CLBLM_R_X3Y147_SLICE_X3Y147_BQ;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_C6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_T1 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_C1 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_C2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_C3 = CLBLM_R_X7Y153_SLICE_X9Y153_DQ;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_C5 = CLBLM_R_X7Y150_SLICE_X9Y150_DO6;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_A1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_A2 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_A3 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_A4 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_A5 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_A6 = 1'b1;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_C5 = CLBLM_R_X11Y153_SLICE_X15Y153_AQ;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_C6 = CLBLM_L_X8Y151_SLICE_X10Y151_AQ;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_B1 = CLBLL_L_X2Y152_SLICE_X1Y152_AO5;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_B2 = LIOB33_X0Y59_IOB_X0Y59_I;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_B3 = CLBLL_L_X2Y154_SLICE_X1Y154_BO5;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_B4 = CLBLM_R_X3Y149_SLICE_X2Y149_CQ;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_B5 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_B6 = CLBLL_L_X2Y151_SLICE_X0Y151_CO5;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_D1 = CLBLM_L_X8Y146_SLICE_X10Y146_BQ;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_D2 = CLBLM_R_X3Y147_SLICE_X3Y147_BQ;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_C1 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_C2 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_C3 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_C4 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_C5 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_C6 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_A1 = CLBLM_R_X5Y152_SLICE_X7Y152_DO5;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_A2 = CLBLM_L_X10Y149_SLICE_X12Y149_AQ;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_A3 = CLBLM_R_X7Y151_SLICE_X8Y151_AQ;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_A4 = CLBLM_R_X5Y149_SLICE_X7Y149_BQ;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_A6 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_AX = CLBLM_R_X7Y151_SLICE_X8Y151_CO6;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_B1 = CLBLM_R_X3Y149_SLICE_X3Y149_AQ;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_D1 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_D2 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_D3 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_D4 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_D5 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_D6 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_B2 = CLBLM_R_X7Y151_SLICE_X8Y151_BQ;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_B3 = CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_B4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_B6 = CLBLM_R_X7Y143_SLICE_X8Y143_CQ;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_C1 = CLBLM_R_X7Y151_SLICE_X8Y151_BQ;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_C2 = CLBLL_L_X4Y145_SLICE_X5Y145_CO6;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_C3 = CLBLM_L_X10Y153_SLICE_X12Y153_CQ;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_C4 = CLBLM_R_X7Y151_SLICE_X8Y151_A5Q;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_C6 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_D1 = CLBLM_L_X10Y149_SLICE_X13Y149_BQ;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_D2 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_D3 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_D4 = CLBLM_R_X5Y152_SLICE_X6Y152_CQ;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_D5 = CLBLM_R_X11Y146_SLICE_X14Y146_DQ;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_D6 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_A1 = CLBLL_L_X2Y154_SLICE_X1Y154_BO6;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_A2 = CLBLM_R_X3Y150_SLICE_X2Y150_AO6;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_A3 = CLBLL_L_X2Y149_SLICE_X1Y149_AO6;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_A4 = CLBLL_L_X2Y150_SLICE_X1Y150_BO6;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_A5 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_A6 = CLBLL_L_X2Y149_SLICE_X0Y149_BO6;
  assign CLBLM_L_X10Y155_SLICE_X12Y155_A6 = CLBLM_L_X8Y153_SLICE_X10Y153_DO6;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_B2 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_B3 = CLBLL_L_X2Y152_SLICE_X1Y152_AO5;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_B4 = CLBLL_L_X2Y154_SLICE_X1Y154_BO5;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_B5 = CLBLL_L_X2Y151_SLICE_X1Y151_AO5;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_B6 = CLBLM_R_X5Y153_SLICE_X6Y153_A5Q;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_C1 = CLBLL_L_X2Y149_SLICE_X1Y149_BO6;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_C2 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_C3 = CLBLM_R_X3Y150_SLICE_X2Y150_CO6;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_C4 = CLBLL_L_X2Y154_SLICE_X1Y154_BO6;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_C5 = CLBLL_L_X2Y149_SLICE_X0Y149_CO6;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_C6 = CLBLL_L_X2Y149_SLICE_X1Y149_CO6;
  assign LIOB33_X0Y177_IOB_X0Y177_O = RIOB33_X105Y129_IOB_X1Y129_I;
  assign LIOB33_X0Y177_IOB_X0Y178_O = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLM_L_X10Y155_SLICE_X12Y155_B1 = CLBLM_L_X10Y156_SLICE_X12Y156_AO5;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_D1 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_D2 = LIOB33_X0Y65_IOB_X0Y65_I;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_D3 = CLBLM_R_X5Y150_SLICE_X6Y150_A5Q;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_D4 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_D5 = CLBLL_L_X2Y152_SLICE_X1Y152_AO5;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_D6 = CLBLL_L_X2Y154_SLICE_X1Y154_BO5;
  assign CLBLM_L_X10Y155_SLICE_X12Y155_B2 = CLBLM_L_X10Y155_SLICE_X13Y155_DO6;
  assign CLBLM_L_X10Y155_SLICE_X12Y155_B3 = CLBLM_L_X10Y153_SLICE_X13Y153_AQ;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_A3 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_A4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X10Y155_SLICE_X12Y155_C6 = CLBLM_L_X10Y155_SLICE_X13Y155_BQ;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_C1 = CLBLM_R_X5Y142_SLICE_X7Y142_AQ;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_C2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_C3 = 1'b1;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_C5 = 1'b1;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign RIOI3_SING_X105Y149_ILOGIC_X1Y149_D = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_A1 = 1'b1;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_A2 = CLBLM_L_X8Y153_SLICE_X10Y153_DO5;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_A4 = CLBLM_R_X5Y152_SLICE_X6Y152_BQ;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_A5 = CLBLM_L_X10Y152_SLICE_X12Y152_BQ;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_A6 = 1'b1;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_B1 = 1'b1;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_B2 = CLBLM_R_X7Y152_SLICE_X9Y152_BQ;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_B4 = 1'b1;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_B6 = CLBLM_R_X7Y152_SLICE_X8Y152_CQ;
  assign CLBLL_L_X2Y151_SLICE_X0Y151_A1 = CLBLL_L_X2Y152_SLICE_X1Y152_AO5;
  assign CLBLL_L_X2Y151_SLICE_X0Y151_A2 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y151_SLICE_X0Y151_A3 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y151_SLICE_X0Y151_A4 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y151_SLICE_X0Y151_A5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y151_SLICE_X0Y151_A6 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_A1 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_A2 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_A3 = 1'b1;
  assign CLBLL_L_X2Y151_SLICE_X0Y151_B1 = CLBLL_L_X2Y152_SLICE_X1Y152_AO5;
  assign CLBLL_L_X2Y151_SLICE_X0Y151_B2 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y151_SLICE_X0Y151_B3 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y151_SLICE_X0Y151_B4 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y151_SLICE_X0Y151_B5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y151_SLICE_X0Y151_B6 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_AX = CLBLM_R_X7Y142_SLICE_X8Y142_AO6;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_B1 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_B2 = 1'b1;
  assign CLBLL_L_X2Y151_SLICE_X0Y151_C1 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y151_SLICE_X0Y151_C2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y151_SLICE_X0Y151_C3 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y151_SLICE_X0Y151_C4 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y151_SLICE_X0Y151_C5 = CLBLL_L_X2Y152_SLICE_X1Y152_AO5;
  assign CLBLL_L_X2Y151_SLICE_X0Y151_C6 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_C3 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_C4 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_C5 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_C6 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_A1 = 1'b1;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_A2 = CLBLM_L_X8Y152_SLICE_X11Y152_BO6;
  assign CLBLL_L_X2Y151_SLICE_X0Y151_D1 = LIOB33_X0Y53_IOB_X0Y54_I;
  assign CLBLL_L_X2Y151_SLICE_X0Y151_D2 = CLBLL_L_X2Y146_SLICE_X1Y146_AQ;
  assign CLBLL_L_X2Y151_SLICE_X0Y151_D3 = CLBLL_L_X2Y151_SLICE_X0Y151_AO5;
  assign CLBLL_L_X2Y151_SLICE_X0Y151_D4 = CLBLL_L_X2Y151_SLICE_X0Y151_CO6;
  assign CLBLL_L_X2Y151_SLICE_X0Y151_D5 = CLBLL_L_X2Y151_SLICE_X0Y151_BO5;
  assign CLBLL_L_X2Y151_SLICE_X0Y151_D6 = CLBLM_R_X5Y146_SLICE_X6Y146_A5Q;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_D1 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_D2 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_D3 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_D4 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_D5 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_D6 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_A1 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_A2 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_A3 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_A4 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_A5 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_A6 = 1'b1;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_C2 = CLBLM_R_X7Y152_SLICE_X8Y152_CQ;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_C3 = CLBLM_R_X7Y153_SLICE_X9Y153_DQ;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_B1 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_B2 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_B3 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_B4 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_B5 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_B6 = 1'b1;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_D2 = CLBLM_R_X7Y153_SLICE_X9Y153_A5Q;
  assign CLBLL_L_X2Y151_SLICE_X1Y151_A1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y151_SLICE_X1Y151_A2 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y151_SLICE_X1Y151_A3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y151_SLICE_X1Y151_A4 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y151_SLICE_X1Y151_A5 = 1'b1;
  assign CLBLL_L_X2Y151_SLICE_X1Y151_A6 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_C1 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_C2 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_C3 = 1'b1;
  assign CLBLL_L_X2Y151_SLICE_X1Y151_B1 = CLBLM_R_X3Y150_SLICE_X2Y150_DO6;
  assign CLBLL_L_X2Y151_SLICE_X1Y151_B2 = CLBLL_L_X2Y151_SLICE_X0Y151_DO6;
  assign CLBLL_L_X2Y151_SLICE_X1Y151_B3 = CLBLM_R_X5Y153_SLICE_X6Y153_DO6;
  assign CLBLL_L_X2Y151_SLICE_X1Y151_B4 = CLBLM_R_X3Y152_SLICE_X3Y152_BO6;
  assign CLBLL_L_X2Y151_SLICE_X1Y151_B5 = CLBLM_R_X3Y155_SLICE_X2Y155_DO6;
  assign CLBLL_L_X2Y151_SLICE_X1Y151_B6 = CLBLL_L_X2Y151_SLICE_X1Y151_CO6;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_D1 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_D2 = 1'b1;
  assign CLBLL_L_X2Y151_SLICE_X1Y151_C1 = CLBLL_L_X2Y154_SLICE_X1Y154_CO5;
  assign CLBLL_L_X2Y151_SLICE_X1Y151_C2 = CLBLM_R_X3Y156_SLICE_X2Y156_CO6;
  assign CLBLL_L_X2Y151_SLICE_X1Y151_C3 = LIOB33_X0Y69_IOB_X0Y70_I;
  assign CLBLL_L_X2Y151_SLICE_X1Y151_C4 = CLBLL_L_X4Y151_SLICE_X4Y151_A5Q;
  assign CLBLL_L_X2Y151_SLICE_X1Y151_C5 = CLBLM_L_X16Y158_SLICE_X22Y158_AO5;
  assign CLBLL_L_X2Y151_SLICE_X1Y151_C6 = CLBLL_L_X2Y150_SLICE_X0Y150_BO6;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_D3 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_D4 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_D5 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_D6 = 1'b1;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_C1 = CLBLM_R_X3Y152_SLICE_X3Y152_CO6;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_C2 = CLBLM_R_X7Y154_SLICE_X9Y154_AQ;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X2Y151_SLICE_X1Y151_D1 = CLBLL_L_X2Y151_SLICE_X1Y151_AO6;
  assign CLBLL_L_X2Y151_SLICE_X1Y151_D2 = LIOB33_X0Y71_IOB_X0Y71_I;
  assign CLBLL_L_X2Y151_SLICE_X1Y151_D3 = CLBLL_L_X2Y152_SLICE_X1Y152_AO5;
  assign CLBLL_L_X2Y151_SLICE_X1Y151_D4 = 1'b1;
  assign CLBLL_L_X2Y151_SLICE_X1Y151_D5 = CLBLL_L_X2Y146_SLICE_X1Y146_CQ;
  assign CLBLL_L_X2Y151_SLICE_X1Y151_D6 = CLBLL_L_X4Y155_SLICE_X4Y155_BO6;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_C5 = CLBLM_R_X7Y153_SLICE_X8Y153_DQ;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I0 = LIOB33_X0Y77_IOB_X0Y78_I;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I1 = 1'b1;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_C6 = 1'b1;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X8Y159_SLICE_X11Y159_A1 = 1'b1;
  assign CLBLM_L_X8Y159_SLICE_X11Y159_A2 = 1'b1;
  assign CLBLM_L_X8Y159_SLICE_X11Y159_A3 = 1'b1;
  assign CLBLM_L_X8Y159_SLICE_X11Y159_A4 = 1'b1;
  assign CLBLM_L_X8Y159_SLICE_X11Y159_A5 = 1'b1;
  assign CLBLM_L_X8Y159_SLICE_X11Y159_A6 = 1'b1;
  assign CLBLM_L_X8Y159_SLICE_X11Y159_B1 = 1'b1;
  assign CLBLM_L_X8Y159_SLICE_X11Y159_B2 = 1'b1;
  assign CLBLM_L_X8Y159_SLICE_X11Y159_B3 = 1'b1;
  assign CLBLM_L_X8Y159_SLICE_X11Y159_B4 = 1'b1;
  assign CLBLM_L_X8Y159_SLICE_X11Y159_B5 = 1'b1;
  assign CLBLM_L_X8Y159_SLICE_X11Y159_B6 = 1'b1;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y159_SLICE_X11Y159_C1 = 1'b1;
  assign CLBLM_L_X8Y159_SLICE_X11Y159_C2 = 1'b1;
  assign CLBLM_L_X8Y159_SLICE_X11Y159_C3 = 1'b1;
  assign CLBLM_L_X8Y159_SLICE_X11Y159_C4 = 1'b1;
  assign CLBLM_L_X8Y159_SLICE_X11Y159_C5 = 1'b1;
  assign CLBLM_L_X8Y159_SLICE_X11Y159_C6 = 1'b1;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_D2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_D3 = CLBLL_L_X4Y147_SLICE_X4Y147_CQ;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_D4 = CLBLM_L_X8Y150_SLICE_X10Y150_DO6;
  assign CLBLM_L_X8Y159_SLICE_X11Y159_D1 = 1'b1;
  assign CLBLM_L_X8Y159_SLICE_X11Y159_D2 = 1'b1;
  assign CLBLM_L_X8Y159_SLICE_X11Y159_D3 = 1'b1;
  assign CLBLM_L_X8Y159_SLICE_X11Y159_D4 = 1'b1;
  assign CLBLM_L_X8Y159_SLICE_X11Y159_D5 = 1'b1;
  assign CLBLM_L_X8Y159_SLICE_X11Y159_D6 = 1'b1;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_D5 = 1'b1;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_D6 = CLBLM_L_X8Y152_SLICE_X10Y152_AQ;
  assign CLBLM_L_X8Y159_SLICE_X10Y159_A1 = CLBLM_L_X8Y151_SLICE_X10Y151_B5Q;
  assign CLBLM_L_X8Y159_SLICE_X10Y159_A2 = 1'b1;
  assign CLBLM_L_X8Y159_SLICE_X10Y159_A3 = 1'b1;
  assign CLBLM_L_X8Y159_SLICE_X10Y159_A4 = 1'b1;
  assign CLBLM_L_X8Y159_SLICE_X10Y159_A5 = 1'b1;
  assign CLBLM_L_X8Y159_SLICE_X10Y159_A6 = 1'b1;
  assign CLBLM_L_X8Y159_SLICE_X10Y159_B1 = 1'b1;
  assign CLBLM_L_X8Y159_SLICE_X10Y159_B2 = 1'b1;
  assign CLBLM_L_X8Y159_SLICE_X10Y159_B3 = 1'b1;
  assign CLBLM_L_X8Y159_SLICE_X10Y159_B4 = 1'b1;
  assign CLBLM_L_X8Y159_SLICE_X10Y159_B5 = 1'b1;
  assign CLBLM_L_X8Y159_SLICE_X10Y159_B6 = 1'b1;
  assign CLBLM_L_X8Y159_SLICE_X10Y159_C1 = 1'b1;
  assign CLBLM_L_X8Y159_SLICE_X10Y159_C2 = 1'b1;
  assign CLBLM_L_X8Y159_SLICE_X10Y159_C3 = 1'b1;
  assign CLBLM_L_X8Y159_SLICE_X10Y159_C4 = 1'b1;
  assign CLBLM_L_X8Y159_SLICE_X10Y159_C5 = 1'b1;
  assign CLBLM_L_X8Y159_SLICE_X10Y159_C6 = 1'b1;
  assign RIOI3_X105Y197_OLOGIC_X1Y198_D1 = CLBLM_L_X16Y158_SLICE_X22Y158_AO6;
  assign RIOI3_SING_X105Y150_OLOGIC_X1Y150_D1 = LIOB33_X0Y75_IOB_X0Y75_I;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_A1 = CLBLM_R_X5Y154_SLICE_X6Y154_BO6;
  assign CLBLM_L_X8Y159_SLICE_X10Y159_D1 = 1'b1;
  assign CLBLM_L_X8Y159_SLICE_X10Y159_D2 = 1'b1;
  assign CLBLM_L_X8Y159_SLICE_X10Y159_D3 = 1'b1;
  assign CLBLM_L_X8Y159_SLICE_X10Y159_D4 = 1'b1;
  assign CLBLM_L_X8Y159_SLICE_X10Y159_D5 = 1'b1;
  assign CLBLM_L_X8Y159_SLICE_X10Y159_D6 = 1'b1;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_A2 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign RIOI3_SING_X105Y150_OLOGIC_X1Y150_T1 = 1'b1;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_A3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_A4 = CLBLM_L_X10Y153_SLICE_X12Y153_DQ;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_A5 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_D4 = CLBLM_L_X8Y146_SLICE_X10Y146_BQ;
  assign CLBLM_R_X5Y155_SLICE_X7Y155_C1 = CLBLM_R_X5Y155_SLICE_X6Y155_AQ;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_D5 = CLBLM_L_X8Y146_SLICE_X11Y146_BQ;
  assign CLBLM_R_X5Y155_SLICE_X7Y155_C2 = CLBLM_R_X5Y152_SLICE_X6Y152_AQ;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_D6 = 1'b1;
  assign CLBLM_R_X5Y155_SLICE_X7Y155_C3 = CLBLM_R_X7Y155_SLICE_X8Y155_AQ;
  assign RIOI3_X105Y197_OLOGIC_X1Y198_T1 = 1'b1;
  assign LIOB33_X0Y181_IOB_X0Y182_O = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_B2 = CLBLM_R_X7Y153_SLICE_X8Y153_BQ;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_A2 = CLBLM_L_X8Y146_SLICE_X10Y146_BQ;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_A3 = CLBLM_R_X7Y155_SLICE_X8Y155_BO5;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_A4 = CLBLM_L_X8Y144_SLICE_X10Y144_BQ;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_B3 = CLBLM_R_X5Y155_SLICE_X7Y155_CO6;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_A5 = CLBLM_R_X5Y146_SLICE_X7Y146_BO6;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_A6 = CLBLM_R_X7Y154_SLICE_X9Y154_CO6;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_SR = CLBLM_R_X11Y151_SLICE_X15Y151_CO6;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_AX = CLBLM_R_X7Y153_SLICE_X9Y153_CO6;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_B1 = CLBLM_L_X8Y152_SLICE_X11Y152_AQ;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_B2 = CLBLM_R_X7Y153_SLICE_X9Y153_BQ;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_B3 = CLBLM_L_X8Y152_SLICE_X11Y152_BO6;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_B4 = 1'b1;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_B5 = CLBLM_R_X7Y155_SLICE_X9Y155_AQ;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_A1 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_A2 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_A3 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_A4 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_A5 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_A6 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_A1 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_A2 = CLBLL_L_X4Y144_SLICE_X4Y144_BQ;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_A3 = CLBLM_R_X5Y143_SLICE_X7Y143_AQ;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_B1 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_B2 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_B3 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_B4 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_B5 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_B6 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_A4 = CLBLM_L_X8Y143_SLICE_X11Y143_AQ;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_A6 = CLBLM_R_X5Y143_SLICE_X7Y143_CO6;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_C1 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_C2 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_C3 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_C4 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_C5 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_C6 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_B3 = CLBLL_L_X2Y153_SLICE_X1Y153_DO6;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_B4 = CLBLM_R_X3Y154_SLICE_X2Y154_BO6;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_B5 = CLBLM_R_X3Y152_SLICE_X3Y152_CO6;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_B6 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_C1 = CLBLM_R_X3Y152_SLICE_X3Y152_CO6;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_C2 = CLBLL_L_X2Y151_SLICE_X1Y151_BO6;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_C3 = CLBLM_R_X5Y145_SLICE_X6Y145_DO6;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_D1 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_D2 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_D3 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_D4 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_D5 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_D6 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_D1 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_D2 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_D3 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_D4 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_D5 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_D6 = 1'b1;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_B1 = CLBLM_R_X7Y155_SLICE_X8Y155_BO5;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_A1 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_A2 = CLBLM_R_X11Y143_SLICE_X14Y143_AQ;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_A3 = CLBLM_R_X5Y143_SLICE_X6Y143_AQ;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_A4 = CLBLM_R_X7Y142_SLICE_X8Y142_DO6;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_A6 = CLBLL_L_X4Y145_SLICE_X4Y145_A5Q;
  assign CLBLM_R_X5Y155_SLICE_X7Y155_D5 = 1'b1;
  assign CLBLM_R_X5Y155_SLICE_X7Y155_D6 = CLBLM_R_X5Y155_SLICE_X6Y155_BQ;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_C1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_B1 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_B2 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_B3 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_B4 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_B5 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_B6 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_A1 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_A2 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_A3 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_A4 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_A5 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_A6 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_C1 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_C2 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_B1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_B2 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_B3 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_B4 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_B5 = CLBLL_L_X2Y152_SLICE_X1Y152_AO6;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_B6 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_C3 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_C4 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_C6 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_C1 = CLBLL_L_X2Y152_SLICE_X1Y152_AO6;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_C2 = CLBLL_L_X4Y155_SLICE_X4Y155_BO6;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_C3 = CLBLL_L_X2Y154_SLICE_X1Y154_BO5;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_C4 = CLBLL_L_X2Y155_SLICE_X1Y155_DO6;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_C5 = CLBLM_R_X3Y145_SLICE_X3Y145_BQ;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_C6 = CLBLL_L_X4Y151_SLICE_X5Y151_AQ;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_D6 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_D1 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_D2 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_D3 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_D4 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_D5 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_D1 = CLBLL_L_X4Y151_SLICE_X5Y151_AQ;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_D2 = CLBLL_L_X4Y155_SLICE_X5Y155_AO6;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_D3 = CLBLL_L_X2Y154_SLICE_X1Y154_BO6;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_D4 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_D5 = CLBLL_L_X2Y152_SLICE_X1Y152_BO5;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_D6 = CLBLM_R_X3Y145_SLICE_X3Y145_BQ;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_D1 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_T1 = 1'b1;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_D2 = CLBLM_L_X10Y153_SLICE_X12Y153_DQ;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_D3 = CLBLM_R_X11Y153_SLICE_X14Y153_AO6;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_D4 = CLBLL_L_X4Y151_SLICE_X5Y151_BQ;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_D5 = 1'b1;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_D6 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE0 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE1 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE0 = 1'b1;
  assign CLBLM_R_X5Y155_SLICE_X6Y155_B5 = CLBLM_R_X5Y155_SLICE_X7Y155_BO6;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE1 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S0 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S1 = 1'b1;
  assign CLBLM_R_X5Y155_SLICE_X6Y155_B6 = CLBLM_R_X5Y152_SLICE_X6Y152_AQ;
  assign CLBLM_R_X5Y155_SLICE_X6Y155_C4 = 1'b1;
  assign CLBLM_R_X5Y155_SLICE_X6Y155_C5 = 1'b1;
  assign CLBLM_R_X5Y155_SLICE_X6Y155_C6 = 1'b1;
  assign LIOI3_X0Y51_ILOGIC_X0Y52_D = LIOB33_X0Y51_IOB_X0Y52_I;
  assign LIOI3_X0Y51_ILOGIC_X0Y51_D = LIOB33_X0Y51_IOB_X0Y51_I;
  assign RIOI3_SING_X105Y199_OLOGIC_X1Y199_D1 = CLBLM_L_X12Y155_SLICE_X17Y155_AQ;
  assign RIOB33_X105Y151_IOB_X1Y152_O = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign RIOB33_X105Y151_IOB_X1Y151_O = LIOB33_X0Y75_IOB_X0Y76_I;
  assign RIOI3_SING_X105Y199_OLOGIC_X1Y199_T1 = 1'b1;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_A1 = CLBLM_L_X8Y154_SLICE_X10Y154_AQ;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_A2 = CLBLM_L_X8Y152_SLICE_X11Y152_AQ;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_C1 = CLBLM_R_X5Y146_SLICE_X6Y146_AQ;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_A3 = 1'b1;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_A6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y58_D = LIOB33_X0Y57_IOB_X0Y58_I;
  assign LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y57_D = LIOB33_X0Y57_IOB_X0Y57_I;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_A1 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_A2 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_A3 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_A4 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_A5 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_A6 = 1'b1;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_B1 = 1'b1;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_B2 = CLBLM_R_X7Y155_SLICE_X9Y155_BO6;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_B3 = CLBLM_R_X7Y151_SLICE_X9Y151_DO5;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_B1 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_B2 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_B3 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_B4 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_B5 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_B6 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_A1 = CLBLM_R_X5Y144_SLICE_X7Y144_AQ;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_A2 = CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_C1 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_C2 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_C3 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_C4 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_C5 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_C6 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_B1 = CLBLM_R_X7Y144_SLICE_X9Y144_A5Q;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_B2 = CLBLM_R_X3Y148_SLICE_X3Y148_AQ;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_B4 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_B5 = CLBLM_R_X5Y152_SLICE_X7Y152_AQ;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_B6 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_D1 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_D2 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_D3 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_D4 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_D5 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_D6 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_C3 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_D2 = CLBLM_L_X10Y144_SLICE_X13Y144_AQ;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_D3 = CLBLM_L_X8Y145_SLICE_X10Y145_CO6;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_D4 = CLBLM_R_X5Y146_SLICE_X7Y146_AO5;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_D5 = CLBLM_R_X5Y144_SLICE_X7Y144_AQ;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_D6 = CLBLM_R_X3Y150_SLICE_X2Y150_BO6;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_A5 = CLBLM_R_X7Y155_SLICE_X8Y155_BO5;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_A6 = CLBLM_R_X7Y153_SLICE_X8Y153_BQ;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_B1 = CLBLM_L_X10Y156_SLICE_X12Y156_CO6;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_B2 = CLBLM_R_X7Y154_SLICE_X8Y154_BQ;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_A1 = CLBLM_R_X7Y147_SLICE_X8Y147_B5Q;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_A2 = CLBLM_R_X5Y147_SLICE_X7Y147_AQ;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_A3 = CLBLM_R_X5Y144_SLICE_X6Y144_AQ;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_A6 = CLBLM_R_X7Y147_SLICE_X8Y147_C5Q;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_C2 = CLBLM_R_X7Y154_SLICE_X8Y154_CQ;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_C3 = CLBLM_R_X5Y152_SLICE_X6Y152_AQ;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_B1 = CLBLM_R_X7Y147_SLICE_X8Y147_B5Q;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_A1 = CLBLL_L_X2Y154_SLICE_X1Y154_BO6;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_A2 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_A3 = CLBLL_L_X2Y152_SLICE_X1Y152_CO6;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_A4 = CLBLL_L_X4Y152_SLICE_X5Y152_BO6;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_A5 = CLBLL_L_X2Y153_SLICE_X1Y153_CO6;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_A6 = CLBLL_L_X4Y153_SLICE_X4Y153_CO6;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_B2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_B3 = CLBLM_R_X7Y147_SLICE_X8Y147_C5Q;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_B4 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_B1 = LIOB33_X0Y67_IOB_X0Y67_I;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_B2 = CLBLL_L_X2Y151_SLICE_X0Y151_BO6;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_B3 = CLBLL_L_X2Y151_SLICE_X0Y151_AO6;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_B4 = CLBLL_L_X4Y152_SLICE_X5Y152_BO6;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_B5 = CLBLM_R_X3Y150_SLICE_X3Y150_BQ;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_B6 = CLBLL_L_X4Y153_SLICE_X4Y153_CO6;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_C1 = CLBLM_R_X3Y149_SLICE_X3Y149_B5Q;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_C2 = CLBLL_L_X4Y145_SLICE_X4Y145_A5Q;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_C1 = CLBLL_L_X2Y151_SLICE_X0Y151_CO5;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_C2 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_C3 = CLBLL_L_X2Y152_SLICE_X1Y152_AO5;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_C4 = CLBLL_L_X2Y154_SLICE_X1Y154_BO5;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_C5 = LIOB33_X0Y67_IOB_X0Y67_I;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_C6 = CLBLM_R_X3Y150_SLICE_X3Y150_BQ;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_D1 = CLBLL_L_X4Y148_SLICE_X4Y148_C5Q;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_D2 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_D3 = CLBLM_R_X5Y152_SLICE_X7Y152_B5Q;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_D4 = CLBLM_R_X5Y144_SLICE_X6Y144_CO6;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_D5 = CLBLM_R_X3Y145_SLICE_X3Y145_A5Q;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_D6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_D1 = CLBLL_L_X2Y155_SLICE_X1Y155_AO6;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_D2 = CLBLL_L_X4Y151_SLICE_X5Y151_CO6;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_D3 = CLBLL_L_X2Y152_SLICE_X1Y152_BO5;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_D4 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_D5 = CLBLL_L_X2Y152_SLICE_X1Y152_DO6;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_D6 = CLBLL_L_X2Y153_SLICE_X1Y153_BO6;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_B5 = CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_B6 = CLBLM_R_X11Y145_SLICE_X14Y145_AQ;
  assign RIOB33_X105Y153_IOB_X1Y154_O = RIOB33_X105Y101_IOB_X1Y102_I;
  assign RIOB33_X105Y153_IOB_X1Y153_O = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_C2 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_C5 = CLBLM_R_X7Y143_SLICE_X8Y143_DO6;
  assign LIOB33_X0Y185_IOB_X0Y186_O = RIOB33_X105Y143_IOB_X1Y143_I;
  assign LIOB33_X0Y185_IOB_X0Y185_O = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_A1 = CLBLM_R_X5Y155_SLICE_X7Y155_CO6;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_A2 = CLBLM_L_X8Y153_SLICE_X10Y153_AQ;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_A3 = CLBLM_R_X7Y155_SLICE_X9Y155_AQ;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_A4 = CLBLM_R_X7Y155_SLICE_X8Y155_BO5;
  assign CLBLL_L_X2Y154_SLICE_X0Y154_A1 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X0Y154_A2 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X0Y154_A3 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X0Y154_A4 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X0Y154_A5 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X0Y154_A6 = 1'b1;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_A6 = CLBLM_R_X5Y152_SLICE_X6Y152_CQ;
  assign CLBLL_L_X2Y154_SLICE_X0Y154_B1 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X0Y154_B2 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X0Y154_B3 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X0Y154_B4 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X0Y154_B5 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X0Y154_B6 = 1'b1;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_A1 = CLBLM_R_X5Y145_SLICE_X7Y145_DO6;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_A2 = CLBLM_R_X5Y148_SLICE_X6Y148_BQ;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_A3 = CLBLM_R_X5Y145_SLICE_X7Y145_AQ;
  assign CLBLL_L_X2Y154_SLICE_X0Y154_C1 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X0Y154_C2 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X0Y154_C3 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X0Y154_C4 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X0Y154_C5 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X0Y154_C6 = 1'b1;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_A4 = CLBLM_R_X11Y146_SLICE_X14Y146_AQ;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_A5 = CLBLM_R_X7Y145_SLICE_X8Y145_AQ;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_B1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_B2 = CLBLM_R_X5Y145_SLICE_X7Y145_BQ;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_B4 = CLBLM_R_X5Y147_SLICE_X7Y147_D5Q;
  assign CLBLL_L_X2Y154_SLICE_X0Y154_D1 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X0Y154_D2 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X0Y154_D3 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X0Y154_D4 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X0Y154_D5 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X0Y154_D6 = 1'b1;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_C2 = CLBLM_L_X8Y148_SLICE_X10Y148_CO6;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_C3 = CLBLM_R_X5Y145_SLICE_X7Y145_BQ;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_C4 = CLBLM_R_X5Y147_SLICE_X7Y147_CQ;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_C5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_C6 = 1'b1;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_D1 = CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_D2 = CLBLM_R_X7Y147_SLICE_X8Y147_AQ;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_D3 = CLBLL_L_X4Y145_SLICE_X4Y145_CQ;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_D4 = 1'b1;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_D5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_D6 = 1'b1;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_A6 = 1'b1;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_B1 = CLBLM_R_X5Y155_SLICE_X7Y155_BO5;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_B2 = CLBLM_R_X7Y155_SLICE_X8Y155_A5Q;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_B3 = CLBLM_R_X7Y153_SLICE_X8Y153_CQ;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_A1 = CLBLM_R_X5Y146_SLICE_X7Y146_AO5;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_A2 = CLBLM_R_X5Y145_SLICE_X7Y145_CQ;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_A4 = 1'b1;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_A6 = CLBLM_R_X5Y145_SLICE_X6Y145_A5Q;
  assign CLBLL_L_X2Y154_SLICE_X1Y154_A1 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y154_SLICE_X1Y154_A2 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y154_SLICE_X1Y154_A3 = CLBLL_L_X2Y152_SLICE_X1Y152_AO6;
  assign CLBLL_L_X2Y154_SLICE_X1Y154_A4 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y154_SLICE_X1Y154_A5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y154_SLICE_X1Y154_A6 = 1'b1;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_AX = CLBLM_R_X5Y145_SLICE_X6Y145_BO6;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_B1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_B2 = CLBLM_L_X10Y146_SLICE_X13Y146_AQ;
  assign CLBLL_L_X2Y154_SLICE_X1Y154_B1 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y154_SLICE_X1Y154_B2 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y154_SLICE_X1Y154_B3 = CLBLL_L_X2Y152_SLICE_X1Y152_AO6;
  assign CLBLL_L_X2Y154_SLICE_X1Y154_B4 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y154_SLICE_X1Y154_B5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y154_SLICE_X1Y154_B6 = 1'b1;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_B4 = CLBLL_L_X4Y145_SLICE_X5Y145_AQ;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_B5 = CLBLL_L_X4Y145_SLICE_X4Y145_BQ;
  assign CLBLL_L_X2Y154_SLICE_X1Y154_C1 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y154_SLICE_X1Y154_C2 = CLBLL_L_X2Y152_SLICE_X1Y152_AO5;
  assign CLBLL_L_X2Y154_SLICE_X1Y154_C3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y154_SLICE_X1Y154_C4 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y154_SLICE_X1Y154_C5 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y154_SLICE_X1Y154_C6 = 1'b1;
  assign CLBLM_L_X12Y154_SLICE_X17Y154_C4 = 1'b1;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_B6 = 1'b1;
  assign CLBLM_L_X12Y154_SLICE_X17Y154_C5 = 1'b1;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_C6 = 1'b1;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_D1 = CLBLM_R_X3Y151_SLICE_X3Y151_AO6;
  assign CLBLM_L_X12Y154_SLICE_X17Y154_C6 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X1Y154_D1 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X1Y154_D2 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X1Y154_D3 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X1Y154_D4 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X1Y154_D5 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X1Y154_D6 = 1'b1;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_D2 = CLBLL_L_X2Y151_SLICE_X1Y151_BO6;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_D3 = CLBLM_R_X3Y154_SLICE_X2Y154_BO6;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_D6 = 1'b1;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_C2 = CLBLM_R_X5Y145_SLICE_X6Y145_CQ;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_C3 = CLBLM_R_X5Y148_SLICE_X7Y148_CQ;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_C4 = CLBLM_R_X5Y147_SLICE_X7Y147_CQ;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_C5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign LIOI3_X0Y175_OLOGIC_X0Y176_D1 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign LIOI3_X0Y175_OLOGIC_X0Y176_T1 = 1'b1;
  assign CLBLM_L_X12Y154_SLICE_X17Y154_D5 = 1'b1;
  assign LIOI3_X0Y115_OLOGIC_X0Y116_D1 = CLBLM_L_X8Y142_SLICE_X10Y142_AQ;
  assign LIOI3_SING_X0Y199_OLOGIC_X0Y199_D1 = LIOB33_X0Y73_IOB_X0Y74_I;
  assign CLBLM_L_X12Y154_SLICE_X17Y154_D6 = 1'b1;
  assign LIOI3_X0Y175_OLOGIC_X0Y175_D1 = RIOB33_X105Y127_IOB_X1Y127_I;
  assign LIOI3_X0Y115_OLOGIC_X0Y116_T1 = 1'b1;
  assign RIOI3_X105Y159_OLOGIC_X1Y160_D1 = CLBLM_R_X11Y151_SLICE_X14Y151_DO5;
  assign LIOI3_X0Y175_OLOGIC_X0Y175_T1 = 1'b1;
  assign LIOI3_X0Y115_OLOGIC_X0Y115_D1 = CLBLM_R_X11Y148_SLICE_X15Y148_BQ;
  assign RIOI3_X105Y159_OLOGIC_X1Y160_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_D1 = RIOB33_X105Y145_IOB_X1Y145_I;
  assign LIOI3_X0Y115_OLOGIC_X0Y115_T1 = 1'b1;
  assign CLBLM_L_X10Y156_SLICE_X13Y156_B3 = 1'b1;
  assign RIOI3_X105Y159_OLOGIC_X1Y159_D1 = CLBLM_R_X11Y151_SLICE_X14Y151_DO6;
  assign CLBLM_L_X10Y156_SLICE_X13Y156_B4 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_T1 = 1'b1;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_D4 = CLBLM_R_X3Y150_SLICE_X2Y150_BO6;
  assign CLBLM_L_X10Y156_SLICE_X13Y156_B5 = 1'b1;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_D5 = CLBLM_R_X5Y147_SLICE_X6Y147_DO6;
  assign RIOI3_X105Y159_OLOGIC_X1Y159_T1 = 1'b1;
  assign CLBLM_L_X10Y156_SLICE_X13Y156_B6 = 1'b1;
  assign RIOB33_X105Y155_IOB_X1Y155_O = RIOB33_X105Y103_IOB_X1Y103_I;
  assign RIOB33_X105Y155_IOB_X1Y156_O = RIOB33_X105Y103_IOB_X1Y104_I;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_D1 = RIOB33_X105Y143_IOB_X1Y144_I;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_T1 = 1'b1;
  assign CLBLM_L_X10Y156_SLICE_X13Y156_C1 = 1'b1;
  assign CLBLM_L_X10Y156_SLICE_X13Y156_C2 = 1'b1;
  assign CLBLM_L_X10Y156_SLICE_X13Y156_C3 = 1'b1;
  assign CLBLM_L_X10Y156_SLICE_X13Y156_C4 = 1'b1;
  assign CLBLM_L_X10Y156_SLICE_X13Y156_C5 = 1'b1;
  assign LIOB33_X0Y187_IOB_X0Y188_O = RIOB33_X105Y145_IOB_X1Y145_I;
  assign LIOB33_X0Y187_IOB_X0Y187_O = RIOB33_X105Y143_IOB_X1Y144_I;
  assign CLBLM_L_X10Y156_SLICE_X13Y156_C6 = 1'b1;
  assign CLBLM_L_X12Y154_SLICE_X16Y154_B5 = CLBLM_R_X11Y154_SLICE_X15Y154_BQ;
  assign CLBLM_L_X12Y154_SLICE_X16Y154_B6 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_A1 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_A2 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_A3 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_A4 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_A5 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_A6 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_B1 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_B2 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_B3 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_B4 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_B5 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_B6 = 1'b1;
  assign CLBLM_L_X10Y156_SLICE_X13Y156_D1 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_C1 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_C2 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_C3 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_C4 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_C5 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_C6 = 1'b1;
  assign CLBLM_L_X10Y156_SLICE_X13Y156_D2 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_A1 = CLBLL_L_X4Y149_SLICE_X5Y149_DQ;
  assign CLBLM_L_X10Y156_SLICE_X13Y156_D3 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_A2 = CLBLM_R_X5Y148_SLICE_X6Y148_BQ;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_A3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_A4 = CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_A5 = CLBLL_L_X4Y148_SLICE_X4Y148_CQ;
  assign CLBLM_L_X10Y156_SLICE_X13Y156_D4 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_D1 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_D2 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_D3 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_D4 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_D5 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_D6 = 1'b1;
  assign CLBLM_L_X10Y156_SLICE_X13Y156_D5 = 1'b1;
  assign CLBLM_L_X12Y154_SLICE_X16Y154_C4 = 1'b1;
  assign CLBLM_L_X10Y156_SLICE_X13Y156_D6 = 1'b1;
  assign CLBLM_L_X12Y154_SLICE_X16Y154_C5 = 1'b1;
  assign CLBLM_L_X12Y154_SLICE_X16Y154_C6 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_C1 = CLBLM_R_X5Y145_SLICE_X7Y145_AQ;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_C2 = CLBLM_L_X10Y147_SLICE_X12Y147_AQ;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_C3 = CLBLM_R_X11Y147_SLICE_X14Y147_BQ;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_C4 = CLBLM_R_X7Y145_SLICE_X8Y145_AQ;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_C5 = CLBLL_L_X4Y146_SLICE_X5Y146_BO5;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_C6 = CLBLM_R_X5Y145_SLICE_X7Y145_DO5;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_D1 = CLBLM_R_X5Y146_SLICE_X7Y146_AO6;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_D2 = CLBLM_R_X3Y153_SLICE_X2Y153_DO6;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_D3 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_D4 = CLBLM_R_X5Y144_SLICE_X7Y144_AQ;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_D5 = CLBLM_L_X10Y144_SLICE_X13Y144_AQ;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_D6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_A1 = CLBLL_L_X4Y149_SLICE_X5Y149_BO5;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_A1 = CLBLL_L_X2Y154_SLICE_X1Y154_CO6;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_A2 = CLBLL_L_X2Y154_SLICE_X1Y154_AO6;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_A3 = CLBLL_L_X2Y154_SLICE_X1Y154_CO5;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_A4 = CLBLM_R_X3Y155_SLICE_X3Y155_AO6;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_A5 = CLBLL_L_X4Y154_SLICE_X5Y154_CO6;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_A6 = CLBLM_L_X16Y158_SLICE_X22Y158_AO5;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_A3 = CLBLM_R_X5Y146_SLICE_X6Y146_AQ;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_A4 = CLBLM_R_X7Y146_SLICE_X9Y146_CQ;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_A5 = CLBLM_R_X3Y151_SLICE_X3Y151_AO6;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_B1 = CLBLL_L_X2Y154_SLICE_X1Y154_CO6;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_B2 = CLBLL_L_X2Y154_SLICE_X1Y154_AO6;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_B3 = CLBLM_R_X3Y156_SLICE_X2Y156_CO6;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_B4 = CLBLM_R_X3Y155_SLICE_X3Y155_AO6;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_B5 = CLBLL_L_X4Y154_SLICE_X5Y154_CO6;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_B6 = CLBLL_L_X2Y155_SLICE_X1Y155_CO6;
  assign CLBLM_L_X10Y156_SLICE_X12Y156_A1 = CLBLM_L_X8Y155_SLICE_X11Y155_DO6;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_B1 = CLBLM_L_X10Y146_SLICE_X12Y146_CQ;
  assign CLBLM_L_X10Y156_SLICE_X12Y156_A2 = CLBLM_L_X8Y155_SLICE_X10Y155_AQ;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_C1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_C2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_C3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_C4 = CLBLL_L_X2Y152_SLICE_X1Y152_AO5;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_C5 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_C6 = CLBLM_L_X16Y158_SLICE_X22Y158_AO5;
  assign CLBLM_L_X10Y156_SLICE_X12Y156_A3 = CLBLM_L_X10Y154_SLICE_X12Y154_DQ;
  assign CLBLM_L_X10Y156_SLICE_X12Y156_A4 = CLBLM_L_X10Y155_SLICE_X13Y155_BQ;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_C2 = CLBLM_R_X7Y146_SLICE_X8Y146_BO5;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_C4 = CLBLM_R_X5Y150_SLICE_X6Y150_BQ;
  assign CLBLM_L_X10Y156_SLICE_X12Y156_A5 = CLBLM_L_X10Y155_SLICE_X13Y155_CQ;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_D1 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_D2 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_D3 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_D4 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_D5 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_D6 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLM_L_X10Y156_SLICE_X12Y156_A6 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_D2 = CLBLM_R_X5Y146_SLICE_X7Y146_AO6;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_D3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_D4 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_D5 = CLBLM_R_X7Y146_SLICE_X9Y146_AQ;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_D6 = CLBLM_R_X5Y151_SLICE_X7Y151_AQ;
  assign LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y70_D = LIOB33_X0Y69_IOB_X0Y70_I;
  assign LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y69_D = LIOB33_X0Y69_IOB_X0Y69_I;
  assign RIOI3_X105Y171_OLOGIC_X1Y171_T1 = 1'b1;
  assign RIOB33_SING_X105Y199_IOB_X1Y199_O = CLBLM_L_X12Y155_SLICE_X17Y155_AQ;
  assign CLBLM_L_X10Y156_SLICE_X12Y156_B4 = CLBLM_L_X8Y155_SLICE_X10Y155_CO6;
  assign CLBLM_L_X10Y156_SLICE_X12Y156_B5 = CLBLM_L_X10Y156_SLICE_X12Y156_AO6;
  assign LIOI3_SING_X0Y199_OLOGIC_X0Y199_T1 = 1'b1;
  assign CLBLM_L_X10Y156_SLICE_X12Y156_B6 = CLBLM_L_X8Y153_SLICE_X10Y153_AQ;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_C3 = CLBLM_L_X10Y156_SLICE_X12Y156_CO6;
  assign RIOB33_X105Y157_IOB_X1Y158_O = CLBLL_L_X36Y146_SLICE_X54Y146_AO6;
  assign RIOB33_X105Y157_IOB_X1Y157_O = RIOB33_X105Y125_IOB_X1Y126_I;
  assign CLBLM_L_X10Y156_SLICE_X12Y156_C4 = CLBLM_L_X10Y155_SLICE_X13Y155_DO6;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_B1 = CLBLL_L_X4Y145_SLICE_X5Y145_AQ;
  assign CLBLM_L_X10Y156_SLICE_X12Y156_C5 = CLBLM_L_X10Y155_SLICE_X12Y155_AQ;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_B2 = CLBLM_R_X11Y152_SLICE_X15Y152_BQ;
  assign CLBLM_L_X10Y156_SLICE_X12Y156_C6 = CLBLM_L_X10Y155_SLICE_X13Y155_BQ;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_A5 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_A6 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_B6 = CLBLM_R_X11Y153_SLICE_X14Y153_CO6;
  assign LIOB33_X0Y189_IOB_X0Y190_O = RIOB33_X105Y147_IOB_X1Y147_I;
  assign LIOB33_X0Y189_IOB_X0Y189_O = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_C1 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_B1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_D1 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_C2 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_C3 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_C4 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_B4 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_C5 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_C6 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_B6 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_C4 = CLBLM_R_X7Y155_SLICE_X8Y155_A5Q;
  assign LIOI3_X0Y61_ILOGIC_X0Y62_D = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y157_SLICE_X9Y157_A1 = 1'b1;
  assign CLBLM_R_X7Y157_SLICE_X9Y157_A2 = 1'b1;
  assign CLBLM_R_X7Y157_SLICE_X9Y157_A3 = 1'b1;
  assign CLBLM_R_X7Y157_SLICE_X9Y157_A4 = 1'b1;
  assign CLBLM_R_X7Y157_SLICE_X9Y157_A5 = 1'b1;
  assign CLBLM_R_X7Y157_SLICE_X9Y157_A6 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_T1 = 1'b1;
  assign CLBLM_R_X7Y157_SLICE_X9Y157_B1 = 1'b1;
  assign CLBLM_R_X7Y157_SLICE_X9Y157_B2 = 1'b1;
  assign CLBLM_R_X7Y157_SLICE_X9Y157_B3 = 1'b1;
  assign CLBLM_R_X7Y157_SLICE_X9Y157_B4 = 1'b1;
  assign CLBLM_R_X7Y157_SLICE_X9Y157_B5 = 1'b1;
  assign CLBLM_R_X7Y157_SLICE_X9Y157_B6 = 1'b1;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_A1 = CLBLL_L_X4Y150_SLICE_X4Y150_B5Q;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_A2 = CLBLM_R_X15Y151_SLICE_X20Y151_AQ;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_A3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_A4 = CLBLM_R_X5Y144_SLICE_X7Y144_BQ;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_A6 = CLBLM_R_X3Y148_SLICE_X3Y148_AQ;
  assign CLBLM_R_X7Y157_SLICE_X9Y157_C1 = 1'b1;
  assign CLBLM_R_X7Y157_SLICE_X9Y157_C2 = 1'b1;
  assign CLBLM_R_X7Y157_SLICE_X9Y157_C3 = 1'b1;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_B1 = CLBLM_R_X5Y152_SLICE_X7Y152_DO5;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_B2 = CLBLM_R_X5Y147_SLICE_X7Y147_BQ;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_B4 = CLBLL_L_X4Y147_SLICE_X4Y147_CQ;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_B5 = CLBLM_L_X8Y143_SLICE_X11Y143_AQ;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_B6 = 1'b1;
  assign CLBLM_R_X7Y157_SLICE_X9Y157_D1 = 1'b1;
  assign CLBLM_R_X7Y157_SLICE_X9Y157_D2 = 1'b1;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_C2 = CLBLM_L_X8Y146_SLICE_X10Y146_BQ;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_C3 = CLBLM_R_X5Y146_SLICE_X6Y146_DQ;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_C4 = 1'b1;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_C5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_C6 = CLBLM_R_X7Y147_SLICE_X9Y147_CO5;
  assign CLBLM_R_X7Y157_SLICE_X9Y157_D3 = 1'b1;
  assign CLBLM_R_X7Y157_SLICE_X9Y157_D4 = 1'b1;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y157_SLICE_X8Y157_A1 = 1'b1;
  assign CLBLM_R_X7Y157_SLICE_X8Y157_A2 = 1'b1;
  assign CLBLM_R_X7Y157_SLICE_X8Y157_A3 = 1'b1;
  assign CLBLM_R_X7Y157_SLICE_X8Y157_A4 = 1'b1;
  assign CLBLM_R_X7Y157_SLICE_X8Y157_A5 = 1'b1;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_D1 = CLBLM_R_X7Y157_SLICE_X8Y157_AQ;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_D2 = CLBLL_L_X2Y147_SLICE_X1Y147_AQ;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_D3 = CLBLM_R_X7Y148_SLICE_X8Y148_D5Q;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_D4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_D5 = CLBLM_L_X8Y153_SLICE_X10Y153_AQ;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_D6 = 1'b1;
  assign CLBLM_R_X7Y157_SLICE_X8Y157_A6 = 1'b1;
  assign CLBLM_R_X7Y157_SLICE_X8Y157_AX = CLBLM_R_X11Y157_SLICE_X14Y157_AO6;
  assign CLBLM_R_X7Y157_SLICE_X8Y157_B1 = 1'b1;
  assign CLBLM_R_X7Y157_SLICE_X8Y157_B2 = 1'b1;
  assign CLBLM_R_X7Y157_SLICE_X8Y157_B3 = 1'b1;
  assign CLBLM_R_X7Y157_SLICE_X8Y157_B4 = 1'b1;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_A1 = CLBLM_L_X10Y147_SLICE_X13Y147_BQ;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_A2 = CLBLM_R_X7Y151_SLICE_X9Y151_CQ;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_A3 = CLBLM_R_X5Y147_SLICE_X6Y147_AQ;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_A5 = CLBLM_R_X5Y152_SLICE_X7Y152_DO6;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_A6 = 1'b1;
  assign CLBLM_R_X7Y157_SLICE_X8Y157_C1 = 1'b1;
  assign CLBLM_R_X7Y157_SLICE_X8Y157_C2 = 1'b1;
  assign CLBLM_R_X7Y157_SLICE_X8Y157_C3 = 1'b1;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_B1 = 1'b1;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_B2 = CLBLM_R_X5Y147_SLICE_X6Y147_BQ;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_B3 = CLBLM_L_X12Y144_SLICE_X16Y144_AQ;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_B4 = CLBLM_R_X5Y152_SLICE_X7Y152_DO5;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_B5 = CLBLL_L_X4Y148_SLICE_X4Y148_BQ;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y157_SLICE_X8Y157_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y157_SLICE_X8Y157_D1 = 1'b1;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_C2 = CLBLM_R_X7Y147_SLICE_X8Y147_B5Q;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_C3 = CLBLM_R_X5Y145_SLICE_X6Y145_BO5;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_C5 = CLBLL_L_X4Y148_SLICE_X4Y148_BQ;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_C6 = 1'b1;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_B5 = CLBLM_R_X7Y155_SLICE_X8Y155_BO5;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_B6 = CLBLM_R_X11Y154_SLICE_X14Y154_AQ;
  assign CLBLM_R_X7Y157_SLICE_X8Y157_D4 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_A6 = 1'b1;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_A2 = CLBLM_R_X11Y152_SLICE_X14Y152_DQ;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_A3 = CLBLM_R_X11Y152_SLICE_X14Y152_AQ;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_D1 = CLBLM_R_X7Y157_SLICE_X8Y157_AQ;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_D2 = CLBLM_L_X16Y158_SLICE_X22Y158_AO5;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_D3 = CLBLM_R_X3Y152_SLICE_X3Y152_CO6;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_D4 = CLBLL_L_X4Y154_SLICE_X4Y154_CO6;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_D5 = CLBLL_L_X2Y153_SLICE_X1Y153_DO6;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_D6 = CLBLM_R_X3Y153_SLICE_X2Y153_DO6;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_A5 = CLBLM_R_X7Y152_SLICE_X8Y152_DQ;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_A6 = CLBLM_R_X11Y153_SLICE_X14Y153_BO5;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_C5 = CLBLM_R_X5Y155_SLICE_X7Y155_BO5;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_C1 = CLBLM_R_X7Y153_SLICE_X9Y153_AQ;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_C2 = CLBLM_R_X7Y153_SLICE_X8Y153_CQ;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_C3 = CLBLM_R_X5Y155_SLICE_X7Y155_BO5;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_C4 = CLBLM_R_X7Y155_SLICE_X8Y155_A5Q;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_C5 = CLBLL_L_X4Y147_SLICE_X5Y147_B5Q;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_C6 = CLBLM_R_X7Y154_SLICE_X8Y154_BQ;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_B4 = CLBLM_R_X11Y154_SLICE_X15Y154_CO6;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_B5 = CLBLM_L_X10Y152_SLICE_X13Y152_BQ;
  assign LIOB33_X0Y183_IOB_X0Y184_O = RIOB33_X105Y135_IOB_X1Y136_I;
  assign LIOB33_X0Y183_IOB_X0Y183_O = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_B6 = CLBLM_R_X11Y152_SLICE_X14Y152_BQ;
  assign RIOB33_X105Y159_IOB_X1Y160_O = CLBLM_R_X11Y151_SLICE_X14Y151_DO5;
  assign RIOB33_X105Y159_IOB_X1Y159_O = CLBLM_R_X11Y151_SLICE_X14Y151_DO6;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_D1 = CLBLM_R_X7Y153_SLICE_X9Y153_AQ;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_D2 = CLBLM_R_X7Y155_SLICE_X8Y155_A5Q;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_D3 = CLBLM_R_X7Y153_SLICE_X9Y153_CO5;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_D4 = CLBLM_R_X7Y153_SLICE_X8Y153_CQ;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_C4 = CLBLM_R_X11Y154_SLICE_X15Y154_CO6;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_D5 = CLBLL_L_X4Y147_SLICE_X5Y147_B5Q;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_C5 = CLBLM_R_X11Y153_SLICE_X14Y153_BO5;
  assign LIOB33_X0Y191_IOB_X0Y191_O = RIOB33_X105Y147_IOB_X1Y148_I;
  assign LIOB33_X0Y191_IOB_X0Y192_O = LIOB33_X0Y51_IOB_X0Y52_I;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_D6 = CLBLM_R_X7Y154_SLICE_X8Y154_BQ;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_C6 = CLBLM_R_X7Y153_SLICE_X9Y153_DQ;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_C6 = CLBLM_R_X5Y153_SLICE_X6Y153_CO6;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_A1 = CLBLM_R_X5Y155_SLICE_X7Y155_CO6;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_A3 = CLBLM_R_X7Y154_SLICE_X8Y154_AQ;
  assign LIOI3_X0Y177_OLOGIC_X0Y178_D1 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_A4 = CLBLM_R_X7Y151_SLICE_X8Y151_A5Q;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_D2 = CLBLM_R_X11Y154_SLICE_X15Y154_CO6;
  assign LIOI3_X0Y177_OLOGIC_X0Y178_T1 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_D3 = CLBLM_R_X11Y152_SLICE_X14Y152_DQ;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_D1 = CLBLM_R_X3Y147_SLICE_X3Y147_CQ;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_D4 = CLBLM_L_X10Y152_SLICE_X12Y152_BQ;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_D5 = CLBLM_R_X11Y153_SLICE_X14Y153_BO5;
  assign LIOI3_X0Y177_OLOGIC_X0Y177_D1 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_D6 = CLBLM_R_X11Y147_SLICE_X14Y147_BQ;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_T1 = 1'b1;
  assign RIOI3_X105Y161_OLOGIC_X1Y162_D1 = CLBLM_L_X10Y152_SLICE_X13Y152_CO5;
  assign LIOI3_X0Y177_OLOGIC_X0Y177_T1 = 1'b1;
  assign LIOI3_X0Y117_OLOGIC_X0Y117_D1 = CLBLM_R_X3Y144_SLICE_X2Y144_B5Q;
  assign RIOI3_X105Y161_OLOGIC_X1Y162_T1 = 1'b1;
  assign LIOI3_X0Y117_OLOGIC_X0Y117_T1 = 1'b1;
  assign RIOI3_X105Y161_OLOGIC_X1Y161_D1 = CLBLM_L_X10Y152_SLICE_X13Y152_CO6;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_B4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_A1 = 1'b1;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_A3 = CLBLM_R_X5Y148_SLICE_X7Y148_AQ;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_A5 = CLBLM_R_X7Y148_SLICE_X8Y148_AQ;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_A6 = CLBLM_R_X5Y150_SLICE_X7Y150_CO6;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_B5 = CLBLM_L_X8Y154_SLICE_X10Y154_BO6;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_B6 = CLBLM_R_X7Y150_SLICE_X8Y150_CQ;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_B1 = 1'b1;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_B2 = CLBLM_R_X7Y147_SLICE_X8Y147_CQ;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_B3 = 1'b1;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_B6 = CLBLM_R_X5Y155_SLICE_X6Y155_BQ;
  assign RIOI3_X105Y161_OLOGIC_X1Y161_T1 = 1'b1;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_C1 = CLBLM_R_X7Y148_SLICE_X8Y148_AQ;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_C2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_C3 = CLBLM_L_X10Y146_SLICE_X12Y146_DQ;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_C4 = CLBLL_L_X4Y150_SLICE_X5Y150_BQ;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_C5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_C6 = 1'b1;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_D1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_D2 = CLBLM_L_X10Y144_SLICE_X13Y144_AQ;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_D3 = 1'b1;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_D4 = CLBLM_R_X5Y144_SLICE_X7Y144_AQ;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_D5 = CLBLM_R_X7Y147_SLICE_X9Y147_CO6;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_D6 = CLBLM_R_X3Y154_SLICE_X2Y154_BO6;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_A1 = CLBLM_R_X7Y147_SLICE_X9Y147_CO6;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_A2 = CLBLM_R_X5Y151_SLICE_X6Y151_CQ;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_A3 = 1'b1;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_A4 = CLBLM_R_X5Y149_SLICE_X7Y149_BQ;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_A6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_C4 = 1'b1;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_B1 = 1'b1;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_B2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_B3 = CLBLM_R_X5Y148_SLICE_X7Y148_C5Q;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_B4 = 1'b1;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_B5 = CLBLM_R_X5Y150_SLICE_X6Y150_CQ;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_C5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_C6 = 1'b1;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_C1 = CLBLM_R_X7Y146_SLICE_X9Y146_AQ;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_C2 = CLBLM_R_X5Y148_SLICE_X6Y148_AQ;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_C4 = CLBLM_R_X5Y147_SLICE_X6Y147_CQ;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_C5 = CLBLM_R_X5Y146_SLICE_X6Y146_DQ;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_C6 = CLBLM_R_X5Y151_SLICE_X6Y151_CQ;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_D1 = CLBLL_L_X4Y148_SLICE_X4Y148_BQ;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_D2 = CLBLM_R_X5Y145_SLICE_X7Y145_CQ;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_D3 = 1'b1;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_D4 = 1'b1;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_D5 = CLBLM_R_X5Y147_SLICE_X7Y147_CQ;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_D6 = CLBLM_R_X5Y149_SLICE_X7Y149_BQ;
  assign RIOB33_X105Y161_IOB_X1Y162_O = CLBLM_L_X10Y152_SLICE_X13Y152_CO5;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_D1 = CLBLM_R_X5Y153_SLICE_X6Y153_CO6;
  assign RIOB33_X105Y161_IOB_X1Y161_O = CLBLM_L_X10Y152_SLICE_X13Y152_CO6;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_D2 = CLBLM_R_X7Y155_SLICE_X8Y155_A5Q;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_D3 = CLBLL_L_X4Y147_SLICE_X5Y147_B5Q;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_D4 = CLBLM_R_X7Y153_SLICE_X8Y153_CQ;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_C1 = 1'b1;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_D5 = CLBLM_L_X10Y156_SLICE_X12Y156_CO6;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_D6 = CLBLM_R_X7Y154_SLICE_X8Y154_BQ;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_C2 = 1'b1;
  assign LIOB33_X0Y193_IOB_X0Y194_O = LIOB33_X0Y59_IOB_X0Y60_I;
  assign LIOB33_X0Y193_IOB_X0Y193_O = LIOB33_X0Y55_IOB_X0Y56_I;
  assign LIOI3_X0Y55_ILOGIC_X0Y56_D = LIOB33_X0Y55_IOB_X0Y56_I;
  assign LIOI3_X0Y55_ILOGIC_X0Y55_D = LIOB33_X0Y55_IOB_X0Y55_I;
  assign RIOI3_X105Y101_ILOGIC_X1Y102_D = RIOB33_X105Y101_IOB_X1Y102_I;
  assign RIOI3_X105Y101_ILOGIC_X1Y101_D = RIOB33_X105Y101_IOB_X1Y101_I;
  assign RIOI3_X105Y151_OLOGIC_X1Y152_T1 = 1'b1;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_A1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_A2 = CLBLM_R_X7Y149_SLICE_X9Y149_BO6;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_A3 = 1'b1;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_A4 = CLBLL_L_X4Y148_SLICE_X5Y148_BQ;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_A6 = CLBLL_L_X4Y147_SLICE_X4Y147_BQ;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_B1 = CLBLL_L_X4Y146_SLICE_X4Y146_CO5;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_B2 = CLBLM_R_X5Y151_SLICE_X7Y151_BQ;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_B3 = 1'b1;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_B4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_B5 = CLBLM_R_X5Y147_SLICE_X6Y147_CQ;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_C2 = CLBLM_R_X5Y149_SLICE_X7Y149_CQ;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_C3 = CLBLM_R_X7Y149_SLICE_X8Y149_DQ;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_C4 = 1'b1;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_C5 = 1'b1;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_C6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_D1 = CLBLL_L_X4Y149_SLICE_X5Y149_A5Q;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_D2 = CLBLM_R_X3Y150_SLICE_X2Y150_BO6;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_D3 = CLBLM_R_X5Y144_SLICE_X7Y144_AQ;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_D4 = 1'b1;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_D5 = CLBLM_L_X10Y144_SLICE_X13Y144_AQ;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_D6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_A1 = CLBLM_R_X5Y149_SLICE_X6Y149_DO6;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_A2 = CLBLM_L_X10Y151_SLICE_X13Y151_AQ;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_A3 = CLBLM_R_X5Y149_SLICE_X6Y149_AQ;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_A6 = CLBLM_R_X5Y148_SLICE_X6Y148_CO6;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_B1 = CLBLM_L_X10Y148_SLICE_X13Y148_BQ;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_B2 = CLBLM_R_X5Y149_SLICE_X6Y149_BQ;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_B3 = CLBLM_L_X10Y149_SLICE_X13Y149_BQ;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_B4 = CLBLM_R_X5Y152_SLICE_X7Y152_DO5;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_B5 = 1'b1;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_C1 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_C2 = CLBLM_R_X5Y154_SLICE_X6Y154_BO6;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_C3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_C4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_C5 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_C6 = 1'b1;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_D1 = CLBLM_R_X5Y145_SLICE_X6Y145_AQ;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_D2 = CLBLM_L_X10Y150_SLICE_X13Y150_CQ;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_D3 = CLBLM_L_X10Y145_SLICE_X12Y145_CQ;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_D4 = CLBLM_R_X5Y148_SLICE_X6Y148_DO6;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_D5 = CLBLM_R_X7Y151_SLICE_X8Y151_DO6;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_D6 = CLBLM_R_X5Y151_SLICE_X6Y151_BQ;
  assign RIOB33_X105Y163_IOB_X1Y163_O = CLBLM_L_X10Y150_SLICE_X13Y150_DO6;
  assign RIOB33_X105Y163_IOB_X1Y164_O = CLBLM_L_X10Y150_SLICE_X13Y150_DO5;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_T1 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_A6 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_B1 = CLBLM_R_X5Y143_SLICE_X7Y143_BO5;
  assign LIOB33_X0Y195_IOB_X0Y196_O = LIOB33_X0Y69_IOB_X0Y69_I;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_B2 = CLBLL_L_X2Y151_SLICE_X1Y151_BO6;
  assign LIOB33_X0Y195_IOB_X0Y195_O = LIOB33_X0Y63_IOB_X0Y64_I;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_B3 = CLBLM_R_X3Y151_SLICE_X3Y151_AO6;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_B4 = CLBLM_R_X3Y150_SLICE_X2Y150_BO6;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_B5 = CLBLM_R_X5Y146_SLICE_X7Y146_CO6;
  assign LIOI3_X0Y53_ILOGIC_X0Y54_D = LIOB33_X0Y53_IOB_X0Y54_I;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_D1 = CLBLM_R_X11Y151_SLICE_X14Y151_DO5;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_B6 = CLBLL_L_X4Y154_SLICE_X4Y154_CO6;
  assign LIOI3_X0Y111_OLOGIC_X0Y112_D1 = CLBLM_R_X11Y148_SLICE_X15Y148_B5Q;
  assign LIOB33_X0Y161_IOB_X0Y162_O = RIOB33_X105Y109_IOB_X1Y109_I;
  assign LIOB33_X0Y161_IOB_X0Y161_O = RIOB33_X105Y107_IOB_X1Y108_I;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_T1 = 1'b1;
  assign LIOI3_X0Y111_OLOGIC_X0Y112_T1 = 1'b1;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_D1 = 1'b0;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_A1 = CLBLM_L_X8Y149_SLICE_X11Y149_B5Q;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_A3 = CLBLM_L_X8Y153_SLICE_X10Y153_DO5;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_A4 = 1'b1;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_A5 = CLBLM_R_X5Y152_SLICE_X6Y152_AQ;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_A6 = 1'b1;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_B2 = 1'b1;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_B3 = 1'b1;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_B4 = CLBLM_R_X7Y147_SLICE_X8Y147_C5Q;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_B5 = CLBLM_R_X3Y150_SLICE_X3Y150_AQ;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_C1 = CLBLM_R_X3Y150_SLICE_X3Y150_AQ;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_C2 = 1'b1;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_C3 = CLBLL_L_X4Y150_SLICE_X5Y150_CO6;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_C4 = CLBLM_R_X7Y153_SLICE_X9Y153_A5Q;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_C5 = CLBLM_R_X7Y152_SLICE_X9Y152_DO6;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_C6 = CLBLM_R_X5Y150_SLICE_X7Y150_DO6;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_T1 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_D1 = CLBLM_R_X5Y149_SLICE_X7Y149_AQ;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_D2 = CLBLM_R_X7Y151_SLICE_X9Y151_CQ;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_D3 = 1'b1;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_D4 = CLBLM_R_X7Y153_SLICE_X9Y153_DQ;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_D5 = CLBLM_R_X7Y149_SLICE_X8Y149_AQ;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_D6 = CLBLL_L_X4Y147_SLICE_X4Y147_CQ;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_A1 = CLBLM_R_X7Y153_SLICE_X8Y153_BQ;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_A2 = CLBLM_R_X3Y150_SLICE_X2Y150_BO6;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_A3 = CLBLM_R_X3Y152_SLICE_X3Y152_CO6;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_A5 = CLBLM_L_X10Y144_SLICE_X13Y144_AQ;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_A6 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_AX = CLBLM_R_X5Y146_SLICE_X6Y146_BO6;
  assign LIOI3_X0Y179_OLOGIC_X0Y180_D1 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign RIOB33_X105Y165_IOB_X1Y165_O = RIOB33_X105Y125_IOB_X1Y125_I;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_B1 = CLBLM_R_X5Y150_SLICE_X6Y150_BQ;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_B2 = CLBLM_R_X3Y147_SLICE_X3Y147_BQ;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_B4 = CLBLM_L_X8Y148_SLICE_X10Y148_A5Q;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_B5 = CLBLM_R_X5Y149_SLICE_X7Y149_CQ;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_B6 = CLBLM_R_X11Y150_SLICE_X14Y150_AO6;
  assign RIOB33_X105Y165_IOB_X1Y166_O = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_B2 = CLBLM_R_X5Y146_SLICE_X6Y146_A5Q;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_C1 = CLBLM_R_X5Y150_SLICE_X7Y150_AQ;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_C2 = 1'b1;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_C3 = 1'b1;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_C4 = CLBLM_R_X7Y142_SLICE_X8Y142_CQ;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_B3 = CLBLM_R_X5Y150_SLICE_X6Y150_AQ;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_C6 = CLBLM_L_X8Y153_SLICE_X10Y153_DO5;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_D1 = CLBLM_R_X3Y144_SLICE_X2Y144_BQ;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_B4 = CLBLL_L_X4Y145_SLICE_X5Y145_CO6;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign LIOI3_X0Y179_OLOGIC_X0Y179_D1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_D1 = CLBLM_R_X5Y145_SLICE_X6Y145_AQ;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_D2 = 1'b1;
  assign CLBLM_L_X12Y155_SLICE_X17Y155_C4 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_B6 = 1'b1;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_D3 = CLBLM_R_X5Y150_SLICE_X6Y150_DQ;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_D4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_D5 = CLBLM_R_X5Y152_SLICE_X7Y152_DO6;
  assign CLBLM_L_X12Y155_SLICE_X17Y155_C5 = 1'b1;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_D6 = CLBLM_R_X5Y147_SLICE_X6Y147_AQ;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_D1 = CLBLM_L_X8Y142_SLICE_X10Y142_A5Q;
  assign LIOI3_X0Y179_OLOGIC_X0Y179_T1 = 1'b1;
  assign CLBLM_L_X12Y155_SLICE_X17Y155_C6 = 1'b1;
  assign RIOI3_X105Y165_OLOGIC_X1Y166_T1 = 1'b1;
  assign LIOB33_X0Y197_IOB_X0Y198_O = LIOB33_X0Y73_IOB_X0Y73_I;
  assign LIOB33_X0Y197_IOB_X0Y197_O = LIOB33_X0Y71_IOB_X0Y72_I;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_T1 = 1'b1;
  assign RIOI3_X105Y165_OLOGIC_X1Y165_D1 = RIOB33_X105Y125_IOB_X1Y125_I;
  assign RIOI3_X105Y165_OLOGIC_X1Y165_T1 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_C5 = CLBLM_L_X8Y146_SLICE_X10Y146_AQ;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_C6 = 1'b1;
  assign CLBLM_L_X12Y155_SLICE_X17Y155_D2 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y155_SLICE_X17Y155_D5 = 1'b1;
  assign CLBLM_L_X12Y155_SLICE_X17Y155_D6 = 1'b1;
  assign CLBLM_L_X12Y155_SLICE_X16Y155_A1 = 1'b1;
  assign LIOI3_X0Y173_OLOGIC_X0Y174_D1 = CLBLM_L_X8Y159_SLICE_X10Y159_AO6;
  assign LIOI3_X0Y59_ILOGIC_X0Y60_D = LIOB33_X0Y59_IOB_X0Y60_I;
  assign CLBLM_L_X12Y155_SLICE_X16Y155_B6 = 1'b1;
  assign LIOI3_X0Y59_ILOGIC_X0Y59_D = LIOB33_X0Y59_IOB_X0Y59_I;
  assign LIOB33_X0Y79_IOB_X0Y80_O = CLBLL_L_X2Y138_SLICE_X0Y138_AO6;
  assign RIOI3_X105Y103_ILOGIC_X1Y104_D = RIOB33_X105Y103_IOB_X1Y104_I;
  assign RIOI3_X105Y103_ILOGIC_X1Y103_D = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_A1 = CLBLM_L_X10Y155_SLICE_X12Y155_AQ;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_A2 = CLBLL_L_X4Y151_SLICE_X4Y151_AQ;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_A3 = CLBLM_R_X5Y151_SLICE_X7Y151_AQ;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_A4 = CLBLM_L_X8Y149_SLICE_X11Y149_AQ;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_A5 = CLBLM_R_X7Y147_SLICE_X8Y147_AQ;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_B1 = 1'b1;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_B2 = CLBLM_R_X5Y151_SLICE_X7Y151_BQ;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_B4 = CLBLM_R_X5Y152_SLICE_X7Y152_DO5;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_B5 = CLBLL_L_X4Y147_SLICE_X4Y147_BQ;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_B6 = CLBLM_R_X7Y153_SLICE_X8Y153_AQ;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_A1 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_A2 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_A3 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_A4 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_A5 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_A6 = 1'b1;
  assign CLBLM_L_X12Y155_SLICE_X16Y155_C4 = 1'b1;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y155_SLICE_X16Y155_C5 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_B1 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_B2 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_B3 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_B4 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_B5 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_B6 = 1'b1;
  assign CLBLM_L_X12Y155_SLICE_X16Y155_C6 = 1'b1;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_C1 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_C2 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_C3 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_C4 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_C5 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_C6 = 1'b1;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_D3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_D4 = CLBLM_R_X5Y152_SLICE_X7Y152_BQ;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_A1 = 1'b1;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_A2 = CLBLM_R_X5Y147_SLICE_X6Y147_BQ;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_A3 = CLBLM_R_X5Y151_SLICE_X6Y151_AQ;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_A4 = CLBLM_R_X5Y152_SLICE_X7Y152_DO5;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_A6 = CLBLM_R_X5Y146_SLICE_X6Y146_DQ;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_D1 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_D2 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_D3 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_D4 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_D5 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_D6 = 1'b1;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_B1 = CLBLM_R_X5Y151_SLICE_X6Y151_CQ;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_B2 = 1'b1;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_B3 = 1'b1;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_B4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_B5 = CLBLL_L_X4Y148_SLICE_X5Y148_AQ;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_A1 = CLBLM_R_X3Y143_SLICE_X3Y143_A5Q;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_A2 = CLBLM_R_X3Y142_SLICE_X2Y142_BQ;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_A3 = CLBLM_R_X3Y142_SLICE_X2Y142_AQ;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_A4 = CLBLM_R_X3Y143_SLICE_X3Y143_BQ;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_A5 = CLBLL_L_X2Y145_SLICE_X1Y145_AQ;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_A6 = CLBLM_R_X3Y143_SLICE_X2Y143_CQ;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_C2 = 1'b1;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_C3 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_B1 = CLBLM_R_X3Y144_SLICE_X3Y144_BO5;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_B2 = CLBLM_R_X3Y150_SLICE_X2Y150_BO6;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_B3 = CLBLM_R_X3Y151_SLICE_X3Y151_AO6;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_B4 = CLBLM_R_X3Y152_SLICE_X3Y152_CO6;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_B5 = LIOB33_X0Y53_IOB_X0Y53_I;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_B6 = CLBLL_L_X4Y142_SLICE_X5Y142_AO5;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_D2 = CLBLL_L_X2Y151_SLICE_X1Y151_BO6;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_C1 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_C2 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_C3 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_C4 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_C5 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_C6 = 1'b1;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_D3 = CLBLM_R_X5Y151_SLICE_X6Y151_DQ;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_D4 = CLBLM_L_X8Y151_SLICE_X11Y151_BQ;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_D5 = CLBLL_L_X4Y149_SLICE_X5Y149_BO5;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_D6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_D1 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_D2 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_D3 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_D4 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_D5 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_D6 = 1'b1;
  assign LIOI3_X0Y173_OLOGIC_X0Y173_T1 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_C4 = CLBLM_R_X13Y152_SLICE_X18Y152_BO6;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_C5 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_C6 = 1'b1;
  assign RIOB33_X105Y169_IOB_X1Y170_O = CLBLM_R_X103Y170_SLICE_X163Y170_AO6;
  assign RIOB33_X105Y169_IOB_X1Y169_O = CLBLM_R_X103Y169_SLICE_X163Y169_AO6;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_A1 = CLBLM_R_X5Y152_SLICE_X7Y152_DO6;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_A2 = CLBLM_R_X5Y144_SLICE_X7Y144_CQ;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_A3 = CLBLM_R_X5Y152_SLICE_X7Y152_AQ;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_A4 = CLBLM_R_X5Y149_SLICE_X7Y149_AQ;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_A6 = 1'b1;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_B1 = CLBLM_R_X7Y153_SLICE_X8Y153_AQ;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_B2 = CLBLM_R_X3Y145_SLICE_X3Y145_CQ;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_B3 = CLBLM_R_X7Y154_SLICE_X8Y154_BQ;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_B5 = CLBLM_R_X7Y143_SLICE_X8Y143_CQ;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_B6 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_D2 = CLBLM_L_X10Y153_SLICE_X12Y153_BQ;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_A1 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_A2 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_A3 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_A4 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_A5 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_A6 = 1'b1;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_C2 = CLBLM_R_X5Y152_SLICE_X7Y152_CQ;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_C3 = CLBLM_L_X10Y153_SLICE_X12Y153_BQ;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_B1 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_B2 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_B3 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_B4 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_B5 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_B6 = 1'b1;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_C1 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_C2 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_C3 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_C4 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_C5 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_C6 = 1'b1;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_D3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_D4 = CLBLM_R_X5Y152_SLICE_X6Y152_CQ;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_A1 = 1'b1;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_A3 = CLBLM_R_X7Y152_SLICE_X9Y152_AQ;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_A4 = CLBLM_R_X3Y150_SLICE_X3Y150_BQ;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_A5 = 1'b1;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_A6 = CLBLM_L_X8Y153_SLICE_X10Y153_DO5;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_D1 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_D2 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_D3 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_D4 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_D5 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_D6 = 1'b1;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_AX = CLBLM_R_X5Y151_SLICE_X7Y151_DO5;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_B1 = 1'b1;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_B3 = 1'b1;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_B4 = CLBLM_R_X5Y150_SLICE_X6Y150_CQ;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_B5 = CLBLM_L_X8Y153_SLICE_X10Y153_DO5;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_A1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_A2 = CLBLM_R_X3Y145_SLICE_X3Y145_D5Q;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_A3 = CLBLM_R_X3Y142_SLICE_X2Y142_AQ;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_A4 = CLBLM_R_X3Y142_SLICE_X2Y142_DO5;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_A6 = CLBLM_R_X5Y149_SLICE_X6Y149_AQ;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_C3 = CLBLM_R_X11Y146_SLICE_X14Y146_DQ;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_C4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_C6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_B1 = CLBLM_R_X3Y143_SLICE_X3Y143_A5Q;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_B2 = CLBLM_R_X3Y142_SLICE_X2Y142_BQ;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_B3 = CLBLM_R_X3Y143_SLICE_X3Y143_CO5;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_B4 = CLBLL_L_X2Y145_SLICE_X1Y145_BQ;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_B6 = CLBLM_R_X3Y143_SLICE_X2Y143_CQ;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_D1 = CLBLL_L_X4Y154_SLICE_X5Y154_CO5;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_D2 = CLBLL_L_X2Y155_SLICE_X1Y155_DO6;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_C2 = CLBLM_R_X3Y142_SLICE_X2Y142_CQ;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_C3 = CLBLM_R_X3Y143_SLICE_X3Y143_DO5;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_C4 = CLBLM_R_X3Y148_SLICE_X3Y148_BQ;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_C5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_C6 = CLBLM_R_X3Y145_SLICE_X3Y145_D5Q;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_D3 = CLBLM_R_X7Y152_SLICE_X8Y152_CQ;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_D4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_D5 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_D6 = CLBLM_R_X7Y152_SLICE_X8Y152_BQ;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_A5 = CLBLM_L_X12Y151_SLICE_X16Y151_DO5;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_A6 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_D1 = CLBLM_R_X3Y142_SLICE_X2Y142_AQ;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_D2 = CLBLM_R_X3Y143_SLICE_X2Y143_CQ;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_D3 = CLBLM_R_X3Y143_SLICE_X3Y143_A5Q;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_D4 = CLBLM_R_X3Y142_SLICE_X2Y142_BQ;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_D5 = CLBLL_L_X2Y145_SLICE_X1Y145_AQ;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_D6 = 1'b1;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_C1 = CLBLM_R_X7Y153_SLICE_X8Y153_CQ;
  assign CLBLM_R_X13Y151_SLICE_X18Y151_D4 = 1'b1;
  assign CLBLM_R_X13Y151_SLICE_X18Y151_D5 = 1'b1;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_C2 = CLBLM_R_X7Y155_SLICE_X8Y155_A5Q;
  assign CLBLM_R_X13Y151_SLICE_X18Y151_D6 = 1'b1;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_C3 = CLBLL_L_X4Y147_SLICE_X5Y147_B5Q;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_C4 = CLBLM_R_X7Y155_SLICE_X8Y155_AQ;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_C5 = CLBLM_R_X7Y154_SLICE_X8Y154_BQ;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_C6 = CLBLM_R_X5Y152_SLICE_X6Y152_BQ;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_B4 = CLBLM_R_X11Y154_SLICE_X15Y154_AQ;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_B5 = CLBLM_L_X12Y151_SLICE_X16Y151_DO5;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_B6 = 1'b1;
  assign LIOI3_X0Y183_OLOGIC_X0Y184_D1 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_BX = CLBLM_R_X11Y154_SLICE_X15Y154_BQ;
  assign LIOI3_X0Y183_OLOGIC_X0Y184_T1 = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_D1 = CLBLM_R_X3Y147_SLICE_X3Y147_C5Q;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_D1 = 1'b1;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_D2 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_C2 = CLBLM_R_X11Y154_SLICE_X15Y154_BQ;
  assign LIOI3_X0Y183_OLOGIC_X0Y183_D1 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_D3 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_C3 = CLBLM_R_X11Y154_SLICE_X14Y154_BO5;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_T1 = 1'b1;
  assign RIOI3_X105Y167_OLOGIC_X1Y168_D1 = CLBLM_L_X8Y159_SLICE_X10Y159_AO6;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_D4 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_C4 = CLBLM_R_X11Y154_SLICE_X14Y154_AQ;
  assign LIOI3_X0Y183_OLOGIC_X0Y183_T1 = 1'b1;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_D5 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_C5 = CLBLM_R_X11Y152_SLICE_X15Y152_BQ;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_D1 = CLBLM_R_X7Y143_SLICE_X8Y143_B5Q;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_D6 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_C6 = 1'b1;
  assign RIOI3_X105Y167_OLOGIC_X1Y168_T1 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_CE = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_T1 = 1'b1;
  assign RIOI3_X105Y167_OLOGIC_X1Y167_D1 = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_D1 = CLBLM_R_X3Y152_SLICE_X2Y152_BO6;
  assign RIOI3_X105Y167_OLOGIC_X1Y167_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_T1 = 1'b1;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_A1 = CLBLM_R_X7Y155_SLICE_X8Y155_DO6;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_D1 = CLBLM_L_X10Y145_SLICE_X13Y145_AQ;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_B4 = 1'b1;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_A2 = CLBLL_L_X4Y154_SLICE_X5Y154_BQ;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_D1 = CLBLL_L_X2Y120_SLICE_X0Y120_AO6;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_CX = CLBLM_R_X5Y150_SLICE_X7Y150_BQ;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_B5 = 1'b1;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_B6 = 1'b1;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_A4 = CLBLM_L_X10Y150_SLICE_X12Y150_A5Q;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_D1 = CLBLM_R_X11Y153_SLICE_X14Y153_AO6;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_T1 = 1'b1;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_A5 = CLBLM_R_X7Y155_SLICE_X8Y155_CO6;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_D2 = CLBLM_R_X11Y154_SLICE_X14Y154_CO6;
  assign RIOB33_X105Y171_IOB_X1Y172_O = CLBLM_R_X103Y170_SLICE_X163Y170_AO5;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_D3 = CLBLM_R_X11Y154_SLICE_X14Y154_DO6;
  assign RIOB33_X105Y171_IOB_X1Y171_O = CLBLM_R_X11Y157_SLICE_X14Y157_AO5;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_D4 = CLBLM_L_X10Y154_SLICE_X13Y154_AQ;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_D5 = CLBLM_R_X7Y153_SLICE_X8Y153_DQ;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_D6 = CLBLM_R_X11Y153_SLICE_X15Y153_BQ;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_C3 = 1'b1;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_C4 = 1'b1;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_C5 = 1'b1;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_A1 = CLBLM_R_X7Y153_SLICE_X8Y153_CQ;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_C6 = 1'b1;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_A3 = CLBLL_L_X4Y142_SLICE_X5Y142_AQ;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_A4 = CLBLM_R_X7Y154_SLICE_X8Y154_BQ;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_A5 = CLBLL_L_X4Y147_SLICE_X5Y147_B5Q;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_A6 = CLBLM_R_X7Y155_SLICE_X8Y155_A5Q;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_B4 = CLBLL_L_X4Y147_SLICE_X5Y147_B5Q;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_B1 = CLBLM_R_X3Y144_SLICE_X2Y144_CO6;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_B2 = CLBLM_R_X5Y153_SLICE_X7Y153_BQ;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_B4 = CLBLM_R_X7Y154_SLICE_X9Y154_BQ;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_B5 = 1'b1;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_B6 = CLBLM_R_X3Y145_SLICE_X3Y145_A5Q;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_B5 = CLBLM_R_X7Y154_SLICE_X8Y154_BQ;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_B6 = 1'b1;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_A1 = CLBLM_L_X8Y155_SLICE_X10Y155_AQ;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_A2 = CLBLM_R_X3Y145_SLICE_X3Y145_D5Q;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_A3 = CLBLM_R_X3Y143_SLICE_X3Y143_AQ;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_A5 = CLBLM_R_X3Y141_SLICE_X2Y141_AO6;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_A6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_C1 = CLBLM_R_X7Y150_SLICE_X9Y150_AQ;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_C2 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_AX = CLBLM_R_X3Y143_SLICE_X3Y143_CO6;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_C3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_B1 = CLBLM_R_X3Y142_SLICE_X2Y142_DO6;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_B4 = CLBLM_R_X3Y145_SLICE_X3Y145_D5Q;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_B5 = CLBLM_R_X3Y143_SLICE_X3Y143_BQ;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_B6 = CLBLM_L_X8Y145_SLICE_X10Y145_A5Q;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_BX = CLBLM_R_X3Y143_SLICE_X3Y143_DO6;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_D1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_C2 = CLBLM_R_X3Y145_SLICE_X3Y145_D5Q;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_C3 = CLBLM_R_X5Y155_SLICE_X7Y155_AQ;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_C4 = CLBLM_R_X3Y143_SLICE_X3Y143_A5Q;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_C5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_C6 = 1'b1;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_D3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_D4 = CLBLL_L_X2Y155_SLICE_X1Y155_DO6;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_A1 = CLBLM_L_X8Y152_SLICE_X11Y152_BO6;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_A2 = 1'b1;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_A3 = CLBLM_R_X5Y153_SLICE_X6Y153_AQ;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_A5 = CLBLM_L_X8Y146_SLICE_X10Y146_AQ;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_D1 = CLBLM_R_X3Y143_SLICE_X3Y143_BQ;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_D2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_D3 = CLBLM_R_X3Y142_SLICE_X2Y142_DO6;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_D4 = CLBLM_R_X3Y146_SLICE_X3Y146_CQ;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_D5 = CLBLM_R_X3Y143_SLICE_X3Y143_AQ;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_D6 = 1'b1;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_A6 = CLBLM_R_X3Y145_SLICE_X3Y145_CQ;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_AX = CLBLM_R_X5Y153_SLICE_X6Y153_CO5;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_B1 = CLBLM_R_X3Y145_SLICE_X3Y145_DQ;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_B2 = CLBLM_R_X5Y153_SLICE_X6Y153_BQ;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_B3 = CLBLM_L_X10Y150_SLICE_X13Y150_CQ;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_A1 = CLBLM_R_X3Y144_SLICE_X2Y144_A5Q;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_A2 = CLBLM_R_X3Y143_SLICE_X3Y143_DO5;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_A3 = CLBLM_R_X3Y143_SLICE_X3Y143_CO5;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_A4 = CLBLM_R_X3Y143_SLICE_X2Y143_AQ;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_A6 = CLBLM_R_X3Y142_SLICE_X2Y142_CQ;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_C2 = CLBLL_L_X4Y145_SLICE_X5Y145_CO6;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_C3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_B1 = CLBLL_L_X4Y145_SLICE_X4Y145_CQ;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_B2 = CLBLM_R_X3Y143_SLICE_X3Y143_DO5;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_B3 = CLBLM_R_X3Y143_SLICE_X2Y143_AQ;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_B4 = CLBLM_R_X3Y145_SLICE_X3Y145_D5Q;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_B6 = CLBLM_R_X3Y142_SLICE_X2Y142_CQ;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_D1 = CLBLM_R_X7Y152_SLICE_X8Y152_AQ;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_D2 = CLBLM_R_X5Y153_SLICE_X7Y153_CO6;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_C2 = CLBLM_R_X3Y143_SLICE_X2Y143_CQ;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_C4 = CLBLM_R_X5Y143_SLICE_X6Y143_AQ;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_C5 = CLBLM_R_X3Y143_SLICE_X3Y143_A5Q;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_C6 = CLBLM_R_X3Y145_SLICE_X3Y145_D5Q;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_D3 = CLBLM_R_X5Y153_SLICE_X7Y153_DO6;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_D4 = CLBLL_L_X2Y154_SLICE_X1Y154_AO5;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_D5 = CLBLM_R_X5Y151_SLICE_X6Y151_DQ;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_D6 = CLBLM_R_X5Y154_SLICE_X7Y154_AO6;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign LIOI3_X0Y61_ILOGIC_X0Y61_D = LIOB33_X0Y61_IOB_X0Y61_I;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_D1 = 1'b1;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_D2 = CLBLM_R_X3Y143_SLICE_X2Y143_CQ;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_D3 = CLBLM_R_X3Y143_SLICE_X2Y143_DQ;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_D4 = CLBLM_R_X3Y144_SLICE_X2Y144_CO6;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_D5 = CLBLM_R_X3Y144_SLICE_X2Y144_A5Q;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_D6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y106_D = RIOB33_X105Y105_IOB_X1Y106_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y105_D = RIOB33_X105Y105_IOB_X1Y105_I;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_T1 = 1'b1;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_D1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_A1 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_A2 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_A3 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_A4 = RIOB33_X105Y123_IOB_X1Y124_I;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_A5 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_A6 = 1'b1;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_D2 = CLBLM_R_X7Y155_SLICE_X8Y155_AQ;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y114_D = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_D3 = CLBLM_L_X8Y153_SLICE_X10Y153_AQ;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_B1 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_B2 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_B3 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_B4 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_B5 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_B6 = 1'b1;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_D4 = CLBLM_R_X5Y155_SLICE_X7Y155_CO6;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_D = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_C1 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_C2 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_C3 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_C4 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_C5 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_C6 = 1'b1;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_D6 = CLBLM_R_X7Y155_SLICE_X8Y155_BO6;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_D1 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_D2 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_D3 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_D4 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_D5 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_D6 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_A1 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_A2 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_A3 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_A4 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_A5 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_A6 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_B1 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_B2 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_B3 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_B4 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_B5 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_B6 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_C1 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_C2 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_C3 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_C4 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_C5 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_C6 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_D1 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_D2 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_D3 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_D4 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_D5 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_D6 = 1'b1;
  assign RIOB33_X105Y173_IOB_X1Y174_O = CLBLM_R_X103Y173_SLICE_X163Y173_AO5;
  assign RIOB33_X105Y173_IOB_X1Y173_O = CLBLM_R_X103Y173_SLICE_X163Y173_AO6;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_C2 = CLBLM_R_X5Y152_SLICE_X6Y152_CQ;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_A1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_A2 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_A3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_A4 = CLBLL_L_X2Y155_SLICE_X1Y155_DO6;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_A5 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_A6 = 1'b1;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_B1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_B2 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_B3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_B4 = CLBLL_L_X4Y148_SLICE_X5Y148_AQ;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_B5 = CLBLM_R_X5Y151_SLICE_X7Y151_CQ;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_B6 = CLBLM_R_X5Y154_SLICE_X7Y154_CO6;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_A1 = CLBLM_R_X11Y146_SLICE_X15Y146_AQ;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_A2 = CLBLM_R_X7Y144_SLICE_X9Y144_DO6;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_A3 = CLBLM_R_X3Y144_SLICE_X3Y144_AQ;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_A4 = CLBLM_R_X3Y144_SLICE_X3Y144_BO6;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_A5 = CLBLL_L_X2Y146_SLICE_X1Y146_CQ;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_C1 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_C2 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_C3 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_B1 = CLBLM_R_X5Y147_SLICE_X7Y147_D5Q;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_B2 = CLBLM_R_X3Y148_SLICE_X3Y148_BQ;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_B3 = CLBLL_L_X2Y147_SLICE_X1Y147_AQ;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_B4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_B5 = CLBLM_L_X8Y145_SLICE_X11Y145_AQ;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_B6 = 1'b1;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_D1 = CLBLM_R_X5Y154_SLICE_X7Y154_AO6;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_D2 = CLBLM_L_X8Y151_SLICE_X11Y151_AQ;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_C1 = CLBLM_R_X3Y146_SLICE_X2Y146_AQ;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_C2 = CLBLM_R_X3Y146_SLICE_X2Y146_BQ;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_C3 = CLBLL_L_X4Y144_SLICE_X4Y144_BQ;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_C4 = CLBLM_R_X3Y146_SLICE_X3Y146_CQ;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_C5 = 1'b1;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_C6 = CLBLL_L_X4Y144_SLICE_X4Y144_AQ;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_D3 = CLBLM_L_X10Y153_SLICE_X12Y153_CQ;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_D4 = CLBLM_R_X5Y154_SLICE_X7Y154_AO5;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_A1 = CLBLM_R_X5Y152_SLICE_X7Y152_DO5;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_A2 = CLBLM_R_X7Y154_SLICE_X9Y154_AQ;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_A3 = CLBLM_R_X5Y154_SLICE_X6Y154_AQ;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_A4 = CLBLM_R_X5Y149_SLICE_X7Y149_BQ;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_A5 = 1'b1;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_D1 = 1'b1;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_D2 = 1'b1;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_D3 = 1'b1;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_D4 = 1'b1;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_D5 = 1'b1;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_D6 = 1'b1;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_B1 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_B2 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_B3 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_B4 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_A1 = CLBLM_R_X3Y144_SLICE_X2Y144_B5Q;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_A2 = CLBLM_R_X3Y145_SLICE_X2Y145_BQ;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_A3 = CLBLL_L_X4Y144_SLICE_X4Y144_BQ;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_A5 = CLBLM_R_X3Y147_SLICE_X3Y147_DQ;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_A6 = 1'b1;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_C1 = 1'b1;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_C2 = 1'b1;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_C3 = 1'b1;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_B1 = 1'b1;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_B3 = CLBLM_R_X3Y146_SLICE_X3Y146_AQ;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_B4 = CLBLM_R_X3Y146_SLICE_X2Y146_BQ;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_B5 = RIOB33_X105Y127_IOB_X1Y127_I;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_B6 = 1'b1;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_D1 = 1'b1;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_D2 = 1'b1;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_D3 = 1'b1;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_C1 = CLBLM_R_X3Y148_SLICE_X3Y148_BQ;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_C2 = CLBLL_L_X4Y143_SLICE_X4Y143_CO6;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_C3 = CLBLM_R_X3Y144_SLICE_X3Y144_BO5;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_C4 = CLBLM_R_X7Y142_SLICE_X8Y142_DO6;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_C5 = CLBLM_L_X8Y144_SLICE_X11Y144_BO6;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_C6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_D4 = 1'b1;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_D5 = 1'b1;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_D6 = 1'b1;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_C1 = CLBLM_L_X12Y145_SLICE_X16Y145_AQ;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_C2 = CLBLM_R_X7Y146_SLICE_X9Y146_CQ;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_C3 = CLBLM_L_X12Y144_SLICE_X16Y144_BQ;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_D1 = CLBLM_R_X3Y144_SLICE_X3Y144_AQ;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_D2 = CLBLL_L_X4Y143_SLICE_X4Y143_CO6;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_D3 = CLBLL_L_X2Y146_SLICE_X1Y146_CQ;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_D4 = CLBLM_R_X7Y142_SLICE_X8Y142_DO6;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_D5 = CLBLM_L_X8Y144_SLICE_X11Y144_BO6;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_D6 = CLBLL_L_X2Y146_SLICE_X1Y146_AQ;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_C5 = CLBLM_L_X12Y144_SLICE_X16Y144_AQ;
  assign LIOI3_X0Y173_OLOGIC_X0Y174_T1 = 1'b1;
  assign RIOB33_X105Y175_IOB_X1Y176_O = CLBLM_R_X103Y176_SLICE_X163Y176_AO6;
  assign RIOB33_X105Y175_IOB_X1Y175_O = CLBLM_R_X15Y153_SLICE_X20Y153_AO6;
  assign LIOI3_X0Y185_OLOGIC_X0Y186_D1 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign LIOI3_X0Y185_OLOGIC_X0Y186_T1 = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_D1 = CLBLM_R_X3Y143_SLICE_X2Y143_BQ;
  assign LIOI3_X0Y185_OLOGIC_X0Y185_D1 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_T1 = 1'b1;
  assign CLBLM_R_X5Y155_SLICE_X7Y155_A1 = CLBLM_R_X5Y155_SLICE_X7Y155_DO6;
  assign CLBLM_R_X5Y155_SLICE_X7Y155_A2 = 1'b1;
  assign CLBLM_R_X5Y155_SLICE_X7Y155_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y155_SLICE_X7Y155_A4 = CLBLM_R_X7Y155_SLICE_X8Y155_BO5;
  assign CLBLM_R_X5Y155_SLICE_X7Y155_A5 = CLBLM_R_X5Y149_SLICE_X7Y149_AQ;
  assign CLBLM_R_X5Y155_SLICE_X7Y155_A6 = CLBLM_R_X5Y155_SLICE_X7Y155_AQ;
  assign LIOI3_X0Y185_OLOGIC_X0Y185_T1 = 1'b1;
  assign RIOI3_X105Y171_OLOGIC_X1Y172_D1 = CLBLM_R_X103Y170_SLICE_X163Y170_AO5;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_D1 = CLBLM_L_X8Y145_SLICE_X11Y145_B5Q;
  assign CLBLM_R_X5Y155_SLICE_X7Y155_B1 = CLBLM_R_X7Y155_SLICE_X8Y155_BO5;
  assign CLBLM_R_X5Y155_SLICE_X7Y155_B2 = CLBLM_R_X5Y152_SLICE_X6Y152_AQ;
  assign CLBLM_R_X5Y155_SLICE_X7Y155_B3 = CLBLM_R_X5Y155_SLICE_X7Y155_AQ;
  assign CLBLM_R_X5Y155_SLICE_X7Y155_B4 = CLBLM_R_X5Y155_SLICE_X6Y155_BQ;
  assign CLBLM_R_X5Y155_SLICE_X7Y155_B5 = CLBLM_R_X5Y155_SLICE_X6Y155_AQ;
  assign CLBLM_R_X5Y155_SLICE_X7Y155_B6 = 1'b1;
  assign RIOI3_X105Y171_OLOGIC_X1Y172_T1 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_A1 = CLBLM_R_X5Y144_SLICE_X6Y144_AQ;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_A2 = CLBLL_L_X4Y154_SLICE_X4Y154_CO6;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_A3 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_A4 = CLBLM_R_X3Y145_SLICE_X3Y145_D5Q;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_A6 = 1'b1;
  assign CLBLM_R_X5Y155_SLICE_X7Y155_C4 = CLBLM_R_X7Y155_SLICE_X8Y155_A5Q;
  assign CLBLM_R_X5Y155_SLICE_X7Y155_C5 = CLBLM_R_X5Y155_SLICE_X7Y155_AQ;
  assign CLBLM_R_X5Y155_SLICE_X7Y155_C6 = CLBLM_R_X5Y155_SLICE_X6Y155_BQ;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_B1 = CLBLM_R_X5Y147_SLICE_X7Y147_CQ;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_B2 = CLBLM_R_X3Y145_SLICE_X3Y145_BQ;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_B3 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_B5 = CLBLM_R_X5Y152_SLICE_X7Y152_DO6;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_B6 = CLBLM_R_X3Y142_SLICE_X2Y142_CQ;
  assign CLBLM_R_X5Y155_SLICE_X7Y155_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X5Y155_SLICE_X7Y155_D1 = CLBLM_R_X5Y155_SLICE_X6Y155_AQ;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_C2 = CLBLM_R_X3Y145_SLICE_X3Y145_CQ;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_C3 = CLBLL_L_X4Y146_SLICE_X4Y146_AQ;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_C4 = CLBLM_R_X5Y144_SLICE_X6Y144_AQ;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_C5 = CLBLM_R_X3Y145_SLICE_X2Y145_A5Q;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_C6 = CLBLM_R_X5Y144_SLICE_X6Y144_BO6;
  assign CLBLM_R_X5Y155_SLICE_X7Y155_D3 = 1'b1;
  assign CLBLM_R_X5Y155_SLICE_X7Y155_D4 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y155_SLICE_X6Y155_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y155_SLICE_X6Y155_A2 = CLBLM_R_X5Y155_SLICE_X6Y155_BQ;
  assign CLBLM_R_X5Y155_SLICE_X6Y155_A3 = CLBLM_R_X5Y155_SLICE_X6Y155_AQ;
  assign CLBLM_R_X5Y155_SLICE_X6Y155_A4 = CLBLM_R_X5Y152_SLICE_X6Y152_AQ;
  assign CLBLM_R_X5Y155_SLICE_X6Y155_A5 = CLBLM_R_X5Y155_SLICE_X7Y155_BO6;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_D2 = CLBLL_L_X4Y146_SLICE_X4Y146_A5Q;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_D3 = CLBLM_R_X11Y146_SLICE_X14Y146_AQ;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_D4 = CLBLM_R_X3Y145_SLICE_X3Y145_BQ;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_D5 = CLBLL_L_X2Y147_SLICE_X1Y147_AQ;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_D6 = 1'b1;
  assign CLBLM_R_X5Y155_SLICE_X6Y155_A6 = CLBLM_R_X7Y152_SLICE_X8Y152_BQ;
  assign CLBLM_R_X5Y155_SLICE_X6Y155_B1 = 1'b1;
  assign CLBLM_R_X5Y155_SLICE_X6Y155_B2 = CLBLM_R_X5Y155_SLICE_X6Y155_BQ;
  assign CLBLM_R_X5Y155_SLICE_X6Y155_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y155_SLICE_X6Y155_B4 = CLBLM_R_X5Y154_SLICE_X6Y154_AQ;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_A1 = CLBLM_R_X5Y152_SLICE_X7Y152_DO6;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_A3 = CLBLM_R_X3Y145_SLICE_X2Y145_AQ;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_A4 = CLBLL_L_X2Y145_SLICE_X1Y145_AQ;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_A5 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_A6 = CLBLM_R_X5Y152_SLICE_X6Y152_A5Q;
  assign CLBLM_R_X5Y155_SLICE_X6Y155_C1 = 1'b1;
  assign CLBLM_R_X5Y155_SLICE_X6Y155_C2 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_AX = CLBLM_R_X3Y145_SLICE_X2Y145_CO6;
  assign CLBLM_R_X5Y155_SLICE_X6Y155_C3 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_B1 = CLBLM_R_X5Y144_SLICE_X6Y144_BO5;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_B2 = CLBLM_R_X3Y145_SLICE_X2Y145_BQ;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_B4 = CLBLM_R_X5Y148_SLICE_X7Y148_CQ;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_B5 = CLBLM_R_X3Y145_SLICE_X2Y145_CO5;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_B6 = CLBLM_R_X3Y145_SLICE_X3Y145_CQ;
  assign CLBLM_R_X5Y155_SLICE_X6Y155_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X5Y155_SLICE_X6Y155_D1 = 1'b1;
  assign CLBLM_R_X5Y155_SLICE_X6Y155_D2 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_C1 = CLBLM_R_X5Y144_SLICE_X6Y144_BO5;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_C2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_C3 = CLBLM_R_X5Y144_SLICE_X6Y144_AQ;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_C4 = CLBLM_R_X3Y145_SLICE_X2Y145_A5Q;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_C5 = CLBLM_L_X12Y147_SLICE_X16Y147_AQ;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_C6 = 1'b1;
  assign CLBLM_R_X5Y155_SLICE_X6Y155_D3 = 1'b1;
  assign CLBLM_R_X5Y155_SLICE_X6Y155_D4 = 1'b1;
  assign CLBLM_R_X5Y155_SLICE_X6Y155_D5 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y155_SLICE_X6Y155_D6 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_D1 = CLBLL_L_X4Y144_SLICE_X4Y144_BQ;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_D2 = CLBLM_R_X5Y144_SLICE_X6Y144_AQ;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_D3 = CLBLM_R_X3Y145_SLICE_X2Y145_A5Q;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_D4 = CLBLM_R_X3Y145_SLICE_X3Y145_CQ;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_D5 = CLBLM_R_X3Y145_SLICE_X2Y145_BQ;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_D6 = CLBLL_L_X4Y144_SLICE_X4Y144_AQ;
  assign RIOB33_X105Y177_IOB_X1Y178_O = CLBLM_R_X103Y178_SLICE_X163Y178_AO6;
  assign RIOB33_X105Y177_IOB_X1Y177_O = CLBLM_R_X103Y176_SLICE_X163Y176_AO5;
  assign LIOI3_X0Y173_OLOGIC_X0Y173_D1 = CLBLM_R_X103Y141_SLICE_X163Y141_AO5;
  assign LIOI3_X0Y65_ILOGIC_X0Y66_D = LIOB33_X0Y65_IOB_X0Y66_I;
  assign LIOI3_X0Y65_ILOGIC_X0Y65_D = LIOB33_X0Y65_IOB_X0Y65_I;
  assign RIOI3_X105Y109_ILOGIC_X1Y110_D = RIOB33_X105Y109_IOB_X1Y110_I;
  assign RIOI3_X105Y109_ILOGIC_X1Y109_D = RIOB33_X105Y109_IOB_X1Y109_I;
  assign RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y138_D = RIOB33_X105Y137_IOB_X1Y138_I;
  assign RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y137_D = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_A1 = CLBLM_L_X8Y149_SLICE_X11Y149_AQ;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_A2 = CLBLM_R_X3Y146_SLICE_X3Y146_BQ;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_A3 = CLBLL_L_X4Y151_SLICE_X4Y151_AQ;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_A5 = CLBLL_L_X4Y143_SLICE_X4Y143_AQ;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_A6 = CLBLM_R_X3Y146_SLICE_X3Y146_AQ;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_B1 = CLBLM_L_X8Y149_SLICE_X11Y149_AQ;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_B3 = CLBLM_R_X11Y146_SLICE_X14Y146_AQ;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_B4 = CLBLM_R_X3Y146_SLICE_X3Y146_DO5;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_B5 = CLBLM_R_X3Y146_SLICE_X2Y146_DO6;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_B6 = CLBLM_R_X3Y146_SLICE_X3Y146_BQ;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_C1 = CLBLM_R_X5Y144_SLICE_X6Y144_BO6;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_C2 = CLBLM_R_X3Y146_SLICE_X2Y146_CO6;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_C3 = 1'b1;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_C4 = CLBLM_R_X3Y147_SLICE_X3Y147_BQ;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_C5 = CLBLM_R_X3Y146_SLICE_X3Y146_CQ;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign RIOI3_X105Y165_OLOGIC_X1Y166_D1 = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_D1 = CLBLL_L_X4Y147_SLICE_X5Y147_BQ;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_D2 = CLBLM_L_X10Y147_SLICE_X12Y147_AQ;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_D3 = CLBLM_R_X3Y146_SLICE_X3Y146_BQ;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_D4 = CLBLL_L_X4Y146_SLICE_X4Y146_DO6;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_D5 = CLBLM_R_X11Y147_SLICE_X14Y147_BQ;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_D6 = 1'b1;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_A2 = CLBLM_R_X3Y149_SLICE_X2Y149_BQ;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_A3 = CLBLM_R_X3Y146_SLICE_X2Y146_AQ;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_A4 = CLBLM_R_X5Y144_SLICE_X6Y144_BO6;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_A5 = 1'b1;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_A6 = CLBLM_R_X3Y145_SLICE_X2Y145_DO6;
  assign LIOB33_X0Y139_IOB_X0Y139_O = CLBLM_R_X3Y143_SLICE_X3Y143_AQ;
  assign LIOB33_X0Y139_IOB_X0Y140_O = CLBLM_R_X3Y142_SLICE_X2Y142_CQ;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_B1 = CLBLM_R_X5Y148_SLICE_X6Y148_AQ;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_B2 = CLBLM_R_X3Y146_SLICE_X2Y146_BQ;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_B3 = CLBLM_R_X3Y146_SLICE_X2Y146_AQ;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_B4 = CLBLM_R_X5Y144_SLICE_X6Y144_BO6;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_B6 = CLBLM_R_X3Y145_SLICE_X2Y145_DO6;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_C1 = 1'b1;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_C2 = CLBLM_R_X3Y146_SLICE_X2Y146_AQ;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_C3 = CLBLM_R_X3Y146_SLICE_X2Y146_BQ;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_C4 = CLBLM_R_X3Y145_SLICE_X2Y145_DO6;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_C5 = 1'b1;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_C6 = 1'b1;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_D1 = 1'b1;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_D2 = 1'b1;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_D3 = CLBLM_R_X11Y147_SLICE_X14Y147_BQ;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_D4 = CLBLL_L_X4Y146_SLICE_X4Y146_DO6;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_D5 = 1'b1;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_D6 = CLBLM_L_X10Y147_SLICE_X12Y147_AQ;
  assign RIOI3_X105Y139_ILOGIC_X1Y140_D = RIOB33_X105Y139_IOB_X1Y140_I;
  assign RIOB33_X105Y179_IOB_X1Y180_O = CLBLM_R_X11Y151_SLICE_X14Y151_DO6;
  assign RIOB33_X105Y179_IOB_X1Y179_O = CLBLM_R_X103Y178_SLICE_X163Y178_AO5;
  assign RIOI3_X105Y139_ILOGIC_X1Y139_D = RIOB33_X105Y139_IOB_X1Y139_I;
  assign CLBLM_R_X11Y154_SLICE_X15Y154_C1 = CLBLM_R_X11Y153_SLICE_X15Y153_CO5;
  assign CLBLM_R_X11Y154_SLICE_X15Y154_C2 = CLBLM_R_X11Y154_SLICE_X14Y154_AQ;
  assign CLBLM_R_X11Y154_SLICE_X15Y154_C6 = 1'b1;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_A1 = CLBLL_L_X4Y144_SLICE_X5Y144_AQ;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_A2 = CLBLM_R_X5Y152_SLICE_X7Y152_DO6;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_A3 = CLBLM_R_X3Y147_SLICE_X3Y147_AQ;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_A4 = 1'b1;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_A5 = CLBLM_R_X3Y150_SLICE_X3Y150_AQ;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y154_SLICE_X15Y154_D2 = CLBLM_R_X11Y154_SLICE_X14Y154_AQ;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_B1 = CLBLM_R_X3Y147_SLICE_X2Y147_DQ;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_B2 = CLBLM_R_X3Y147_SLICE_X3Y147_BQ;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_B4 = CLBLM_R_X11Y146_SLICE_X14Y146_AQ;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_B5 = 1'b1;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_B6 = CLBLM_R_X3Y146_SLICE_X3Y146_DO6;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_C1 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_C2 = CLBLL_L_X4Y147_SLICE_X4Y147_BQ;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_C3 = 1'b1;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_C4 = CLBLM_R_X3Y147_SLICE_X2Y147_CQ;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_C6 = 1'b1;
  assign CLBLM_R_X11Y154_SLICE_X15Y154_D5 = CLBLM_R_X11Y154_SLICE_X15Y154_AQ;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y154_SLICE_X15Y154_D6 = CLBLM_L_X10Y154_SLICE_X13Y154_AQ;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_D1 = CLBLL_L_X4Y147_SLICE_X5Y147_BQ;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_D2 = CLBLM_L_X8Y148_SLICE_X10Y148_A5Q;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_D3 = CLBLM_R_X3Y147_SLICE_X3Y147_DQ;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_D4 = CLBLM_R_X11Y150_SLICE_X14Y150_BO6;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_D5 = CLBLM_R_X5Y142_SLICE_X7Y142_AQ;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_D6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_A1 = 1'b1;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_A2 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_A3 = CLBLM_R_X3Y147_SLICE_X2Y147_AQ;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_A4 = CLBLM_R_X5Y152_SLICE_X7Y152_BQ;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_A6 = 1'b1;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_AX = CLBLM_R_X3Y147_SLICE_X2Y147_BO6;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_B1 = CLBLM_L_X8Y149_SLICE_X11Y149_AQ;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_B2 = CLBLM_R_X3Y147_SLICE_X3Y147_AQ;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_B3 = CLBLL_L_X4Y151_SLICE_X4Y151_AQ;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_B4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_B6 = 1'b1;
  assign LIOI3_X0Y189_OLOGIC_X0Y190_D1 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_C1 = CLBLL_L_X4Y151_SLICE_X4Y151_AQ;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_C2 = CLBLM_R_X3Y147_SLICE_X2Y147_CQ;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_C4 = CLBLL_L_X4Y146_SLICE_X4Y146_A5Q;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_C5 = CLBLM_L_X8Y149_SLICE_X11Y149_AQ;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_C6 = CLBLM_R_X11Y147_SLICE_X14Y147_BQ;
  assign LIOI3_X0Y189_OLOGIC_X0Y190_T1 = 1'b1;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_D1 = CLBLL_L_X2Y147_SLICE_X1Y147_AQ;
  assign CLBLM_R_X13Y152_SLICE_X18Y152_D1 = 1'b1;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_D2 = CLBLM_L_X8Y152_SLICE_X11Y152_BO6;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_D3 = CLBLM_R_X3Y147_SLICE_X2Y147_DQ;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_D4 = CLBLM_R_X5Y146_SLICE_X6Y146_CQ;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_D5 = 1'b1;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_D6 = CLBLM_R_X3Y148_SLICE_X2Y148_AQ;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_T1 = 1'b1;
  assign LIOI3_X0Y189_OLOGIC_X0Y189_D1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign RIOI3_X105Y173_OLOGIC_X1Y174_D1 = CLBLM_R_X103Y173_SLICE_X163Y173_AO5;
  assign LIOI3_X0Y189_OLOGIC_X0Y189_T1 = 1'b1;
  assign CLBLM_R_X13Y152_SLICE_X18Y152_D4 = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_D1 = CLBLL_L_X4Y147_SLICE_X5Y147_CQ;
  assign RIOB33_X105Y181_IOB_X1Y182_O = CLBLM_L_X10Y152_SLICE_X13Y152_CO6;
  assign RIOB33_X105Y181_IOB_X1Y181_O = CLBLM_R_X11Y151_SLICE_X14Y151_DO5;
  assign RIOI3_X105Y173_OLOGIC_X1Y174_T1 = 1'b1;
  assign CLBLM_R_X13Y152_SLICE_X18Y152_D6 = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_T1 = 1'b1;
  assign RIOI3_X105Y173_OLOGIC_X1Y173_D1 = CLBLM_R_X103Y173_SLICE_X163Y173_AO6;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_D1 = CLBLM_R_X5Y142_SLICE_X7Y142_AQ;
  assign RIOI3_X105Y173_OLOGIC_X1Y173_T1 = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_D1 = CLBLM_L_X10Y150_SLICE_X13Y150_DO5;
  assign CLBLM_R_X11Y154_SLICE_X14Y154_B5 = CLBLM_R_X11Y154_SLICE_X15Y154_AQ;
  assign CLBLM_R_X11Y154_SLICE_X14Y154_B6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_D1 = CLBLM_R_X7Y142_SLICE_X8Y142_AO5;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_D1 = CLBLM_L_X10Y150_SLICE_X13Y150_DO6;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_T1 = 1'b1;
  assign CLBLM_R_X11Y154_SLICE_X14Y154_C3 = CLBLM_R_X11Y154_SLICE_X15Y154_BQ;
  assign CLBLM_R_X11Y154_SLICE_X14Y154_C4 = 1'b1;
  assign CLBLM_R_X11Y154_SLICE_X14Y154_C5 = CLBLM_L_X10Y153_SLICE_X13Y153_BQ;
  assign CLBLM_R_X11Y154_SLICE_X14Y154_C6 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_D3 = CLBLM_L_X12Y153_SLICE_X16Y153_DO6;
  assign LIOI3_X0Y67_ILOGIC_X0Y68_D = LIOB33_X0Y67_IOB_X0Y68_I;
  assign LIOI3_X0Y67_ILOGIC_X0Y67_D = LIOB33_X0Y67_IOB_X0Y67_I;
  assign RIOI3_X105Y111_ILOGIC_X1Y112_D = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_A1 = CLBLM_R_X3Y148_SLICE_X3Y148_B5Q;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_A2 = CLBLM_R_X3Y148_SLICE_X2Y148_CQ;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_A4 = CLBLM_R_X5Y148_SLICE_X7Y148_C5Q;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_A5 = CLBLM_R_X3Y148_SLICE_X2Y148_AQ;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_A6 = CLBLM_R_X3Y148_SLICE_X2Y148_BQ;
  assign RIOI3_X105Y111_ILOGIC_X1Y111_D = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_D4 = CLBLM_L_X10Y154_SLICE_X13Y154_CO5;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_B1 = CLBLL_L_X4Y149_SLICE_X4Y149_CQ;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_B3 = CLBLL_L_X4Y144_SLICE_X4Y144_DO6;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_B4 = CLBLM_R_X3Y148_SLICE_X3Y148_DO6;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_B5 = CLBLM_R_X7Y149_SLICE_X8Y149_AQ;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_B6 = 1'b1;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_C1 = CLBLL_L_X4Y148_SLICE_X4Y148_C5Q;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_C2 = CLBLM_R_X3Y148_SLICE_X3Y148_CQ;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_C3 = CLBLM_R_X3Y144_SLICE_X2Y144_CO6;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_C4 = CLBLL_L_X4Y146_SLICE_X5Y146_A5Q;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_C6 = 1'b1;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_D5 = CLBLM_R_X11Y153_SLICE_X15Y153_AQ;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_D1 = CLBLM_R_X3Y148_SLICE_X2Y148_AQ;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_D2 = CLBLL_L_X2Y148_SLICE_X1Y148_BO6;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_D3 = CLBLM_R_X11Y150_SLICE_X14Y150_BO6;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_D4 = CLBLM_R_X3Y148_SLICE_X2Y148_CQ;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_D5 = CLBLM_R_X3Y148_SLICE_X3Y148_B5Q;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_D6 = CLBLM_R_X3Y148_SLICE_X2Y148_BQ;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_A2 = CLBLL_L_X4Y148_SLICE_X4Y148_C5Q;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_A3 = CLBLM_R_X3Y148_SLICE_X2Y148_AQ;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_A4 = CLBLM_R_X11Y150_SLICE_X14Y150_BO6;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_A5 = CLBLL_L_X2Y148_SLICE_X1Y148_BO6;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_A6 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_D6 = CLBLM_R_X11Y153_SLICE_X14Y153_CO5;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_B1 = CLBLM_L_X8Y150_SLICE_X11Y150_AQ;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_B2 = CLBLM_R_X3Y148_SLICE_X2Y148_BQ;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_B3 = CLBLL_L_X2Y147_SLICE_X1Y147_AO6;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_B4 = CLBLM_R_X3Y148_SLICE_X2Y148_CQ;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_B6 = CLBLM_R_X3Y148_SLICE_X2Y148_AO5;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_C1 = CLBLL_L_X2Y147_SLICE_X1Y147_AO6;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_C2 = CLBLM_R_X3Y148_SLICE_X2Y148_CQ;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_C4 = CLBLM_R_X3Y148_SLICE_X2Y148_AO5;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_C5 = 1'b1;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_C6 = CLBLM_R_X7Y144_SLICE_X9Y144_CQ;
  assign RIOB33_X105Y183_IOB_X1Y183_O = CLBLM_L_X10Y152_SLICE_X13Y152_CO5;
  assign RIOB33_X105Y183_IOB_X1Y184_O = CLBLM_L_X10Y150_SLICE_X13Y150_DO6;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_D1 = 1'b1;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_D2 = CLBLM_L_X10Y145_SLICE_X12Y145_CQ;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_D3 = CLBLM_R_X3Y148_SLICE_X2Y148_DQ;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_D4 = CLBLM_R_X3Y147_SLICE_X3Y147_CQ;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_D5 = CLBLM_R_X5Y152_SLICE_X7Y152_DO6;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_D6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_B1 = CLBLM_R_X7Y154_SLICE_X9Y154_DO6;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_B2 = CLBLL_L_X4Y147_SLICE_X5Y147_B5Q;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_B3 = CLBLM_R_X7Y154_SLICE_X8Y154_BQ;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_B4 = CLBLM_R_X7Y154_SLICE_X9Y154_BQ;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_B5 = CLBLM_R_X7Y153_SLICE_X8Y153_CQ;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_B6 = CLBLM_R_X7Y155_SLICE_X9Y155_CO6;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_A6 = 1'b1;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_A1 = CLBLM_R_X5Y152_SLICE_X7Y152_DO6;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_A2 = CLBLM_R_X11Y148_SLICE_X15Y148_B5Q;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_A3 = CLBLM_R_X7Y149_SLICE_X8Y149_AQ;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_A4 = CLBLM_R_X3Y149_SLICE_X3Y149_AQ;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_A6 = 1'b1;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_B2 = CLBLM_R_X3Y149_SLICE_X3Y149_BQ;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_B3 = CLBLM_R_X3Y146_SLICE_X2Y146_BQ;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_B4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_B5 = CLBLM_R_X3Y149_SLICE_X2Y149_CQ;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_B6 = 1'b1;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_C2 = CLBLM_R_X3Y149_SLICE_X3Y149_CQ;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_C3 = CLBLL_L_X4Y145_SLICE_X4Y145_CQ;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_C4 = CLBLM_R_X11Y150_SLICE_X14Y150_BO6;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_C5 = CLBLM_L_X8Y148_SLICE_X10Y148_A5Q;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_C6 = CLBLM_R_X11Y150_SLICE_X15Y150_AQ;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_D1 = CLBLM_R_X5Y153_SLICE_X6Y153_A5Q;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_D2 = CLBLM_R_X11Y150_SLICE_X14Y150_BO6;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_D3 = CLBLM_R_X3Y149_SLICE_X3Y149_DQ;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_D4 = CLBLM_L_X8Y148_SLICE_X10Y148_A5Q;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_D6 = CLBLM_R_X7Y145_SLICE_X8Y145_AQ;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_B3 = CLBLM_R_X11Y144_SLICE_X14Y144_AQ;
  assign RIOB33_X105Y185_IOB_X1Y186_O = CLBLM_L_X12Y151_SLICE_X16Y151_AQ;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_B4 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign RIOB33_X105Y185_IOB_X1Y185_O = CLBLM_L_X10Y150_SLICE_X13Y150_DO5;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_A1 = CLBLM_R_X3Y148_SLICE_X2Y148_DQ;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_A2 = CLBLL_L_X4Y151_SLICE_X4Y151_AQ;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_A3 = CLBLM_R_X3Y149_SLICE_X2Y149_AQ;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_A4 = CLBLL_L_X4Y145_SLICE_X4Y145_CQ;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_A5 = CLBLM_L_X8Y149_SLICE_X11Y149_AQ;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_B5 = CLBLM_R_X5Y142_SLICE_X7Y142_AQ;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_B6 = CLBLM_R_X11Y144_SLICE_X14Y144_CO6;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_B1 = CLBLM_R_X5Y150_SLICE_X7Y150_AQ;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_B2 = CLBLM_R_X3Y149_SLICE_X2Y149_BQ;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_B4 = CLBLM_R_X7Y150_SLICE_X9Y150_A5Q;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_B5 = CLBLM_L_X8Y152_SLICE_X11Y152_BO6;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_B6 = 1'b1;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_C1 = CLBLM_R_X7Y150_SLICE_X9Y150_A5Q;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_C2 = CLBLM_R_X5Y152_SLICE_X7Y152_B5Q;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_C4 = 1'b1;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_C5 = CLBLM_R_X3Y144_SLICE_X2Y144_CO6;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_C6 = CLBLM_R_X3Y149_SLICE_X2Y149_CQ;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_D1 = CLBLM_R_X7Y145_SLICE_X9Y145_AQ;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_D2 = 1'b1;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_D3 = 1'b1;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_D4 = CLBLM_R_X3Y147_SLICE_X2Y147_CQ;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_D5 = CLBLL_L_X2Y152_SLICE_X1Y152_BO6;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_D6 = CLBLL_L_X4Y152_SLICE_X5Y152_AO6;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_A1 = 1'b1;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_A2 = 1'b1;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_A3 = 1'b1;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_A4 = 1'b1;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_A5 = 1'b1;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_A6 = 1'b1;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_B1 = 1'b1;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_B2 = 1'b1;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_B3 = 1'b1;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_B4 = 1'b1;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_B5 = 1'b1;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_B6 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_C6 = CLBLM_R_X3Y145_SLICE_X3Y145_DQ;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_C1 = 1'b1;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_C2 = 1'b1;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_C3 = 1'b1;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_C4 = 1'b1;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_C5 = 1'b1;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_C6 = 1'b1;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_D1 = 1'b1;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_D2 = 1'b1;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_D3 = 1'b1;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_D4 = 1'b1;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_D5 = 1'b1;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_D6 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_A1 = CLBLM_R_X3Y145_SLICE_X2Y145_AQ;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_A2 = CLBLM_L_X10Y152_SLICE_X12Y152_DQ;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_A5 = CLBLM_L_X12Y145_SLICE_X16Y145_CO5;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_A6 = 1'b1;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_B1 = CLBLM_L_X12Y144_SLICE_X16Y144_DO6;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_B2 = CLBLM_L_X12Y144_SLICE_X16Y144_BQ;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_B3 = CLBLM_R_X7Y142_SLICE_X8Y142_DO6;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_B5 = CLBLM_L_X10Y144_SLICE_X12Y144_AQ;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_B6 = CLBLM_L_X12Y144_SLICE_X16Y144_AO5;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_C1 = CLBLM_L_X10Y152_SLICE_X12Y152_DQ;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_C2 = CLBLM_L_X12Y144_SLICE_X16Y144_CQ;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_C5 = CLBLM_L_X12Y144_SLICE_X16Y144_DO6;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_C6 = CLBLM_L_X12Y154_SLICE_X16Y154_AQ;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_A6 = CLBLL_L_X4Y149_SLICE_X5Y149_CQ;
  assign LIOI3_X0Y191_OLOGIC_X0Y192_D1 = LIOB33_X0Y51_IOB_X0Y52_I;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_D1 = CLBLM_L_X12Y145_SLICE_X16Y145_AQ;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_D2 = CLBLM_L_X12Y144_SLICE_X16Y144_CQ;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_D3 = CLBLM_R_X7Y142_SLICE_X8Y142_DO6;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_D4 = CLBLM_L_X12Y144_SLICE_X16Y144_AQ;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_D5 = CLBLM_L_X12Y144_SLICE_X16Y144_BQ;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_D6 = 1'b1;
  assign LIOI3_X0Y191_OLOGIC_X0Y192_T1 = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_D1 = CLBLL_L_X52Y126_SLICE_X78Y126_AO6;
  assign LIOI3_X0Y191_OLOGIC_X0Y191_D1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_T1 = 1'b1;
  assign RIOI3_X105Y175_OLOGIC_X1Y176_D1 = CLBLM_R_X103Y176_SLICE_X163Y176_AO6;
  assign LIOI3_X0Y191_OLOGIC_X0Y191_T1 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_B3 = CLBLM_R_X11Y148_SLICE_X15Y148_AQ;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_D1 = CLBLM_R_X3Y148_SLICE_X3Y148_AQ;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_B4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign RIOI3_X105Y175_OLOGIC_X1Y176_T1 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_B5 = CLBLM_R_X7Y152_SLICE_X9Y152_CQ;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_B6 = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_T1 = 1'b1;
  assign RIOI3_X105Y175_OLOGIC_X1Y175_D1 = CLBLM_R_X15Y153_SLICE_X20Y153_AO6;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_D1 = LIOB33_X0Y57_IOB_X0Y57_I;
  assign RIOI3_X105Y175_OLOGIC_X1Y175_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_D1 = CLBLM_L_X10Y155_SLICE_X13Y155_AQ;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_D1 = LIOB33_X0Y55_IOB_X0Y55_I;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_D1 = CLBLM_R_X11Y151_SLICE_X14Y151_BQ;
  assign LIOB33_X0Y101_IOB_X0Y102_O = CLBLL_L_X2Y138_SLICE_X0Y138_BO5;
  assign LIOB33_X0Y101_IOB_X0Y101_O = CLBLL_L_X2Y138_SLICE_X0Y138_BO6;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_T1 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_A1 = CLBLL_L_X4Y151_SLICE_X4Y151_A5Q;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_A2 = CLBLM_R_X5Y152_SLICE_X6Y152_A5Q;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_A4 = CLBLM_R_X3Y147_SLICE_X2Y147_A5Q;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_A6 = 1'b1;
  assign RIOB33_X105Y167_IOB_X1Y168_O = CLBLM_L_X8Y159_SLICE_X10Y159_AO6;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_B2 = CLBLM_R_X3Y150_SLICE_X3Y150_BQ;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_B3 = CLBLM_R_X3Y144_SLICE_X2Y144_CO6;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_B4 = CLBLM_R_X3Y143_SLICE_X3Y143_B5Q;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_B5 = 1'b1;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_B6 = CLBLM_R_X5Y150_SLICE_X6Y150_A5Q;
  assign RIOB33_X105Y187_IOB_X1Y187_O = CLBLM_R_X11Y151_SLICE_X14Y151_BQ;
  assign RIOB33_X105Y187_IOB_X1Y188_O = CLBLM_L_X10Y155_SLICE_X13Y155_AQ;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_C1 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_C2 = CLBLL_L_X2Y150_SLICE_X1Y150_DO6;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_C3 = CLBLL_L_X2Y154_SLICE_X1Y154_BO6;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_C4 = CLBLL_L_X4Y149_SLICE_X4Y149_AQ;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_C5 = CLBLL_L_X2Y149_SLICE_X1Y149_DO6;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_C6 = CLBLL_L_X4Y152_SLICE_X4Y152_AO6;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign RIOB33_X105Y167_IOB_X1Y167_O = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_D1 = CLBLL_L_X4Y145_SLICE_X4Y145_AQ;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_D2 = CLBLL_L_X4Y155_SLICE_X4Y155_AO5;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_D3 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_D4 = CLBLM_R_X3Y147_SLICE_X3Y147_DQ;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_D5 = CLBLL_L_X2Y151_SLICE_X0Y151_CO5;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_D6 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_A1 = CLBLL_L_X2Y155_SLICE_X1Y155_DO6;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_A2 = CLBLM_L_X8Y153_SLICE_X11Y153_DQ;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_A3 = CLBLM_R_X3Y156_SLICE_X2Y156_AO6;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_A4 = CLBLM_L_X8Y150_SLICE_X11Y150_AQ;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_A5 = CLBLL_L_X2Y150_SLICE_X0Y150_AO6;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_A6 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_B1 = CLBLM_R_X3Y151_SLICE_X2Y151_DO6;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_B2 = CLBLL_L_X4Y150_SLICE_X4Y150_DO6;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_B3 = CLBLM_R_X3Y149_SLICE_X2Y149_DO6;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_B4 = CLBLL_L_X2Y150_SLICE_X1Y150_AO6;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_B5 = CLBLM_R_X3Y155_SLICE_X2Y155_DO6;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_B6 = CLBLL_L_X4Y150_SLICE_X5Y150_DO6;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_C1 = CLBLM_R_X3Y156_SLICE_X2Y156_AO6;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_C2 = CLBLL_L_X2Y155_SLICE_X1Y155_DO6;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_C3 = CLBLM_R_X3Y147_SLICE_X2Y147_DQ;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_C4 = CLBLM_L_X10Y146_SLICE_X12Y146_C5Q;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_C5 = CLBLL_L_X2Y150_SLICE_X0Y150_AO6;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_C6 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_D1 = CLBLM_R_X3Y149_SLICE_X2Y149_BQ;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_D2 = 1'b1;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_D3 = CLBLM_R_X7Y150_SLICE_X8Y150_AQ;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_D4 = 1'b1;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_D5 = CLBLL_L_X4Y152_SLICE_X5Y152_AO6;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_D6 = CLBLL_L_X2Y152_SLICE_X1Y152_BO6;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_A1 = 1'b1;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_A2 = 1'b1;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_A3 = 1'b1;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_A4 = 1'b1;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_A5 = 1'b1;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_A6 = 1'b1;
  assign LIOI3_X0Y71_ILOGIC_X0Y72_D = LIOB33_X0Y71_IOB_X0Y72_I;
  assign LIOI3_X0Y71_ILOGIC_X0Y71_D = LIOB33_X0Y71_IOB_X0Y71_I;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_B1 = 1'b1;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_B2 = 1'b1;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_B3 = 1'b1;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_B4 = 1'b1;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_B5 = 1'b1;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_B6 = 1'b1;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_B5 = CLBLM_R_X5Y153_SLICE_X7Y153_AQ;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_C1 = 1'b1;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_C2 = 1'b1;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_C3 = 1'b1;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_C4 = 1'b1;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_C5 = 1'b1;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_C6 = 1'b1;
  assign RIOI3_X105Y115_ILOGIC_X1Y116_D = RIOB33_X105Y115_IOB_X1Y116_I;
  assign RIOI3_X105Y115_ILOGIC_X1Y115_D = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_D1 = 1'b1;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_D2 = 1'b1;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_D3 = 1'b1;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_D4 = 1'b1;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_D5 = 1'b1;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_D6 = 1'b1;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_A3 = CLBLM_L_X12Y145_SLICE_X16Y145_AQ;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_A4 = CLBLM_R_X7Y142_SLICE_X8Y142_BQ;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_A5 = CLBLM_L_X10Y152_SLICE_X12Y152_DQ;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_A6 = CLBLM_L_X12Y145_SLICE_X16Y145_CO6;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_B1 = CLBLL_L_X4Y145_SLICE_X5Y145_DO6;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_B2 = CLBLM_L_X12Y145_SLICE_X16Y145_BQ;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_B3 = CLBLM_R_X11Y152_SLICE_X14Y152_AQ;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_B5 = CLBLM_R_X11Y145_SLICE_X14Y145_BQ;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_B6 = 1'b1;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_C1 = CLBLM_L_X12Y144_SLICE_X16Y144_BQ;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_C2 = CLBLM_L_X12Y145_SLICE_X16Y145_AQ;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_C3 = CLBLM_R_X7Y142_SLICE_X8Y142_DO6;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_C4 = CLBLM_L_X12Y144_SLICE_X16Y144_CQ;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_C5 = CLBLM_L_X12Y144_SLICE_X16Y144_AQ;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_C6 = 1'b1;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_D1 = 1'b1;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_D2 = 1'b1;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_D3 = 1'b1;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_D4 = 1'b1;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_D5 = 1'b1;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_D6 = 1'b1;
  assign LIOB33_X0Y141_IOB_X0Y142_O = LIOB33_X0Y53_IOB_X0Y54_I;
  assign LIOB33_X0Y141_IOB_X0Y141_O = CLBLM_R_X3Y143_SLICE_X2Y143_AQ;
  assign LIOB33_X0Y103_IOB_X0Y104_O = CLBLL_L_X2Y141_SLICE_X0Y141_AO5;
  assign LIOB33_X0Y103_IOB_X0Y103_O = CLBLL_L_X2Y141_SLICE_X0Y141_AO6;
  assign RIOB33_X105Y189_IOB_X1Y190_O = CLBLM_L_X12Y152_SLICE_X17Y152_AQ;
  assign RIOB33_X105Y189_IOB_X1Y189_O = CLBLM_R_X11Y153_SLICE_X14Y153_CQ;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_A1 = CLBLM_R_X3Y152_SLICE_X2Y152_DO6;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_A2 = CLBLL_L_X4Y150_SLICE_X4Y150_CO6;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_A3 = CLBLM_R_X3Y151_SLICE_X2Y151_CO6;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_A4 = CLBLM_R_X3Y151_SLICE_X3Y151_BO6;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_A5 = CLBLM_R_X3Y155_SLICE_X2Y155_DO6;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_A6 = CLBLL_L_X4Y151_SLICE_X4Y151_BO6;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_B1 = CLBLL_L_X4Y149_SLICE_X4Y149_CQ;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_B2 = CLBLM_L_X8Y151_SLICE_X10Y151_DQ;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_B3 = CLBLL_L_X2Y154_SLICE_X1Y154_BO6;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_B4 = CLBLL_L_X4Y152_SLICE_X4Y152_AO6;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_B5 = CLBLL_L_X4Y155_SLICE_X5Y155_AO6;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_B6 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_C1 = 1'b1;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_C2 = CLBLL_L_X2Y151_SLICE_X0Y151_CO5;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_C3 = CLBLL_L_X2Y154_SLICE_X1Y154_BO5;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_C4 = CLBLM_R_X3Y149_SLICE_X3Y149_AQ;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_C5 = CLBLM_R_X5Y150_SLICE_X6Y150_DQ;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_C6 = CLBLL_L_X2Y155_SLICE_X1Y155_DO6;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_D1 = CLBLM_R_X3Y147_SLICE_X3Y147_AQ;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_D2 = CLBLL_L_X4Y155_SLICE_X5Y155_AO5;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_D3 = CLBLM_R_X3Y152_SLICE_X2Y152_AO5;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_D4 = CLBLM_R_X3Y151_SLICE_X3Y151_CO6;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_D5 = 1'b1;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_D6 = CLBLM_R_X5Y147_SLICE_X6Y147_BQ;
  assign RIOI3_X105Y153_OLOGIC_X1Y153_T1 = 1'b1;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_A1 = CLBLL_L_X2Y151_SLICE_X1Y151_BO6;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_A2 = CLBLM_R_X3Y153_SLICE_X2Y153_AO6;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_A3 = CLBLM_R_X3Y151_SLICE_X3Y151_AO6;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_A4 = CLBLM_R_X3Y154_SLICE_X3Y154_AO6;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_A5 = CLBLM_R_X3Y150_SLICE_X2Y150_BO6;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_A6 = CLBLM_R_X3Y152_SLICE_X3Y152_CO6;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_B1 = CLBLL_L_X2Y151_SLICE_X1Y151_AO5;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_B2 = CLBLM_L_X8Y149_SLICE_X11Y149_B5Q;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_B3 = CLBLM_R_X7Y151_SLICE_X8Y151_A5Q;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_B4 = CLBLM_L_X16Y158_SLICE_X22Y158_AO5;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_B5 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_B6 = CLBLL_L_X2Y152_SLICE_X1Y152_AO5;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_C1 = CLBLM_R_X3Y148_SLICE_X2Y148_CQ;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_C2 = CLBLL_L_X4Y148_SLICE_X4Y148_AQ;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_C3 = CLBLL_L_X2Y152_SLICE_X1Y152_BO5;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_C4 = CLBLL_L_X4Y155_SLICE_X5Y155_AO5;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_C5 = CLBLM_R_X3Y152_SLICE_X2Y152_CO6;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_C6 = CLBLM_R_X3Y151_SLICE_X2Y151_BO6;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_D1 = 1'b1;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_D2 = CLBLL_L_X4Y155_SLICE_X5Y155_AO5;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_D3 = CLBLL_L_X2Y152_SLICE_X1Y152_BO5;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_D4 = CLBLM_R_X7Y151_SLICE_X8Y151_AQ;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_D5 = CLBLM_R_X5Y152_SLICE_X6Y152_DO6;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_D6 = CLBLM_R_X3Y148_SLICE_X2Y148_BQ;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_A1 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_A2 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_A3 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_A4 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_A5 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_A6 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_B1 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_B2 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_B3 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_B4 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_B5 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_B6 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_C1 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_C2 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_C3 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_C4 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_C5 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_C6 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_D1 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_D2 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_D3 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_D4 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_D5 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_D6 = 1'b1;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_D4 = CLBLM_L_X12Y149_SLICE_X17Y149_BQ;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_A1 = CLBLM_R_X11Y146_SLICE_X15Y146_CQ;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_A2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_A3 = CLBLM_L_X12Y146_SLICE_X16Y146_AQ;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_A4 = CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_A5 = CLBLM_L_X10Y143_SLICE_X13Y143_AQ;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_B1 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_B2 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_B3 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_B4 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_B5 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_B6 = 1'b1;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_D5 = CLBLM_L_X10Y150_SLICE_X12Y150_AQ;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_C1 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_C2 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_C3 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_C4 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_C5 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_C6 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_D1 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_D2 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_D3 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_D4 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_D5 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_D6 = 1'b1;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_D6 = CLBLM_L_X12Y149_SLICE_X17Y149_CQ;
  assign LIOB33_X0Y105_IOB_X0Y106_O = CLBLL_L_X2Y138_SLICE_X0Y138_CO5;
  assign LIOB33_X0Y105_IOB_X0Y105_O = CLBLL_L_X2Y138_SLICE_X0Y138_CO6;
  assign CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_CE = 1'b1;
  assign CLBLM_R_X7Y157_SLICE_X8Y157_C6 = 1'b1;
  assign RIOB33_X105Y191_IOB_X1Y192_O = CLBLM_R_X11Y151_SLICE_X15Y151_AQ;
  assign RIOB33_X105Y191_IOB_X1Y191_O = CLBLM_L_X10Y149_SLICE_X12Y149_AQ;
  assign LIOI3_X0Y195_OLOGIC_X0Y196_D1 = LIOB33_X0Y69_IOB_X0Y69_I;
  assign CLBLL_L_X2Y134_SLICE_X0Y134_A3 = CLBLL_L_X2Y147_SLICE_X0Y147_AO6;
  assign LIOI3_X0Y195_OLOGIC_X0Y196_T1 = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_D1 = CLBLM_R_X3Y143_SLICE_X2Y143_CQ;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_A1 = CLBLL_L_X4Y155_SLICE_X4Y155_BO6;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_A2 = CLBLL_L_X2Y152_SLICE_X1Y152_AO6;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_A3 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_A4 = CLBLL_L_X2Y155_SLICE_X1Y155_DO6;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_A5 = CLBLL_L_X2Y151_SLICE_X1Y151_AO6;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_A6 = CLBLM_R_X7Y152_SLICE_X8Y152_DQ;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_T1 = 1'b1;
  assign LIOI3_X0Y195_OLOGIC_X0Y195_D1 = LIOB33_X0Y63_IOB_X0Y64_I;
  assign RIOI3_X105Y177_OLOGIC_X1Y178_D1 = CLBLM_R_X103Y178_SLICE_X163Y178_AO6;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_B1 = CLBLM_R_X3Y152_SLICE_X3Y152_DO6;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_B2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_B3 = CLBLL_L_X4Y152_SLICE_X4Y152_CO6;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_B4 = CLBLL_L_X4Y152_SLICE_X5Y152_CO6;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_B5 = CLBLM_R_X3Y152_SLICE_X3Y152_AO6;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_B6 = CLBLL_L_X2Y154_SLICE_X1Y154_BO6;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_D1 = CLBLM_R_X3Y143_SLICE_X3Y143_A5Q;
  assign LIOI3_X0Y195_OLOGIC_X0Y195_T1 = 1'b1;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_C1 = CLBLL_L_X4Y153_SLICE_X5Y153_CO6;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_C2 = CLBLM_R_X3Y151_SLICE_X3Y151_DO6;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_C3 = CLBLL_L_X4Y152_SLICE_X4Y152_DO6;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_C4 = CLBLM_R_X3Y150_SLICE_X3Y150_CO6;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_C5 = CLBLM_R_X3Y155_SLICE_X3Y155_AO5;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_C6 = CLBLL_L_X2Y155_SLICE_X1Y155_BO6;
  assign RIOI3_X105Y177_OLOGIC_X1Y178_T1 = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_T1 = 1'b1;
  assign RIOI3_X105Y177_OLOGIC_X1Y177_D1 = CLBLM_R_X103Y176_SLICE_X163Y176_AO5;
  assign CLBLL_L_X2Y134_SLICE_X0Y134_B2 = 1'b1;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_D1 = CLBLL_L_X4Y154_SLICE_X5Y154_CO5;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_D2 = CLBLM_R_X3Y149_SLICE_X3Y149_DQ;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_D3 = CLBLM_R_X3Y148_SLICE_X2Y148_AQ;
  assign CLBLL_L_X2Y134_SLICE_X0Y134_B3 = 1'b1;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_D4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_D5 = 1'b1;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_D6 = CLBLL_L_X2Y152_SLICE_X1Y152_AO6;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_D1 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLL_L_X2Y134_SLICE_X0Y134_B4 = 1'b1;
  assign RIOI3_X105Y177_OLOGIC_X1Y177_T1 = 1'b1;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_A1 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_A2 = CLBLL_L_X2Y155_SLICE_X1Y155_DO6;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_A3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_A4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_A5 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y134_SLICE_X0Y134_B6 = 1'b1;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_A6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_T1 = 1'b1;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_B1 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_B2 = CLBLL_L_X4Y151_SLICE_X5Y151_BQ;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_B3 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_B4 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_B5 = CLBLM_R_X5Y145_SLICE_X6Y145_DO5;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_B6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_D1 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_C1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_C2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_C3 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_C4 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_C5 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_C6 = CLBLL_L_X2Y152_SLICE_X1Y152_AO6;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_T1 = 1'b1;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_D1 = CLBLM_R_X3Y152_SLICE_X2Y152_AO6;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_D2 = CLBLL_L_X2Y151_SLICE_X0Y151_BO6;
  assign CLBLL_L_X2Y134_SLICE_X0Y134_C3 = 1'b1;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_D3 = LIOB33_X0Y61_IOB_X0Y61_I;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_D4 = CLBLM_R_X3Y152_SLICE_X2Y152_AO5;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_D5 = CLBLM_R_X5Y154_SLICE_X6Y154_AQ;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_D6 = CLBLM_R_X5Y147_SLICE_X6Y147_AQ;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_A1 = 1'b1;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_A2 = 1'b1;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_A3 = 1'b1;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_A4 = 1'b1;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_A5 = 1'b1;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_A6 = 1'b1;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_B1 = 1'b1;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_B2 = 1'b1;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_B3 = 1'b1;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_B4 = 1'b1;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_B5 = 1'b1;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_B6 = 1'b1;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_C1 = 1'b1;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_C2 = 1'b1;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_C3 = 1'b1;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_C4 = 1'b1;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_C5 = 1'b1;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_C6 = 1'b1;
  assign CLBLM_R_X7Y157_SLICE_X9Y157_C4 = 1'b1;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_D1 = 1'b1;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_D2 = 1'b1;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_D3 = 1'b1;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_D4 = 1'b1;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_D5 = 1'b1;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_D6 = 1'b1;
  assign CLBLM_R_X7Y157_SLICE_X9Y157_C5 = 1'b1;
  assign CLBLM_R_X7Y157_SLICE_X9Y157_C6 = 1'b1;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_A2 = CLBLM_L_X10Y151_SLICE_X13Y151_CQ;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_A3 = CLBLM_L_X12Y147_SLICE_X16Y147_AQ;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_A4 = CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_A5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_A6 = CLBLM_L_X12Y146_SLICE_X16Y146_AQ;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_B1 = 1'b1;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_B2 = 1'b1;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_B3 = 1'b1;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_B4 = 1'b1;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_B5 = 1'b1;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_B6 = 1'b1;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_C1 = 1'b1;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_C2 = 1'b1;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_C3 = 1'b1;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_C4 = 1'b1;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_C5 = 1'b1;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_C6 = 1'b1;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_D1 = 1'b1;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_D2 = 1'b1;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_D3 = 1'b1;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_D4 = 1'b1;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_D5 = 1'b1;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_D6 = 1'b1;
  assign LIOB33_X0Y107_IOB_X0Y108_O = CLBLM_R_X3Y152_SLICE_X2Y152_BO6;
  assign LIOB33_X0Y107_IOB_X0Y107_O = CLBLL_L_X2Y120_SLICE_X0Y120_AO6;
  assign CLBLM_R_X7Y157_SLICE_X9Y157_D5 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_SR = CLBLM_R_X11Y151_SLICE_X15Y151_CO6;
  assign LIOI3_X0Y73_ILOGIC_X0Y74_D = LIOB33_X0Y73_IOB_X0Y74_I;
  assign CLBLM_R_X7Y157_SLICE_X9Y157_D6 = 1'b1;
  assign LIOI3_X0Y73_ILOGIC_X0Y73_D = LIOB33_X0Y73_IOB_X0Y73_I;
  assign CLBLM_R_X15Y151_SLICE_X21Y151_A1 = 1'b1;
  assign CLBLM_R_X15Y151_SLICE_X21Y151_A2 = 1'b1;
  assign CLBLM_R_X15Y151_SLICE_X21Y151_A3 = 1'b1;
  assign CLBLM_R_X15Y151_SLICE_X21Y151_A4 = 1'b1;
  assign CLBLM_R_X15Y151_SLICE_X21Y151_A5 = 1'b1;
  assign CLBLM_R_X15Y151_SLICE_X21Y151_A6 = 1'b1;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_AX = CLBLM_L_X10Y147_SLICE_X12Y147_BO6;
  assign CLBLM_R_X15Y151_SLICE_X21Y151_B2 = 1'b1;
  assign CLBLM_R_X15Y151_SLICE_X21Y151_B3 = 1'b1;
  assign CLBLM_R_X15Y151_SLICE_X21Y151_B4 = 1'b1;
  assign CLBLM_R_X15Y151_SLICE_X21Y151_B5 = 1'b1;
  assign CLBLM_R_X15Y151_SLICE_X21Y151_B6 = 1'b1;
  assign CLBLM_R_X15Y151_SLICE_X21Y151_B1 = 1'b1;
  assign RIOB33_X105Y193_IOB_X1Y193_O = CLBLM_R_X11Y153_SLICE_X14Y153_AQ;
  assign RIOB33_X105Y193_IOB_X1Y194_O = CLBLM_L_X12Y155_SLICE_X17Y155_AQ;
  assign CLBLM_R_X15Y151_SLICE_X21Y151_C1 = 1'b1;
  assign CLBLM_R_X15Y151_SLICE_X21Y151_C2 = 1'b1;
  assign CLBLM_R_X15Y151_SLICE_X21Y151_C3 = 1'b1;
  assign CLBLM_R_X15Y151_SLICE_X21Y151_C4 = 1'b1;
  assign CLBLM_R_X7Y157_SLICE_X8Y157_D2 = 1'b1;
  assign CLBLM_R_X15Y151_SLICE_X21Y151_C5 = 1'b1;
  assign CLBLM_R_X15Y151_SLICE_X21Y151_C6 = 1'b1;
  assign CLBLM_R_X15Y151_SLICE_X21Y151_D1 = 1'b1;
  assign CLBLM_R_X15Y151_SLICE_X21Y151_D2 = 1'b1;
  assign CLBLM_R_X15Y151_SLICE_X21Y151_D3 = 1'b1;
  assign CLBLM_R_X15Y151_SLICE_X21Y151_D4 = 1'b1;
  assign CLBLM_R_X15Y151_SLICE_X21Y151_D5 = 1'b1;
  assign CLBLM_R_X15Y151_SLICE_X21Y151_D6 = 1'b1;
  assign CLBLM_R_X15Y151_SLICE_X20Y151_A1 = 1'b1;
  assign CLBLM_R_X7Y157_SLICE_X8Y157_D3 = 1'b1;
  assign CLBLM_R_X15Y151_SLICE_X20Y151_A2 = 1'b1;
  assign CLBLM_R_X15Y151_SLICE_X20Y151_A3 = 1'b1;
  assign CLBLM_R_X15Y151_SLICE_X20Y151_A4 = 1'b1;
  assign CLBLM_R_X15Y151_SLICE_X20Y151_A5 = 1'b1;
  assign CLBLM_R_X15Y151_SLICE_X20Y151_A6 = 1'b1;
  assign CLBLM_R_X15Y151_SLICE_X20Y151_AX = CLBLM_R_X15Y153_SLICE_X20Y153_AO5;
  assign CLBLM_R_X15Y151_SLICE_X20Y151_B1 = 1'b1;
  assign CLBLM_R_X15Y151_SLICE_X20Y151_B2 = 1'b1;
  assign CLBLM_R_X15Y151_SLICE_X20Y151_B3 = 1'b1;
  assign CLBLM_R_X15Y151_SLICE_X20Y151_B4 = 1'b1;
  assign CLBLM_R_X15Y151_SLICE_X20Y151_B5 = 1'b1;
  assign CLBLM_R_X15Y151_SLICE_X20Y151_B6 = 1'b1;
  assign CLBLM_R_X15Y151_SLICE_X20Y151_C1 = 1'b1;
  assign CLBLM_R_X15Y151_SLICE_X20Y151_C2 = 1'b1;
  assign CLBLM_R_X15Y151_SLICE_X20Y151_C3 = 1'b1;
  assign CLBLM_R_X15Y151_SLICE_X20Y151_C4 = 1'b1;
  assign CLBLM_R_X15Y151_SLICE_X20Y151_C5 = 1'b1;
  assign CLBLM_R_X15Y151_SLICE_X20Y151_C6 = 1'b1;
  assign CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_I = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLM_R_X15Y151_SLICE_X20Y151_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X15Y151_SLICE_X20Y151_D1 = 1'b1;
  assign CLBLM_R_X15Y151_SLICE_X20Y151_D2 = 1'b1;
  assign CLBLM_R_X15Y151_SLICE_X20Y151_D3 = 1'b1;
  assign CLBLM_R_X15Y151_SLICE_X20Y151_D4 = 1'b1;
  assign CLBLM_R_X15Y151_SLICE_X20Y151_D5 = 1'b1;
  assign CLBLM_R_X15Y151_SLICE_X20Y151_D6 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_A1 = CLBLM_R_X3Y153_SLICE_X3Y153_DO6;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_A2 = CLBLM_R_X3Y155_SLICE_X3Y155_BO6;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_A3 = CLBLL_L_X4Y154_SLICE_X5Y154_DO6;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_A4 = CLBLM_R_X3Y153_SLICE_X3Y153_BO6;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_A5 = CLBLL_L_X4Y153_SLICE_X4Y153_BO6;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_A6 = CLBLM_R_X3Y150_SLICE_X3Y150_DO6;
  assign CLBLM_R_X7Y157_SLICE_X8Y157_D5 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_B1 = CLBLL_L_X2Y154_SLICE_X1Y154_BO5;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_B2 = CLBLM_R_X5Y152_SLICE_X7Y152_CQ;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_B3 = CLBLL_L_X2Y151_SLICE_X0Y151_CO5;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_B4 = CLBLL_L_X2Y152_SLICE_X1Y152_AO5;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_B5 = LIOB33_X0Y65_IOB_X0Y66_I;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_B6 = CLBLM_R_X3Y152_SLICE_X2Y152_BO5;
  assign CLBLM_R_X7Y157_SLICE_X8Y157_B5 = 1'b1;
  assign CLBLM_R_X7Y157_SLICE_X8Y157_B6 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_C1 = LIOB33_X0Y65_IOB_X0Y66_I;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_C2 = CLBLL_L_X4Y151_SLICE_X5Y151_BQ;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_C3 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_C4 = CLBLL_L_X2Y152_SLICE_X1Y152_AO5;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_C5 = CLBLL_L_X2Y154_SLICE_X1Y154_BO5;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_C6 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X7Y157_SLICE_X8Y157_D6 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X1Y134_A4 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X1Y134_A5 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_D1 = CLBLL_L_X2Y151_SLICE_X1Y151_AO6;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_D2 = CLBLM_R_X3Y148_SLICE_X2Y148_DQ;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_D3 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_D4 = CLBLL_L_X2Y155_SLICE_X1Y155_DO6;
  assign CLBLL_L_X2Y134_SLICE_X1Y134_A6 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_D5 = CLBLM_R_X3Y145_SLICE_X2Y145_AQ;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_D6 = CLBLL_L_X4Y155_SLICE_X4Y155_BO6;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_C1 = CLBLM_R_X7Y154_SLICE_X8Y154_BQ;
  assign LIOI3_X0Y155_OLOGIC_X0Y155_D1 = LIOB33_X0Y69_IOB_X0Y70_I;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_A1 = CLBLL_L_X2Y152_SLICE_X1Y152_BO5;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_A2 = CLBLL_L_X4Y151_SLICE_X5Y151_CO6;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_A3 = CLBLM_R_X3Y153_SLICE_X3Y153_AO6;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_A4 = CLBLL_L_X2Y153_SLICE_X1Y153_AO6;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_A5 = CLBLL_L_X2Y155_SLICE_X1Y155_AO6;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_A6 = CLBLM_R_X3Y156_SLICE_X2Y156_CO6;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_B1 = CLBLL_L_X2Y151_SLICE_X0Y151_AO6;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_B2 = CLBLM_R_X3Y152_SLICE_X2Y152_AO5;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_B3 = CLBLM_R_X3Y153_SLICE_X3Y153_CO6;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_B4 = CLBLM_R_X5Y152_SLICE_X7Y152_CQ;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_B5 = CLBLM_R_X3Y145_SLICE_X2Y145_AQ;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_B6 = CLBLM_R_X3Y153_SLICE_X2Y153_CO6;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_C2 = CLBLM_R_X7Y155_SLICE_X8Y155_AQ;
  assign CLBLM_R_X7Y157_SLICE_X8Y157_C4 = 1'b1;
  assign CLBLM_R_X7Y157_SLICE_X8Y157_C5 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_C1 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_C2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_C3 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_L_X16Y158_SLICE_X23Y158_A1 = 1'b1;
  assign CLBLM_L_X16Y158_SLICE_X23Y158_A2 = 1'b1;
  assign CLBLM_L_X16Y158_SLICE_X23Y158_A3 = 1'b1;
  assign CLBLM_L_X16Y158_SLICE_X23Y158_A4 = 1'b1;
  assign CLBLM_L_X16Y158_SLICE_X23Y158_A5 = 1'b1;
  assign CLBLM_L_X16Y158_SLICE_X23Y158_A6 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X1Y134_B3 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X1Y134_B4 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_C4 = CLBLL_L_X2Y155_SLICE_X1Y155_DO6;
  assign CLBLM_L_X16Y158_SLICE_X23Y158_B1 = 1'b1;
  assign CLBLM_L_X16Y158_SLICE_X23Y158_B2 = 1'b1;
  assign CLBLM_L_X16Y158_SLICE_X23Y158_B3 = 1'b1;
  assign CLBLM_L_X16Y158_SLICE_X23Y158_B4 = 1'b1;
  assign CLBLM_L_X16Y158_SLICE_X23Y158_B5 = 1'b1;
  assign CLBLM_L_X16Y158_SLICE_X23Y158_B6 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X1Y134_B5 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X1Y134_B6 = 1'b1;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_A1 = 1'b1;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_A2 = 1'b1;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_A3 = 1'b1;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_A4 = 1'b1;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_A5 = 1'b1;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_A6 = 1'b1;
  assign CLBLM_L_X16Y158_SLICE_X23Y158_C1 = 1'b1;
  assign CLBLM_L_X16Y158_SLICE_X23Y158_C2 = 1'b1;
  assign CLBLM_L_X16Y158_SLICE_X23Y158_C3 = 1'b1;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_B1 = 1'b1;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_B2 = 1'b1;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_B3 = 1'b1;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_B4 = 1'b1;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_B5 = 1'b1;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_B6 = 1'b1;
  assign CLBLM_L_X16Y158_SLICE_X23Y158_D1 = 1'b1;
  assign CLBLM_L_X16Y158_SLICE_X23Y158_D2 = 1'b1;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_C1 = 1'b1;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_C2 = 1'b1;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_C3 = 1'b1;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_C4 = 1'b1;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_C5 = 1'b1;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_C6 = 1'b1;
  assign CLBLM_L_X16Y158_SLICE_X23Y158_D3 = 1'b1;
  assign CLBLM_L_X16Y158_SLICE_X23Y158_D4 = 1'b1;
  assign CLBLM_L_X16Y158_SLICE_X22Y158_A1 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_L_X16Y158_SLICE_X23Y158_D6 = 1'b1;
  assign CLBLM_L_X16Y158_SLICE_X22Y158_A2 = 1'b1;
  assign CLBLM_L_X16Y158_SLICE_X22Y158_A3 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLM_L_X16Y158_SLICE_X22Y158_A4 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_D1 = 1'b1;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_D2 = 1'b1;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_D3 = 1'b1;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_D4 = 1'b1;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_D5 = 1'b1;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_D6 = 1'b1;
  assign CLBLM_L_X16Y158_SLICE_X22Y158_A5 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLM_L_X16Y158_SLICE_X22Y158_A6 = 1'b1;
  assign CLBLM_L_X16Y158_SLICE_X22Y158_B1 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_A1 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_A2 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_A3 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_A4 = CLBLL_L_X2Y141_SLICE_X0Y141_BO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_A5 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_A6 = 1'b1;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_A1 = CLBLM_L_X10Y151_SLICE_X12Y151_BQ;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_A2 = CLBLM_L_X10Y152_SLICE_X12Y152_DQ;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_A3 = CLBLM_L_X12Y148_SLICE_X16Y148_AQ;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_B1 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_B2 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_B3 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_B4 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_B5 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_B6 = 1'b1;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_A6 = CLBLM_R_X11Y147_SLICE_X14Y147_CO6;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_C1 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_C2 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_C3 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_C4 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_C5 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_C6 = 1'b1;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_B5 = CLBLM_L_X12Y149_SLICE_X16Y149_AQ;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_C1 = CLBLM_L_X8Y144_SLICE_X10Y144_AQ;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_C2 = 1'b1;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_C3 = 1'b1;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_C4 = CLBLM_L_X8Y151_SLICE_X11Y151_CQ;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_C5 = CLBLM_L_X10Y145_SLICE_X12Y145_BQ;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_D1 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_D2 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_D3 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_D4 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_D5 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_D6 = 1'b1;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_D1 = 1'b1;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_D2 = 1'b1;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_D3 = 1'b1;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_D4 = 1'b1;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_D5 = 1'b1;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_D6 = 1'b1;
  assign RIOB33_X105Y195_IOB_X1Y196_O = CLBLM_R_X11Y153_SLICE_X14Y153_BQ;
  assign RIOB33_X105Y195_IOB_X1Y195_O = CLBLM_R_X11Y151_SLICE_X14Y151_AQ;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_A1 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_A2 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_A3 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_A4 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_A5 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_A6 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_B1 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_B2 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_B3 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_B4 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_B5 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_B6 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_C1 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_C2 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_C3 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_C4 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_C5 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_C6 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_D1 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_D2 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_D3 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_D4 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_D5 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_D6 = 1'b1;
  assign LIOI3_X0Y53_ILOGIC_X0Y53_D = LIOB33_X0Y53_IOB_X0Y53_I;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_D3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOB33_SING_X0Y149_IOB_X0Y149_O = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_D4 = CLBLL_L_X2Y151_SLICE_X1Y151_BO6;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_A4 = CLBLM_R_X11Y148_SLICE_X14Y148_AQ;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_A1 = CLBLL_L_X2Y150_SLICE_X1Y150_CO6;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_A2 = CLBLM_R_X5Y154_SLICE_X7Y154_DO6;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_A3 = CLBLM_R_X3Y155_SLICE_X2Y155_DO6;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_A4 = CLBLM_R_X3Y154_SLICE_X3Y154_BO6;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_A5 = CLBLL_L_X4Y154_SLICE_X4Y154_BO6;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_A6 = CLBLM_R_X3Y155_SLICE_X2Y155_AO6;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_T1 = 1'b1;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_B1 = CLBLL_L_X4Y155_SLICE_X4Y155_CO6;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_B2 = CLBLL_L_X2Y154_SLICE_X1Y154_AO5;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_B3 = CLBLM_R_X3Y154_SLICE_X2Y154_AO6;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_B4 = CLBLM_R_X3Y149_SLICE_X2Y149_AQ;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_B5 = CLBLM_R_X3Y154_SLICE_X3Y154_CO6;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_B6 = CLBLL_L_X4Y151_SLICE_X4Y151_DO6;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_C1 = CLBLL_L_X2Y154_SLICE_X1Y154_BO5;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_C2 = CLBLL_L_X4Y155_SLICE_X4Y155_BO6;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_C3 = 1'b1;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_C4 = CLBLM_R_X3Y149_SLICE_X3Y149_CQ;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_C5 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_C6 = CLBLL_L_X2Y152_SLICE_X1Y152_AO6;
  assign LIOI3_X0Y155_OLOGIC_X0Y155_T1 = 1'b1;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_D1 = CLBLM_R_X3Y150_SLICE_X3Y150_DO6;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_D2 = CLBLL_L_X2Y154_SLICE_X1Y154_BO6;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_D3 = 1'b1;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_D4 = CLBLL_L_X4Y150_SLICE_X5Y150_BQ;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_D5 = CLBLL_L_X4Y155_SLICE_X5Y155_AO6;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_D6 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_B1 = CLBLM_R_X11Y143_SLICE_X14Y143_BQ;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_B2 = CLBLM_R_X11Y145_SLICE_X14Y145_BQ;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_A1 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_A2 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_A3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_A4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_A5 = CLBLM_R_X7Y153_SLICE_X9Y153_BQ;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_A6 = CLBLL_L_X2Y155_SLICE_X1Y155_DO6;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_B3 = CLBLL_L_X4Y145_SLICE_X5Y145_DO6;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_B1 = CLBLM_R_X3Y154_SLICE_X2Y154_DO6;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_B2 = CLBLM_R_X3Y155_SLICE_X2Y155_BO6;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_B3 = CLBLL_L_X4Y152_SLICE_X5Y152_AO6;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_B4 = CLBLM_R_X3Y156_SLICE_X2Y156_BO6;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_B5 = CLBLM_R_X7Y153_SLICE_X9Y153_BQ;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_B6 = CLBLM_R_X3Y154_SLICE_X2Y154_CO6;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_B6 = 1'b1;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_C1 = LIOB33_X0Y67_IOB_X0Y68_I;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_C2 = CLBLL_L_X2Y154_SLICE_X1Y154_AO5;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_C3 = CLBLM_R_X3Y149_SLICE_X2Y149_AQ;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_C4 = 1'b1;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_C5 = CLBLL_L_X4Y155_SLICE_X4Y155_DO6;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_C6 = CLBLL_L_X2Y151_SLICE_X0Y151_BO6;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_D1 = CLBLL_L_X4Y151_SLICE_X4Y151_DO6;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_D2 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_D3 = CLBLM_R_X3Y149_SLICE_X3Y149_CQ;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_D4 = CLBLL_L_X2Y154_SLICE_X1Y154_BO6;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_D5 = 1'b1;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_D6 = CLBLL_L_X2Y152_SLICE_X1Y152_BO5;
  assign LIOI3_X0Y197_OLOGIC_X0Y198_D1 = LIOB33_X0Y73_IOB_X0Y73_I;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_A1 = CLBLM_R_X11Y152_SLICE_X14Y152_DQ;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_A2 = CLBLM_L_X12Y148_SLICE_X16Y148_BQ;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_A5 = CLBLM_R_X11Y147_SLICE_X14Y147_CO6;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_A6 = CLBLM_L_X12Y149_SLICE_X17Y149_AQ;
  assign LIOI3_X0Y197_OLOGIC_X0Y198_T1 = 1'b1;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_B1 = CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_B2 = CLBLM_L_X12Y149_SLICE_X17Y149_BQ;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_B4 = CLBLM_R_X11Y147_SLICE_X14Y147_CO6;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_B6 = CLBLM_L_X12Y149_SLICE_X17Y149_AQ;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_B6 = CLBLM_R_X3Y146_SLICE_X3Y146_CQ;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_D1 = CLBLL_L_X2Y145_SLICE_X1Y145_AQ;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_C1 = CLBLM_L_X12Y150_SLICE_X16Y150_BQ;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_C2 = CLBLM_L_X12Y149_SLICE_X17Y149_CQ;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_C4 = CLBLM_R_X7Y151_SLICE_X9Y151_AQ;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_C5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_C6 = CLBLM_R_X11Y147_SLICE_X14Y147_CO6;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_C5 = CLBLM_L_X10Y145_SLICE_X13Y145_A5Q;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_C6 = CLBLM_R_X7Y142_SLICE_X8Y142_DO6;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_T1 = 1'b1;
  assign RIOI3_X105Y179_OLOGIC_X1Y180_D1 = CLBLM_R_X11Y151_SLICE_X14Y151_DO6;
  assign LIOI3_X0Y197_OLOGIC_X0Y197_T1 = 1'b1;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_D1 = 1'b1;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_D2 = 1'b1;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_D3 = 1'b1;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_D4 = 1'b1;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_D5 = 1'b1;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_D6 = 1'b1;
  assign LIOB33_X0Y111_IOB_X0Y111_O = 1'b0;
  assign LIOB33_X0Y111_IOB_X0Y112_O = CLBLM_R_X11Y148_SLICE_X15Y148_B5Q;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_D1 = CLBLM_R_X3Y142_SLICE_X2Y142_BQ;
  assign RIOI3_X105Y179_OLOGIC_X1Y180_T1 = 1'b1;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_A1 = CLBLL_L_X4Y143_SLICE_X4Y143_BQ;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_A2 = CLBLM_R_X11Y147_SLICE_X14Y147_CO6;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_A3 = CLBLM_L_X12Y149_SLICE_X16Y149_AQ;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_A6 = CLBLM_L_X12Y149_SLICE_X17Y149_CQ;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_T1 = 1'b1;
  assign RIOI3_X105Y179_OLOGIC_X1Y179_D1 = CLBLM_R_X103Y178_SLICE_X163Y178_AO5;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_B1 = CLBLM_L_X12Y149_SLICE_X16Y149_DO6;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_B2 = 1'b1;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_B3 = 1'b1;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_B4 = CLBLM_R_X11Y149_SLICE_X14Y149_AQ;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_B5 = CLBLM_L_X10Y145_SLICE_X12Y145_BQ;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_B6 = CLBLM_L_X12Y149_SLICE_X16Y149_CO6;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_D1 = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign RIOI3_X105Y179_OLOGIC_X1Y179_T1 = 1'b1;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_C1 = CLBLM_L_X12Y150_SLICE_X16Y150_BQ;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_C2 = 1'b1;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_C3 = CLBLM_L_X8Y151_SLICE_X11Y151_CQ;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_C4 = CLBLM_L_X10Y150_SLICE_X12Y150_AQ;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_C5 = 1'b1;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_C6 = CLBLM_L_X8Y144_SLICE_X10Y144_AQ;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_T1 = 1'b1;
  assign RIOB33_X105Y197_IOB_X1Y198_O = CLBLM_L_X16Y158_SLICE_X22Y158_AO6;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOB33_X105Y197_IOB_X1Y197_O = CLBLM_L_X16Y158_SLICE_X22Y158_AO6;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_D1 = RIOB33_X105Y121_IOB_X1Y122_I;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_D1 = CLBLM_R_X7Y146_SLICE_X9Y146_BQ;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_D2 = CLBLL_L_X4Y148_SLICE_X5Y148_BQ;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_D3 = CLBLM_L_X10Y151_SLICE_X12Y151_BQ;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_D4 = CLBLM_L_X12Y149_SLICE_X17Y149_CQ;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_D5 = 1'b1;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_D6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_T1 = 1'b1;
  assign CLBLM_R_X5Y155_SLICE_X7Y155_D2 = CLBLM_R_X5Y152_SLICE_X6Y152_AQ;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_B1 = CLBLM_R_X7Y147_SLICE_X8Y147_CQ;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_B2 = CLBLM_R_X7Y153_SLICE_X8Y153_DQ;
  assign CLBLM_R_X15Y153_SLICE_X21Y153_A1 = 1'b1;
  assign CLBLM_R_X15Y153_SLICE_X21Y153_A2 = 1'b1;
  assign CLBLM_R_X15Y153_SLICE_X21Y153_A3 = 1'b1;
  assign CLBLM_R_X15Y153_SLICE_X21Y153_A4 = 1'b1;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_B3 = CLBLM_R_X11Y153_SLICE_X14Y153_AO6;
  assign CLBLM_R_X15Y153_SLICE_X21Y153_A5 = 1'b1;
  assign CLBLM_R_X15Y153_SLICE_X21Y153_A6 = 1'b1;
  assign CLBLM_R_X15Y153_SLICE_X21Y153_B1 = 1'b1;
  assign CLBLM_R_X15Y153_SLICE_X21Y153_B2 = 1'b1;
  assign CLBLM_R_X15Y153_SLICE_X21Y153_B3 = 1'b1;
  assign CLBLM_R_X15Y153_SLICE_X21Y153_B4 = 1'b1;
  assign CLBLM_R_X15Y153_SLICE_X21Y153_B5 = 1'b1;
  assign CLBLM_R_X15Y153_SLICE_X21Y153_B6 = 1'b1;
  assign CLBLM_R_X15Y153_SLICE_X21Y153_C1 = 1'b1;
  assign CLBLM_R_X15Y153_SLICE_X21Y153_C2 = 1'b1;
  assign CLBLM_R_X15Y153_SLICE_X21Y153_C3 = 1'b1;
  assign CLBLM_R_X15Y153_SLICE_X21Y153_C4 = 1'b1;
  assign CLBLM_R_X15Y153_SLICE_X21Y153_C5 = 1'b1;
  assign CLBLM_R_X15Y153_SLICE_X21Y153_C6 = 1'b1;
  assign CLBLM_R_X15Y153_SLICE_X21Y153_D1 = 1'b1;
  assign CLBLM_R_X15Y153_SLICE_X21Y153_D2 = 1'b1;
  assign CLBLM_R_X15Y153_SLICE_X21Y153_D3 = 1'b1;
  assign CLBLM_R_X15Y153_SLICE_X21Y153_D4 = 1'b1;
  assign CLBLM_R_X15Y153_SLICE_X21Y153_D5 = 1'b1;
  assign CLBLM_R_X15Y153_SLICE_X21Y153_D6 = 1'b1;
  assign CLBLM_R_X15Y153_SLICE_X20Y153_A1 = 1'b1;
  assign CLBLM_R_X15Y153_SLICE_X20Y153_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X15Y153_SLICE_X20Y153_A3 = CLBLM_L_X10Y150_SLICE_X12Y150_C5Q;
  assign CLBLM_R_X15Y153_SLICE_X20Y153_A4 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_R_X15Y153_SLICE_X20Y153_A5 = CLBLM_R_X11Y153_SLICE_X14Y153_AQ;
  assign CLBLM_R_X15Y153_SLICE_X20Y153_A6 = 1'b1;
  assign CLBLM_R_X15Y153_SLICE_X20Y153_B1 = 1'b1;
  assign CLBLM_R_X15Y153_SLICE_X20Y153_B2 = 1'b1;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_C2 = CLBLM_R_X7Y153_SLICE_X8Y153_CQ;
  assign CLBLM_R_X15Y153_SLICE_X20Y153_B3 = 1'b1;
  assign CLBLM_R_X15Y153_SLICE_X20Y153_B4 = 1'b1;
  assign CLBLM_R_X15Y153_SLICE_X20Y153_B5 = 1'b1;
  assign CLBLM_R_X15Y153_SLICE_X20Y153_B6 = 1'b1;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_C5 = CLBLM_R_X7Y147_SLICE_X8Y147_B5Q;
  assign CLBLM_R_X15Y153_SLICE_X20Y153_C1 = 1'b1;
  assign CLBLM_R_X15Y153_SLICE_X20Y153_C2 = 1'b1;
  assign CLBLM_R_X15Y153_SLICE_X20Y153_C3 = 1'b1;
  assign CLBLM_R_X15Y153_SLICE_X20Y153_C4 = 1'b1;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_C6 = 1'b1;
  assign CLBLM_R_X15Y153_SLICE_X20Y153_C5 = 1'b1;
  assign CLBLM_R_X15Y153_SLICE_X20Y153_C6 = 1'b1;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_C3 = CLBLM_R_X3Y143_SLICE_X3Y143_AQ;
  assign CLBLM_R_X15Y153_SLICE_X20Y153_D1 = 1'b1;
  assign CLBLM_R_X15Y153_SLICE_X20Y153_D2 = 1'b1;
  assign CLBLM_R_X15Y153_SLICE_X20Y153_D3 = 1'b1;
  assign CLBLM_R_X15Y153_SLICE_X20Y153_D4 = 1'b1;
  assign CLBLM_R_X15Y153_SLICE_X20Y153_D5 = 1'b1;
  assign CLBLM_R_X15Y153_SLICE_X20Y153_D6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_D1 = CLBLM_L_X10Y146_SLICE_X13Y146_BQ;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_A1 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_A2 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_A3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_A4 = CLBLL_L_X2Y155_SLICE_X1Y155_DO6;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_A5 = 1'b1;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_A6 = 1'b1;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_B1 = CLBLL_L_X4Y150_SLICE_X5Y150_BQ;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_B2 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_B3 = CLBLL_L_X2Y154_SLICE_X1Y154_BO5;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_B4 = CLBLL_L_X4Y155_SLICE_X4Y155_AO5;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_B5 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_B6 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_C4 = CLBLM_L_X10Y156_SLICE_X12Y156_CO6;
  assign LIOI3_X0Y75_ILOGIC_X0Y76_D = LIOB33_X0Y75_IOB_X0Y76_I;
  assign LIOI3_X0Y75_ILOGIC_X0Y75_D = LIOB33_X0Y75_IOB_X0Y75_I;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_C1 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_C2 = CLBLL_L_X2Y152_SLICE_X1Y152_AO5;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_C3 = CLBLL_L_X2Y155_SLICE_X1Y155_DO6;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_C4 = CLBLM_L_X16Y158_SLICE_X22Y158_AO5;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_C5 = CLBLM_R_X3Y155_SLICE_X3Y155_DO6;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_C6 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign RIOI3_X105Y121_ILOGIC_X1Y122_D = RIOB33_X105Y121_IOB_X1Y122_I;
  assign RIOI3_X105Y121_ILOGIC_X1Y121_D = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_D1 = 1'b1;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_D2 = 1'b1;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_D3 = 1'b1;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_D4 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_D5 = 1'b1;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_D6 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_A1 = CLBLM_R_X3Y156_SLICE_X2Y156_CO6;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_A2 = CLBLL_L_X4Y155_SLICE_X4Y155_BO5;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_A3 = CLBLM_R_X3Y155_SLICE_X3Y155_CO6;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_A4 = CLBLL_L_X4Y154_SLICE_X5Y154_CO6;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_A5 = CLBLL_L_X2Y152_SLICE_X1Y152_BO5;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_A6 = CLBLL_L_X2Y154_SLICE_X1Y154_CO6;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_B1 = CLBLL_L_X2Y154_SLICE_X1Y154_CO6;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_B2 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_B3 = CLBLM_R_X3Y155_SLICE_X3Y155_AO6;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_B4 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_B5 = CLBLL_L_X2Y154_SLICE_X1Y154_CO5;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_B6 = CLBLL_L_X4Y154_SLICE_X5Y154_CO6;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_C6 = CLBLL_L_X4Y147_SLICE_X5Y147_B5Q;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_C1 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_C2 = CLBLL_L_X2Y150_SLICE_X0Y150_AO6;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_C3 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_C4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_C5 = CLBLM_R_X3Y156_SLICE_X2Y156_AO5;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_C6 = CLBLL_L_X4Y155_SLICE_X4Y155_AO5;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_D1 = CLBLL_L_X2Y152_SLICE_X1Y152_BO5;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_D2 = CLBLM_R_X3Y155_SLICE_X3Y155_CO6;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_D3 = CLBLL_L_X2Y154_SLICE_X1Y154_AO6;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_D4 = CLBLM_R_X3Y155_SLICE_X2Y155_CO6;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_D5 = CLBLL_L_X2Y154_SLICE_X1Y154_CO6;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_D6 = CLBLL_L_X4Y154_SLICE_X5Y154_CO6;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_A1 = 1'b1;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_A2 = 1'b1;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_A3 = 1'b1;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_A4 = 1'b1;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_A5 = 1'b1;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_A6 = 1'b1;
  assign LIOB33_X0Y113_IOB_X0Y113_O = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_B1 = 1'b1;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_B2 = 1'b1;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_B3 = 1'b1;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_B4 = 1'b1;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_B5 = 1'b1;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_B6 = 1'b1;
  assign LIOB33_X0Y113_IOB_X0Y114_O = CLBLM_R_X7Y143_SLICE_X8Y143_BQ;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_C1 = 1'b1;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_C2 = 1'b1;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_C3 = 1'b1;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_C4 = 1'b1;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_C5 = 1'b1;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_C6 = 1'b1;
  assign RIOI3_X105Y117_ILOGIC_X1Y118_D = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_D1 = 1'b1;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_D2 = 1'b1;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_D3 = 1'b1;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_D4 = 1'b1;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_D5 = 1'b1;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_D6 = 1'b1;
  assign RIOI3_X105Y117_ILOGIC_X1Y117_D = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_A1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_A2 = CLBLM_R_X11Y150_SLICE_X15Y150_CQ;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_A3 = CLBLM_L_X12Y150_SLICE_X16Y150_AQ;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_A4 = CLBLM_L_X12Y151_SLICE_X16Y151_AQ;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_A5 = CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_B2 = CLBLM_L_X12Y150_SLICE_X16Y150_BQ;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_B3 = CLBLM_L_X12Y148_SLICE_X16Y148_AQ;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_B4 = CLBLM_L_X12Y152_SLICE_X17Y152_BQ;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_B6 = CLBLM_R_X11Y147_SLICE_X14Y147_CO6;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_C1 = CLBLM_R_X11Y150_SLICE_X15Y150_CQ;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_C2 = CLBLM_L_X12Y150_SLICE_X16Y150_CQ;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_C3 = CLBLM_R_X11Y154_SLICE_X15Y154_CO6;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_C5 = CLBLM_L_X12Y151_SLICE_X16Y151_CQ;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_C6 = CLBLM_L_X12Y150_SLICE_X16Y150_DO5;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_D1 = CLBLM_L_X10Y149_SLICE_X13Y149_A5Q;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_D2 = CLBLM_R_X11Y151_SLICE_X15Y151_A5Q;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_D3 = CLBLM_L_X12Y151_SLICE_X16Y151_BQ;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_D4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_D5 = CLBLM_R_X7Y147_SLICE_X9Y147_AQ;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_D6 = 1'b1;
  assign LIOB33_X0Y181_IOB_X0Y181_O = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_A1 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_A2 = CLBLM_R_X11Y151_SLICE_X14Y151_BQ;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_A3 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_A4 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_A5 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_A6 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_B1 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_B2 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_B3 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_B4 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_B5 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_B6 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_C1 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_C2 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_C3 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_C4 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_C5 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_C6 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_D1 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_D2 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_D3 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_D4 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_D5 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_D6 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_A1 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_A2 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_A3 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_A4 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_A5 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_A6 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_B1 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_B2 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_B3 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_B4 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_B5 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_B6 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_C1 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_C2 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_C3 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_C4 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_C5 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_C6 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_D1 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_D2 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_D3 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_D4 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_D5 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_D6 = 1'b1;
  assign LIOB33_SING_X0Y100_IOB_X0Y100_O = CLBLL_L_X2Y138_SLICE_X0Y138_AO5;
  assign CLBLM_R_X3Y156_SLICE_X3Y156_A1 = 1'b1;
  assign CLBLM_R_X3Y156_SLICE_X3Y156_A2 = 1'b1;
  assign CLBLM_R_X3Y156_SLICE_X3Y156_A3 = 1'b1;
  assign CLBLM_R_X3Y156_SLICE_X3Y156_A4 = 1'b1;
  assign CLBLM_R_X3Y156_SLICE_X3Y156_A5 = 1'b1;
  assign CLBLM_R_X3Y156_SLICE_X3Y156_A6 = 1'b1;
  assign LIOI3_X0Y103_OLOGIC_X0Y104_T1 = 1'b1;
  assign CLBLM_R_X3Y156_SLICE_X3Y156_B1 = 1'b1;
  assign CLBLM_R_X3Y156_SLICE_X3Y156_B2 = 1'b1;
  assign CLBLM_R_X3Y156_SLICE_X3Y156_B3 = 1'b1;
  assign CLBLM_R_X3Y156_SLICE_X3Y156_B4 = 1'b1;
  assign CLBLM_R_X3Y156_SLICE_X3Y156_B5 = 1'b1;
  assign CLBLM_R_X3Y156_SLICE_X3Y156_B6 = 1'b1;
  assign CLBLM_R_X3Y156_SLICE_X3Y156_C1 = 1'b1;
  assign CLBLM_R_X3Y156_SLICE_X3Y156_C2 = 1'b1;
  assign CLBLM_R_X3Y156_SLICE_X3Y156_C3 = 1'b1;
  assign CLBLM_R_X3Y156_SLICE_X3Y156_C4 = 1'b1;
  assign CLBLM_R_X3Y156_SLICE_X3Y156_C5 = 1'b1;
  assign CLBLM_R_X3Y156_SLICE_X3Y156_C6 = 1'b1;
  assign CLBLM_R_X3Y156_SLICE_X3Y156_D1 = 1'b1;
  assign CLBLM_R_X3Y156_SLICE_X3Y156_D2 = 1'b1;
  assign CLBLM_R_X3Y156_SLICE_X3Y156_D3 = 1'b1;
  assign CLBLM_R_X3Y156_SLICE_X3Y156_D4 = 1'b1;
  assign CLBLM_R_X3Y156_SLICE_X3Y156_D5 = 1'b1;
  assign CLBLM_R_X3Y156_SLICE_X3Y156_D6 = 1'b1;
  assign LIOI3_X0Y77_ILOGIC_X0Y78_D = LIOB33_X0Y77_IOB_X0Y78_I;
  assign CLBLM_R_X3Y156_SLICE_X2Y156_A1 = 1'b1;
  assign CLBLM_R_X3Y156_SLICE_X2Y156_A2 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y156_SLICE_X2Y156_A3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y156_SLICE_X2Y156_A4 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y156_SLICE_X2Y156_A5 = 1'b1;
  assign CLBLM_R_X3Y156_SLICE_X2Y156_A6 = 1'b1;
  assign CLBLM_R_X3Y156_SLICE_X2Y156_B1 = CLBLL_L_X2Y152_SLICE_X1Y152_AO6;
  assign CLBLM_R_X3Y156_SLICE_X2Y156_B2 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y156_SLICE_X2Y156_B3 = CLBLM_R_X3Y156_SLICE_X2Y156_CO6;
  assign CLBLM_R_X3Y156_SLICE_X2Y156_B4 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y156_SLICE_X2Y156_B5 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y156_SLICE_X2Y156_B6 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign LIOI3_X0Y103_OLOGIC_X0Y103_D1 = CLBLL_L_X2Y141_SLICE_X0Y141_AO6;
  assign LIOI3_X0Y77_ILOGIC_X0Y77_D = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y156_SLICE_X2Y156_C1 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X3Y156_SLICE_X2Y156_C2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y156_SLICE_X2Y156_C3 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X3Y156_SLICE_X2Y156_C4 = CLBLM_R_X3Y156_SLICE_X2Y156_AO5;
  assign CLBLM_R_X3Y156_SLICE_X2Y156_C5 = CLBLM_L_X16Y158_SLICE_X22Y158_AO5;
  assign CLBLM_R_X3Y156_SLICE_X2Y156_C6 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign LIOB33_X0Y115_IOB_X0Y115_O = CLBLM_R_X11Y148_SLICE_X15Y148_BQ;
  assign LIOB33_X0Y115_IOB_X0Y116_O = CLBLM_L_X8Y142_SLICE_X10Y142_AQ;
  assign CLBLM_R_X3Y156_SLICE_X2Y156_D1 = 1'b1;
  assign CLBLM_R_X3Y156_SLICE_X2Y156_D2 = 1'b1;
  assign CLBLM_R_X3Y156_SLICE_X2Y156_D3 = 1'b1;
  assign CLBLM_R_X3Y156_SLICE_X2Y156_D4 = 1'b1;
  assign CLBLM_R_X3Y156_SLICE_X2Y156_D5 = 1'b1;
  assign CLBLM_R_X3Y156_SLICE_X2Y156_D6 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_A1 = CLBLM_R_X13Y151_SLICE_X18Y151_AO6;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_A2 = CLBLM_L_X12Y153_SLICE_X16Y153_DO6;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_A3 = CLBLM_R_X11Y153_SLICE_X14Y153_CO5;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_A4 = CLBLM_L_X12Y152_SLICE_X17Y152_BQ;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_A5 = CLBLM_R_X13Y151_SLICE_X18Y151_BO6;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_A6 = CLBLM_R_X11Y152_SLICE_X14Y152_CQ;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_B1 = CLBLM_R_X13Y151_SLICE_X18Y151_AO6;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_B2 = CLBLM_L_X12Y152_SLICE_X17Y152_BQ;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_B3 = CLBLM_R_X11Y153_SLICE_X14Y153_CO5;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_B4 = CLBLM_R_X11Y152_SLICE_X14Y152_BQ;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_B5 = CLBLM_R_X13Y151_SLICE_X18Y151_BO6;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_B6 = CLBLM_L_X12Y153_SLICE_X16Y153_DO6;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_A1 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_A2 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_C3 = CLBLM_L_X12Y152_SLICE_X17Y152_CQ;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_C4 = CLBLM_L_X10Y151_SLICE_X13Y151_CQ;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_C5 = CLBLM_L_X12Y151_SLICE_X17Y151_DO6;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_C6 = CLBLM_R_X13Y151_SLICE_X18Y151_CO6;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_A3 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_A4 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_A5 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_A6 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_B1 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_B2 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_B3 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_B4 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_B5 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_B6 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_D1 = CLBLM_L_X12Y154_SLICE_X16Y154_AQ;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_D5 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_D6 = CLBLM_L_X12Y152_SLICE_X17Y152_BQ;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_D2 = CLBLM_L_X12Y152_SLICE_X16Y152_AQ;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_C1 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_C2 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_C3 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_C4 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_C5 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_C6 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_A1 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_A2 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_A3 = CLBLM_L_X12Y151_SLICE_X16Y151_AQ;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_A5 = CLBLM_R_X5Y142_SLICE_X7Y142_AQ;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_A6 = CLBLM_L_X8Y152_SLICE_X10Y152_CQ;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_D1 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_D2 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_D3 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_D4 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_D5 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_D6 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_B1 = CLBLM_R_X11Y154_SLICE_X15Y154_CO6;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_B2 = CLBLM_R_X11Y151_SLICE_X14Y151_AO5;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_B3 = CLBLM_R_X11Y151_SLICE_X14Y151_BQ;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_B4 = CLBLM_L_X12Y151_SLICE_X16Y151_DO5;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_B5 = CLBLM_L_X12Y151_SLICE_X16Y151_BQ;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_A1 = CLBLM_R_X7Y144_SLICE_X8Y144_DQ;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_A2 = CLBLM_L_X12Y145_SLICE_X16Y145_AQ;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_C4 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_A3 = CLBLM_L_X12Y144_SLICE_X16Y144_CQ;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_A4 = CLBLM_L_X12Y144_SLICE_X16Y144_AQ;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_A5 = CLBLM_L_X12Y144_SLICE_X16Y144_BQ;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_A6 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_C1 = CLBLL_L_X4Y149_SLICE_X4Y149_AQ;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_C2 = CLBLM_L_X12Y151_SLICE_X16Y151_CQ;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_B1 = CLBLM_L_X12Y144_SLICE_X16Y144_AQ;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_B2 = CLBLM_R_X7Y142_SLICE_X8Y142_BQ;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_B3 = CLBLM_L_X12Y144_SLICE_X16Y144_CQ;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_B4 = CLBLM_L_X12Y145_SLICE_X16Y145_AQ;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_B5 = CLBLM_L_X12Y144_SLICE_X16Y144_BQ;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_B6 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_D1 = CLBLM_L_X12Y151_SLICE_X16Y151_BQ;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_D2 = CLBLM_R_X11Y151_SLICE_X15Y151_A5Q;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_C1 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_C2 = CLBLM_L_X12Y144_SLICE_X16Y144_CQ;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_C3 = CLBLM_L_X12Y144_SLICE_X16Y144_BQ;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_C4 = CLBLM_L_X12Y144_SLICE_X16Y144_AQ;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_C5 = CLBLM_R_X11Y146_SLICE_X15Y146_AQ;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_C6 = CLBLM_L_X12Y145_SLICE_X16Y145_AQ;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_D5 = CLBLM_L_X12Y151_SLICE_X16Y151_CQ;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_D6 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_D1 = CLBLM_L_X12Y144_SLICE_X16Y144_BQ;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_D2 = CLBLM_R_X7Y142_SLICE_X8Y142_CQ;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_D3 = CLBLM_L_X12Y144_SLICE_X16Y144_CQ;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_D4 = CLBLM_L_X12Y144_SLICE_X16Y144_AQ;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_D5 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_D6 = CLBLM_L_X12Y145_SLICE_X16Y145_AQ;
  assign CLBLM_R_X103Y170_SLICE_X163Y170_A1 = CLBLM_L_X12Y152_SLICE_X17Y152_AQ;
  assign CLBLM_R_X103Y170_SLICE_X163Y170_A2 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X163Y170_A3 = CLBLM_L_X10Y155_SLICE_X13Y155_AQ;
  assign CLBLM_R_X103Y170_SLICE_X163Y170_A4 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X163Y170_A5 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_R_X103Y170_SLICE_X163Y170_A6 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X163Y170_B1 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X163Y170_B2 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X163Y170_B3 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X163Y170_B4 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X163Y170_B5 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X163Y170_B6 = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_D1 = CLBLM_R_X3Y142_SLICE_X2Y142_CQ;
  assign CLBLM_R_X103Y170_SLICE_X163Y170_C1 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X163Y170_C2 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X163Y170_C3 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X163Y170_C4 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X163Y170_C5 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X163Y170_C6 = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_T1 = 1'b1;
  assign RIOI3_X105Y183_OLOGIC_X1Y184_D1 = CLBLM_L_X10Y150_SLICE_X13Y150_DO6;
  assign CLBLM_R_X103Y170_SLICE_X163Y170_D1 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X163Y170_D2 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X163Y170_D3 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X163Y170_D4 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X163Y170_D5 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X163Y170_D6 = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_D1 = CLBLM_R_X3Y143_SLICE_X3Y143_AQ;
  assign RIOI3_X105Y183_OLOGIC_X1Y184_T1 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X162Y170_A1 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X162Y170_A2 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X162Y170_A3 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X162Y170_A4 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X162Y170_A5 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X162Y170_A6 = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_T1 = 1'b1;
  assign RIOI3_X105Y183_OLOGIC_X1Y183_D1 = CLBLM_L_X10Y152_SLICE_X13Y152_CO5;
  assign LIOB33_SING_X0Y150_IOB_X0Y150_O = LIOB33_X0Y63_IOB_X0Y63_I;
  assign CLBLM_R_X103Y170_SLICE_X162Y170_B1 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X162Y170_B2 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X162Y170_B3 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X162Y170_B4 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X162Y170_B5 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X162Y170_B6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_D1 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign RIOI3_X105Y183_OLOGIC_X1Y183_T1 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X162Y170_C1 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X162Y170_C2 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X162Y170_C3 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X162Y170_C4 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X162Y170_C5 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X162Y170_C6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_T1 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X162Y170_D1 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X162Y170_D2 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X162Y170_D3 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X162Y170_D4 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X162Y170_D5 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X162Y170_D6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_D1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_T1 = 1'b1;
  assign LIOB33_X0Y117_IOB_X0Y118_O = CLBLM_R_X3Y147_SLICE_X3Y147_CQ;
  assign LIOB33_X0Y117_IOB_X0Y117_O = CLBLM_R_X3Y144_SLICE_X2Y144_B5Q;
  assign LIOB33_SING_X0Y199_IOB_X0Y199_O = LIOB33_X0Y73_IOB_X0Y74_I;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_A2 = 1'b1;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_A3 = CLBLM_L_X12Y152_SLICE_X17Y152_CQ;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_A4 = CLBLM_L_X12Y152_SLICE_X17Y152_AQ;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_A5 = CLBLM_R_X5Y142_SLICE_X7Y142_AQ;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_A6 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_B1 = CLBLM_R_X11Y154_SLICE_X15Y154_CO5;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_B2 = 1'b1;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_B4 = CLBLM_L_X12Y151_SLICE_X17Y151_BO6;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_B5 = CLBLM_L_X10Y154_SLICE_X13Y154_CO5;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_B6 = CLBLM_R_X7Y144_SLICE_X8Y144_CQ;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_A1 = 1'b1;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_C2 = 1'b1;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_C4 = CLBLM_R_X11Y154_SLICE_X15Y154_CO5;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_C5 = CLBLM_R_X11Y148_SLICE_X14Y148_DQ;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_C6 = CLBLM_L_X12Y151_SLICE_X17Y151_CO6;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_A3 = CLBLM_L_X10Y142_SLICE_X13Y142_AQ;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_A4 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_A5 = CLBLM_L_X10Y145_SLICE_X12Y145_C5Q;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_B1 = CLBLM_L_X10Y143_SLICE_X13Y143_BQ;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_B2 = CLBLM_L_X12Y145_SLICE_X16Y145_AQ;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_B3 = CLBLM_L_X12Y144_SLICE_X16Y144_BQ;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_D1 = CLBLM_L_X12Y153_SLICE_X16Y153_DO6;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_D2 = CLBLM_R_X11Y152_SLICE_X14Y152_DQ;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_D3 = CLBLM_L_X12Y154_SLICE_X16Y154_BO5;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_D4 = CLBLM_R_X11Y153_SLICE_X15Y153_AQ;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_D5 = CLBLM_L_X12Y152_SLICE_X16Y152_BQ;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_D6 = CLBLM_R_X11Y153_SLICE_X14Y153_CO5;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_B4 = CLBLM_L_X12Y144_SLICE_X16Y144_CQ;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_B5 = CLBLM_L_X12Y144_SLICE_X16Y144_AQ;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_B6 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_C1 = CLBLM_L_X8Y145_SLICE_X11Y145_BQ;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_C2 = CLBLM_R_X5Y143_SLICE_X7Y143_BO6;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_C3 = CLBLM_R_X5Y145_SLICE_X6Y145_DO6;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_C4 = CLBLM_R_X5Y144_SLICE_X6Y144_DO6;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_C5 = CLBLM_R_X11Y143_SLICE_X14Y143_CO6;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_C6 = CLBLM_R_X7Y142_SLICE_X9Y142_AO6;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_A2 = CLBLM_L_X10Y154_SLICE_X13Y154_CO5;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_A3 = CLBLM_L_X12Y152_SLICE_X16Y152_AQ;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_D1 = CLBLM_L_X10Y145_SLICE_X12Y145_C5Q;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_D2 = CLBLM_R_X5Y144_SLICE_X6Y144_DO6;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_D3 = CLBLM_L_X10Y143_SLICE_X13Y143_CO6;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_B2 = CLBLM_R_X11Y154_SLICE_X15Y154_CO5;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_B3 = CLBLM_L_X10Y154_SLICE_X13Y154_CO5;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_B5 = 1'b1;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_B6 = CLBLM_R_X11Y147_SLICE_X15Y147_CQ;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_D4 = CLBLM_R_X3Y151_SLICE_X2Y151_AO6;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_D5 = CLBLM_R_X3Y145_SLICE_X3Y145_DQ;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_D6 = CLBLM_L_X10Y141_SLICE_X12Y141_AO6;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_A1 = CLBLM_R_X5Y145_SLICE_X6Y145_DO6;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_A2 = CLBLM_R_X15Y151_SLICE_X20Y151_AQ;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_C2 = CLBLM_R_X11Y153_SLICE_X14Y153_CO5;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_C3 = CLBLM_L_X12Y153_SLICE_X17Y153_DO6;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_C4 = CLBLM_L_X12Y153_SLICE_X16Y153_AQ;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_C5 = CLBLM_L_X12Y153_SLICE_X17Y153_CO6;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_C6 = CLBLM_L_X10Y152_SLICE_X13Y152_BQ;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_A3 = CLBLM_L_X10Y141_SLICE_X12Y141_BO5;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_A4 = CLBLM_R_X7Y142_SLICE_X9Y142_AO6;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_A5 = CLBLM_R_X5Y144_SLICE_X6Y144_DO6;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_A6 = CLBLM_R_X5Y143_SLICE_X7Y143_BO6;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_B1 = CLBLM_L_X10Y142_SLICE_X12Y142_DO6;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_B2 = CLBLM_L_X10Y142_SLICE_X13Y142_DO6;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_B3 = CLBLM_L_X10Y142_SLICE_X13Y142_CO6;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_B4 = CLBLM_L_X10Y143_SLICE_X13Y143_DO6;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_B5 = CLBLM_L_X10Y142_SLICE_X12Y142_AO6;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_B6 = CLBLM_L_X10Y142_SLICE_X12Y142_CO6;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_D2 = CLBLM_R_X11Y153_SLICE_X15Y153_AQ;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_D3 = CLBLM_L_X10Y152_SLICE_X12Y152_BQ;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_D1 = CLBLM_L_X12Y153_SLICE_X16Y153_DO6;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_C1 = CLBLM_R_X5Y144_SLICE_X6Y144_DO6;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_C2 = CLBLM_R_X5Y143_SLICE_X7Y143_BO6;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_C3 = CLBLM_R_X5Y145_SLICE_X6Y145_DO6;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_C4 = CLBLM_L_X10Y141_SLICE_X12Y141_CO6;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_C5 = CLBLM_R_X5Y144_SLICE_X7Y144_B5Q;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_C6 = CLBLM_R_X7Y142_SLICE_X9Y142_AO6;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_B2 = CLBLM_L_X12Y148_SLICE_X16Y148_BQ;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_D5 = CLBLM_L_X12Y154_SLICE_X16Y154_BO5;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_D6 = CLBLM_R_X11Y153_SLICE_X14Y153_CO5;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_B3 = CLBLM_L_X12Y150_SLICE_X16Y150_AQ;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_D = RIOB33_X105Y107_IOB_X1Y108_I;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_D = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_D1 = CLBLM_R_X5Y144_SLICE_X6Y144_DO6;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_D2 = CLBLM_R_X3Y151_SLICE_X2Y151_AO6;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_D3 = CLBLM_L_X10Y142_SLICE_X13Y142_BO5;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_D4 = CLBLM_L_X10Y145_SLICE_X13Y145_A5Q;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_D5 = CLBLM_L_X10Y141_SLICE_X12Y141_DO6;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_D6 = CLBLM_L_X8Y148_SLICE_X10Y148_BQ;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_B4 = CLBLM_R_X11Y147_SLICE_X14Y147_CO6;
  assign LIOB33_X0Y169_IOB_X0Y169_O = RIOB33_X105Y121_IOB_X1Y122_I;
  assign LIOI3_X0Y165_OLOGIC_X0Y165_T1 = 1'b1;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_C6 = CLBLL_L_X4Y148_SLICE_X5Y148_BQ;
  assign CLBLM_R_X103Y141_SLICE_X163Y141_B5 = 1'b1;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOB33_X0Y119_IOB_X0Y120_O = CLBLM_L_X10Y145_SLICE_X13Y145_AQ;
  assign LIOB33_X0Y119_IOB_X0Y119_O = CLBLM_L_X10Y146_SLICE_X13Y146_BQ;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_B2 = CLBLM_R_X11Y143_SLICE_X14Y143_BQ;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_A1 = CLBLM_R_X11Y154_SLICE_X15Y154_CO5;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_A3 = 1'b1;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_A4 = CLBLM_L_X12Y153_SLICE_X17Y153_BO6;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_A5 = CLBLM_R_X11Y154_SLICE_X15Y154_AQ;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_A6 = CLBLM_L_X10Y154_SLICE_X13Y154_CO5;
  assign RIOI3_X105Y141_ILOGIC_X1Y142_D = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_B1 = CLBLM_L_X12Y153_SLICE_X17Y153_AQ;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_B2 = CLBLM_R_X11Y153_SLICE_X14Y153_CO5;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_B3 = CLBLM_R_X13Y152_SLICE_X18Y152_AO6;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_B4 = CLBLM_L_X12Y153_SLICE_X16Y153_DO6;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_B5 = CLBLM_R_X13Y152_SLICE_X18Y152_BO6;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_B6 = CLBLM_L_X10Y154_SLICE_X13Y154_BQ;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_B3 = CLBLM_R_X11Y143_SLICE_X14Y143_AQ;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_A2 = CLBLM_L_X10Y143_SLICE_X12Y143_BO6;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_A3 = CLBLM_R_X5Y142_SLICE_X7Y142_AQ;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_C4 = CLBLM_R_X11Y154_SLICE_X15Y154_BQ;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_C5 = CLBLM_R_X11Y152_SLICE_X15Y152_AQ;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_C6 = CLBLM_L_X12Y152_SLICE_X16Y152_BQ;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_A4 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_A5 = 1'b1;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_A6 = CLBLM_L_X8Y148_SLICE_X10Y148_A5Q;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_C1 = CLBLM_R_X11Y154_SLICE_X15Y154_AQ;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_C2 = CLBLM_R_X11Y153_SLICE_X15Y153_AQ;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_B1 = CLBLM_L_X10Y145_SLICE_X13Y145_CQ;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_B2 = CLBLM_L_X10Y143_SLICE_X13Y143_BQ;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_B3 = 1'b1;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_B4 = CLBLM_R_X7Y142_SLICE_X8Y142_DO6;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_B5 = CLBLM_R_X7Y143_SLICE_X9Y143_CQ;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_D3 = CLBLM_R_X11Y154_SLICE_X15Y154_BQ;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_C1 = CLBLM_L_X12Y145_SLICE_X16Y145_AQ;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_C2 = CLBLM_L_X10Y148_SLICE_X12Y148_BQ;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_C4 = CLBLM_L_X12Y144_SLICE_X16Y144_AQ;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_C5 = CLBLM_L_X12Y144_SLICE_X16Y144_BQ;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_C3 = CLBLM_L_X12Y144_SLICE_X16Y144_CQ;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_C6 = 1'b1;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_D6 = CLBLM_L_X12Y152_SLICE_X16Y152_BQ;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_A3 = 1'b1;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_A4 = CLBLM_L_X12Y153_SLICE_X16Y153_BO6;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_A5 = 1'b1;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_A6 = CLBLM_R_X11Y154_SLICE_X15Y154_CO5;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_D1 = CLBLM_R_X11Y144_SLICE_X15Y144_AO6;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_D2 = CLBLM_R_X11Y144_SLICE_X15Y144_CO6;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_D3 = CLBLM_R_X11Y148_SLICE_X15Y148_A5Q;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_D5 = CLBLM_R_X7Y145_SLICE_X9Y145_CQ;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_D6 = CLBLM_R_X3Y151_SLICE_X2Y151_AO6;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_B1 = CLBLM_L_X12Y153_SLICE_X16Y153_DO6;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_B2 = CLBLM_L_X10Y154_SLICE_X13Y154_CO5;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_B3 = CLBLM_L_X12Y153_SLICE_X16Y153_AQ;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_B4 = CLBLM_R_X11Y153_SLICE_X14Y153_CO5;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_B5 = CLBLM_R_X11Y152_SLICE_X14Y152_AQ;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_B6 = CLBLM_L_X12Y153_SLICE_X16Y153_CO6;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_A1 = CLBLM_R_X7Y145_SLICE_X9Y145_CQ;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_C1 = CLBLM_R_X11Y154_SLICE_X15Y154_AQ;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_C2 = CLBLM_R_X11Y152_SLICE_X15Y152_AQ;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_C3 = CLBLM_R_X11Y154_SLICE_X14Y154_AQ;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_C4 = CLBLM_R_X11Y154_SLICE_X15Y154_BQ;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_A2 = CLBLM_R_X7Y142_SLICE_X8Y142_DO6;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_C6 = CLBLM_L_X12Y152_SLICE_X16Y152_BQ;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_A3 = CLBLM_L_X10Y143_SLICE_X13Y143_CO5;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_A4 = CLBLM_L_X10Y141_SLICE_X12Y141_BO6;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_A5 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_A6 = CLBLM_L_X10Y145_SLICE_X13Y145_CQ;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_B4 = CLBLM_R_X7Y142_SLICE_X8Y142_DO6;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_B1 = CLBLM_R_X5Y144_SLICE_X7Y144_B5Q;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_B2 = CLBLM_L_X10Y141_SLICE_X12Y141_BO6;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_D1 = CLBLM_L_X12Y151_SLICE_X16Y151_DO5;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_D2 = CLBLM_L_X10Y153_SLICE_X13Y153_CQ;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_D3 = CLBLM_L_X10Y153_SLICE_X13Y153_BQ;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_D4 = CLBLM_R_X11Y154_SLICE_X15Y154_BQ;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_D5 = CLBLM_R_X11Y154_SLICE_X14Y154_AQ;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_C2 = CLBLM_L_X10Y145_SLICE_X12Y145_DQ;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_C3 = CLBLM_L_X8Y144_SLICE_X11Y144_AQ;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_C4 = 1'b1;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_D6 = CLBLM_R_X11Y154_SLICE_X15Y154_AQ;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_C1 = CLBLM_L_X10Y145_SLICE_X12Y145_C5Q;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_C5 = CLBLM_L_X10Y143_SLICE_X12Y143_DO6;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_C6 = CLBLM_L_X8Y145_SLICE_X11Y145_BQ;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_B6 = 1'b1;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_D1 = 1'b1;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_D2 = CLBLM_L_X10Y144_SLICE_X12Y144_BQ;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_D3 = CLBLM_R_X5Y144_SLICE_X7Y144_B5Q;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_D4 = 1'b1;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_D5 = CLBLM_R_X11Y148_SLICE_X15Y148_A5Q;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_D6 = CLBLM_L_X8Y144_SLICE_X10Y144_BQ;
  assign CLBLM_R_X103Y141_SLICE_X162Y141_B5 = 1'b1;
  assign CLBLM_R_X103Y141_SLICE_X162Y141_B6 = 1'b1;
  assign RIOI3_X105Y197_OLOGIC_X1Y197_D1 = CLBLM_L_X16Y158_SLICE_X22Y158_AO6;
  assign CLBLM_R_X103Y141_SLICE_X162Y141_C1 = 1'b1;
  assign CLBLM_R_X103Y141_SLICE_X162Y141_C2 = 1'b1;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_A4 = 1'b1;
  assign CLBLM_R_X103Y141_SLICE_X162Y141_C3 = 1'b1;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_A5 = CLBLM_R_X7Y148_SLICE_X9Y148_DQ;
  assign CLBLM_R_X103Y141_SLICE_X162Y141_C4 = 1'b1;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_A6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X103Y141_SLICE_X162Y141_C5 = 1'b1;
  assign CLBLM_R_X103Y141_SLICE_X162Y141_C6 = 1'b1;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOB33_X0Y121_IOB_X0Y121_O = CLBLM_L_X8Y142_SLICE_X10Y142_A5Q;
  assign LIOB33_X0Y121_IOB_X0Y122_O = CLBLM_R_X3Y144_SLICE_X2Y144_BQ;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_B2 = CLBLL_L_X4Y150_SLICE_X4Y150_B5Q;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_B3 = CLBLM_R_X11Y153_SLICE_X14Y153_AO6;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_B4 = 1'b1;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_B5 = CLBLM_R_X7Y147_SLICE_X9Y147_AQ;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_B6 = 1'b1;
  assign CLBLM_R_X103Y141_SLICE_X162Y141_D1 = 1'b1;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_A5 = CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  assign CLBLM_R_X103Y141_SLICE_X162Y141_D2 = 1'b1;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_A6 = CLBLM_L_X8Y146_SLICE_X10Y146_B5Q;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_D1 = LIOB33_X0Y53_IOB_X0Y54_I;
  assign CLBLM_R_X103Y141_SLICE_X162Y141_D3 = 1'b1;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X103Y141_SLICE_X162Y141_D4 = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_T1 = 1'b1;
  assign CLBLM_R_X103Y141_SLICE_X162Y141_D5 = 1'b1;
  assign RIOI3_X105Y185_OLOGIC_X1Y186_D1 = CLBLM_L_X12Y151_SLICE_X16Y151_AQ;
  assign LIOI3_X0Y79_OLOGIC_X0Y80_D1 = CLBLL_L_X2Y138_SLICE_X0Y138_AO6;
  assign CLBLM_R_X103Y141_SLICE_X162Y141_D6 = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_D1 = CLBLM_R_X3Y143_SLICE_X2Y143_AQ;
  assign RIOI3_X105Y185_OLOGIC_X1Y186_T1 = 1'b1;
  assign LIOI3_X0Y79_OLOGIC_X0Y80_T1 = 1'b1;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_T1 = 1'b1;
  assign RIOI3_X105Y185_OLOGIC_X1Y185_D1 = CLBLM_L_X10Y150_SLICE_X13Y150_DO5;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_D1 = LIOB33_X0Y59_IOB_X0Y60_I;
  assign RIOI3_X105Y185_OLOGIC_X1Y185_T1 = 1'b1;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_B6 = CLBLM_L_X8Y146_SLICE_X10Y146_B5Q;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_D1 = LIOB33_X0Y55_IOB_X0Y56_I;
  assign CLBLM_L_X12Y154_SLICE_X17Y154_A1 = 1'b1;
  assign CLBLM_L_X12Y154_SLICE_X17Y154_A2 = 1'b1;
  assign CLBLM_L_X12Y154_SLICE_X17Y154_A3 = 1'b1;
  assign CLBLM_L_X12Y154_SLICE_X17Y154_A4 = 1'b1;
  assign CLBLM_L_X12Y154_SLICE_X17Y154_A5 = 1'b1;
  assign CLBLM_L_X12Y154_SLICE_X17Y154_A6 = 1'b1;
  assign CLBLM_L_X12Y154_SLICE_X17Y154_B1 = 1'b1;
  assign CLBLM_L_X12Y154_SLICE_X17Y154_B2 = 1'b1;
  assign CLBLM_L_X12Y154_SLICE_X17Y154_B3 = 1'b1;
  assign CLBLM_L_X12Y154_SLICE_X17Y154_B4 = 1'b1;
  assign CLBLM_L_X12Y154_SLICE_X17Y154_B5 = 1'b1;
  assign CLBLM_L_X12Y154_SLICE_X17Y154_B6 = 1'b1;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_D2 = CLBLM_R_X7Y145_SLICE_X8Y145_AQ;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_C1 = CLBLM_R_X7Y146_SLICE_X9Y146_AQ;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_A1 = CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_A2 = 1'b1;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_A3 = CLBLM_L_X10Y144_SLICE_X13Y144_AQ;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_A4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_A5 = CLBLM_L_X10Y142_SLICE_X13Y142_AQ;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y154_SLICE_X17Y154_C1 = 1'b1;
  assign CLBLM_L_X12Y154_SLICE_X17Y154_C2 = 1'b1;
  assign CLBLM_L_X12Y154_SLICE_X17Y154_C3 = 1'b1;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_B1 = CLBLM_L_X10Y144_SLICE_X13Y144_DO6;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_B2 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_B3 = CLBLM_R_X5Y142_SLICE_X7Y142_AQ;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_B4 = CLBLM_L_X10Y145_SLICE_X12Y145_CQ;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_B5 = 1'b1;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y154_SLICE_X17Y154_D1 = 1'b1;
  assign CLBLM_L_X12Y154_SLICE_X17Y154_D2 = 1'b1;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_C1 = 1'b1;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_C2 = CLBLM_L_X10Y144_SLICE_X13Y144_CQ;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_C4 = CLBLM_L_X10Y147_SLICE_X12Y147_A5Q;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_C5 = CLBLM_R_X11Y145_SLICE_X15Y145_AQ;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_C6 = CLBLM_R_X7Y142_SLICE_X8Y142_DO6;
  assign CLBLM_L_X12Y154_SLICE_X17Y154_D3 = 1'b1;
  assign CLBLM_L_X12Y154_SLICE_X17Y154_D4 = 1'b1;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y154_SLICE_X16Y154_A1 = CLBLM_L_X10Y154_SLICE_X13Y154_CO5;
  assign CLBLM_L_X12Y154_SLICE_X16Y154_A2 = CLBLL_L_X4Y150_SLICE_X5Y150_AQ;
  assign CLBLM_L_X12Y154_SLICE_X16Y154_A3 = CLBLM_L_X12Y154_SLICE_X16Y154_AQ;
  assign CLBLM_L_X12Y154_SLICE_X16Y154_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y154_SLICE_X16Y154_A5 = CLBLM_R_X11Y154_SLICE_X15Y154_CO5;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_D1 = CLBLM_L_X10Y145_SLICE_X12Y145_C5Q;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_D2 = CLBLM_L_X12Y144_SLICE_X16Y144_DO5;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_D3 = CLBLM_L_X10Y144_SLICE_X13Y144_BQ;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_D4 = CLBLM_R_X7Y142_SLICE_X8Y142_DO6;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_D5 = 1'b1;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_D6 = CLBLM_L_X10Y148_SLICE_X12Y148_BQ;
  assign CLBLM_L_X12Y154_SLICE_X16Y154_A6 = CLBLM_L_X12Y152_SLICE_X16Y152_CO6;
  assign CLBLM_L_X12Y154_SLICE_X16Y154_B1 = CLBLM_L_X10Y153_SLICE_X13Y153_BQ;
  assign CLBLM_L_X12Y154_SLICE_X16Y154_B2 = CLBLM_L_X10Y153_SLICE_X13Y153_CQ;
  assign CLBLM_L_X12Y154_SLICE_X16Y154_B3 = CLBLM_R_X11Y154_SLICE_X15Y154_AQ;
  assign CLBLM_L_X12Y154_SLICE_X16Y154_B4 = CLBLM_R_X11Y154_SLICE_X14Y154_AQ;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_A1 = CLBLM_R_X11Y151_SLICE_X15Y151_CO6;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_A2 = CLBLM_R_X7Y151_SLICE_X8Y151_CO5;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_A3 = CLBLM_L_X10Y144_SLICE_X12Y144_AQ;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_A4 = CLBLM_L_X10Y142_SLICE_X12Y142_BO6;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_A5 = CLBLM_R_X7Y144_SLICE_X9Y144_DO5;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_A6 = CLBLM_L_X8Y147_SLICE_X11Y147_BO5;
  assign CLBLM_L_X12Y154_SLICE_X16Y154_C1 = 1'b1;
  assign CLBLM_L_X12Y154_SLICE_X16Y154_C2 = 1'b1;
  assign CLBLM_L_X12Y154_SLICE_X16Y154_C3 = 1'b1;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_B1 = CLBLM_R_X5Y144_SLICE_X7Y144_AQ;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_B2 = CLBLM_L_X10Y144_SLICE_X12Y144_BQ;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_B3 = CLBLM_R_X5Y143_SLICE_X7Y143_AQ;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_B4 = CLBLM_R_X7Y142_SLICE_X8Y142_DO6;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_B5 = 1'b1;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y154_SLICE_X16Y154_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X12Y154_SLICE_X16Y154_D1 = 1'b1;
  assign CLBLM_L_X12Y154_SLICE_X16Y154_D2 = 1'b1;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_C1 = CLBLM_R_X7Y144_SLICE_X9Y144_DO5;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_C2 = CLBLM_L_X10Y144_SLICE_X12Y144_CQ;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_C3 = CLBLM_R_X5Y146_SLICE_X6Y146_BO5;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_C4 = CLBLM_R_X11Y151_SLICE_X15Y151_CO6;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_C5 = CLBLM_L_X8Y144_SLICE_X11Y144_DO6;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_C6 = CLBLM_L_X10Y142_SLICE_X12Y142_BO6;
  assign CLBLM_L_X12Y154_SLICE_X16Y154_D3 = 1'b1;
  assign CLBLM_L_X12Y154_SLICE_X16Y154_D4 = 1'b1;
  assign CLBLM_L_X12Y154_SLICE_X16Y154_D5 = 1'b1;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y154_SLICE_X16Y154_D6 = 1'b1;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_A5 = CLBLM_R_X7Y148_SLICE_X9Y148_AQ;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_A6 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_D1 = CLBLM_L_X12Y145_SLICE_X16Y145_AQ;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_D2 = CLBLM_R_X11Y144_SLICE_X15Y144_DO6;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_D3 = CLBLM_L_X12Y144_SLICE_X16Y144_BQ;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_D4 = CLBLM_L_X10Y146_SLICE_X12Y146_CQ;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_D5 = CLBLM_L_X12Y144_SLICE_X16Y144_CQ;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_D6 = CLBLM_L_X12Y144_SLICE_X16Y144_AQ;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_A1 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_A2 = CLBLM_L_X10Y149_SLICE_X12Y149_AQ;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_A3 = CLBLM_R_X11Y151_SLICE_X15Y151_AQ;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_A4 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_A5 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_A6 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_B1 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_B2 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_B3 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_B4 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_B5 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_B6 = 1'b1;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_B1 = CLBLM_R_X7Y148_SLICE_X9Y148_DQ;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_C1 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_C2 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_C3 = 1'b1;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_B2 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_C4 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_C5 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_C6 = 1'b1;
  assign CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_I = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_B3 = CLBLM_R_X7Y147_SLICE_X8Y147_CQ;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_B4 = CLBLM_R_X5Y146_SLICE_X6Y146_A5Q;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_D1 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_D2 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_D3 = 1'b1;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_D4 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_D5 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_D6 = 1'b1;
  assign LIOI3_X0Y79_ILOGIC_X0Y79_D = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_B6 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_A1 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_A2 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_A3 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_A4 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_A5 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_A6 = 1'b1;
  assign RIOI3_X105Y125_ILOGIC_X1Y126_D = RIOB33_X105Y125_IOB_X1Y126_I;
  assign LIOB33_X0Y123_IOB_X0Y124_O = CLBLM_R_X3Y147_SLICE_X3Y147_C5Q;
  assign LIOB33_X0Y123_IOB_X0Y123_O = CLBLM_R_X7Y143_SLICE_X8Y143_B5Q;
  assign RIOI3_X105Y125_ILOGIC_X1Y125_D = RIOB33_X105Y125_IOB_X1Y125_I;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_B1 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_B2 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_B3 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_B4 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_B5 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_B6 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_C1 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_C2 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_C3 = 1'b1;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_C1 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_C4 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_C5 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_C6 = 1'b1;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_C2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_D1 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_D2 = 1'b1;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_C4 = CLBLM_R_X7Y150_SLICE_X8Y150_CQ;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_D3 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_D4 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_D5 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_D6 = 1'b1;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_C5 = 1'b1;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_C6 = CLBLM_R_X5Y147_SLICE_X7Y147_BQ;
  assign RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_D = RIOB33_X105Y119_IOB_X1Y119_I;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_D1 = CLBLM_R_X7Y143_SLICE_X8Y143_BQ;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_D5 = RIOB33_X105Y143_IOB_X1Y144_I;
  assign LIOI3_X0Y197_OLOGIC_X0Y197_D1 = LIOB33_X0Y71_IOB_X0Y72_I;
  assign CLBLM_L_X12Y155_SLICE_X17Y155_A1 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_L_X12Y155_SLICE_X17Y155_A2 = CLBLM_R_X7Y155_SLICE_X9Y155_AQ;
  assign CLBLM_L_X12Y155_SLICE_X17Y155_A3 = CLBLM_L_X12Y155_SLICE_X17Y155_AQ;
  assign CLBLM_L_X12Y155_SLICE_X17Y155_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y155_SLICE_X17Y155_A5 = CLBLM_R_X5Y142_SLICE_X7Y142_AQ;
  assign CLBLM_L_X12Y155_SLICE_X17Y155_A6 = 1'b1;
  assign CLBLM_L_X12Y155_SLICE_X17Y155_B1 = 1'b1;
  assign CLBLM_L_X12Y155_SLICE_X17Y155_B2 = 1'b1;
  assign CLBLM_L_X12Y155_SLICE_X17Y155_B3 = 1'b1;
  assign CLBLM_L_X12Y155_SLICE_X17Y155_B4 = 1'b1;
  assign CLBLM_L_X12Y155_SLICE_X17Y155_B5 = 1'b1;
  assign CLBLM_L_X12Y155_SLICE_X17Y155_B6 = 1'b1;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_A1 = CLBLM_L_X10Y147_SLICE_X12Y147_A5Q;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_A2 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_A3 = CLBLM_R_X11Y145_SLICE_X15Y145_AQ;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_A5 = CLBLL_L_X4Y145_SLICE_X4Y145_AQ;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_A6 = 1'b1;
  assign CLBLM_L_X12Y155_SLICE_X17Y155_C1 = 1'b1;
  assign CLBLM_L_X12Y155_SLICE_X17Y155_C2 = 1'b1;
  assign CLBLM_L_X12Y155_SLICE_X17Y155_C3 = 1'b1;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_B1 = 1'b1;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_B2 = CLBLM_L_X10Y146_SLICE_X13Y146_AQ;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_B3 = CLBLM_L_X12Y145_SLICE_X16Y145_AQ;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_B6 = 1'b1;
  assign CLBLM_L_X12Y155_SLICE_X17Y155_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X12Y155_SLICE_X17Y155_D1 = 1'b1;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_C2 = CLBLM_L_X10Y145_SLICE_X13Y145_CQ;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_C3 = CLBLM_L_X10Y146_SLICE_X12Y146_A5Q;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_C4 = CLBLM_R_X7Y146_SLICE_X9Y146_CQ;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_C5 = CLBLL_L_X4Y145_SLICE_X5Y145_DO6;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_C6 = 1'b1;
  assign CLBLM_L_X12Y155_SLICE_X17Y155_D3 = 1'b1;
  assign CLBLM_L_X12Y155_SLICE_X17Y155_D4 = 1'b1;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y155_SLICE_X16Y155_A2 = 1'b1;
  assign CLBLM_L_X12Y155_SLICE_X16Y155_A3 = 1'b1;
  assign CLBLM_L_X12Y155_SLICE_X16Y155_A4 = 1'b1;
  assign CLBLM_L_X12Y155_SLICE_X16Y155_A5 = 1'b1;
  assign CLBLM_L_X12Y155_SLICE_X16Y155_A6 = 1'b1;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_D1 = CLBLM_L_X8Y148_SLICE_X10Y148_BQ;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_D2 = CLBLM_R_X7Y142_SLICE_X8Y142_DO6;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_D3 = CLBLM_R_X11Y146_SLICE_X15Y146_DQ;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_D4 = CLBLM_L_X10Y142_SLICE_X13Y142_BO6;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_D5 = CLBLM_L_X10Y143_SLICE_X13Y143_BQ;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_D6 = CLBLM_L_X12Y144_SLICE_X16Y144_CQ;
  assign CLBLM_L_X12Y155_SLICE_X16Y155_B1 = 1'b1;
  assign CLBLM_L_X12Y155_SLICE_X16Y155_B2 = 1'b1;
  assign CLBLM_L_X12Y155_SLICE_X16Y155_B3 = 1'b1;
  assign CLBLM_L_X12Y155_SLICE_X16Y155_B4 = 1'b1;
  assign CLBLM_L_X12Y155_SLICE_X16Y155_B5 = 1'b1;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_A1 = CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_A2 = CLBLM_L_X8Y145_SLICE_X10Y145_DO6;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_A3 = CLBLM_L_X10Y145_SLICE_X12Y145_AQ;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_A4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_A5 = CLBLM_R_X11Y143_SLICE_X14Y143_BQ;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y155_SLICE_X16Y155_C1 = 1'b1;
  assign CLBLM_L_X12Y155_SLICE_X16Y155_C2 = 1'b1;
  assign CLBLM_L_X12Y155_SLICE_X16Y155_C3 = 1'b1;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_B1 = CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_B2 = CLBLM_L_X10Y145_SLICE_X12Y145_BQ;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_B3 = CLBLM_R_X7Y145_SLICE_X9Y145_BQ;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_B4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_B5 = CLBLM_R_X5Y145_SLICE_X7Y145_BQ;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y155_SLICE_X16Y155_D1 = 1'b1;
  assign CLBLM_L_X12Y155_SLICE_X16Y155_D2 = 1'b1;
  assign CLBLM_L_X12Y155_SLICE_X16Y155_D3 = 1'b1;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_C1 = CLBLM_L_X10Y144_SLICE_X13Y144_BQ;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_C2 = CLBLM_R_X7Y151_SLICE_X9Y151_CQ;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_C3 = CLBLM_L_X10Y149_SLICE_X12Y149_CO6;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_C5 = CLBLM_L_X10Y146_SLICE_X12Y146_A5Q;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_C6 = 1'b1;
  assign CLBLM_L_X12Y155_SLICE_X16Y155_D4 = 1'b1;
  assign CLBLM_L_X12Y155_SLICE_X16Y155_D5 = 1'b1;
  assign CLBLM_L_X12Y155_SLICE_X16Y155_D6 = 1'b1;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_D1 = 1'b1;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_D2 = CLBLM_R_X7Y142_SLICE_X8Y142_DO6;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_D3 = CLBLM_L_X10Y145_SLICE_X12Y145_DQ;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_D4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_D5 = CLBLM_L_X8Y144_SLICE_X10Y144_BQ;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_D6 = CLBLM_L_X10Y151_SLICE_X13Y151_BQ;
  assign LIOB33_X0Y125_IOB_X0Y126_O = CLBLM_R_X3Y143_SLICE_X2Y143_BQ;
  assign LIOB33_X0Y125_IOB_X0Y125_O = CLBLM_L_X8Y145_SLICE_X11Y145_B5Q;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_A1 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_A2 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_A3 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_A4 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_A5 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_A6 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_B1 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_B2 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_B3 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_B4 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_B5 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_B6 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_C1 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_C2 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_C3 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_C4 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_C5 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_C6 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_D1 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_D2 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_D3 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_D4 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_D5 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_D6 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_A1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_A2 = CLBLL_L_X4Y147_SLICE_X5Y147_CQ;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_A3 = CLBLL_L_X4Y142_SLICE_X5Y142_AQ;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_A5 = CLBLM_R_X5Y151_SLICE_X6Y151_DQ;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_A6 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_B1 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_B2 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_B3 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_B4 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_B5 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_B6 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_C1 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_C2 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_C3 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_C4 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_C5 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_C6 = 1'b1;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_A1 = CLBLM_R_X7Y149_SLICE_X8Y149_CQ;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_A2 = CLBLM_R_X11Y149_SLICE_X14Y149_CQ;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_A3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_A4 = CLBLM_L_X10Y146_SLICE_X13Y146_CQ;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_A6 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_D1 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_D2 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_D3 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_D4 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_D5 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_D6 = 1'b1;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_B2 = CLBLM_L_X10Y145_SLICE_X13Y145_BQ;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_B3 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_B5 = CLBLM_L_X10Y147_SLICE_X12Y147_AQ;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_B6 = 1'b1;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_C2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_C3 = 1'b1;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_C4 = CLBLM_R_X11Y148_SLICE_X15Y148_A5Q;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_C5 = CLBLM_L_X10Y147_SLICE_X13Y147_BQ;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_C6 = 1'b1;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_T1 = 1'b1;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_D1 = CLBLM_L_X10Y148_SLICE_X13Y148_BQ;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_D2 = CLBLM_L_X10Y146_SLICE_X13Y146_CQ;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_D3 = 1'b1;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_D4 = CLBLM_L_X10Y146_SLICE_X13Y146_A5Q;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_D5 = 1'b1;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_D6 = CLBLM_L_X10Y145_SLICE_X13Y145_BQ;
  assign RIOI3_X105Y189_OLOGIC_X1Y190_D1 = CLBLM_L_X12Y152_SLICE_X17Y152_AQ;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_D1 = LIOB33_X0Y57_IOB_X0Y58_I;
  assign RIOI3_X105Y189_OLOGIC_X1Y190_T1 = 1'b1;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_A1 = CLBLM_L_X10Y146_SLICE_X12Y146_B5Q;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_A2 = CLBLM_R_X5Y154_SLICE_X6Y154_BO6;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_A3 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_A4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_A5 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_T1 = 1'b1;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_AX = CLBLM_R_X7Y148_SLICE_X8Y148_BO6;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_B1 = 1'b1;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_B2 = CLBLM_L_X10Y146_SLICE_X12Y146_BQ;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_B4 = CLBLM_R_X7Y142_SLICE_X8Y142_DO6;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_B5 = CLBLM_R_X11Y146_SLICE_X15Y146_AQ;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_B6 = CLBLM_R_X7Y148_SLICE_X8Y148_CQ;
  assign RIOI3_X105Y189_OLOGIC_X1Y189_D1 = CLBLM_R_X11Y153_SLICE_X14Y153_CQ;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_BX = CLBLM_L_X10Y148_SLICE_X12Y148_AO6;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_C1 = CLBLM_R_X11Y153_SLICE_X15Y153_BQ;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_C2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_C3 = CLBLM_L_X12Y144_SLICE_X16Y144_BQ;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_C4 = CLBLM_L_X10Y144_SLICE_X12Y144_CQ;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_C5 = CLBLM_L_X10Y146_SLICE_X12Y146_B5Q;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_C6 = 1'b1;
  assign RIOI3_X105Y189_OLOGIC_X1Y189_T1 = 1'b1;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_D1 = CLBLM_L_X8Y145_SLICE_X10Y145_BQ;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_D2 = CLBLM_L_X10Y146_SLICE_X13Y146_A5Q;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_D3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_D4 = CLBLM_R_X7Y148_SLICE_X8Y148_DQ;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_D6 = 1'b1;
  assign LIOB33_X0Y127_IOB_X0Y127_O = CLBLL_L_X4Y147_SLICE_X5Y147_CQ;
  assign LIOB33_X0Y127_IOB_X0Y128_O = CLBLL_L_X2Y147_SLICE_X1Y147_AQ;
  assign LIOI3_X0Y153_OLOGIC_X0Y154_D1 = LIOB33_X0Y67_IOB_X0Y68_I;
  assign LIOI3_X0Y153_OLOGIC_X0Y154_T1 = 1'b1;
  assign CLBLM_R_X11Y157_SLICE_X15Y157_C3 = 1'b1;
  assign CLBLM_R_X11Y157_SLICE_X15Y157_C4 = 1'b1;
  assign CLBLM_R_X11Y157_SLICE_X15Y157_C5 = 1'b1;
  assign CLBLM_R_X11Y157_SLICE_X15Y157_C6 = 1'b1;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_A1 = CLBLM_L_X8Y145_SLICE_X11Y145_AQ;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_A3 = CLBLL_L_X4Y143_SLICE_X4Y143_AQ;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_A5 = CLBLL_L_X4Y143_SLICE_X4Y143_CO5;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_A6 = CLBLM_R_X3Y143_SLICE_X2Y143_DQ;
  assign LIOI3_X0Y153_OLOGIC_X0Y153_D1 = LIOB33_X0Y67_IOB_X0Y67_I;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_B1 = 1'b1;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_B2 = CLBLL_L_X4Y143_SLICE_X4Y143_BQ;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_B5 = CLBLM_R_X3Y142_SLICE_X2Y142_AQ;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_B6 = CLBLM_R_X5Y148_SLICE_X7Y148_CQ;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_C1 = CLBLM_R_X7Y142_SLICE_X8Y142_DO6;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_C2 = CLBLL_L_X4Y143_SLICE_X4Y143_AQ;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_C3 = CLBLL_L_X4Y144_SLICE_X5Y144_BQ;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_C4 = CLBLL_L_X4Y144_SLICE_X5Y144_AQ;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_C5 = CLBLL_L_X4Y144_SLICE_X5Y144_A5Q;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_C6 = 1'b1;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y157_SLICE_X15Y157_D3 = 1'b1;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_D1 = 1'b1;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_D2 = 1'b1;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_D3 = 1'b1;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_D4 = 1'b1;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_D5 = 1'b1;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_D6 = 1'b1;
  assign CLBLM_R_X11Y157_SLICE_X15Y157_D5 = 1'b1;
  assign RIOI3_X105Y127_ILOGIC_X1Y128_D = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLM_R_X11Y157_SLICE_X15Y157_D6 = 1'b1;
  assign RIOI3_X105Y127_ILOGIC_X1Y127_D = RIOB33_X105Y127_IOB_X1Y127_I;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_B4 = CLBLL_L_X4Y145_SLICE_X5Y145_DO6;
  assign LIOI3_X0Y153_OLOGIC_X0Y153_T1 = 1'b1;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_A1 = CLBLL_L_X4Y144_SLICE_X5Y144_BQ;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_A2 = CLBLL_L_X4Y144_SLICE_X5Y144_AQ;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_A3 = 1'b1;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_A4 = CLBLL_L_X4Y145_SLICE_X5Y145_DO6;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_A5 = CLBLL_L_X4Y143_SLICE_X4Y143_AQ;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_A6 = CLBLL_L_X4Y144_SLICE_X5Y144_A5Q;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_B1 = 1'b1;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_B2 = 1'b1;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_B3 = 1'b1;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_B4 = 1'b1;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_B5 = 1'b1;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_B6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y132_D = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_C1 = 1'b1;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_C2 = 1'b1;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_C3 = 1'b1;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_C4 = 1'b1;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_C5 = 1'b1;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_C6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y131_D = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_A1 = CLBLM_L_X10Y147_SLICE_X13Y147_DO6;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_A2 = CLBLM_L_X10Y147_SLICE_X13Y147_BQ;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_A3 = CLBLM_L_X10Y147_SLICE_X13Y147_AQ;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_D1 = 1'b1;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_D2 = 1'b1;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_D3 = 1'b1;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_D4 = 1'b1;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_D5 = 1'b1;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_D6 = 1'b1;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_A6 = CLBLM_L_X8Y145_SLICE_X11Y145_A5Q;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_B3 = CLBLM_L_X8Y146_SLICE_X11Y146_BQ;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_B4 = 1'b1;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_B5 = CLBLM_L_X8Y145_SLICE_X10Y145_AQ;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_B6 = 1'b1;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_C2 = CLBLM_L_X10Y144_SLICE_X13Y144_AQ;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_C3 = CLBLM_R_X3Y151_SLICE_X3Y151_AO6;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_C4 = CLBLM_R_X5Y145_SLICE_X6Y145_BO5;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_C5 = CLBLM_R_X5Y144_SLICE_X7Y144_AQ;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_C6 = 1'b1;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_X105Y155_OLOGIC_X1Y156_D1 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_D1 = 1'b1;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_D2 = CLBLM_L_X8Y147_SLICE_X11Y147_CO6;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_D3 = CLBLM_L_X10Y149_SLICE_X13Y149_DQ;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_D4 = CLBLM_L_X10Y146_SLICE_X13Y146_CQ;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_D5 = CLBLM_L_X10Y147_SLICE_X13Y147_AQ;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_D6 = 1'b1;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_B5 = CLBLM_R_X5Y152_SLICE_X7Y152_DO5;
  assign CLBLM_R_X11Y157_SLICE_X14Y157_B1 = 1'b1;
  assign CLBLM_R_X11Y157_SLICE_X14Y157_B2 = 1'b1;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_A2 = CLBLM_R_X11Y147_SLICE_X14Y147_BQ;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_A3 = CLBLM_L_X10Y147_SLICE_X12Y147_AQ;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_A4 = CLBLL_L_X4Y146_SLICE_X4Y146_DO6;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_A5 = CLBLM_R_X11Y146_SLICE_X14Y146_AQ;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_A6 = CLBLM_L_X10Y148_SLICE_X13Y148_AQ;
  assign CLBLM_R_X11Y157_SLICE_X14Y157_B3 = 1'b1;
  assign CLBLM_R_X11Y157_SLICE_X14Y157_B4 = 1'b1;
  assign LIOB33_X0Y129_IOB_X0Y129_O = CLBLM_R_X3Y148_SLICE_X3Y148_AQ;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_AX = CLBLM_L_X10Y152_SLICE_X12Y152_CO6;
  assign LIOB33_X0Y129_IOB_X0Y130_O = CLBLL_L_X52Y126_SLICE_X78Y126_AO6;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_B1 = CLBLM_R_X11Y148_SLICE_X15Y148_CQ;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_B2 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_B4 = CLBLM_L_X10Y146_SLICE_X13Y146_B5Q;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_B5 = CLBLM_L_X10Y145_SLICE_X13Y145_CQ;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_B6 = 1'b1;
  assign CLBLM_R_X11Y157_SLICE_X14Y157_B5 = 1'b1;
  assign CLBLM_R_X11Y157_SLICE_X14Y157_B6 = 1'b1;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_C2 = CLBLM_R_X11Y146_SLICE_X14Y146_DQ;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_C3 = CLBLM_L_X10Y150_SLICE_X12Y150_DQ;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_C5 = CLBLM_L_X10Y147_SLICE_X12Y147_BO5;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_C6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_T1 = 1'b1;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_D1 = CLBLM_R_X3Y143_SLICE_X2Y143_BQ;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_D2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_D3 = CLBLM_L_X10Y146_SLICE_X13Y146_AQ;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_D4 = CLBLM_R_X11Y147_SLICE_X15Y147_BQ;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_D5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_D6 = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y156_T1 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X163Y176_A1 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X163Y176_A2 = 1'b1;
  assign CLBLM_R_X11Y157_SLICE_X14Y157_C1 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X163Y176_A3 = CLBLM_L_X12Y155_SLICE_X17Y155_AQ;
  assign CLBLM_R_X103Y176_SLICE_X163Y176_A4 = CLBLM_L_X12Y151_SLICE_X16Y151_AQ;
  assign CLBLM_R_X103Y176_SLICE_X163Y176_A5 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_R_X103Y176_SLICE_X163Y176_A6 = 1'b1;
  assign CLBLM_R_X11Y157_SLICE_X14Y157_C2 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X163Y176_B1 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X163Y176_B2 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X163Y176_B3 = 1'b1;
  assign CLBLM_R_X11Y157_SLICE_X14Y157_C3 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X163Y176_B4 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X163Y176_B5 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X163Y176_B6 = 1'b1;
  assign CLBLM_R_X11Y157_SLICE_X14Y157_C4 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X163Y176_C1 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X163Y176_C2 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X163Y176_C3 = 1'b1;
  assign CLBLM_R_X11Y157_SLICE_X14Y157_C5 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X163Y176_C4 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X163Y176_C5 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X163Y176_C6 = 1'b1;
  assign CLBLM_R_X11Y157_SLICE_X14Y157_C6 = 1'b1;
  assign CLBLM_R_X13Y151_SLICE_X19Y151_A1 = 1'b1;
  assign CLBLM_R_X13Y151_SLICE_X19Y151_A2 = 1'b1;
  assign CLBLM_R_X13Y151_SLICE_X19Y151_A3 = 1'b1;
  assign CLBLM_R_X13Y151_SLICE_X19Y151_A4 = 1'b1;
  assign CLBLM_R_X13Y151_SLICE_X19Y151_A5 = 1'b1;
  assign CLBLM_R_X13Y151_SLICE_X19Y151_A6 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X163Y176_D1 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X163Y176_D2 = 1'b1;
  assign CLBLM_R_X13Y151_SLICE_X19Y151_B1 = 1'b1;
  assign CLBLM_R_X13Y151_SLICE_X19Y151_B2 = 1'b1;
  assign CLBLM_R_X13Y151_SLICE_X19Y151_B3 = 1'b1;
  assign CLBLM_R_X13Y151_SLICE_X19Y151_B4 = 1'b1;
  assign CLBLM_R_X13Y151_SLICE_X19Y151_B5 = 1'b1;
  assign CLBLM_R_X13Y151_SLICE_X19Y151_B6 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X162Y176_A1 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X162Y176_A2 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X162Y176_A3 = 1'b1;
  assign CLBLM_R_X13Y151_SLICE_X19Y151_C1 = 1'b1;
  assign CLBLM_R_X13Y151_SLICE_X19Y151_C2 = 1'b1;
  assign CLBLM_R_X13Y151_SLICE_X19Y151_C3 = 1'b1;
  assign CLBLM_R_X13Y151_SLICE_X19Y151_C4 = 1'b1;
  assign CLBLM_R_X13Y151_SLICE_X19Y151_C5 = 1'b1;
  assign CLBLM_R_X13Y151_SLICE_X19Y151_C6 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X162Y176_A4 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X162Y176_A5 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X162Y176_A6 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X162Y176_B1 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X162Y176_B2 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X162Y176_B3 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X162Y176_B4 = 1'b1;
  assign CLBLM_R_X13Y151_SLICE_X19Y151_D1 = 1'b1;
  assign CLBLM_R_X13Y151_SLICE_X19Y151_D2 = 1'b1;
  assign CLBLM_R_X13Y151_SLICE_X19Y151_D3 = 1'b1;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_B6 = 1'b1;
  assign CLBLM_R_X13Y151_SLICE_X19Y151_D4 = 1'b1;
  assign CLBLM_R_X13Y151_SLICE_X19Y151_D5 = 1'b1;
  assign CLBLM_R_X13Y151_SLICE_X19Y151_D6 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X162Y176_C5 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X162Y176_C6 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X162Y176_C1 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X162Y176_C2 = 1'b1;
  assign CLBLM_R_X13Y151_SLICE_X18Y151_A1 = CLBLM_L_X12Y154_SLICE_X16Y154_BO5;
  assign CLBLM_R_X13Y151_SLICE_X18Y151_A2 = CLBLM_L_X12Y152_SLICE_X16Y152_BQ;
  assign CLBLM_R_X11Y157_SLICE_X14Y157_D1 = 1'b1;
  assign CLBLM_R_X13Y151_SLICE_X18Y151_A3 = CLBLM_R_X11Y153_SLICE_X15Y153_AQ;
  assign CLBLM_R_X13Y151_SLICE_X18Y151_A4 = CLBLM_L_X12Y153_SLICE_X16Y153_AQ;
  assign CLBLM_R_X13Y151_SLICE_X18Y151_A5 = CLBLM_L_X12Y154_SLICE_X16Y154_AQ;
  assign CLBLM_R_X13Y151_SLICE_X18Y151_A6 = CLBLM_R_X11Y152_SLICE_X15Y152_AQ;
  assign CLBLM_R_X11Y157_SLICE_X14Y157_D2 = 1'b1;
  assign CLBLM_R_X103Y176_SLICE_X162Y176_D1 = 1'b1;
  assign CLBLM_R_X13Y151_SLICE_X18Y151_B1 = CLBLM_L_X12Y154_SLICE_X16Y154_BO5;
  assign CLBLM_R_X11Y157_SLICE_X14Y157_D3 = 1'b1;
  assign CLBLM_R_X13Y151_SLICE_X18Y151_B2 = CLBLM_L_X12Y152_SLICE_X16Y152_BQ;
  assign CLBLM_R_X13Y151_SLICE_X18Y151_B3 = CLBLM_R_X11Y153_SLICE_X15Y153_AQ;
  assign CLBLM_R_X13Y151_SLICE_X18Y151_B4 = CLBLM_L_X12Y153_SLICE_X16Y153_AQ;
  assign CLBLM_R_X13Y151_SLICE_X18Y151_B5 = CLBLM_L_X12Y154_SLICE_X16Y154_AQ;
  assign CLBLM_R_X11Y157_SLICE_X14Y157_D4 = 1'b1;
  assign CLBLM_R_X13Y151_SLICE_X18Y151_B6 = CLBLM_R_X11Y152_SLICE_X15Y152_AQ;
  assign CLBLM_R_X103Y176_SLICE_X162Y176_D6 = 1'b1;
  assign CLBLM_R_X11Y157_SLICE_X14Y157_D5 = 1'b1;
  assign CLBLM_R_X13Y151_SLICE_X18Y151_C1 = CLBLM_L_X12Y154_SLICE_X16Y154_AQ;
  assign CLBLM_R_X13Y151_SLICE_X18Y151_C2 = CLBLM_L_X12Y152_SLICE_X17Y152_BQ;
  assign CLBLM_R_X13Y151_SLICE_X18Y151_C3 = CLBLM_L_X12Y152_SLICE_X16Y152_AQ;
  assign CLBLM_R_X13Y151_SLICE_X18Y151_C4 = CLBLM_L_X12Y153_SLICE_X17Y153_CO6;
  assign CLBLM_R_X11Y157_SLICE_X14Y157_D6 = 1'b1;
  assign CLBLM_R_X13Y151_SLICE_X18Y151_C5 = CLBLM_L_X12Y153_SLICE_X16Y153_AQ;
  assign CLBLM_R_X13Y151_SLICE_X18Y151_C6 = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y155_T1 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_A1 = CLBLM_R_X7Y145_SLICE_X9Y145_CQ;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_A2 = CLBLL_L_X4Y144_SLICE_X4Y144_BQ;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_A3 = CLBLL_L_X4Y144_SLICE_X4Y144_AQ;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_A5 = CLBLL_L_X4Y144_SLICE_X4Y144_CO5;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_A6 = CLBLM_R_X5Y144_SLICE_X6Y144_BO5;
  assign CLBLM_R_X13Y151_SLICE_X18Y151_D1 = 1'b1;
  assign CLBLM_R_X13Y151_SLICE_X18Y151_D2 = 1'b1;
  assign CLBLM_R_X13Y151_SLICE_X18Y151_D3 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_B1 = CLBLL_L_X4Y154_SLICE_X5Y154_AQ;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_B2 = CLBLL_L_X4Y144_SLICE_X4Y144_BQ;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_B3 = CLBLM_R_X5Y144_SLICE_X6Y144_BO6;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_B5 = CLBLL_L_X4Y144_SLICE_X4Y144_CO5;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_B6 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_C1 = CLBLM_R_X3Y145_SLICE_X2Y145_BQ;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_C2 = CLBLM_R_X5Y144_SLICE_X6Y144_AQ;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_C3 = CLBLM_R_X3Y145_SLICE_X2Y145_A5Q;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_C4 = CLBLM_R_X3Y145_SLICE_X3Y145_CQ;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_C5 = CLBLM_R_X3Y144_SLICE_X3Y144_CO6;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_C6 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_D1 = CLBLL_L_X4Y144_SLICE_X5Y144_AQ;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_D2 = CLBLL_L_X4Y144_SLICE_X5Y144_A5Q;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_D3 = CLBLM_L_X8Y144_SLICE_X11Y144_BO6;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_D4 = CLBLM_R_X7Y142_SLICE_X8Y142_DO6;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_D5 = CLBLL_L_X4Y143_SLICE_X4Y143_AQ;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_D6 = CLBLL_L_X4Y144_SLICE_X5Y144_BQ;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_A1 = CLBLM_R_X5Y155_SLICE_X6Y155_AQ;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_A3 = CLBLL_L_X4Y144_SLICE_X5Y144_AQ;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_A4 = CLBLM_R_X7Y142_SLICE_X8Y142_DO6;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_A5 = CLBLL_L_X4Y144_SLICE_X5Y144_CO5;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_A6 = CLBLL_L_X4Y143_SLICE_X4Y143_CO6;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_AX = CLBLL_L_X4Y144_SLICE_X5Y144_CO6;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_B1 = CLBLL_L_X4Y143_SLICE_X4Y143_AQ;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_B2 = CLBLL_L_X4Y144_SLICE_X5Y144_BQ;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_B3 = CLBLL_L_X4Y143_SLICE_X4Y143_CO5;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_B5 = CLBLL_L_X4Y144_SLICE_X5Y144_CO5;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_B6 = CLBLL_L_X4Y149_SLICE_X5Y149_DQ;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_C1 = CLBLL_L_X4Y143_SLICE_X5Y143_AO6;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_C2 = CLBLM_L_X10Y145_SLICE_X12Y145_AQ;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_C3 = CLBLM_L_X8Y145_SLICE_X11Y145_AQ;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_C5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_C6 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_A1 = CLBLM_L_X8Y148_SLICE_X10Y148_DO6;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_D1 = CLBLM_R_X3Y144_SLICE_X2Y144_A5Q;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_D2 = CLBLM_R_X3Y145_SLICE_X3Y145_A5Q;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_D3 = CLBLL_L_X4Y145_SLICE_X5Y145_BO5;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_D4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_D5 = CLBLM_R_X3Y149_SLICE_X3Y149_B5Q;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_D6 = CLBLM_R_X7Y145_SLICE_X8Y145_C5Q;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_A2 = CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_A3 = CLBLM_L_X10Y148_SLICE_X13Y148_AQ;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_A5 = CLBLM_L_X10Y150_SLICE_X13Y150_AQ;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_A6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_B1 = 1'b1;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_B4 = 1'b1;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_B5 = CLBLL_L_X4Y148_SLICE_X4Y148_CQ;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_B6 = CLBLM_L_X10Y150_SLICE_X13Y150_A5Q;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_C1 = CLBLL_L_X4Y146_SLICE_X5Y146_A5Q;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_C2 = CLBLM_L_X10Y148_SLICE_X13Y148_AQ;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_C3 = CLBLM_R_X7Y152_SLICE_X9Y152_CQ;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_C4 = CLBLM_L_X8Y149_SLICE_X11Y149_CQ;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_C5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_C6 = 1'b1;
  assign LIOB33_X0Y131_IOB_X0Y131_O = CLBLM_R_X7Y142_SLICE_X8Y142_AO5;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOB33_X0Y131_IOB_X0Y132_O = CLBLM_R_X5Y142_SLICE_X7Y142_AQ;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_D1 = CLBLM_L_X8Y145_SLICE_X10Y145_CO5;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_D2 = CLBLM_R_X3Y151_SLICE_X3Y151_AO6;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_D3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_D4 = CLBLM_R_X5Y144_SLICE_X7Y144_AQ;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_D5 = CLBLM_L_X10Y148_SLICE_X13Y148_CO5;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_D6 = CLBLM_L_X10Y144_SLICE_X13Y144_AQ;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_A1 = CLBLM_L_X10Y149_SLICE_X13Y149_DQ;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_A3 = CLBLL_L_X4Y146_SLICE_X5Y146_A5Q;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_A4 = CLBLM_L_X10Y148_SLICE_X12Y148_CQ;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_A5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_A6 = 1'b1;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_B1 = CLBLL_L_X4Y145_SLICE_X5Y145_DO6;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_B2 = CLBLM_L_X10Y148_SLICE_X12Y148_BQ;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_B3 = CLBLM_L_X10Y146_SLICE_X12Y146_BQ;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_B5 = 1'b1;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_B6 = CLBLM_L_X8Y151_SLICE_X10Y151_CQ;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_C2 = CLBLM_L_X10Y148_SLICE_X12Y148_CQ;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_C3 = CLBLM_L_X10Y148_SLICE_X12Y148_BQ;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_C4 = CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_C5 = CLBLM_L_X10Y148_SLICE_X12Y148_DO6;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_C6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_D1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_D2 = CLBLM_L_X10Y148_SLICE_X13Y148_CO6;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_D3 = CLBLM_R_X5Y144_SLICE_X7Y144_AQ;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_D4 = CLBLL_L_X2Y151_SLICE_X1Y151_BO6;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_D5 = 1'b1;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_D6 = CLBLM_L_X10Y144_SLICE_X13Y144_AQ;
  assign CLBLM_R_X13Y152_SLICE_X19Y152_A1 = 1'b1;
  assign CLBLM_R_X13Y152_SLICE_X19Y152_A2 = 1'b1;
  assign CLBLM_R_X13Y152_SLICE_X19Y152_A3 = 1'b1;
  assign CLBLM_R_X13Y152_SLICE_X19Y152_A4 = 1'b1;
  assign CLBLM_R_X13Y152_SLICE_X19Y152_A5 = 1'b1;
  assign CLBLM_R_X13Y152_SLICE_X19Y152_A6 = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_D1 = LIOB33_X0Y61_IOB_X0Y61_I;
  assign CLBLM_R_X13Y152_SLICE_X19Y152_B1 = 1'b1;
  assign CLBLM_R_X13Y152_SLICE_X19Y152_B2 = 1'b1;
  assign CLBLM_R_X13Y152_SLICE_X19Y152_B3 = 1'b1;
  assign CLBLM_R_X13Y152_SLICE_X19Y152_B4 = 1'b1;
  assign CLBLM_R_X13Y152_SLICE_X19Y152_B5 = 1'b1;
  assign CLBLM_R_X13Y152_SLICE_X19Y152_B6 = 1'b1;
  assign CLBLM_R_X13Y152_SLICE_X19Y152_C1 = 1'b1;
  assign CLBLM_R_X13Y152_SLICE_X19Y152_C2 = 1'b1;
  assign CLBLM_R_X13Y152_SLICE_X19Y152_C3 = 1'b1;
  assign CLBLM_R_X13Y152_SLICE_X19Y152_C4 = 1'b1;
  assign CLBLM_R_X13Y152_SLICE_X19Y152_C5 = 1'b1;
  assign CLBLM_R_X13Y152_SLICE_X19Y152_C6 = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_T1 = 1'b1;
  assign RIOI3_X105Y191_OLOGIC_X1Y192_D1 = CLBLM_R_X11Y151_SLICE_X15Y151_AQ;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_D4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_D1 = LIOB33_X0Y71_IOB_X0Y71_I;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_D5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X13Y152_SLICE_X19Y152_D1 = 1'b1;
  assign CLBLM_R_X13Y152_SLICE_X19Y152_D2 = 1'b1;
  assign CLBLM_R_X13Y152_SLICE_X19Y152_D3 = 1'b1;
  assign CLBLM_R_X13Y152_SLICE_X19Y152_D4 = 1'b1;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_D6 = CLBLM_L_X12Y152_SLICE_X17Y152_AQ;
  assign CLBLM_R_X13Y152_SLICE_X19Y152_D5 = 1'b1;
  assign CLBLM_R_X13Y152_SLICE_X19Y152_D6 = 1'b1;
  assign RIOI3_X105Y191_OLOGIC_X1Y192_T1 = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_T1 = 1'b1;
  assign RIOI3_X105Y191_OLOGIC_X1Y191_D1 = CLBLM_L_X10Y149_SLICE_X12Y149_AQ;
  assign CLBLM_R_X13Y152_SLICE_X18Y152_A1 = CLBLM_L_X12Y153_SLICE_X17Y153_DO6;
  assign CLBLM_R_X13Y152_SLICE_X18Y152_A2 = CLBLM_L_X12Y152_SLICE_X17Y152_CQ;
  assign CLBLM_R_X13Y152_SLICE_X18Y152_A3 = CLBLM_L_X12Y154_SLICE_X16Y154_AQ;
  assign CLBLM_R_X13Y152_SLICE_X18Y152_A4 = CLBLM_L_X12Y152_SLICE_X16Y152_AQ;
  assign CLBLM_R_X13Y152_SLICE_X18Y152_A5 = CLBLM_L_X12Y153_SLICE_X16Y153_AQ;
  assign CLBLM_R_X13Y152_SLICE_X18Y152_A6 = CLBLM_L_X12Y152_SLICE_X17Y152_BQ;
  assign CLBLM_R_X13Y152_SLICE_X18Y152_B1 = CLBLM_L_X12Y153_SLICE_X16Y153_AQ;
  assign CLBLM_R_X13Y152_SLICE_X18Y152_B2 = CLBLM_L_X12Y152_SLICE_X17Y152_CQ;
  assign CLBLM_R_X13Y152_SLICE_X18Y152_B3 = CLBLM_L_X12Y154_SLICE_X16Y154_AQ;
  assign CLBLM_R_X13Y152_SLICE_X18Y152_B4 = CLBLM_L_X12Y152_SLICE_X16Y152_AQ;
  assign CLBLM_R_X13Y152_SLICE_X18Y152_B5 = CLBLM_L_X12Y152_SLICE_X17Y152_BQ;
  assign CLBLM_R_X13Y152_SLICE_X18Y152_B6 = CLBLM_L_X12Y153_SLICE_X17Y153_CO6;
  assign RIOI3_X105Y191_OLOGIC_X1Y191_T1 = 1'b1;
  assign CLBLM_R_X13Y152_SLICE_X18Y152_C1 = 1'b1;
  assign CLBLM_R_X13Y152_SLICE_X18Y152_C2 = 1'b1;
  assign CLBLM_R_X13Y152_SLICE_X18Y152_C3 = 1'b1;
  assign CLBLM_R_X13Y152_SLICE_X18Y152_C4 = 1'b1;
  assign CLBLM_R_X13Y152_SLICE_X18Y152_C5 = 1'b1;
  assign CLBLM_R_X13Y152_SLICE_X18Y152_C6 = 1'b1;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_A1 = CLBLM_R_X7Y151_SLICE_X8Y151_AQ;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_A1 = 1'b1;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_A3 = CLBLL_L_X4Y145_SLICE_X4Y145_AQ;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_A4 = CLBLM_R_X5Y152_SLICE_X7Y152_DO6;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_A5 = CLBLM_L_X10Y145_SLICE_X13Y145_AQ;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_A6 = CLBLM_R_X7Y149_SLICE_X8Y149_DQ;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_AX = CLBLL_L_X4Y146_SLICE_X4Y146_CO6;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_A3 = CLBLM_R_X11Y146_SLICE_X14Y146_CQ;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_B1 = CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_B2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_B3 = CLBLM_R_X7Y145_SLICE_X8Y145_DO6;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_B4 = CLBLM_R_X3Y143_SLICE_X2Y143_AQ;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_B6 = 1'b1;
  assign CLBLM_R_X13Y152_SLICE_X18Y152_D2 = 1'b1;
  assign CLBLM_R_X13Y152_SLICE_X18Y152_D3 = 1'b1;
  assign CLBLM_R_X13Y152_SLICE_X18Y152_D5 = 1'b1;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_C1 = CLBLM_R_X7Y147_SLICE_X8Y147_AQ;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_C2 = CLBLL_L_X4Y145_SLICE_X4Y145_CQ;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_C3 = CLBLM_R_X11Y146_SLICE_X14Y146_AQ;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_C5 = CLBLL_L_X4Y145_SLICE_X4Y145_BO5;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_C6 = CLBLM_L_X10Y146_SLICE_X12Y146_C5Q;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_D1 = CLBLM_R_X3Y149_SLICE_X3Y149_B5Q;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_D2 = 1'b1;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_D3 = CLBLM_R_X3Y145_SLICE_X3Y145_A5Q;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_D4 = 1'b1;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_D5 = 1'b1;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_D6 = 1'b1;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_A1 = CLBLL_L_X4Y147_SLICE_X5Y147_CQ;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_A3 = CLBLL_L_X4Y142_SLICE_X5Y142_AQ;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_A5 = CLBLM_R_X11Y145_SLICE_X14Y145_AQ;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_A6 = LIOB33_X0Y53_IOB_X0Y53_I;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_B1 = CLBLM_R_X3Y143_SLICE_X3Y143_B5Q;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_B2 = CLBLM_R_X3Y144_SLICE_X2Y144_A5Q;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_B3 = CLBLM_R_X3Y144_SLICE_X2Y144_AQ;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_B4 = CLBLL_L_X4Y145_SLICE_X4Y145_A5Q;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_B5 = CLBLL_L_X4Y148_SLICE_X4Y148_C5Q;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_B6 = 1'b1;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_C2 = LIOB33_X0Y53_IOB_X0Y53_I;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_C3 = CLBLL_L_X4Y147_SLICE_X5Y147_CQ;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_C4 = CLBLL_L_X4Y142_SLICE_X5Y142_AQ;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_C5 = CLBLM_R_X5Y145_SLICE_X6Y145_A5Q;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_C6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign LIOB33_X0Y147_IOB_X0Y147_O = LIOB33_X0Y71_IOB_X0Y71_I;
  assign LIOB33_X0Y147_IOB_X0Y148_O = LIOB33_X0Y61_IOB_X0Y61_I;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOB33_X0Y133_IOB_X0Y134_O = CLBLM_R_X3Y143_SLICE_X2Y143_CQ;
  assign LIOB33_X0Y133_IOB_X0Y133_O = CLBLM_R_X3Y143_SLICE_X3Y143_A5Q;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_D1 = CLBLM_R_X7Y145_SLICE_X8Y145_C5Q;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_D2 = CLBLM_R_X3Y151_SLICE_X2Y151_AO6;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_D3 = CLBLL_L_X4Y145_SLICE_X4Y145_DO6;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_D4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_D5 = CLBLM_R_X5Y152_SLICE_X7Y152_B5Q;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_D6 = CLBLL_L_X4Y145_SLICE_X5Y145_BO6;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_A1 = CLBLM_R_X11Y147_SLICE_X14Y147_CO6;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_A3 = CLBLM_L_X10Y149_SLICE_X13Y149_AQ;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_A4 = CLBLM_R_X11Y150_SLICE_X15Y150_AQ;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_A6 = CLBLM_L_X8Y149_SLICE_X11Y149_CQ;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_AX = CLBLM_L_X10Y149_SLICE_X13Y149_CO6;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_B1 = 1'b1;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_B3 = CLBLM_R_X7Y145_SLICE_X9Y145_C5Q;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_B4 = CLBLM_L_X10Y150_SLICE_X13Y150_CQ;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_B6 = CLBLM_L_X10Y148_SLICE_X13Y148_CO6;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_D4 = CLBLM_R_X7Y147_SLICE_X9Y147_CO5;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_C1 = CLBLL_L_X4Y148_SLICE_X4Y148_CQ;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_C2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_C3 = CLBLM_L_X12Y148_SLICE_X16Y148_AQ;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_C4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_C5 = CLBLM_R_X11Y147_SLICE_X15Y147_DQ;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_C6 = 1'b1;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_D5 = 1'b1;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_D6 = CLBLM_L_X10Y144_SLICE_X13Y144_AQ;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_D1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_D2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_D3 = CLBLL_L_X4Y146_SLICE_X5Y146_A5Q;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_D4 = 1'b1;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_D5 = 1'b1;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_D6 = CLBLM_R_X11Y153_SLICE_X15Y153_AQ;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_A1 = CLBLM_L_X10Y149_SLICE_X12Y149_DO6;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_A2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_A3 = CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_A4 = CLBLM_R_X11Y147_SLICE_X15Y147_AQ;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_A6 = 1'b1;
  assign RIOI3_X105Y129_ILOGIC_X1Y130_D = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_AX = CLBLM_L_X8Y144_SLICE_X10Y144_CQ;
  assign RIOI3_X105Y129_ILOGIC_X1Y129_D = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_B1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_B3 = CLBLM_R_X7Y145_SLICE_X9Y145_C5Q;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_B4 = CLBLM_L_X8Y148_SLICE_X11Y148_AQ;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_B5 = CLBLM_L_X10Y146_SLICE_X12Y146_BQ;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_B6 = 1'b1;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_C1 = CLBLM_R_X5Y151_SLICE_X6Y151_BQ;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_C2 = CLBLM_L_X10Y150_SLICE_X13Y150_CQ;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_C3 = 1'b1;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_C4 = CLBLM_L_X10Y145_SLICE_X12Y145_CQ;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_C5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_C6 = CLBLM_L_X10Y149_SLICE_X13Y149_BQ;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_CE = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_A4 = CLBLM_L_X8Y148_SLICE_X11Y148_CO6;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_D1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_D2 = CLBLM_R_X5Y144_SLICE_X7Y144_AQ;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_D3 = CLBLM_L_X10Y150_SLICE_X13Y150_A5Q;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_D4 = CLBLL_L_X4Y154_SLICE_X4Y154_CO6;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_D5 = 1'b1;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_D6 = CLBLM_L_X10Y144_SLICE_X13Y144_AQ;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_A1 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_A2 = CLBLM_R_X11Y153_SLICE_X14Y153_BQ;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_SR = CLBLM_R_X11Y151_SLICE_X15Y151_CO6;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_A3 = CLBLM_R_X11Y151_SLICE_X14Y151_AQ;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_A4 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_A5 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_A6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y144_D = RIOB33_X105Y143_IOB_X1Y144_I;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_B1 = 1'b1;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_C2 = CLBLM_R_X5Y151_SLICE_X7Y151_CQ;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_B2 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_B3 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_B4 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_B5 = 1'b1;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_B6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y143_D = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_C1 = 1'b1;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_C4 = CLBLL_L_X4Y154_SLICE_X4Y154_CO6;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_C2 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_C3 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_C4 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_C5 = 1'b1;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_C5 = CLBLL_L_X4Y149_SLICE_X5Y149_BO5;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_C6 = 1'b1;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_C6 = CLBLM_R_X5Y145_SLICE_X7Y145_CQ;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_D1 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_D2 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_D3 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_D4 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_D5 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_D6 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_A1 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_A2 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_A3 = 1'b1;
  assign CLBLM_L_X16Y158_SLICE_X23Y158_C4 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_A4 = 1'b1;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_B6 = CLBLM_L_X10Y150_SLICE_X12Y150_CQ;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_A1 = 1'b1;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_A2 = 1'b1;
  assign CLBLM_L_X16Y158_SLICE_X23Y158_C5 = 1'b1;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_A3 = 1'b1;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_A4 = 1'b1;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_A5 = 1'b1;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_A6 = 1'b1;
  assign CLBLM_L_X16Y158_SLICE_X23Y158_C6 = 1'b1;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_B1 = 1'b1;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_B2 = 1'b1;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_B3 = 1'b1;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_B4 = 1'b1;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_B5 = 1'b1;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_B6 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_B2 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_B3 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_B5 = 1'b1;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_C1 = 1'b1;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_C2 = 1'b1;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_C3 = 1'b1;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_C4 = 1'b1;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_C5 = 1'b1;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_C6 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_C1 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_C2 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_C3 = 1'b1;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_D1 = CLBLM_R_X5Y149_SLICE_X7Y149_AQ;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_C5 = 1'b1;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_D2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_D1 = 1'b1;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_D2 = 1'b1;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_D3 = 1'b1;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_D4 = 1'b1;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_D5 = 1'b1;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_D6 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_D1 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_D2 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_D3 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_D4 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_D5 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_D6 = 1'b1;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_D5 = CLBLL_L_X4Y150_SLICE_X4Y150_AQ;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_A2 = CLBLM_R_X7Y142_SLICE_X8Y142_DO6;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_A3 = CLBLM_R_X11Y143_SLICE_X14Y143_AQ;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_A4 = CLBLM_L_X8Y144_SLICE_X11Y144_AQ;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_A5 = 1'b1;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_D6 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_A1 = CLBLM_L_X8Y149_SLICE_X11Y149_AQ;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_A2 = CLBLM_R_X5Y145_SLICE_X7Y145_AQ;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_A3 = CLBLL_L_X4Y146_SLICE_X4Y146_AQ;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_A5 = CLBLL_L_X4Y151_SLICE_X4Y151_AQ;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_A6 = CLBLM_R_X3Y146_SLICE_X2Y146_AQ;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_A6 = CLBLM_R_X11Y145_SLICE_X14Y145_BQ;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_AX = CLBLM_R_X7Y146_SLICE_X8Y146_BO6;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_B1 = CLBLL_L_X4Y147_SLICE_X5Y147_CQ;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_B2 = CLBLL_L_X4Y146_SLICE_X4Y146_BQ;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_B3 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_B5 = CLBLM_R_X11Y146_SLICE_X15Y146_DQ;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_B6 = CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_B5 = CLBLM_L_X10Y143_SLICE_X13Y143_BQ;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_C2 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_C3 = CLBLM_L_X8Y147_SLICE_X10Y147_CQ;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_C4 = CLBLM_L_X10Y146_SLICE_X13Y146_B5Q;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_C5 = CLBLM_R_X3Y146_SLICE_X2Y146_AQ;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_C6 = 1'b1;
  assign CLBLM_L_X16Y158_SLICE_X23Y158_D5 = 1'b1;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_C4 = CLBLM_L_X12Y144_SLICE_X16Y144_CQ;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_C6 = 1'b1;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_D1 = 1'b1;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_D2 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_D1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_D2 = CLBLL_L_X4Y145_SLICE_X4Y145_CQ;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_D3 = CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_D4 = CLBLM_R_X7Y147_SLICE_X8Y147_AQ;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_D5 = CLBLM_R_X5Y145_SLICE_X7Y145_AQ;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_D6 = CLBLM_R_X7Y145_SLICE_X8Y145_AQ;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_D3 = 1'b1;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_D4 = 1'b1;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_D5 = 1'b1;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_D6 = 1'b1;
  assign CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_CE = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_A1 = CLBLM_L_X8Y149_SLICE_X11Y149_AQ;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_A2 = CLBLL_L_X4Y147_SLICE_X5Y147_BQ;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_A3 = CLBLL_L_X4Y146_SLICE_X5Y146_AQ;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_A4 = CLBLM_R_X7Y146_SLICE_X8Y146_C5Q;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_A5 = CLBLL_L_X4Y151_SLICE_X4Y151_AQ;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOB33_X0Y135_IOB_X0Y136_O = CLBLL_L_X2Y145_SLICE_X1Y145_AQ;
  assign LIOB33_X0Y135_IOB_X0Y135_O = CLBLM_R_X3Y142_SLICE_X2Y142_BQ;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_AX = CLBLL_L_X4Y146_SLICE_X5Y146_BO6;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_B1 = CLBLM_R_X7Y146_SLICE_X8Y146_DQ;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_B2 = CLBLL_L_X4Y147_SLICE_X5Y147_BQ;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_B4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_B5 = CLBLM_R_X3Y146_SLICE_X3Y146_BQ;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_B6 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_C1 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_C2 = CLBLL_L_X4Y146_SLICE_X5Y146_CQ;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_C3 = CLBLL_L_X4Y145_SLICE_X5Y145_CO6;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_C4 = CLBLM_L_X12Y144_SLICE_X16Y144_CQ;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_C5 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_D1 = CLBLM_R_X7Y146_SLICE_X8Y146_C5Q;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_D2 = CLBLM_R_X11Y147_SLICE_X14Y147_BQ;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_D3 = CLBLM_R_X3Y147_SLICE_X3Y147_BQ;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_D4 = CLBLM_L_X8Y146_SLICE_X10Y146_BQ;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_D5 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_D6 = CLBLL_L_X4Y147_SLICE_X5Y147_BQ;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_A1 = CLBLM_L_X10Y150_SLICE_X13Y150_AQ;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_A2 = CLBLM_R_X11Y152_SLICE_X15Y152_BQ;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_A3 = CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_A5 = CLBLM_R_X7Y149_SLICE_X9Y149_DO6;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_A6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_AX = CLBLM_L_X10Y149_SLICE_X12Y149_AO6;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_B2 = CLBLM_L_X10Y150_SLICE_X13Y150_BQ;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_B3 = CLBLM_L_X12Y149_SLICE_X17Y149_BQ;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_B4 = CLBLM_R_X11Y147_SLICE_X14Y147_CO6;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_B5 = CLBLM_L_X8Y147_SLICE_X10Y147_BQ;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X16Y158_SLICE_X22Y158_B2 = 1'b1;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_C2 = CLBLM_R_X5Y145_SLICE_X6Y145_AQ;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_C4 = CLBLM_R_X11Y151_SLICE_X15Y151_A5Q;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_C5 = CLBLM_L_X10Y148_SLICE_X13Y148_CO5;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_C6 = 1'b1;
  assign CLBLM_L_X16Y158_SLICE_X22Y158_B3 = 1'b1;
  assign CLBLM_L_X16Y158_SLICE_X22Y158_B4 = 1'b1;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X16Y158_SLICE_X22Y158_B5 = 1'b1;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_D1 = CLBLL_L_X4Y149_SLICE_X5Y149_A5Q;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_D2 = CLBLM_L_X8Y146_SLICE_X10Y146_BQ;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_D3 = CLBLM_R_X5Y144_SLICE_X7Y144_CQ;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_D4 = CLBLM_L_X10Y150_SLICE_X13Y150_A5Q;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_D5 = CLBLM_L_X10Y150_SLICE_X13Y150_AQ;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_D6 = 1'b1;
  assign CLBLM_L_X16Y158_SLICE_X22Y158_B6 = 1'b1;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_A1 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_A2 = CLBLM_R_X11Y149_SLICE_X14Y149_BQ;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_A3 = CLBLM_L_X10Y150_SLICE_X12Y150_AQ;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_A6 = CLBLM_R_X11Y147_SLICE_X14Y147_CO6;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_C4 = CLBLM_R_X5Y151_SLICE_X7Y151_CQ;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_AX = CLBLM_L_X10Y149_SLICE_X12Y149_BO6;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_C5 = CLBLM_L_X10Y149_SLICE_X13Y149_BQ;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_B1 = 1'b1;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_B2 = 1'b1;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_B3 = CLBLM_R_X5Y148_SLICE_X6Y148_BQ;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_B4 = CLBLM_L_X10Y150_SLICE_X13Y150_BQ;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_C6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X16Y158_SLICE_X22Y158_C1 = 1'b1;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_BX = CLBLM_L_X10Y147_SLICE_X12Y147_DO6;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_C2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_C3 = CLBLM_L_X10Y149_SLICE_X13Y149_A5Q;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_C4 = CLBLM_L_X10Y147_SLICE_X12Y147_CQ;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_C5 = 1'b1;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_C6 = CLBLM_L_X10Y149_SLICE_X12Y149_BO5;
  assign CLBLM_L_X16Y158_SLICE_X22Y158_C2 = 1'b1;
  assign CLBLM_L_X16Y158_SLICE_X22Y158_C3 = 1'b1;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X16Y158_SLICE_X22Y158_C4 = 1'b1;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_CX = CLBLM_L_X8Y147_SLICE_X11Y147_AO6;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_D1 = CLBLM_L_X10Y147_SLICE_X12Y147_DO5;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_D2 = CLBLM_R_X7Y148_SLICE_X8Y148_CQ;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_D3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_D4 = CLBLM_L_X12Y152_SLICE_X16Y152_BQ;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_D5 = 1'b1;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_D6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X16Y158_SLICE_X22Y158_C5 = 1'b1;
  assign CLBLM_L_X16Y158_SLICE_X22Y158_C6 = 1'b1;
  assign CLBLM_L_X16Y158_SLICE_X22Y158_D1 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_A1 = CLBLM_L_X10Y145_SLICE_X13Y145_CQ;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_A2 = CLBLM_L_X12Y144_SLICE_X16Y144_CQ;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_A3 = CLBLM_L_X12Y144_SLICE_X16Y144_BQ;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_A4 = CLBLM_L_X12Y144_SLICE_X16Y144_AQ;
  assign CLBLM_L_X16Y158_SLICE_X22Y158_D2 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_A5 = CLBLM_L_X12Y145_SLICE_X16Y145_AQ;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_A6 = 1'b1;
  assign CLBLM_L_X16Y158_SLICE_X22Y158_D3 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_B1 = CLBLM_L_X10Y145_SLICE_X13Y145_CQ;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_B2 = CLBLM_L_X10Y146_SLICE_X12Y146_BQ;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_B3 = CLBLM_L_X10Y143_SLICE_X13Y143_BQ;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_B4 = CLBLM_R_X7Y142_SLICE_X8Y142_BQ;
  assign CLBLM_L_X16Y158_SLICE_X22Y158_D4 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_B5 = CLBLM_R_X11Y146_SLICE_X15Y146_AQ;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_B6 = CLBLM_R_X7Y142_SLICE_X8Y142_CQ;
  assign CLBLM_L_X16Y158_SLICE_X22Y158_D5 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_C1 = CLBLM_L_X12Y144_SLICE_X16Y144_AQ;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_C2 = CLBLM_L_X12Y144_SLICE_X16Y144_BQ;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_C3 = CLBLM_L_X12Y144_SLICE_X16Y144_CQ;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_C4 = 1'b1;
  assign CLBLM_L_X16Y158_SLICE_X22Y158_D6 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_C5 = CLBLM_L_X12Y145_SLICE_X16Y145_AQ;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_C6 = CLBLM_L_X10Y146_SLICE_X12Y146_BQ;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_D1 = CLBLM_R_X11Y145_SLICE_X15Y145_AQ;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_D2 = CLBLM_L_X10Y144_SLICE_X13Y144_CQ;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_D3 = CLBLM_R_X11Y144_SLICE_X14Y144_DO6;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_D4 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_D5 = CLBLM_R_X11Y145_SLICE_X15Y145_DO6;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_D6 = CLBLM_R_X11Y144_SLICE_X15Y144_BO6;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_A1 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_A1 = CLBLL_L_X4Y147_SLICE_X4Y147_DO6;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_A2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_A3 = CLBLL_L_X4Y147_SLICE_X4Y147_AQ;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_A4 = CLBLM_R_X3Y148_SLICE_X2Y148_BQ;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_A6 = CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_A3 = CLBLM_R_X11Y144_SLICE_X14Y144_AQ;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_A5 = CLBLM_R_X5Y145_SLICE_X6Y145_AQ;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_B2 = CLBLM_L_X8Y148_SLICE_X11Y148_BO6;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_B3 = 1'b1;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_B4 = CLBLM_R_X3Y145_SLICE_X2Y145_BQ;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_B5 = CLBLM_L_X8Y150_SLICE_X10Y150_BQ;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_B1 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_C1 = CLBLM_R_X7Y149_SLICE_X8Y149_AQ;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_C2 = 1'b1;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_C5 = CLBLL_L_X4Y147_SLICE_X4Y147_DO6;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_C6 = CLBLM_R_X3Y147_SLICE_X3Y147_C5Q;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_C1 = CLBLM_L_X12Y144_SLICE_X16Y144_BQ;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_C2 = CLBLM_R_X11Y144_SLICE_X15Y144_AO5;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_C3 = CLBLM_R_X7Y144_SLICE_X8Y144_DQ;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_C4 = CLBLM_R_X7Y142_SLICE_X8Y142_DO6;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_C5 = CLBLM_R_X11Y144_SLICE_X14Y144_BQ;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_C5 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_D1 = CLBLL_L_X4Y143_SLICE_X4Y143_BQ;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_D2 = CLBLL_L_X4Y148_SLICE_X4Y148_CQ;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_D3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_D4 = CLBLM_L_X8Y148_SLICE_X10Y148_DO5;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_D5 = 1'b1;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_D6 = CLBLM_R_X7Y144_SLICE_X9Y144_CQ;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_C6 = CLBLM_R_X3Y148_SLICE_X2Y148_DQ;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_D1 = CLBLM_R_X11Y143_SLICE_X14Y143_BQ;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_D2 = CLBLM_R_X7Y144_SLICE_X8Y144_DQ;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_D3 = CLBLM_R_X11Y145_SLICE_X14Y145_BQ;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_D4 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_D5 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_D6 = CLBLM_L_X12Y145_SLICE_X16Y145_BQ;
  assign LIOB33_X0Y137_IOB_X0Y137_O = CLBLM_R_X3Y142_SLICE_X2Y142_AQ;
  assign LIOB33_X0Y137_IOB_X0Y138_O = CLBLM_R_X3Y143_SLICE_X3Y143_BQ;
  assign LIOB33_X0Y159_IOB_X0Y160_O = RIOB33_X105Y107_IOB_X1Y107_I;
  assign LIOI3_X0Y151_OLOGIC_X0Y152_D1 = LIOB33_X0Y65_IOB_X0Y66_I;
  assign LIOI3_SING_X0Y50_ILOGIC_X0Y50_D = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign LIOI3_X0Y151_OLOGIC_X0Y152_T1 = 1'b1;
  assign RIOI3_X105Y195_OLOGIC_X1Y196_D1 = CLBLM_R_X11Y153_SLICE_X14Y153_BQ;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_A1 = CLBLM_R_X5Y152_SLICE_X7Y152_DO5;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_A3 = CLBLL_L_X4Y147_SLICE_X5Y147_AQ;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_A4 = CLBLM_L_X8Y146_SLICE_X10Y146_CQ;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_A5 = 1'b1;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_A6 = CLBLM_R_X7Y146_SLICE_X9Y146_AQ;
  assign LIOB33_X0Y159_IOB_X0Y159_O = RIOB33_X105Y117_IOB_X1Y117_I;
  assign LIOI3_X0Y151_OLOGIC_X0Y151_D1 = LIOB33_X0Y65_IOB_X0Y65_I;
  assign RIOI3_X105Y195_OLOGIC_X1Y196_T1 = 1'b1;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_B1 = CLBLL_L_X4Y147_SLICE_X5Y147_DO6;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_B2 = CLBLM_R_X7Y143_SLICE_X9Y143_BQ;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_B4 = CLBLM_R_X7Y147_SLICE_X8Y147_AQ;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_B5 = CLBLM_R_X7Y154_SLICE_X8Y154_DO6;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_B6 = 1'b1;
  assign LIOI3_X0Y151_OLOGIC_X0Y151_T1 = 1'b1;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_C2 = CLBLM_R_X5Y146_SLICE_X6Y146_A5Q;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_C3 = CLBLM_R_X5Y153_SLICE_X6Y153_A5Q;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_C4 = CLBLL_L_X4Y146_SLICE_X5Y146_CQ;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_C5 = CLBLM_R_X7Y151_SLICE_X8Y151_A5Q;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_C6 = CLBLM_L_X12Y146_SLICE_X16Y146_AQ;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_D1 = CLBLL_L_X2Y155_SLICE_X1Y155_AO6;
  assign RIOI3_X105Y195_OLOGIC_X1Y195_D1 = CLBLM_R_X11Y151_SLICE_X14Y151_AQ;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_D2 = CLBLM_R_X3Y156_SLICE_X2Y156_CO6;
  assign RIOI3_X105Y195_OLOGIC_X1Y195_T1 = 1'b1;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_D1 = CLBLL_L_X4Y147_SLICE_X5Y147_BQ;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_D2 = CLBLM_L_X10Y147_SLICE_X12Y147_AQ;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_D3 = CLBLL_L_X4Y146_SLICE_X4Y146_DO6;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_D4 = CLBLM_R_X3Y146_SLICE_X3Y146_BQ;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_D5 = CLBLM_R_X11Y146_SLICE_X14Y146_AQ;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_D6 = CLBLM_R_X11Y147_SLICE_X14Y147_BQ;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_D3 = CLBLM_R_X3Y154_SLICE_X3Y154_DO6;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_D4 = CLBLL_L_X4Y153_SLICE_X5Y153_DO6;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_D5 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_A1 = CLBLM_R_X5Y152_SLICE_X7Y152_BQ;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_A3 = CLBLM_L_X10Y151_SLICE_X13Y151_AQ;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_A5 = CLBLM_R_X11Y151_SLICE_X14Y151_BO6;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_A6 = CLBLM_L_X10Y151_SLICE_X12Y151_CQ;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_D6 = CLBLM_R_X3Y153_SLICE_X2Y153_BO6;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_B1 = CLBLM_R_X5Y152_SLICE_X7Y152_BQ;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_B2 = CLBLM_L_X10Y151_SLICE_X13Y151_BQ;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_B3 = CLBLM_R_X7Y143_SLICE_X8Y143_AQ;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_B4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_B5 = CLBLM_R_X11Y151_SLICE_X14Y151_CO5;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_D1 = CLBLL_L_X36Y146_SLICE_X54Y146_AO6;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_C1 = CLBLM_R_X5Y150_SLICE_X6Y150_DQ;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_C2 = CLBLM_L_X10Y151_SLICE_X13Y151_CQ;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_C3 = CLBLM_R_X11Y153_SLICE_X14Y153_BO5;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_C4 = CLBLM_R_X11Y152_SLICE_X14Y152_CQ;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_C5 = CLBLM_R_X11Y154_SLICE_X15Y154_CO6;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_T1 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_D1 = CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_D2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_D3 = CLBLM_L_X10Y151_SLICE_X13Y151_DQ;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_D4 = CLBLM_R_X11Y149_SLICE_X14Y149_CQ;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_D6 = CLBLM_R_X11Y152_SLICE_X14Y152_BQ;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_D1 = RIOB33_X105Y125_IOB_X1Y126_I;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_A1 = CLBLM_R_X7Y151_SLICE_X8Y151_BQ;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_A3 = CLBLM_L_X10Y151_SLICE_X12Y151_AQ;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_A4 = CLBLM_L_X10Y154_SLICE_X13Y154_BQ;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_A5 = CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_A6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_T1 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_B2 = CLBLM_L_X10Y151_SLICE_X12Y151_BQ;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_B3 = CLBLM_L_X10Y150_SLICE_X12Y150_AQ;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_B5 = CLBLM_R_X11Y147_SLICE_X14Y147_CO6;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_B6 = CLBLM_L_X8Y153_SLICE_X11Y153_CQ;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_C1 = CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_C2 = CLBLM_L_X10Y144_SLICE_X12Y144_CQ;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_C3 = CLBLM_L_X10Y151_SLICE_X12Y151_DQ;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_C4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_C5 = CLBLM_L_X10Y151_SLICE_X12Y151_CQ;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_D1 = CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_D2 = CLBLM_R_X3Y150_SLICE_X3Y150_A5Q;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_D3 = CLBLM_L_X10Y151_SLICE_X12Y151_DQ;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_D4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_D6 = CLBLM_L_X10Y148_SLICE_X12Y148_DO6;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_A2 = CLBLM_R_X11Y145_SLICE_X15Y145_BQ;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_A3 = CLBLM_R_X11Y145_SLICE_X15Y145_AQ;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_A4 = CLBLL_L_X4Y145_SLICE_X5Y145_DO6;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_A5 = 1'b1;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_A6 = CLBLM_L_X10Y147_SLICE_X12Y147_CQ;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_B2 = CLBLM_R_X11Y145_SLICE_X15Y145_BQ;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_B3 = CLBLM_L_X10Y154_SLICE_X12Y154_AQ;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_B4 = CLBLL_L_X4Y145_SLICE_X5Y145_DO6;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_B5 = CLBLM_L_X12Y145_SLICE_X16Y145_BQ;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_B6 = 1'b1;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_C1 = CLBLM_R_X11Y144_SLICE_X15Y144_AO5;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_C2 = CLBLM_R_X7Y142_SLICE_X8Y142_DO6;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_C3 = CLBLM_L_X12Y144_SLICE_X16Y144_BQ;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_C4 = CLBLM_R_X15Y151_SLICE_X20Y151_AQ;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_C5 = CLBLM_R_X11Y146_SLICE_X15Y146_BQ;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_C6 = CLBLM_R_X7Y142_SLICE_X8Y142_BQ;
  assign RIOI3_X105Y133_ILOGIC_X1Y134_D = RIOB33_X105Y133_IOB_X1Y134_I;
  assign RIOI3_X105Y133_ILOGIC_X1Y133_D = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_D1 = CLBLM_R_X7Y146_SLICE_X9Y146_CQ;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_D2 = CLBLM_L_X10Y148_SLICE_X12Y148_BQ;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_D3 = 1'b1;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_D4 = CLBLM_R_X11Y145_SLICE_X15Y145_BQ;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_D5 = 1'b1;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_D6 = 1'b1;
  assign RIOI3_X105Y123_ILOGIC_X1Y124_D = RIOB33_X105Y123_IOB_X1Y124_I;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_A1 = 1'b1;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_A2 = CLBLM_R_X7Y148_SLICE_X8Y148_D5Q;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_A3 = CLBLL_L_X4Y148_SLICE_X4Y148_AQ;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_A5 = CLBLM_R_X5Y148_SLICE_X6Y148_AQ;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_A6 = CLBLM_R_X5Y152_SLICE_X7Y152_DO5;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_A2 = 1'b1;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_A3 = CLBLM_R_X5Y142_SLICE_X7Y142_AQ;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_B1 = CLBLM_L_X10Y145_SLICE_X12Y145_CQ;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_B3 = 1'b1;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_B4 = 1'b1;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_B6 = CLBLM_R_X5Y149_SLICE_X6Y149_BQ;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_A5 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_A6 = CLBLM_R_X11Y145_SLICE_X14Y145_CO6;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_C2 = CLBLL_L_X4Y144_SLICE_X4Y144_AQ;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_C3 = CLBLM_R_X3Y149_SLICE_X3Y149_DQ;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_C4 = CLBLM_R_X5Y148_SLICE_X7Y148_BQ;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_C6 = 1'b1;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_B5 = CLBLM_R_X11Y149_SLICE_X14Y149_AQ;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_C1 = CLBLM_R_X11Y143_SLICE_X14Y143_CO5;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_C2 = CLBLM_R_X11Y145_SLICE_X14Y145_AQ;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_C3 = CLBLM_L_X12Y144_SLICE_X16Y144_CQ;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_C4 = CLBLM_R_X7Y142_SLICE_X8Y142_CQ;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_D1 = CLBLM_R_X3Y146_SLICE_X3Y146_BQ;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_D2 = CLBLM_L_X8Y148_SLICE_X10Y148_A5Q;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_D3 = CLBLL_L_X4Y148_SLICE_X4Y148_DQ;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_D4 = CLBLM_R_X11Y150_SLICE_X14Y150_BO6;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_D6 = CLBLM_L_X10Y147_SLICE_X12Y147_AQ;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_D1 = CLBLM_R_X11Y143_SLICE_X14Y143_CO5;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_D2 = CLBLM_R_X11Y149_SLICE_X14Y149_CQ;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_D3 = CLBLM_L_X12Y144_SLICE_X16Y144_CQ;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_D4 = CLBLM_R_X11Y148_SLICE_X15Y148_A5Q;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_D5 = CLBLM_R_X7Y142_SLICE_X8Y142_DO6;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_D6 = CLBLM_L_X10Y146_SLICE_X12Y146_BQ;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_A1 = CLBLM_L_X10Y147_SLICE_X12Y147_AQ;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_A2 = CLBLM_L_X8Y149_SLICE_X11Y149_AQ;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_A3 = CLBLL_L_X4Y148_SLICE_X5Y148_AQ;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_A4 = CLBLL_L_X4Y151_SLICE_X4Y151_AQ;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_A5 = CLBLL_L_X4Y147_SLICE_X4Y147_AQ;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_B1 = CLBLM_R_X3Y148_SLICE_X3Y148_CQ;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_B2 = CLBLL_L_X4Y148_SLICE_X5Y148_BQ;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_B3 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X2Y134_SLICE_X0Y134_A4 = CLBLM_R_X5Y145_SLICE_X6Y145_DO5;
  assign CLBLL_L_X2Y134_SLICE_X0Y134_A5 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X0Y134_A6 = 1'b1;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_B4 = CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_B6 = CLBLM_R_X7Y144_SLICE_X8Y144_CQ;
  assign CLBLL_L_X2Y134_SLICE_X0Y134_A1 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X0Y134_A2 = CLBLL_L_X2Y141_SLICE_X0Y141_BO6;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_C1 = CLBLL_L_X2Y148_SLICE_X1Y148_AQ;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_C2 = 1'b1;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_C3 = CLBLL_L_X4Y146_SLICE_X5Y146_DO6;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_C4 = 1'b1;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_C5 = CLBLL_L_X4Y148_SLICE_X5Y148_DO6;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X2Y134_SLICE_X0Y134_B1 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X0Y134_C1 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X0Y134_C2 = 1'b1;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y134_SLICE_X0Y134_B5 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X0Y134_C5 = 1'b1;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_D1 = CLBLM_R_X3Y146_SLICE_X3Y146_BQ;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_D2 = CLBLL_L_X4Y145_SLICE_X4Y145_CQ;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_D3 = CLBLM_R_X7Y145_SLICE_X8Y145_AQ;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_D4 = CLBLM_R_X5Y145_SLICE_X7Y145_AQ;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_D5 = CLBLM_R_X7Y147_SLICE_X8Y147_AQ;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_D6 = CLBLM_L_X10Y147_SLICE_X12Y147_AQ;
  assign CLBLL_L_X2Y134_SLICE_X0Y134_C4 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X0Y134_C6 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X0Y134_D1 = 1'b1;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X2Y134_SLICE_X0Y134_D2 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X0Y134_D3 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X0Y134_D4 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X0Y134_D5 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X0Y134_D6 = 1'b1;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_A1 = CLBLM_L_X10Y147_SLICE_X13Y147_CO6;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_A3 = CLBLM_L_X10Y152_SLICE_X13Y152_AQ;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_A4 = CLBLM_L_X8Y151_SLICE_X11Y151_AQ;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_A5 = CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_A6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_B2 = CLBLM_L_X10Y152_SLICE_X13Y152_BQ;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_B3 = CLBLM_L_X10Y152_SLICE_X13Y152_AQ;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_B4 = CLBLM_R_X11Y154_SLICE_X15Y154_CO6;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_B5 = CLBLM_R_X11Y152_SLICE_X14Y152_AQ;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_B6 = CLBLM_R_X11Y153_SLICE_X14Y153_BO5;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_C1 = CLBLM_L_X10Y145_SLICE_X12Y145_AQ;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_C2 = CLBLM_L_X10Y152_SLICE_X13Y152_AQ;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_C3 = CLBLM_L_X10Y153_SLICE_X13Y153_DQ;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_C4 = CLBLM_L_X8Y146_SLICE_X10Y146_BQ;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_C5 = CLBLM_R_X7Y144_SLICE_X8Y144_AQ;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_A1 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_A2 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_A3 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_A4 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_A5 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_A6 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X1Y134_A1 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X1Y134_A2 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_B4 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_B5 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X1Y134_A3 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_B1 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_B2 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_B3 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_B6 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X1Y134_B1 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_C5 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_C6 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X1Y134_B2 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_C1 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_C2 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_C3 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_C4 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X1Y134_C1 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X1Y134_C2 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X1Y134_C3 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X1Y134_C4 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X1Y134_C5 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X1Y134_C6 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_D5 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_D1 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_D2 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_D3 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_D6 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_D4 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X1Y134_D1 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X1Y134_D2 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X1Y134_D3 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X1Y134_D4 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X1Y134_D5 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X1Y134_D6 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_A2 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_A3 = CLBLM_R_X3Y142_SLICE_X2Y142_BQ;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_A4 = RIOB33_X105Y125_IOB_X1Y126_I;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_A5 = CLBLM_R_X11Y152_SLICE_X15Y152_AQ;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_A6 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_B1 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_B2 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_B3 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_B4 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_B5 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_B6 = 1'b1;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_D1 = CLBLM_L_X10Y153_SLICE_X12Y153_AQ;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_D2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_C1 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_C2 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_C3 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_C4 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_C5 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_C6 = 1'b1;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_D4 = CLBLM_R_X11Y144_SLICE_X14Y144_BQ;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_D5 = CLBLM_R_X7Y154_SLICE_X9Y154_BQ;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_C6 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_D1 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_D2 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_D3 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_D4 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_D5 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_D6 = 1'b1;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign RIOI3_X105Y141_ILOGIC_X1Y141_D = RIOB33_X105Y141_IOB_X1Y141_I;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_D1 = 1'b1;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_A1 = 1'b1;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_A3 = CLBLM_R_X11Y146_SLICE_X15Y146_AQ;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_A4 = CLBLM_R_X11Y148_SLICE_X15Y148_AQ;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_D2 = CLBLM_R_X11Y153_SLICE_X14Y153_BO5;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_A5 = CLBLM_R_X7Y142_SLICE_X8Y142_DO6;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_A6 = CLBLM_R_X7Y142_SLICE_X8Y142_CQ;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_D3 = 1'b1;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_B1 = 1'b1;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_B2 = CLBLL_L_X4Y146_SLICE_X5Y146_AQ;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_B3 = CLBLM_R_X5Y142_SLICE_X7Y142_AQ;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_B4 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_D4 = 1'b1;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_B5 = CLBLM_R_X11Y145_SLICE_X15Y145_CO6;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_D5 = 1'b1;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_C2 = CLBLM_R_X11Y146_SLICE_X15Y146_CQ;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_C3 = CLBLM_R_X11Y147_SLICE_X15Y147_DQ;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_D6 = CLBLM_L_X10Y154_SLICE_X13Y154_BQ;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_C5 = CLBLM_R_X11Y146_SLICE_X14Y146_DQ;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_C6 = CLBLM_L_X8Y146_SLICE_X10Y146_CQ;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_D1 = CLBLM_R_X5Y142_SLICE_X7Y142_AQ;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_D2 = CLBLM_L_X12Y148_SLICE_X16Y148_BQ;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_D3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_D4 = CLBLM_L_X10Y145_SLICE_X13Y145_DO6;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_A2 = CLBLM_L_X8Y148_SLICE_X10Y148_A5Q;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_A3 = CLBLL_L_X4Y149_SLICE_X4Y149_AQ;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_A4 = CLBLM_R_X11Y150_SLICE_X14Y150_AO6;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_A5 = CLBLM_R_X5Y144_SLICE_X7Y144_BQ;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_A6 = CLBLM_R_X3Y146_SLICE_X3Y146_BQ;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_D5 = 1'b1;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_D6 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_A1 = CLBLM_R_X11Y146_SLICE_X14Y146_CQ;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_B1 = CLBLM_R_X3Y145_SLICE_X3Y145_AQ;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_B2 = CLBLL_L_X4Y149_SLICE_X4Y149_BQ;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_B4 = 1'b1;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_B5 = CLBLM_R_X7Y150_SLICE_X8Y150_CQ;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_B6 = CLBLM_L_X8Y152_SLICE_X11Y152_BO6;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_A2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_A3 = CLBLM_R_X11Y146_SLICE_X14Y146_AQ;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_C1 = CLBLM_R_X5Y152_SLICE_X7Y152_DO5;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_C2 = CLBLL_L_X4Y149_SLICE_X4Y149_CQ;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_C3 = 1'b1;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_C5 = CLBLM_R_X5Y151_SLICE_X6Y151_CQ;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_C6 = CLBLL_L_X4Y149_SLICE_X5Y149_A5Q;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_A1 = CLBLM_L_X8Y145_SLICE_X10Y145_DO6;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_B1 = 1'b1;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_B3 = CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_B4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_B5 = CLBLM_R_X11Y146_SLICE_X14Y146_BQ;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_A3 = CLBLM_L_X10Y152_SLICE_X12Y152_AQ;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_D2 = CLBLM_R_X3Y148_SLICE_X3Y148_B5Q;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_D3 = CLBLL_L_X4Y149_SLICE_X4Y149_DQ;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_D4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_D5 = 1'b1;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_D6 = CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_A4 = CLBLM_R_X7Y152_SLICE_X8Y152_AQ;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_A5 = CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_D1 = CLBLM_R_X11Y146_SLICE_X14Y146_BQ;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_D2 = CLBLM_L_X8Y147_SLICE_X11Y147_CO6;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_A6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_D3 = CLBLM_L_X10Y147_SLICE_X13Y147_AQ;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_D4 = CLBLM_R_X11Y146_SLICE_X15Y146_CQ;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_D6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign LIOI3_SING_X0Y100_OLOGIC_X0Y100_D1 = CLBLL_L_X2Y138_SLICE_X0Y138_AO5;
  assign LIOI3_SING_X0Y100_OLOGIC_X0Y100_T1 = 1'b1;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_A1 = CLBLL_L_X4Y149_SLICE_X5Y149_BO5;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_A2 = CLBLM_R_X3Y150_SLICE_X2Y150_BO6;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_A3 = CLBLL_L_X4Y149_SLICE_X5Y149_AQ;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_A4 = CLBLL_L_X4Y147_SLICE_X5Y147_B5Q;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_A6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_AX = CLBLL_L_X4Y149_SLICE_X5Y149_BO6;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_B1 = CLBLM_L_X10Y152_SLICE_X12Y152_BQ;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_B1 = CLBLM_R_X5Y149_SLICE_X7Y149_DO6;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_B2 = CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_B4 = CLBLL_L_X4Y147_SLICE_X4Y147_CQ;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_B5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_B6 = 1'b1;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_B2 = CLBLM_L_X10Y150_SLICE_X12Y150_BQ;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_B3 = CLBLM_L_X10Y153_SLICE_X12Y153_BQ;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_C1 = 1'b1;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_C2 = CLBLL_L_X4Y149_SLICE_X5Y149_CQ;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_C3 = CLBLM_R_X5Y152_SLICE_X7Y152_DO6;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_C5 = CLBLL_L_X4Y149_SLICE_X5Y149_AQ;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_C6 = CLBLM_L_X8Y150_SLICE_X10Y150_BQ;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_B4 = CLBLM_R_X11Y154_SLICE_X15Y154_CO6;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_B5 = CLBLM_R_X11Y153_SLICE_X14Y153_BO5;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_D1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_D2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_D3 = CLBLL_L_X4Y149_SLICE_X5Y149_DQ;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_D4 = CLBLM_R_X7Y149_SLICE_X9Y149_BO6;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_D5 = CLBLM_R_X3Y149_SLICE_X3Y149_CQ;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_D6 = CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_A1 = CLBLM_R_X7Y155_SLICE_X8Y155_BO5;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_A3 = CLBLM_L_X10Y153_SLICE_X13Y153_AQ;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_A4 = CLBLM_R_X5Y155_SLICE_X7Y155_CO6;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_A5 = CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_A6 = CLBLM_L_X10Y154_SLICE_X12Y154_BQ;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_C1 = CLBLM_L_X10Y146_SLICE_X12Y146_DQ;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_B1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_C2 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_B2 = CLBLM_L_X10Y153_SLICE_X13Y153_BQ;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_B3 = CLBLL_L_X4Y151_SLICE_X5Y151_AQ;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_B4 = CLBLM_R_X11Y154_SLICE_X14Y154_BO6;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_C3 = CLBLM_L_X10Y152_SLICE_X12Y152_AQ;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_B6 = CLBLM_R_X11Y153_SLICE_X14Y153_BO6;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_C2 = CLBLM_L_X10Y153_SLICE_X13Y153_CQ;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_C4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_C5 = CLBLM_L_X10Y152_SLICE_X13Y152_DO6;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_C6 = CLBLM_R_X11Y153_SLICE_X14Y153_AO5;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_A2 = CLBLM_L_X8Y145_SLICE_X10Y145_BQ;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_A3 = CLBLM_L_X8Y143_SLICE_X11Y143_AQ;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_A4 = CLBLM_R_X5Y143_SLICE_X7Y143_CO6;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_A5 = 1'b1;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_A6 = CLBLM_L_X10Y143_SLICE_X13Y143_AQ;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_C5 = CLBLM_L_X10Y152_SLICE_X12Y152_D5Q;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_B1 = CLBLM_L_X8Y144_SLICE_X10Y144_BQ;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_B2 = CLBLM_R_X5Y143_SLICE_X6Y143_AQ;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_D1 = CLBLM_R_X7Y149_SLICE_X9Y149_CO6;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_D2 = CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_D3 = CLBLM_L_X10Y153_SLICE_X13Y153_DQ;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_B3 = CLBLM_L_X8Y144_SLICE_X11Y144_AQ;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_D6 = CLBLM_L_X10Y155_SLICE_X13Y155_BQ;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_B4 = CLBLM_L_X10Y145_SLICE_X12Y145_DQ;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_B5 = CLBLM_L_X10Y144_SLICE_X12Y144_BQ;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_B6 = CLBLM_R_X11Y143_SLICE_X14Y143_AQ;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_C1 = 1'b1;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_C2 = CLBLM_L_X8Y145_SLICE_X10Y145_BQ;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_C3 = CLBLM_R_X3Y145_SLICE_X3Y145_DQ;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_C4 = CLBLM_R_X15Y151_SLICE_X20Y151_AQ;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_C5 = CLBLM_L_X8Y143_SLICE_X11Y143_DO6;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_C6 = CLBLM_L_X8Y143_SLICE_X11Y143_AQ;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_A1 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_A2 = CLBLM_L_X10Y150_SLICE_X12Y150_C5Q;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_A4 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_A5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_D1 = CLBLM_L_X8Y148_SLICE_X10Y148_BQ;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_D2 = CLBLM_R_X11Y143_SLICE_X14Y143_AQ;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_D3 = CLBLM_R_X7Y145_SLICE_X9Y145_CQ;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_D4 = 1'b1;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_B6 = CLBLM_R_X11Y154_SLICE_X15Y154_CO6;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_D5 = 1'b1;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_D6 = CLBLM_R_X5Y143_SLICE_X6Y143_AQ;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_B2 = CLBLM_L_X10Y153_SLICE_X12Y153_BQ;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_B3 = CLBLM_R_X11Y153_SLICE_X14Y153_BO5;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_B4 = CLBLM_L_X10Y154_SLICE_X13Y154_BQ;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_A1 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_A2 = CLBLM_L_X10Y143_SLICE_X12Y143_AO6;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_C6 = CLBLM_L_X10Y153_SLICE_X13Y153_BQ;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_A3 = CLBLM_R_X5Y142_SLICE_X7Y142_AQ;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_A4 = CLBLL_L_X4Y149_SLICE_X4Y149_BQ;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_A5 = 1'b1;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_C2 = CLBLM_R_X11Y154_SLICE_X14Y154_AQ;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_C3 = CLBLM_R_X11Y154_SLICE_X15Y154_BQ;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_B1 = CLBLM_R_X5Y143_SLICE_X7Y143_CO6;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_B2 = CLBLM_L_X8Y148_SLICE_X10Y148_BQ;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_B3 = 1'b1;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_B4 = CLBLM_R_X5Y143_SLICE_X6Y143_AQ;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_B5 = CLBLM_L_X8Y143_SLICE_X10Y143_BQ;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_D1 = CLBLM_R_X11Y154_SLICE_X15Y154_AQ;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_D2 = CLBLM_R_X11Y154_SLICE_X14Y154_AQ;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_C1 = CLBLM_L_X8Y143_SLICE_X10Y143_BQ;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_C2 = CLBLM_R_X7Y143_SLICE_X9Y143_CQ;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_C3 = CLBLM_L_X8Y143_SLICE_X11Y143_BO6;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_D3 = CLBLM_L_X10Y150_SLICE_X12Y150_CQ;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_C4 = CLBLM_R_X7Y143_SLICE_X9Y143_DO6;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_C5 = 1'b1;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_C6 = CLBLM_L_X8Y145_SLICE_X10Y145_BQ;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_X105Y197_OLOGIC_X1Y197_T1 = 1'b1;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_D1 = 1'b1;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_D2 = 1'b1;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_D3 = 1'b1;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_D4 = 1'b1;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_D5 = 1'b1;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_D6 = 1'b1;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_D6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_D1 = CLBLM_R_X103Y170_SLICE_X163Y170_AO6;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_T1 = 1'b1;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_A1 = CLBLM_R_X11Y148_SLICE_X15Y148_DO6;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_A2 = CLBLM_R_X11Y147_SLICE_X15Y147_BQ;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_A3 = CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_A5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_A6 = CLBLM_L_X8Y147_SLICE_X11Y147_BO5;
  assign LIOB33_X0Y151_IOB_X0Y152_O = LIOB33_X0Y65_IOB_X0Y66_I;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_D1 = CLBLM_R_X103Y169_SLICE_X163Y169_AO6;
  assign LIOB33_X0Y143_IOB_X0Y143_O = LIOB33_X0Y55_IOB_X0Y55_I;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_B1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_B2 = CLBLM_R_X11Y147_SLICE_X15Y147_BQ;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_B3 = CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_B4 = CLBLM_R_X7Y145_SLICE_X8Y145_BQ;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_B5 = CLBLM_L_X10Y147_SLICE_X13Y147_CO6;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_D3 = CLBLM_R_X11Y147_SLICE_X14Y147_DO6;
  assign LIOB33_X0Y151_IOB_X0Y151_O = LIOB33_X0Y65_IOB_X0Y65_I;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_T1 = 1'b1;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_C2 = CLBLM_R_X11Y147_SLICE_X15Y147_CQ;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_C3 = CLBLM_R_X11Y146_SLICE_X14Y146_DQ;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_C4 = CLBLM_L_X10Y143_SLICE_X13Y143_BQ;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_C5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_C6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_D5 = CLBLM_L_X12Y150_SLICE_X16Y150_AQ;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_D6 = CLBLM_L_X12Y148_SLICE_X16Y148_CO6;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_A1 = 1'b1;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_A2 = CLBLL_L_X4Y150_SLICE_X4Y150_BQ;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_A3 = CLBLL_L_X4Y150_SLICE_X4Y150_AQ;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_A4 = CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_A5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_D1 = CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_D2 = CLBLM_R_X5Y146_SLICE_X7Y146_DO6;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_D3 = CLBLM_R_X11Y147_SLICE_X15Y147_DQ;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_B1 = CLBLM_R_X11Y150_SLICE_X14Y150_AO6;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_B3 = CLBLM_R_X11Y149_SLICE_X14Y149_BQ;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_B4 = CLBLL_L_X2Y153_SLICE_X1Y153_DO6;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_B5 = CLBLM_R_X3Y147_SLICE_X2Y147_A5Q;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_B6 = 1'b1;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_A4 = CLBLM_R_X11Y147_SLICE_X14Y147_AQ;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_A5 = CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_A6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_C1 = CLBLL_L_X4Y146_SLICE_X4Y146_AQ;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_C2 = CLBLL_L_X4Y152_SLICE_X5Y152_AO5;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_C3 = CLBLM_R_X5Y149_SLICE_X6Y149_AQ;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_C4 = CLBLL_L_X4Y152_SLICE_X5Y152_AO6;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_C5 = CLBLM_L_X8Y147_SLICE_X10Y147_BQ;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_C6 = CLBLL_L_X2Y152_SLICE_X1Y152_BO6;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_B1 = CLBLM_L_X12Y150_SLICE_X16Y150_BQ;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_B2 = CLBLM_R_X11Y147_SLICE_X14Y147_BQ;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_B3 = CLBLM_R_X11Y146_SLICE_X14Y146_AQ;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_B4 = 1'b1;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_B5 = CLBLL_L_X4Y146_SLICE_X4Y146_DO6;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_D1 = CLBLL_L_X4Y155_SLICE_X5Y155_AO6;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_D2 = CLBLL_L_X4Y152_SLICE_X4Y152_AO5;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_D3 = CLBLM_R_X5Y149_SLICE_X6Y149_BQ;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_D4 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_D5 = CLBLL_L_X4Y152_SLICE_X4Y152_AO6;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_D6 = CLBLM_L_X8Y151_SLICE_X10Y151_CQ;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_C1 = CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_C2 = 1'b1;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_C3 = CLBLM_R_X3Y147_SLICE_X2Y147_AQ;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_C4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_C5 = CLBLM_R_X11Y146_SLICE_X14Y146_AQ;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_C6 = 1'b1;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_D1 = CLBLM_R_X7Y145_SLICE_X9Y145_BQ;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_D2 = CLBLM_R_X11Y147_SLICE_X14Y147_AQ;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_D3 = 1'b1;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_D4 = 1'b1;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_D5 = CLBLM_L_X12Y147_SLICE_X16Y147_AQ;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_D6 = CLBLM_R_X7Y146_SLICE_X9Y146_BQ;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_A4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_A1 = 1'b1;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_A2 = CLBLM_R_X5Y152_SLICE_X7Y152_DO5;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_A3 = CLBLL_L_X4Y150_SLICE_X5Y150_AQ;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_A4 = CLBLM_R_X5Y147_SLICE_X6Y147_CQ;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_A5 = CLBLM_R_X7Y150_SLICE_X8Y150_AQ;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_B1 = 1'b1;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_B2 = CLBLM_R_X5Y145_SLICE_X7Y145_CQ;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_B3 = CLBLL_L_X4Y148_SLICE_X4Y148_DQ;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_B4 = CLBLM_R_X5Y152_SLICE_X7Y152_DO5;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_B5 = CLBLL_L_X4Y150_SLICE_X5Y150_BQ;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_C1 = CLBLM_R_X5Y150_SLICE_X7Y150_BQ;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_C2 = CLBLL_L_X4Y147_SLICE_X4Y147_BQ;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_C3 = 1'b1;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_C4 = CLBLM_R_X5Y152_SLICE_X6Y152_A5Q;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_C5 = CLBLM_R_X7Y149_SLICE_X8Y149_DQ;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_C6 = 1'b1;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_B1 = CLBLM_R_X11Y148_SLICE_X14Y148_BQ;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_B2 = CLBLM_R_X11Y147_SLICE_X14Y147_AQ;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_D1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_B3 = CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  assign LIOI3_SING_X0Y150_OLOGIC_X0Y150_T1 = 1'b1;
  assign RIOI3_X105Y135_ILOGIC_X1Y136_D = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_D1 = 1'b1;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_D2 = CLBLL_L_X4Y152_SLICE_X5Y152_AO5;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_D3 = CLBLL_L_X4Y149_SLICE_X5Y149_AQ;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_D4 = 1'b1;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_D5 = CLBLL_L_X2Y154_SLICE_X1Y154_AO5;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_D6 = CLBLM_R_X5Y148_SLICE_X7Y148_AQ;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_T1 = 1'b1;
  assign RIOI3_X105Y135_ILOGIC_X1Y135_D = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_B6 = CLBLM_L_X8Y148_SLICE_X11Y148_BO6;
  assign CLBLM_L_X10Y154_SLICE_X13Y154_A1 = CLBLM_L_X10Y154_SLICE_X13Y154_AQ;
  assign CLBLM_L_X10Y154_SLICE_X13Y154_A2 = CLBLM_R_X5Y153_SLICE_X6Y153_BQ;
  assign CLBLM_L_X10Y154_SLICE_X13Y154_A3 = CLBLM_R_X11Y154_SLICE_X15Y154_CO5;
  assign CLBLM_L_X10Y154_SLICE_X13Y154_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y154_SLICE_X13Y154_A5 = CLBLM_R_X11Y154_SLICE_X14Y154_BO6;
  assign CLBLM_L_X10Y154_SLICE_X13Y154_A6 = CLBLM_L_X10Y154_SLICE_X13Y154_CO6;
  assign CLBLM_L_X10Y154_SLICE_X13Y154_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y154_SLICE_X13Y154_B2 = CLBLM_R_X7Y154_SLICE_X8Y154_AQ;
  assign CLBLM_L_X10Y154_SLICE_X13Y154_B3 = CLBLM_R_X11Y153_SLICE_X14Y153_BO5;
  assign CLBLM_L_X10Y154_SLICE_X13Y154_B4 = CLBLM_R_X11Y154_SLICE_X15Y154_CO6;
  assign CLBLM_L_X10Y154_SLICE_X13Y154_B5 = CLBLM_L_X10Y151_SLICE_X13Y151_CQ;
  assign CLBLM_L_X10Y154_SLICE_X13Y154_B6 = CLBLM_L_X10Y154_SLICE_X13Y154_BQ;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_D1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_D2 = CLBLM_L_X8Y149_SLICE_X10Y149_AO5;
  assign LIOI3_X0Y103_OLOGIC_X0Y103_T1 = 1'b1;
  assign CLBLM_L_X10Y154_SLICE_X13Y154_C1 = CLBLM_R_X11Y154_SLICE_X14Y154_AQ;
  assign CLBLM_L_X10Y154_SLICE_X13Y154_C2 = CLBLM_L_X10Y153_SLICE_X13Y153_BQ;
  assign CLBLM_L_X10Y154_SLICE_X13Y154_C3 = CLBLM_R_X11Y154_SLICE_X15Y154_AQ;
  assign CLBLM_L_X10Y154_SLICE_X13Y154_C4 = CLBLM_L_X10Y153_SLICE_X13Y153_CQ;
  assign CLBLM_L_X10Y154_SLICE_X13Y154_C5 = CLBLM_R_X11Y154_SLICE_X15Y154_BQ;
  assign CLBLM_L_X10Y154_SLICE_X13Y154_C6 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_A2 = 1'b1;
  assign CLBLM_L_X10Y154_SLICE_X13Y154_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_A3 = CLBLM_L_X10Y145_SLICE_X12Y145_DQ;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_A4 = CLBLM_R_X7Y142_SLICE_X8Y142_DO6;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_A5 = CLBLM_L_X8Y152_SLICE_X10Y152_DQ;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_B2 = CLBLM_L_X10Y143_SLICE_X12Y143_CO6;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_B3 = CLBLM_R_X5Y143_SLICE_X7Y143_AQ;
  assign CLBLM_L_X10Y154_SLICE_X13Y154_D1 = 1'b1;
  assign CLBLM_L_X10Y154_SLICE_X13Y154_D2 = 1'b1;
  assign CLBLM_L_X10Y154_SLICE_X13Y154_D3 = 1'b1;
  assign CLBLM_L_X10Y154_SLICE_X13Y154_D4 = CLBLM_L_X10Y150_SLICE_X12Y150_B5Q;
  assign CLBLM_L_X10Y154_SLICE_X13Y154_D5 = CLBLM_L_X10Y154_SLICE_X13Y154_AQ;
  assign CLBLM_L_X10Y154_SLICE_X13Y154_D6 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_B6 = CLBLM_L_X10Y146_SLICE_X12Y146_CQ;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_C1 = CLBLM_R_X11Y144_SLICE_X14Y144_AQ;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_C2 = CLBLM_L_X10Y142_SLICE_X13Y142_AQ;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_C3 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_C4 = CLBLM_L_X8Y147_SLICE_X10Y147_DQ;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_C5 = CLBLM_R_X7Y144_SLICE_X9Y144_CQ;
  assign CLBLM_L_X10Y154_SLICE_X12Y154_A2 = CLBLM_R_X5Y155_SLICE_X7Y155_CO6;
  assign CLBLM_L_X10Y154_SLICE_X12Y154_A3 = CLBLM_L_X10Y154_SLICE_X12Y154_AQ;
  assign CLBLM_L_X10Y154_SLICE_X12Y154_A4 = CLBLM_L_X10Y154_SLICE_X12Y154_CQ;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_C6 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y154_SLICE_X12Y154_A1 = CLBLM_R_X7Y155_SLICE_X8Y155_BO5;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_D1 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_D2 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_D3 = CLBLM_L_X10Y144_SLICE_X12Y144_DO6;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_D4 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_D5 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_D6 = CLBLM_R_X5Y143_SLICE_X7Y143_CO6;
  assign CLBLM_L_X10Y154_SLICE_X12Y154_B4 = CLBLM_R_X5Y155_SLICE_X7Y155_CO6;
  assign CLBLM_L_X10Y154_SLICE_X12Y154_B5 = CLBLM_R_X7Y145_SLICE_X8Y145_C5Q;
  assign CLBLM_L_X10Y154_SLICE_X12Y154_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y154_SLICE_X12Y154_B1 = CLBLM_R_X7Y155_SLICE_X8Y155_BO5;
  assign CLBLM_L_X10Y154_SLICE_X12Y154_B2 = CLBLM_L_X10Y154_SLICE_X12Y154_BQ;
  assign CLBLM_L_X10Y154_SLICE_X12Y154_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y154_SLICE_X12Y154_C2 = CLBLM_L_X10Y154_SLICE_X12Y154_CQ;
  assign CLBLM_L_X10Y154_SLICE_X12Y154_C3 = CLBLM_L_X8Y145_SLICE_X11Y145_CQ;
  assign CLBLM_L_X10Y154_SLICE_X12Y154_C4 = CLBLM_R_X5Y155_SLICE_X7Y155_CO6;
  assign CLBLM_L_X10Y154_SLICE_X12Y154_C5 = CLBLM_R_X7Y155_SLICE_X8Y155_BO5;
  assign CLBLM_L_X10Y154_SLICE_X12Y154_C6 = CLBLM_R_X7Y154_SLICE_X8Y154_AQ;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_A6 = CLBLM_L_X8Y144_SLICE_X11Y144_AQ;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_A1 = CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y154_SLICE_X12Y154_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_A4 = CLBLM_R_X7Y144_SLICE_X9Y144_AQ;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_B1 = CLBLM_R_X7Y145_SLICE_X9Y145_AQ;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_B2 = CLBLM_L_X8Y144_SLICE_X10Y144_BQ;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y154_SLICE_X12Y154_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y154_SLICE_X12Y154_D2 = CLBLM_L_X8Y153_SLICE_X10Y153_DO6;
  assign CLBLM_L_X10Y154_SLICE_X12Y154_D3 = CLBLM_L_X10Y154_SLICE_X12Y154_DQ;
  assign CLBLM_L_X10Y154_SLICE_X12Y154_D4 = CLBLM_L_X8Y153_SLICE_X10Y153_CO5;
  assign CLBLM_L_X10Y154_SLICE_X12Y154_D5 = CLBLM_L_X10Y155_SLICE_X12Y155_DO6;
  assign CLBLM_L_X10Y154_SLICE_X12Y154_D6 = CLBLM_L_X10Y148_SLICE_X12Y148_CQ;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_C1 = CLBLM_L_X8Y150_SLICE_X11Y150_BQ;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_C2 = CLBLM_L_X8Y144_SLICE_X10Y144_CQ;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_C4 = CLBLM_R_X7Y143_SLICE_X9Y143_CQ;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_B1 = CLBLM_L_X10Y145_SLICE_X13Y145_A5Q;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_C5 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_C6 = CLBLM_R_X5Y143_SLICE_X7Y143_CO6;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_D1 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_D2 = CLBLM_L_X8Y144_SLICE_X10Y144_CQ;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_D3 = CLBLM_L_X10Y146_SLICE_X12Y146_CQ;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_D4 = CLBLM_L_X8Y143_SLICE_X10Y143_CO6;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_D5 = CLBLM_L_X8Y145_SLICE_X11Y145_CQ;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_D6 = CLBLL_L_X4Y143_SLICE_X4Y143_CO6;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_B4 = CLBLM_L_X8Y144_SLICE_X10Y144_DO6;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_B5 = CLBLM_L_X8Y143_SLICE_X11Y143_CO6;
  assign LIOB33_X0Y145_IOB_X0Y146_O = LIOB33_X0Y59_IOB_X0Y59_I;
  assign LIOB33_X0Y145_IOB_X0Y145_O = LIOB33_X0Y57_IOB_X0Y58_I;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_C4 = 1'b1;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_C5 = CLBLM_R_X3Y149_SLICE_X3Y149_B5Q;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_B1 = CLBLM_L_X8Y150_SLICE_X10Y150_CQ;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_C6 = CLBLM_R_X3Y144_SLICE_X2Y144_CO6;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_B2 = CLBLM_R_X7Y150_SLICE_X8Y150_BQ;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_B3 = CLBLM_R_X7Y149_SLICE_X8Y149_CQ;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_A1 = CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_A3 = CLBLM_R_X11Y148_SLICE_X15Y148_AQ;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_A4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_A5 = CLBLM_R_X11Y151_SLICE_X14Y151_AQ;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_A6 = CLBLM_L_X10Y148_SLICE_X13Y148_DO6;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_AX = CLBLM_L_X12Y150_SLICE_X16Y150_DO6;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_B6 = CLBLM_L_X8Y152_SLICE_X11Y152_BO6;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_B1 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_B2 = CLBLM_L_X10Y146_SLICE_X12Y146_D5Q;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_B4 = CLBLM_R_X11Y146_SLICE_X15Y146_BQ;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_B5 = CLBLM_L_X12Y149_SLICE_X17Y149_AQ;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_B6 = 1'b1;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_C1 = CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_C2 = CLBLM_R_X11Y148_SLICE_X15Y148_CQ;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_C3 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_C4 = CLBLM_R_X7Y149_SLICE_X9Y149_CO6;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_C6 = CLBLM_R_X11Y145_SLICE_X15Y145_BQ;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_A1 = 1'b1;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_A2 = CLBLL_L_X4Y151_SLICE_X5Y151_B5Q;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_A4 = 1'b1;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_A5 = CLBLM_L_X8Y149_SLICE_X11Y149_AQ;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_A6 = CLBLM_R_X3Y150_SLICE_X3Y150_A5Q;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_D1 = CLBLM_L_X10Y151_SLICE_X12Y151_AQ;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_AX = CLBLM_R_X7Y151_SLICE_X9Y151_DO6;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_D2 = CLBLM_R_X11Y147_SLICE_X15Y147_AQ;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_B1 = CLBLL_L_X2Y151_SLICE_X1Y151_DO6;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_B2 = CLBLL_L_X4Y151_SLICE_X5Y151_DO6;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_B3 = CLBLL_L_X2Y149_SLICE_X0Y149_AO6;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_B4 = CLBLL_L_X2Y154_SLICE_X1Y154_AO5;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_B5 = CLBLM_R_X5Y146_SLICE_X6Y146_AQ;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_B6 = CLBLL_L_X4Y151_SLICE_X4Y151_CO6;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_D2 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_D4 = 1'b1;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_C1 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_C2 = CLBLM_R_X5Y152_SLICE_X6Y152_CQ;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_C3 = CLBLL_L_X2Y155_SLICE_X1Y155_DO6;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_C4 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_C5 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_C6 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_A2 = CLBLM_L_X10Y146_SLICE_X12Y146_D5Q;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_A3 = CLBLM_R_X11Y148_SLICE_X14Y148_AQ;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_C6 = 1'b1;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_D5 = CLBLM_R_X11Y146_SLICE_X14Y146_DQ;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_A5 = CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_A6 = CLBLM_L_X10Y148_SLICE_X13Y148_DO6;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_D6 = 1'b1;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_D1 = 1'b1;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_D2 = CLBLL_L_X2Y155_SLICE_X1Y155_DO6;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_D3 = CLBLM_R_X5Y151_SLICE_X6Y151_AQ;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_D4 = CLBLM_R_X5Y151_SLICE_X7Y151_BQ;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_D5 = CLBLL_L_X2Y154_SLICE_X1Y154_BO5;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_D6 = CLBLL_L_X4Y155_SLICE_X4Y155_BO6;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_B4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_C2 = CLBLM_R_X11Y148_SLICE_X14Y148_CQ;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_C4 = CLBLM_R_X11Y148_SLICE_X14Y148_BQ;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_C5 = 1'b1;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_C6 = 1'b1;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_D2 = CLBLM_L_X10Y146_SLICE_X13Y146_AQ;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_D3 = CLBLM_R_X11Y148_SLICE_X14Y148_DQ;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_D4 = CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_D5 = CLBLM_R_X5Y148_SLICE_X7Y148_DO6;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_D6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_A1 = CLBLM_R_X11Y150_SLICE_X14Y150_BO6;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_A2 = CLBLM_L_X8Y148_SLICE_X10Y148_A5Q;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_A3 = CLBLL_L_X4Y151_SLICE_X5Y151_AQ;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_A5 = CLBLM_R_X7Y150_SLICE_X8Y150_BQ;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_A6 = CLBLM_R_X7Y147_SLICE_X8Y147_AQ;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_B1 = CLBLM_R_X3Y153_SLICE_X2Y153_DO6;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_B2 = CLBLM_R_X3Y154_SLICE_X2Y154_BO6;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_B3 = CLBLM_L_X8Y144_SLICE_X10Y144_AQ;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_B5 = CLBLL_L_X4Y148_SLICE_X5Y148_CQ;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_B6 = 1'b1;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_C1 = CLBLL_L_X4Y152_SLICE_X5Y152_AO6;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_C2 = CLBLM_R_X7Y151_SLICE_X9Y151_BQ;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_C3 = CLBLM_R_X5Y151_SLICE_X7Y151_AQ;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_C4 = CLBLL_L_X2Y152_SLICE_X1Y152_BO6;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_C5 = CLBLL_L_X2Y154_SLICE_X1Y154_AO5;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_C6 = CLBLM_R_X7Y150_SLICE_X8Y150_BQ;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign RIOI3_X105Y171_OLOGIC_X1Y171_D1 = CLBLM_R_X11Y157_SLICE_X14Y157_AO5;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_D1 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_D2 = CLBLM_L_X8Y152_SLICE_X10Y152_BQ;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_D3 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_D4 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_D5 = CLBLL_L_X2Y155_SLICE_X1Y155_DO6;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_D6 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_A3 = CLBLM_L_X8Y144_SLICE_X10Y144_AQ;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_A5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_A6 = CLBLM_L_X10Y144_SLICE_X12Y144_BQ;
  assign CLBLM_L_X10Y155_SLICE_X13Y155_A1 = CLBLM_L_X10Y155_SLICE_X13Y155_CQ;
  assign CLBLM_L_X10Y155_SLICE_X13Y155_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y155_SLICE_X13Y155_A3 = CLBLM_L_X10Y155_SLICE_X13Y155_AQ;
  assign CLBLM_L_X10Y155_SLICE_X13Y155_A4 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_L_X10Y155_SLICE_X13Y155_A5 = 1'b1;
  assign CLBLM_L_X10Y155_SLICE_X13Y155_A6 = CLBLM_R_X5Y142_SLICE_X7Y142_AQ;
  assign CLBLM_L_X10Y155_SLICE_X13Y155_B1 = 1'b1;
  assign CLBLM_L_X10Y155_SLICE_X13Y155_B2 = CLBLM_L_X10Y155_SLICE_X12Y155_BO6;
  assign CLBLM_L_X10Y155_SLICE_X13Y155_B3 = CLBLM_L_X10Y154_SLICE_X13Y154_AQ;
  assign CLBLM_L_X10Y155_SLICE_X13Y155_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y155_SLICE_X13Y155_B5 = CLBLM_L_X8Y153_SLICE_X10Y153_CO5;
  assign CLBLM_L_X10Y155_SLICE_X13Y155_B6 = CLBLM_L_X8Y153_SLICE_X10Y153_DO6;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_B6 = CLBLM_L_X8Y152_SLICE_X10Y152_BQ;
  assign LIOI3_SING_X0Y150_OLOGIC_X0Y150_D1 = LIOB33_X0Y63_IOB_X0Y63_I;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_A1 = CLBLM_L_X8Y145_SLICE_X11Y145_B5Q;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_A2 = CLBLM_L_X10Y146_SLICE_X12Y146_AQ;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y155_SLICE_X13Y155_C4 = CLBLM_L_X8Y153_SLICE_X10Y153_DO6;
  assign CLBLM_L_X10Y155_SLICE_X13Y155_C5 = CLBLM_L_X10Y155_SLICE_X13Y155_CQ;
  assign CLBLM_L_X10Y155_SLICE_X13Y155_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_A5 = CLBLM_L_X8Y145_SLICE_X11Y145_A5Q;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_A6 = 1'b1;
  assign CLBLM_L_X10Y155_SLICE_X13Y155_C1 = CLBLM_L_X8Y153_SLICE_X10Y153_CO5;
  assign CLBLM_L_X10Y155_SLICE_X13Y155_C2 = CLBLM_L_X10Y155_SLICE_X12Y155_CO6;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_B1 = CLBLM_R_X11Y146_SLICE_X14Y146_AQ;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_B2 = CLBLM_R_X7Y144_SLICE_X8Y144_BQ;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_B3 = CLBLM_L_X10Y150_SLICE_X12Y150_A5Q;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y155_SLICE_X13Y155_D2 = CLBLM_L_X10Y154_SLICE_X12Y154_DQ;
  assign CLBLM_L_X10Y155_SLICE_X13Y155_D3 = CLBLM_L_X8Y153_SLICE_X11Y153_BQ;
  assign CLBLM_L_X10Y155_SLICE_X13Y155_D4 = CLBLM_L_X8Y155_SLICE_X10Y155_AQ;
  assign CLBLM_L_X10Y155_SLICE_X13Y155_D5 = 1'b1;
  assign CLBLM_L_X10Y155_SLICE_X13Y155_D6 = CLBLM_L_X8Y155_SLICE_X11Y155_CO6;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_B5 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_B6 = 1'b1;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_C1 = CLBLM_L_X8Y144_SLICE_X10Y144_CQ;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_C2 = CLBLM_L_X8Y145_SLICE_X11Y145_CQ;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_C3 = CLBLM_L_X8Y144_SLICE_X11Y144_AQ;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_C4 = CLBLM_R_X7Y142_SLICE_X8Y142_DO6;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_C5 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_B4 = CLBLM_L_X10Y144_SLICE_X12Y144_BQ;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y155_SLICE_X12Y155_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y155_SLICE_X12Y155_A1 = CLBLM_L_X10Y150_SLICE_X12Y150_B5Q;
  assign CLBLM_L_X10Y155_SLICE_X12Y155_A2 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_B5 = 1'b1;
  assign CLBLM_L_X10Y155_SLICE_X12Y155_A3 = CLBLM_L_X8Y153_SLICE_X10Y153_CO5;
  assign CLBLM_L_X10Y155_SLICE_X12Y155_A4 = CLBLM_L_X10Y156_SLICE_X12Y156_BO6;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_D1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_B6 = CLBLM_R_X7Y142_SLICE_X8Y142_DO6;
  assign CLBLM_L_X10Y155_SLICE_X12Y155_B4 = CLBLM_L_X10Y155_SLICE_X13Y155_BQ;
  assign CLBLM_L_X10Y155_SLICE_X12Y155_B5 = CLBLM_L_X8Y155_SLICE_X10Y155_CO6;
  assign CLBLM_L_X10Y155_SLICE_X12Y155_B6 = CLBLM_L_X8Y154_SLICE_X11Y154_DO6;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_D2 = CLBLM_R_X7Y145_SLICE_X9Y145_DO6;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_D3 = CLBLM_L_X8Y145_SLICE_X11Y145_DQ;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_D4 = CLBLM_L_X10Y145_SLICE_X12Y145_DQ;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_D5 = CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_D6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y155_SLICE_X12Y155_C1 = CLBLM_L_X8Y155_SLICE_X10Y155_CO6;
  assign CLBLM_L_X10Y155_SLICE_X12Y155_C2 = CLBLM_L_X8Y153_SLICE_X10Y153_BQ;
  assign CLBLM_L_X10Y155_SLICE_X12Y155_C3 = CLBLM_L_X10Y155_SLICE_X13Y155_DO6;
  assign CLBLM_L_X10Y155_SLICE_X12Y155_C4 = CLBLM_L_X10Y156_SLICE_X12Y156_AO5;
  assign CLBLM_L_X10Y155_SLICE_X12Y155_C5 = CLBLM_L_X8Y154_SLICE_X11Y154_DO6;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_A1 = CLBLM_L_X10Y147_SLICE_X13Y147_AQ;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
endmodule
