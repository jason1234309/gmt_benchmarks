module top(
  input LIOB33_SING_X0Y100_IOB_X0Y100_IPAD,
  input LIOB33_X0Y101_IOB_X0Y101_IPAD,
  input LIOB33_X0Y101_IOB_X0Y102_IPAD,
  input LIOB33_X0Y103_IOB_X0Y103_IPAD,
  input LIOB33_X0Y103_IOB_X0Y104_IPAD,
  input LIOB33_X0Y105_IOB_X0Y105_IPAD,
  input LIOB33_X0Y105_IOB_X0Y106_IPAD,
  input LIOB33_X0Y107_IOB_X0Y107_IPAD,
  input LIOB33_X0Y107_IOB_X0Y108_IPAD,
  input LIOB33_X0Y109_IOB_X0Y109_IPAD,
  input LIOB33_X0Y109_IOB_X0Y110_IPAD,
  input LIOB33_X0Y111_IOB_X0Y111_IPAD,
  input LIOB33_X0Y111_IOB_X0Y112_IPAD,
  input LIOB33_X0Y113_IOB_X0Y113_IPAD,
  input LIOB33_X0Y113_IOB_X0Y114_IPAD,
  input LIOB33_X0Y115_IOB_X0Y115_IPAD,
  input LIOB33_X0Y115_IOB_X0Y116_IPAD,
  input LIOB33_X0Y117_IOB_X0Y117_IPAD,
  input RIOB33_SING_X105Y100_IOB_X1Y100_IPAD,
  input RIOB33_X105Y101_IOB_X1Y101_IPAD,
  input RIOB33_X105Y101_IOB_X1Y102_IPAD,
  input RIOB33_X105Y103_IOB_X1Y103_IPAD,
  input RIOB33_X105Y103_IOB_X1Y104_IPAD,
  input RIOB33_X105Y105_IOB_X1Y105_IPAD,
  input RIOB33_X105Y105_IOB_X1Y106_IPAD,
  input RIOB33_X105Y107_IOB_X1Y107_IPAD,
  input RIOB33_X105Y107_IOB_X1Y108_IPAD,
  input RIOB33_X105Y109_IOB_X1Y109_IPAD,
  input RIOB33_X105Y109_IOB_X1Y110_IPAD,
  input RIOB33_X105Y111_IOB_X1Y111_IPAD,
  input RIOB33_X105Y111_IOB_X1Y112_IPAD,
  input RIOB33_X105Y113_IOB_X1Y113_IPAD,
  output LIOB33_SING_X0Y149_IOB_X0Y149_OPAD,
  output LIOB33_X0Y117_IOB_X0Y118_OPAD,
  output LIOB33_X0Y119_IOB_X0Y119_OPAD,
  output LIOB33_X0Y119_IOB_X0Y120_OPAD,
  output LIOB33_X0Y121_IOB_X0Y121_OPAD,
  output LIOB33_X0Y121_IOB_X0Y122_OPAD,
  output LIOB33_X0Y123_IOB_X0Y123_OPAD,
  output LIOB33_X0Y123_IOB_X0Y124_OPAD,
  output LIOB33_X0Y125_IOB_X0Y125_OPAD,
  output LIOB33_X0Y125_IOB_X0Y126_OPAD,
  output LIOB33_X0Y127_IOB_X0Y127_OPAD,
  output LIOB33_X0Y127_IOB_X0Y128_OPAD,
  output LIOB33_X0Y129_IOB_X0Y129_OPAD,
  output LIOB33_X0Y129_IOB_X0Y130_OPAD,
  output LIOB33_X0Y131_IOB_X0Y131_OPAD,
  output LIOB33_X0Y131_IOB_X0Y132_OPAD,
  output LIOB33_X0Y133_IOB_X0Y133_OPAD,
  output LIOB33_X0Y133_IOB_X0Y134_OPAD,
  output LIOB33_X0Y135_IOB_X0Y135_OPAD,
  output LIOB33_X0Y135_IOB_X0Y136_OPAD,
  output LIOB33_X0Y137_IOB_X0Y137_OPAD,
  output LIOB33_X0Y137_IOB_X0Y138_OPAD,
  output LIOB33_X0Y139_IOB_X0Y139_OPAD,
  output LIOB33_X0Y139_IOB_X0Y140_OPAD,
  output LIOB33_X0Y141_IOB_X0Y141_OPAD,
  output LIOB33_X0Y141_IOB_X0Y142_OPAD,
  output LIOB33_X0Y143_IOB_X0Y143_OPAD,
  output LIOB33_X0Y145_IOB_X0Y145_OPAD,
  output LIOB33_X0Y145_IOB_X0Y146_OPAD,
  output LIOB33_X0Y147_IOB_X0Y147_OPAD,
  output LIOB33_X0Y147_IOB_X0Y148_OPAD
  );
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_A;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_A1;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_A2;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_A3;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_A4;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_A5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_A6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_AMUX;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_AO5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_AO6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_A_CY;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_A_XOR;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_B;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_B1;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_B2;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_B3;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_B4;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_B5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_B6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_BMUX;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_BO5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_BO6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_B_CY;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_B_XOR;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_C;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_C1;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_C2;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_C3;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_C4;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_C5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_C6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_CO5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_CO6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_C_CY;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_C_XOR;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_D;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_D1;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_D2;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_D3;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_D4;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_D5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_D6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_DO5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_DO6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_D_CY;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_D_XOR;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_A;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_A1;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_A2;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_A3;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_A4;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_A5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_A6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_AMUX;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_AO5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_AO6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_A_CY;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_A_XOR;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_B;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_B1;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_B2;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_B3;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_B4;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_B5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_B6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_BO5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_BO6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_B_CY;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_B_XOR;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_C;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_C1;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_C2;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_C3;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_C4;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_C5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_C6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_CO5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_CO6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_C_CY;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_C_XOR;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_D;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_D1;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_D2;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_D3;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_D4;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_D5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_D6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_DO5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_DO6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_D_CY;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_D_XOR;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_A;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_A1;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_A2;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_A3;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_A4;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_A5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_A6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_AMUX;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_AO5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_AO6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_A_CY;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_A_XOR;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_B;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_B1;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_B2;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_B3;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_B4;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_B5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_B6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_BO5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_BO6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_B_CY;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_B_XOR;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_C;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_C1;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_C2;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_C3;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_C4;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_C5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_C6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_CO5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_CO6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_C_CY;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_C_XOR;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_D;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_D1;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_D2;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_D3;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_D4;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_D5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_D6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_DO5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_DO6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_D_CY;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_D_XOR;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_A;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_A1;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_A2;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_A3;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_A4;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_A5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_A6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_AMUX;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_AO5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_AO6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_A_CY;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_A_XOR;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_B;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_B1;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_B2;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_B3;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_B4;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_B5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_B6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_BO5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_BO6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_B_CY;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_B_XOR;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_C;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_C1;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_C2;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_C3;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_C4;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_C5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_C6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_CMUX;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_CO5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_CO6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_C_CY;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_C_XOR;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_D;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_D1;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_D2;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_D3;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_D4;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_D5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_D6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_DO5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_DO6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_D_CY;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_D_XOR;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_A;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_A1;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_A2;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_A3;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_A4;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_A5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_A6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_AMUX;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_AO5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_AO6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_A_CY;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_A_XOR;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_B;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_B1;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_B2;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_B3;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_B4;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_B5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_B6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_BO5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_BO6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_B_CY;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_B_XOR;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_C;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_C1;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_C2;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_C3;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_C4;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_C5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_C6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_CO5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_CO6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_C_CY;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_C_XOR;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_D;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_D1;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_D2;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_D3;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_D4;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_D5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_D6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_DO5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_DO6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_D_CY;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_D_XOR;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_A;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_A1;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_A2;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_A3;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_A4;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_A5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_A6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_AMUX;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_AO5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_AO6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_A_CY;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_A_XOR;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_B;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_B1;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_B2;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_B3;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_B4;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_B5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_B6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_BMUX;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_BO5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_BO6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_B_CY;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_B_XOR;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_C;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_C1;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_C2;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_C3;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_C4;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_C5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_C6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_CMUX;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_CO5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_CO6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_C_CY;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_C_XOR;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_D;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_D1;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_D2;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_D3;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_D4;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_D5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_D6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_DO5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_DO6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_D_CY;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_D_XOR;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A1;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A2;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A3;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A4;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_AMUX;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_AO5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_AO6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A_CY;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A_XOR;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B1;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B2;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B3;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B4;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_BMUX;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_BO5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_BO6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B_CY;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B_XOR;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C1;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C2;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C3;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C4;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_CMUX;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_CO5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_CO6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C_CY;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C_XOR;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D1;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D2;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D3;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D4;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_DO5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_DO6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D_CY;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D_XOR;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A1;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A2;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A3;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A4;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_AO5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_AO6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A_CY;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A_XOR;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B1;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B2;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B3;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B4;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_BO5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_BO6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B_CY;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B_XOR;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C1;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C2;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C3;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C4;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_CO5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_CO6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C_CY;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C_XOR;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D1;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D2;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D3;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D4;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_DO5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_DO6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D_CY;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D_XOR;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A1;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A2;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A3;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A4;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_AO5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_AO6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A_CY;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A_XOR;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B1;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B2;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B3;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B4;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_BO5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_BO6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B_CY;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B_XOR;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C1;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C2;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C3;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C4;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_CO5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_CO6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C_CY;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C_XOR;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D1;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D2;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D3;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D4;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_DO5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_DO6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D_CY;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D_XOR;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A1;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A2;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A3;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A4;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_AO5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_AO6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A_CY;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A_XOR;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B1;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B2;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B3;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B4;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_BO5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_BO6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B_CY;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B_XOR;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C1;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C2;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C3;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C4;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_CO5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_CO6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C_CY;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C_XOR;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D1;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D2;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D3;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D4;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_DO5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_DO6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D_CY;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D_XOR;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_A;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_A1;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_A2;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_A3;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_A4;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_A5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_A6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_AO5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_AO6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_A_CY;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_A_XOR;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_B;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_B1;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_B2;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_B3;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_B4;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_B5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_B6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_BO5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_BO6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_B_CY;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_B_XOR;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_C;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_C1;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_C2;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_C3;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_C4;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_C5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_C6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_CO5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_CO6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_C_CY;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_C_XOR;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_D;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_D1;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_D2;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_D3;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_D4;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_D5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_D6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_DO5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_DO6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_D_CY;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_D_XOR;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_A;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_A1;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_A2;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_A3;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_A4;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_A5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_A6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_AO5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_AO6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_A_CY;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_A_XOR;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_B;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_B1;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_B2;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_B3;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_B4;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_B5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_B6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_BO5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_BO6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_B_CY;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_B_XOR;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_C;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_C1;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_C2;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_C3;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_C4;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_C5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_C6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_CO5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_CO6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_C_CY;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_C_XOR;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_D;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_D1;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_D2;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_D3;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_D4;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_D5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_D6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_DO5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_DO6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_D_CY;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_D_XOR;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_A;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_A1;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_A2;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_A3;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_A4;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_A5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_A6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_AMUX;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_AO5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_AO6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_A_CY;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_A_XOR;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_B;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_B1;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_B2;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_B3;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_B4;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_B5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_B6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_BO5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_BO6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_B_CY;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_B_XOR;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_C;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_C1;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_C2;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_C3;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_C4;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_C5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_C6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_CO5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_CO6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_C_CY;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_C_XOR;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_D;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_D1;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_D2;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_D3;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_D4;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_D5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_D6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_DO5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_DO6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_D_CY;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_D_XOR;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_A;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_A1;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_A2;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_A3;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_A4;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_A5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_A6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_AO5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_AO6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_A_CY;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_A_XOR;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_B;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_B1;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_B2;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_B3;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_B4;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_B5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_B6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_BO5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_BO6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_B_CY;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_B_XOR;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_C;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_C1;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_C2;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_C3;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_C4;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_C5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_C6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_CO5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_CO6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_C_CY;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_C_XOR;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_D;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_D1;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_D2;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_D3;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_D4;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_D5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_D6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_DO5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_DO6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_D_CY;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_D_XOR;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_A;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_A1;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_A2;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_A3;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_A4;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_A5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_A6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_AMUX;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_AO5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_AO6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_A_CY;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_A_XOR;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_B;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_B1;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_B2;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_B3;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_B4;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_B5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_B6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_BO5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_BO6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_B_CY;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_B_XOR;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_C;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_C1;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_C2;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_C3;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_C4;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_C5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_C6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_CO5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_CO6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_C_CY;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_C_XOR;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_D;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_D1;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_D2;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_D3;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_D4;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_D5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_D6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_DO5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_DO6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_D_CY;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_D_XOR;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_A;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_A1;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_A2;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_A3;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_A4;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_A5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_A6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_AO5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_AO6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_A_CY;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_A_XOR;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_B;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_B1;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_B2;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_B3;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_B4;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_B5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_B6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_BO5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_BO6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_B_CY;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_B_XOR;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_C;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_C1;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_C2;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_C3;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_C4;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_C5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_C6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_CO5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_CO6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_C_CY;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_C_XOR;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_D;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_D1;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_D2;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_D3;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_D4;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_D5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_D6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_DO5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_DO6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_D_CY;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_D_XOR;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_A;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_A1;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_A2;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_A3;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_A4;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_A5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_A6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_AMUX;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_AO5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_AO6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_A_CY;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_A_XOR;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_B;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_B1;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_B2;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_B3;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_B4;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_B5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_B6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_BO5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_BO6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_B_CY;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_B_XOR;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_C;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_C1;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_C2;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_C3;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_C4;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_C5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_C6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_CO5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_CO6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_C_CY;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_C_XOR;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_D;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_D1;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_D2;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_D3;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_D4;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_D5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_D6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_DO5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_DO6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_D_CY;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_D_XOR;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_A;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_A1;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_A2;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_A3;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_A4;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_A5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_A6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_AO5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_AO6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_A_CY;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_A_XOR;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_B;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_B1;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_B2;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_B3;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_B4;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_B5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_B6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_BO5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_BO6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_B_CY;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_B_XOR;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_C;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_C1;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_C2;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_C3;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_C4;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_C5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_C6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_CO5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_CO6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_C_CY;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_C_XOR;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_D;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_D1;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_D2;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_D3;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_D4;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_D5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_D6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_DO5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_DO6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_D_CY;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_D_XOR;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A1;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A2;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A3;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A4;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_AO5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_AO6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A_CY;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A_XOR;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B1;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B2;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B3;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B4;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_BO5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_BO6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B_CY;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B_XOR;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C1;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C2;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C3;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C4;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_CO5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_CO6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C_CY;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C_XOR;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D1;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D2;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D3;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D4;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_DO5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_DO6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D_CY;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D_XOR;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A1;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A2;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A3;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A4;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_AO5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_AO6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A_CY;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A_XOR;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B1;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B2;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B3;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B4;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_BO5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_BO6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B_CY;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B_XOR;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C1;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C2;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C3;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C4;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_CO5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_CO6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C_CY;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C_XOR;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D1;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D2;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D3;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D4;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_DO5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_DO6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D_CY;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D_XOR;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A1;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A2;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A3;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A4;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_AO5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_AO6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A_CY;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A_XOR;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B1;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B2;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B3;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B4;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_BO5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_BO6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B_CY;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B_XOR;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C1;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C2;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C3;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C4;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_CO5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_CO6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C_CY;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C_XOR;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D1;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D2;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D3;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D4;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_DO5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_DO6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D_CY;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D_XOR;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A1;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A2;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A3;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A4;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_AMUX;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_AO5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_AO6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A_CY;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A_XOR;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B1;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B2;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B3;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B4;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_BO5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_BO6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B_CY;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B_XOR;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C1;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C2;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C3;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C4;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_CO5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_CO6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C_CY;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C_XOR;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D1;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D2;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D3;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D4;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_DO5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_DO6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D_CY;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_AMUX;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_AO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_AO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_BO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_BO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_CO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_CO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_DO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_DO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_AO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_AO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_BO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_BO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_CO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_CO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_DO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_DO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D_XOR;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A1;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A2;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A3;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A4;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_AMUX;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_AO5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_AO6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A_CY;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A_XOR;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B1;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B2;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B3;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B4;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_BMUX;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_BO5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_BO6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B_CY;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B_XOR;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C1;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C2;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C3;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C4;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_CO5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_CO6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C_CY;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C_XOR;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D1;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D2;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D3;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D4;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_DO5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_DO6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D_CY;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D_XOR;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A1;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A2;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A3;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A4;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_AO5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_AO6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A_CY;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A_XOR;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B1;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B2;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B3;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B4;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_BO5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_BO6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B_CY;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B_XOR;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C1;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C2;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C3;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C4;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_CO5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_CO6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C_CY;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C_XOR;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D1;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D2;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D3;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D4;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_DO5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_DO6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D_CY;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D_XOR;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A1;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A2;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A3;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A4;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_AMUX;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_AO5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_AO6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A_CY;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A_XOR;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B1;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B2;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B3;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B4;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_BO5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_BO6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B_CY;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B_XOR;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C1;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C2;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C3;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C4;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_CO5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_CO6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C_CY;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C_XOR;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D1;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D2;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D3;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D4;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_DO5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_DO6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D_CY;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D_XOR;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A1;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A2;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A3;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A4;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_AO5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_AO6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A_CY;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A_XOR;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B1;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B2;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B3;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B4;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_BMUX;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_BO5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_BO6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B_CY;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B_XOR;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C1;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C2;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C3;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C4;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_CO5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_CO6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C_CY;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C_XOR;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D1;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D2;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D3;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D4;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_DO5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_DO6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D_CY;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_AO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_AO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_BO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_BO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_CO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_CO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_DO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_DO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_AMUX;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_AO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_AO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_BMUX;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_BO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_BO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_CO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_CO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_DO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_DO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_AMUX;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_AO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_AO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_BO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_BO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_CO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_CO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_DO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_DO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_AMUX;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_AO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_AO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_BMUX;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_BO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_BO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_CMUX;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_CO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_CO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_DO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_DO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D_XOR;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A1;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A2;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A3;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A4;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_AO5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_AO6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A_CY;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A_XOR;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B1;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B2;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B3;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B4;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_BO5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_BO6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B_CY;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B_XOR;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C1;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C2;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C3;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C4;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_CO5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_CO6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C_CY;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C_XOR;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D1;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D2;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D3;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D4;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_DO5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_DO6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D_CY;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D_XOR;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A1;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A2;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A3;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A4;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_AMUX;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_AO5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_AO6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A_CY;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A_XOR;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B1;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B2;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B3;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B4;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_BO5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_BO6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B_CY;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B_XOR;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C1;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C2;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C3;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C4;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_CO5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_CO6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C_CY;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C_XOR;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D1;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D2;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D3;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D4;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_DO5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_DO6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D_CY;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_AMUX;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_AO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_AO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_BO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_BO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_CO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_CO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_DO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_DO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_AMUX;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_AO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_AO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_BO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_BO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_CO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_CO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_DO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_DO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D_XOR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A1;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A2;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A3;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A4;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_AMUX;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_AO5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_AO6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A_CY;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A_XOR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B1;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B2;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B3;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B4;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_BO5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_BO6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B_CY;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B_XOR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C1;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C2;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C3;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C4;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_CO5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_CO6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C_CY;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C_XOR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D1;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D2;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D3;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D4;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_DO5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_DO6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D_CY;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D_XOR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A1;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A2;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A3;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A4;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_AMUX;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_AO5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_AO6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A_CY;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A_XOR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B1;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B2;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B3;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B4;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_BMUX;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_BO5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_BO6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B_CY;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B_XOR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C1;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C2;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C3;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C4;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_CMUX;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_CO5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_CO6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C_CY;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C_XOR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D1;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D2;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D3;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D4;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_DMUX;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_DO5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_DO6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D_CY;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D_XOR;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_A;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_A1;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_A2;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_A3;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_A4;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_A5;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_A6;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_AO5;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_AO6;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_A_CY;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_A_XOR;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_B;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_B1;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_B2;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_B3;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_B4;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_B5;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_B6;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_BO5;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_BO6;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_B_CY;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_B_XOR;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_C;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_C1;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_C2;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_C3;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_C4;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_C5;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_C6;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_CMUX;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_CO5;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_CO6;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_C_CY;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_C_XOR;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_D;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_D1;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_D2;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_D3;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_D4;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_D5;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_D6;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_DO5;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_DO6;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_D_CY;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_D_XOR;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_A;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_A1;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_A2;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_A3;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_A4;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_A5;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_A6;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_AMUX;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_AO5;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_AO6;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_A_CY;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_A_XOR;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_B;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_B1;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_B2;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_B3;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_B4;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_B5;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_B6;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_BO5;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_BO6;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_B_CY;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_B_XOR;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_C;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_C1;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_C2;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_C3;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_C4;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_C5;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_C6;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_CO5;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_CO6;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_C_CY;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_C_XOR;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_D;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_D1;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_D2;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_D3;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_D4;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_D5;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_D6;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_DO5;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_DO6;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_D_CY;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_D_XOR;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_A;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_A1;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_A2;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_A3;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_A4;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_A5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_A6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_AMUX;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_AO5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_AO6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_A_CY;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_A_XOR;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_B;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_B1;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_B2;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_B3;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_B4;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_B5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_B6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_BO5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_BO6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_B_CY;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_B_XOR;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_C;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_C1;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_C2;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_C3;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_C4;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_C5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_C6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_CO5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_CO6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_C_CY;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_C_XOR;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_D;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_D1;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_D2;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_D3;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_D4;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_D5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_D6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_DO5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_DO6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_D_CY;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_D_XOR;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_A;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_A1;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_A2;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_A3;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_A4;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_A5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_A6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_AMUX;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_AO5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_AO6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_A_CY;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_A_XOR;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_B;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_B1;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_B2;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_B3;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_B4;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_B5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_B6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_BO5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_BO6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_B_CY;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_B_XOR;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_C;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_C1;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_C2;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_C3;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_C4;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_C5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_C6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_CO5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_CO6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_C_CY;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_C_XOR;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_D;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_D1;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_D2;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_D3;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_D4;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_D5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_D6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_DO5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_DO6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_D_CY;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_D_XOR;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_A;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_A1;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_A2;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_A3;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_A4;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_A5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_A6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_AO5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_AO6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_A_CY;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_A_XOR;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_B;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_B1;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_B2;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_B3;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_B4;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_B5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_B6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_BO5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_BO6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_B_CY;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_B_XOR;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_C;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_C1;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_C2;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_C3;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_C4;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_C5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_C6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_CO5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_CO6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_C_CY;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_C_XOR;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_D;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_D1;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_D2;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_D3;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_D4;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_D5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_D6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_DO5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_DO6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_D_CY;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_D_XOR;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_A;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_A1;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_A2;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_A3;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_A4;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_A5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_A6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_AO5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_AO6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_A_CY;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_A_XOR;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_B;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_B1;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_B2;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_B3;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_B4;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_B5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_B6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_BMUX;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_BO5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_BO6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_B_CY;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_B_XOR;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_C;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_C1;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_C2;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_C3;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_C4;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_C5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_C6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_CMUX;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_CO5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_CO6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_C_CY;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_C_XOR;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_D;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_D1;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_D2;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_D3;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_D4;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_D5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_D6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_DO5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_DO6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_D_CY;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_D_XOR;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_A;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_A1;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_A2;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_A3;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_A4;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_A5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_A6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_AMUX;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_AO5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_AO6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_A_CY;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_A_XOR;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_B;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_B1;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_B2;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_B3;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_B4;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_B5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_B6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_BO5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_BO6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_B_CY;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_B_XOR;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_C;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_C1;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_C2;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_C3;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_C4;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_C5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_C6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_CO5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_CO6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_C_CY;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_C_XOR;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_D;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_D1;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_D2;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_D3;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_D4;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_D5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_D6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_DO5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_DO6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_D_CY;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_D_XOR;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_A;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_A1;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_A2;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_A3;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_A4;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_A5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_A6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_AMUX;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_AO5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_AO6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_A_CY;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_A_XOR;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_B;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_B1;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_B2;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_B3;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_B4;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_B5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_B6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_BO5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_BO6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_B_CY;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_B_XOR;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_C;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_C1;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_C2;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_C3;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_C4;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_C5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_C6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_CMUX;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_CO5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_CO6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_C_CY;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_C_XOR;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_D;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_D1;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_D2;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_D3;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_D4;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_D5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_D6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_DO5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_DO6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_D_CY;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_D_XOR;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_A;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_A1;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_A2;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_A3;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_A4;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_A5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_A6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_AO5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_AO6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_A_CY;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_A_XOR;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_B;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_B1;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_B2;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_B3;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_B4;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_B5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_B6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_BO5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_BO6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_B_CY;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_B_XOR;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_C;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_C1;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_C2;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_C3;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_C4;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_C5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_C6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_CO5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_CO6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_C_CY;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_C_XOR;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_D;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_D1;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_D2;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_D3;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_D4;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_D5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_D6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_DO5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_DO6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_D_CY;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_D_XOR;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_A;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_A1;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_A2;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_A3;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_A4;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_A5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_A6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_AO5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_AO6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_A_CY;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_A_XOR;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_B;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_B1;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_B2;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_B3;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_B4;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_B5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_B6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_BO5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_BO6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_B_CY;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_B_XOR;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_C;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_C1;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_C2;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_C3;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_C4;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_C5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_C6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_CO5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_CO6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_C_CY;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_C_XOR;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_D;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_D1;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_D2;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_D3;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_D4;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_D5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_D6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_DO5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_DO6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_D_CY;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_D_XOR;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_A;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_A1;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_A2;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_A3;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_A4;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_A5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_A6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_AMUX;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_AO5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_AO6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_A_CY;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_A_XOR;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_B;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_B1;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_B2;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_B3;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_B4;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_B5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_B6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_BMUX;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_BO5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_BO6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_B_CY;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_B_XOR;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_C;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_C1;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_C2;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_C3;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_C4;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_C5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_C6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_CO5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_CO6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_C_CY;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_C_XOR;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_D;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_D1;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_D2;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_D3;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_D4;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_D5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_D6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_DO5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_DO6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_D_CY;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_D_XOR;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_A;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_A1;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_A2;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_A3;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_A4;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_A5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_A6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_AMUX;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_AO5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_AO6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_A_CY;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_A_XOR;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_B;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_B1;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_B2;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_B3;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_B4;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_B5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_B6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_BO5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_BO6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_B_CY;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_B_XOR;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_C;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_C1;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_C2;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_C3;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_C4;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_C5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_C6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_CO5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_CO6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_C_CY;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_C_XOR;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_D;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_D1;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_D2;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_D3;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_D4;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_D5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_D6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_DO5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_DO6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_D_CY;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_D_XOR;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_A;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_A1;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_A2;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_A3;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_A4;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_A5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_A6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_AMUX;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_AO5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_AO6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_A_CY;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_A_XOR;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_B;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_B1;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_B2;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_B3;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_B4;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_B5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_B6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_BO5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_BO6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_B_CY;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_B_XOR;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_C;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_C1;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_C2;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_C3;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_C4;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_C5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_C6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_CO5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_CO6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_C_CY;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_C_XOR;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_D;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_D1;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_D2;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_D3;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_D4;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_D5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_D6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_DO5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_DO6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_D_CY;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_D_XOR;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_A;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_A1;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_A2;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_A3;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_A4;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_A5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_A6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_AMUX;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_AO5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_AO6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_A_CY;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_A_XOR;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_B;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_B1;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_B2;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_B3;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_B4;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_B5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_B6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_BO5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_BO6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_B_CY;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_B_XOR;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_C;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_C1;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_C2;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_C3;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_C4;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_C5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_C6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_CO5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_CO6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_C_CY;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_C_XOR;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_D;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_D1;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_D2;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_D3;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_D4;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_D5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_D6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_DO5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_DO6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_D_CY;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_D_XOR;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_A;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_A1;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_A2;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_A3;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_A4;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_A5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_A6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_AMUX;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_AO5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_AO6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_A_CY;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_A_XOR;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_B;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_B1;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_B2;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_B3;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_B4;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_B5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_B6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_BO5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_BO6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_B_CY;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_B_XOR;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_C;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_C1;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_C2;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_C3;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_C4;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_C5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_C6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_CO5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_CO6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_C_CY;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_C_XOR;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_D;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_D1;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_D2;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_D3;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_D4;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_D5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_D6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_DO5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_DO6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_D_CY;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_D_XOR;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_A;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_A1;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_A2;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_A3;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_A4;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_A5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_A6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_AMUX;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_AO5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_AO6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_A_CY;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_A_XOR;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_B;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_B1;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_B2;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_B3;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_B4;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_B5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_B6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_BO5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_BO6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_B_CY;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_B_XOR;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_C;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_C1;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_C2;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_C3;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_C4;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_C5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_C6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_CO5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_CO6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_C_CY;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_C_XOR;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_D;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_D1;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_D2;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_D3;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_D4;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_D5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_D6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_DMUX;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_DO5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_DO6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_D_CY;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_D_XOR;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_A;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_A1;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_A2;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_A3;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_A4;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_A5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_A6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_AO5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_AO6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_A_CY;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_A_XOR;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_B;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_B1;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_B2;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_B3;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_B4;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_B5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_B6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_BO5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_BO6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_B_CY;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_B_XOR;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_C;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_C1;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_C2;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_C3;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_C4;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_C5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_C6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_CO5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_CO6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_C_CY;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_C_XOR;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_D;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_D1;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_D2;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_D3;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_D4;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_D5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_D6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_DO5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_DO6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_D_CY;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_D_XOR;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_A;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_A1;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_A2;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_A3;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_A4;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_A5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_A6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_AMUX;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_AO5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_AO6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_A_CY;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_A_XOR;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_B;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_B1;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_B2;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_B3;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_B4;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_B5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_B6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_BO5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_BO6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_B_CY;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_B_XOR;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_C;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_C1;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_C2;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_C3;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_C4;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_C5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_C6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_CO5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_CO6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_C_CY;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_C_XOR;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_D;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_D1;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_D2;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_D3;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_D4;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_D5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_D6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_DO5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_DO6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_D_CY;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_D_XOR;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_A;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_A1;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_A2;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_A3;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_A4;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_A5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_A6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_AO5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_AO6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_A_CY;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_A_XOR;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_B;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_B1;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_B2;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_B3;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_B4;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_B5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_B6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_BO5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_BO6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_B_CY;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_B_XOR;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_C;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_C1;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_C2;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_C3;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_C4;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_C5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_C6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_CO5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_CO6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_C_CY;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_C_XOR;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_D;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_D1;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_D2;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_D3;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_D4;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_D5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_D6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_DO5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_DO6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_D_CY;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_D_XOR;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_A;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_A1;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_A2;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_A3;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_A4;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_A5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_A6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_AO5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_AO6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_A_CY;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_A_XOR;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_B;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_B1;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_B2;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_B3;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_B4;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_B5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_B6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_BO5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_BO6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_B_CY;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_B_XOR;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_C;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_C1;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_C2;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_C3;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_C4;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_C5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_C6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_CO5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_CO6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_C_CY;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_C_XOR;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_D;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_D1;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_D2;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_D3;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_D4;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_D5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_D6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_DO5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_DO6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_D_CY;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_D_XOR;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_A;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_A1;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_A2;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_A3;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_A4;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_A5;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_A6;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_AMUX;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_AO5;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_AO6;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_A_CY;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_A_XOR;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_B;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_B1;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_B2;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_B3;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_B4;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_B5;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_B6;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_BO5;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_BO6;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_B_CY;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_B_XOR;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_C;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_C1;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_C2;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_C3;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_C4;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_C5;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_C6;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_CO5;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_CO6;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_C_CY;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_C_XOR;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_D;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_D1;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_D2;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_D3;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_D4;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_D5;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_D6;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_DO5;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_DO6;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_D_CY;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_D_XOR;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_A;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_A1;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_A2;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_A3;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_A4;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_A5;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_A6;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_AO5;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_AO6;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_A_CY;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_A_XOR;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_B;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_B1;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_B2;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_B3;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_B4;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_B5;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_B6;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_BO5;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_BO6;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_B_CY;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_B_XOR;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_C;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_C1;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_C2;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_C3;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_C4;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_C5;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_C6;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_CO5;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_CO6;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_C_CY;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_C_XOR;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_D;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_D1;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_D2;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_D3;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_D4;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_D5;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_D6;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_DO5;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_DO6;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_D_CY;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_D_XOR;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_A;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_A1;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_A2;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_A3;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_A4;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_A5;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_A6;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_AMUX;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_AO5;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_AO6;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_A_CY;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_A_XOR;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_B;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_B1;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_B2;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_B3;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_B4;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_B5;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_B6;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_BO5;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_BO6;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_B_CY;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_B_XOR;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_C;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_C1;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_C2;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_C3;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_C4;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_C5;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_C6;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_CO5;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_CO6;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_C_CY;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_C_XOR;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_D;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_D1;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_D2;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_D3;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_D4;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_D5;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_D6;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_DO5;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_DO6;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_D_CY;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_D_XOR;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_A;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_A1;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_A2;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_A3;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_A4;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_A5;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_A6;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_AO5;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_AO6;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_A_CY;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_A_XOR;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_B;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_B1;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_B2;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_B3;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_B4;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_B5;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_B6;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_BO5;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_BO6;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_B_CY;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_B_XOR;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_C;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_C1;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_C2;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_C3;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_C4;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_C5;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_C6;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_CO5;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_CO6;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_C_CY;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_C_XOR;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_D;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_D1;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_D2;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_D3;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_D4;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_D5;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_D6;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_DO5;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_DO6;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_D_CY;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_D_XOR;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_A;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_A1;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_A2;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_A3;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_A4;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_A5;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_A6;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_AMUX;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_AO5;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_AO6;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_A_CY;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_A_XOR;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_B;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_B1;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_B2;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_B3;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_B4;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_B5;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_B6;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_BO5;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_BO6;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_B_CY;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_B_XOR;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_C;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_C1;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_C2;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_C3;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_C4;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_C5;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_C6;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_CMUX;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_CO5;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_CO6;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_C_CY;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_C_XOR;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_D;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_D1;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_D2;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_D3;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_D4;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_D5;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_D6;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_DO5;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_DO6;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_D_CY;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_D_XOR;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_A;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_A1;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_A2;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_A3;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_A4;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_A5;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_A6;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_AO5;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_AO6;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_A_CY;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_A_XOR;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_B;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_B1;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_B2;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_B3;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_B4;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_B5;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_B6;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_BO5;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_BO6;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_B_CY;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_B_XOR;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_C;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_C1;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_C2;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_C3;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_C4;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_C5;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_C6;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_CO5;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_CO6;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_C_CY;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_C_XOR;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_D;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_D1;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_D2;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_D3;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_D4;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_D5;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_D6;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_DO5;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_DO6;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_D_CY;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_D_XOR;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_A;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_A1;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_A2;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_A3;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_A4;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_A5;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_A6;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_AMUX;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_AO5;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_AO6;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_A_CY;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_A_XOR;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_B;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_B1;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_B2;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_B3;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_B4;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_B5;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_B6;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_BMUX;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_BO5;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_BO6;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_B_CY;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_B_XOR;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_C;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_C1;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_C2;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_C3;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_C4;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_C5;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_C6;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_CO5;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_CO6;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_C_CY;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_C_XOR;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_D;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_D1;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_D2;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_D3;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_D4;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_D5;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_D6;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_DO5;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_DO6;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_D_CY;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_D_XOR;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_A;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_A1;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_A2;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_A3;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_A4;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_A5;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_A6;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_AMUX;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_AO5;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_AO6;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_A_CY;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_A_XOR;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_B;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_B1;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_B2;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_B3;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_B4;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_B5;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_B6;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_BO5;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_BO6;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_B_CY;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_B_XOR;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_C;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_C1;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_C2;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_C3;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_C4;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_C5;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_C6;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_CO5;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_CO6;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_C_CY;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_C_XOR;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_D;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_D1;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_D2;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_D3;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_D4;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_D5;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_D6;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_DO5;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_DO6;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_D_CY;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_D_XOR;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_A;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_A1;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_A2;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_A3;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_A4;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_A5;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_A6;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_AMUX;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_AO5;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_AO6;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_A_CY;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_A_XOR;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_B;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_B1;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_B2;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_B3;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_B4;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_B5;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_B6;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_BO5;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_BO6;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_B_CY;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_B_XOR;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_C;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_C1;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_C2;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_C3;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_C4;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_C5;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_C6;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_CO5;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_CO6;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_C_CY;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_C_XOR;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_D;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_D1;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_D2;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_D3;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_D4;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_D5;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_D6;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_DO5;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_DO6;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_D_CY;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_D_XOR;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_A;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_A1;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_A2;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_A3;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_A4;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_A5;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_A6;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_AMUX;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_AO5;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_AO6;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_A_CY;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_A_XOR;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_B;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_B1;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_B2;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_B3;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_B4;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_B5;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_B6;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_BO5;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_BO6;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_B_CY;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_B_XOR;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_C;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_C1;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_C2;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_C3;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_C4;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_C5;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_C6;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_CO5;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_CO6;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_C_CY;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_C_XOR;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_D;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_D1;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_D2;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_D3;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_D4;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_D5;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_D6;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_DO5;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_DO6;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_D_CY;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_D_XOR;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_A;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_A1;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_A2;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_A3;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_A4;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_A5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_A6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_AMUX;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_AO5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_AO6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_A_CY;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_A_XOR;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_B;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_B1;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_B2;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_B3;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_B4;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_B5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_B6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_BO5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_BO6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_B_CY;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_B_XOR;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_C;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_C1;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_C2;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_C3;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_C4;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_C5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_C6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_CO5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_CO6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_C_CY;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_C_XOR;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_D;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_D1;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_D2;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_D3;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_D4;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_D5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_D6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_DO5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_DO6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_D_CY;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_D_XOR;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_A;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_A1;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_A2;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_A3;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_A4;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_A5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_A6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_AO5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_AO6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_A_CY;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_A_XOR;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_B;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_B1;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_B2;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_B3;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_B4;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_B5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_B6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_BO5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_BO6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_B_CY;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_B_XOR;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_C;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_C1;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_C2;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_C3;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_C4;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_C5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_C6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_CO5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_CO6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_C_CY;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_C_XOR;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_D;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_D1;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_D2;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_D3;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_D4;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_D5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_D6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_DO5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_DO6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_D_CY;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_D_XOR;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_A;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_A1;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_A2;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_A3;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_A4;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_A5;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_A6;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_AO5;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_AO6;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_A_CY;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_A_XOR;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_B;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_B1;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_B2;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_B3;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_B4;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_B5;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_B6;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_BO5;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_BO6;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_B_CY;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_B_XOR;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_C;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_C1;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_C2;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_C3;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_C4;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_C5;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_C6;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_CO5;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_CO6;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_C_CY;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_C_XOR;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_D;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_D1;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_D2;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_D3;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_D4;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_D5;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_D6;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_DO5;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_DO6;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_D_CY;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_D_XOR;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_A;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_A1;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_A2;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_A3;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_A4;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_A5;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_A6;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_AO5;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_AO6;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_A_CY;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_A_XOR;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_B;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_B1;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_B2;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_B3;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_B4;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_B5;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_B6;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_BO5;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_BO6;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_B_CY;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_B_XOR;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_C;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_C1;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_C2;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_C3;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_C4;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_C5;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_C6;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_CO5;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_CO6;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_C_CY;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_C_XOR;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_D;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_D1;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_D2;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_D3;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_D4;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_D5;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_D6;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_DO5;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_DO6;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_D_CY;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_D_XOR;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_A;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_A1;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_A2;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_A3;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_A4;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_A5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_A6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_AO5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_AO6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_A_CY;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_A_XOR;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_B;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_B1;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_B2;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_B3;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_B4;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_B5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_B6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_BO5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_BO6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_B_CY;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_B_XOR;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_C;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_C1;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_C2;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_C3;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_C4;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_C5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_C6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_CO5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_CO6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_C_CY;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_C_XOR;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_D;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_D1;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_D2;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_D3;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_D4;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_D5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_D6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_DO5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_DO6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_D_CY;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_D_XOR;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_A;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_A1;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_A2;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_A3;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_A4;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_A5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_A6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_AO5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_AO6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_A_CY;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_A_XOR;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_B;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_B1;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_B2;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_B3;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_B4;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_B5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_B6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_BO5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_BO6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_B_CY;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_B_XOR;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_C;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_C1;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_C2;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_C3;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_C4;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_C5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_C6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_CO5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_CO6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_C_CY;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_C_XOR;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_D;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_D1;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_D2;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_D3;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_D4;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_D5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_D6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_DO5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_DO6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_D_CY;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_D_XOR;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_A;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_A1;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_A2;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_A3;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_A4;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_A5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_A6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_AMUX;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_AO5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_AO6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_A_CY;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_A_XOR;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_B;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_B1;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_B2;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_B3;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_B4;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_B5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_B6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_BMUX;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_BO5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_BO6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_B_CY;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_B_XOR;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_C;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_C1;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_C2;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_C3;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_C4;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_C5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_C6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_CO5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_CO6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_C_CY;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_C_XOR;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_D;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_D1;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_D2;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_D3;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_D4;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_D5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_D6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_DO5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_DO6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_D_CY;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_D_XOR;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_A;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_A1;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_A2;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_A3;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_A4;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_A5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_A6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_AO5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_AO6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_A_CY;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_A_XOR;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_B;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_B1;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_B2;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_B3;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_B4;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_B5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_B6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_BO5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_BO6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_B_CY;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_B_XOR;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_C;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_C1;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_C2;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_C3;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_C4;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_C5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_C6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_CO5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_CO6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_C_CY;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_C_XOR;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_D;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_D1;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_D2;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_D3;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_D4;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_D5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_D6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_DO5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_DO6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_D_CY;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_D_XOR;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_A;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_A1;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_A2;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_A3;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_A4;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_A5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_A6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_AO5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_AO6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_A_CY;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_A_XOR;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_B;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_B1;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_B2;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_B3;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_B4;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_B5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_B6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_BO5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_BO6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_B_CY;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_B_XOR;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_C;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_C1;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_C2;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_C3;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_C4;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_C5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_C6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_CO5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_CO6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_C_CY;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_C_XOR;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_D;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_D1;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_D2;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_D3;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_D4;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_D5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_D6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_DO5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_DO6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_D_CY;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_D_XOR;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_A;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_A1;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_A2;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_A3;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_A4;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_A5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_A6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_AO5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_AO6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_A_CY;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_A_XOR;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_B;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_B1;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_B2;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_B3;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_B4;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_B5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_B6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_BO5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_BO6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_B_CY;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_B_XOR;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_C;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_C1;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_C2;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_C3;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_C4;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_C5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_C6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_CO5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_CO6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_C_CY;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_C_XOR;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_D;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_D1;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_D2;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_D3;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_D4;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_D5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_D6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_DO5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_DO6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_D_CY;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_D_XOR;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_A;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_A1;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_A2;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_A3;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_A4;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_A5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_A6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_AMUX;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_AO5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_AO6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_A_CY;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_A_XOR;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_B;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_B1;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_B2;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_B3;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_B4;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_B5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_B6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_BO5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_BO6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_B_CY;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_B_XOR;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_C;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_C1;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_C2;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_C3;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_C4;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_C5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_C6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_CO5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_CO6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_C_CY;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_C_XOR;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_D;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_D1;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_D2;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_D3;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_D4;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_D5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_D6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_DO5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_DO6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_D_CY;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_D_XOR;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_A;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_A1;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_A2;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_A3;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_A4;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_A5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_A6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_AMUX;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_AO5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_AO6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_A_CY;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_A_XOR;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_B;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_B1;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_B2;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_B3;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_B4;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_B5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_B6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_BO5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_BO6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_B_CY;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_B_XOR;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_C;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_C1;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_C2;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_C3;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_C4;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_C5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_C6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_CO5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_CO6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_C_CY;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_C_XOR;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_D;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_D1;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_D2;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_D3;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_D4;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_D5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_D6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_DO5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_DO6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_D_CY;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_D_XOR;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_A;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_A1;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_A2;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_A3;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_A4;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_A5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_A6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_AO5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_AO6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_A_CY;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_A_XOR;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_B;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_B1;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_B2;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_B3;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_B4;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_B5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_B6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_BO5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_BO6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_B_CY;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_B_XOR;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_C;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_C1;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_C2;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_C3;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_C4;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_C5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_C6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_CO5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_CO6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_C_CY;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_C_XOR;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_D;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_D1;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_D2;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_D3;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_D4;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_D5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_D6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_DO5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_DO6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_D_CY;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_D_XOR;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_A;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_A1;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_A2;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_A3;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_A4;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_A5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_A6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_AMUX;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_AO5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_AO6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_A_CY;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_A_XOR;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_B;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_B1;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_B2;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_B3;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_B4;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_B5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_B6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_BO5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_BO6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_B_CY;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_B_XOR;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_C;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_C1;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_C2;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_C3;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_C4;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_C5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_C6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_CO5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_CO6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_C_CY;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_C_XOR;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_D;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_D1;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_D2;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_D3;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_D4;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_D5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_D6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_DO5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_DO6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_D_CY;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_D_XOR;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_A;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_A1;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_A2;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_A3;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_A4;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_A5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_A6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_AO5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_AO6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_A_CY;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_A_XOR;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_B;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_B1;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_B2;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_B3;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_B4;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_B5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_B6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_BO5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_BO6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_B_CY;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_B_XOR;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_C;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_C1;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_C2;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_C3;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_C4;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_C5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_C6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_CO5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_CO6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_C_CY;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_C_XOR;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_D;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_D1;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_D2;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_D3;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_D4;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_D5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_D6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_DO5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_DO6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_D_CY;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_D_XOR;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_A;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_A1;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_A2;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_A3;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_A4;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_A5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_A6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_AMUX;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_AO5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_AO6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_A_CY;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_A_XOR;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_B;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_B1;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_B2;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_B3;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_B4;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_B5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_B6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_BO5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_BO6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_B_CY;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_B_XOR;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_C;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_C1;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_C2;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_C3;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_C4;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_C5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_C6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_CO5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_CO6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_C_CY;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_C_XOR;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_D;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_D1;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_D2;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_D3;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_D4;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_D5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_D6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_DO5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_DO6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_D_CY;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_D_XOR;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A1;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A2;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A3;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A4;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_AMUX;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_AO5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_AO6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A_CY;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A_XOR;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B1;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B2;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B3;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B4;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_BO5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_BO6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B_CY;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B_XOR;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C1;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C2;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C3;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C4;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_CO5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_CO6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C_CY;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C_XOR;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D1;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D2;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D3;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D4;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_DO5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_DO6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D_CY;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D_XOR;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A1;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A2;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A3;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A4;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_AO5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_AO6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A_CY;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A_XOR;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B1;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B2;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B3;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B4;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_BMUX;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_BO5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_BO6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B_CY;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B_XOR;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C1;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C2;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C3;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C4;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_CO5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_CO6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C_CY;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C_XOR;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D1;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D2;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D3;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D4;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_DO5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_DO6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D_CY;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D_XOR;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A1;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A2;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A3;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A4;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_AMUX;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_AO5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_AO6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A_CY;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A_XOR;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B1;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B2;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B3;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B4;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_BO5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_BO6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B_CY;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B_XOR;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C1;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C2;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C3;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C4;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_CO5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_CO6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C_CY;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C_XOR;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D1;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D2;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D3;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D4;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_DO5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_DO6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D_CY;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D_XOR;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A1;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A2;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A3;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A4;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_AO5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_AO6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A_CY;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A_XOR;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B1;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B2;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B3;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B4;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_BO5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_BO6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B_CY;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B_XOR;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C1;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C2;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C3;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C4;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_CO5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_CO6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C_CY;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C_XOR;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D1;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D2;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D3;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D4;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_DO5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_DO6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D_CY;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D_XOR;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A1;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A2;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A3;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A4;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_AMUX;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_AO5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_AO6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A_CY;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A_XOR;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B1;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B2;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B3;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B4;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_BO5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_BO6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B_CY;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B_XOR;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C1;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C2;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C3;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C4;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_CO5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_CO6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C_CY;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C_XOR;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D1;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D2;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D3;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D4;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_DO5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_DO6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D_CY;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D_XOR;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A1;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A2;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A3;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A4;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_AO5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_AO6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A_CY;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A_XOR;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B1;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B2;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B3;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B4;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_BO5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_BO6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B_CY;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B_XOR;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C1;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C2;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C3;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C4;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_CO5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_CO6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C_CY;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C_XOR;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D1;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D2;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D3;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D4;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_DO5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_DO6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D_CY;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D_XOR;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A1;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A2;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A3;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A4;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_AMUX;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_AO5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_AO6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A_CY;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A_XOR;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B1;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B2;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B3;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B4;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_BO5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_BO6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B_CY;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B_XOR;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C1;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C2;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C3;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C4;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_CO5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_CO6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C_CY;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C_XOR;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D1;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D2;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D3;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D4;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_DO5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_DO6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D_CY;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D_XOR;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A1;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A2;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A3;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A4;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_AO5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_AO6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A_CY;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A_XOR;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B1;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B2;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B3;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B4;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_BO5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_BO6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B_CY;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B_XOR;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C1;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C2;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C3;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C4;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_CO5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_CO6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C_CY;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C_XOR;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D1;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D2;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D3;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D4;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_DO5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_DO6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D_CY;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D_XOR;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_A;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_A1;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_A2;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_A3;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_A4;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_A5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_A6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_AO5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_AO6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_A_CY;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_A_XOR;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_B;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_B1;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_B2;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_B3;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_B4;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_B5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_B6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_BO5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_BO6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_B_CY;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_B_XOR;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_C;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_C1;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_C2;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_C3;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_C4;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_C5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_C6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_CO5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_CO6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_C_CY;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_C_XOR;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_D;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_D1;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_D2;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_D3;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_D4;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_D5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_D6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_DO5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_DO6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_D_CY;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_D_XOR;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_A;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_A1;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_A2;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_A3;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_A4;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_A5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_A6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_AO5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_AO6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_A_CY;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_A_XOR;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_B;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_B1;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_B2;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_B3;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_B4;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_B5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_B6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_BO5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_BO6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_B_CY;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_B_XOR;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_C;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_C1;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_C2;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_C3;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_C4;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_C5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_C6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_CO5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_CO6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_C_CY;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_C_XOR;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_D;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_D1;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_D2;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_D3;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_D4;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_D5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_D6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_DO5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_DO6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_D_CY;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_D_XOR;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_A;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_A1;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_A2;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_A3;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_A4;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_A5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_A6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_AMUX;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_AO5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_AO6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_A_CY;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_A_XOR;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_B;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_B1;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_B2;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_B3;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_B4;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_B5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_B6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_BO5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_BO6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_B_CY;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_B_XOR;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_C;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_C1;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_C2;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_C3;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_C4;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_C5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_C6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_CMUX;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_CO5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_CO6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_C_CY;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_C_XOR;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_D;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_D1;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_D2;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_D3;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_D4;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_D5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_D6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_DO5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_DO6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_D_CY;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_D_XOR;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_A;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_A1;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_A2;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_A3;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_A4;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_A5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_A6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_AO5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_AO6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_A_CY;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_A_XOR;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_B;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_B1;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_B2;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_B3;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_B4;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_B5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_B6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_BO5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_BO6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_B_CY;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_B_XOR;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_C;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_C1;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_C2;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_C3;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_C4;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_C5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_C6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_CO5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_CO6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_C_CY;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_C_XOR;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_D;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_D1;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_D2;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_D3;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_D4;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_D5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_D6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_DO5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_DO6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_D_CY;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_D_XOR;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_A;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_A1;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_A2;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_A3;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_A4;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_A5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_A6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_AMUX;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_AO5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_AO6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_A_CY;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_A_XOR;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_B;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_B1;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_B2;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_B3;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_B4;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_B5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_B6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_BO5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_BO6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_B_CY;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_B_XOR;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_C;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_C1;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_C2;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_C3;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_C4;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_C5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_C6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_CO5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_CO6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_C_CY;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_C_XOR;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_D;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_D1;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_D2;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_D3;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_D4;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_D5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_D6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_DO5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_DO6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_D_CY;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_D_XOR;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_A;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_A1;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_A2;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_A3;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_A4;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_A5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_A6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_AO5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_AO6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_A_CY;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_A_XOR;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_B;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_B1;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_B2;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_B3;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_B4;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_B5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_B6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_BO5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_BO6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_B_CY;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_B_XOR;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_C;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_C1;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_C2;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_C3;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_C4;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_C5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_C6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_CO5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_CO6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_C_CY;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_C_XOR;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_D;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_D1;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_D2;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_D3;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_D4;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_D5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_D6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_DO5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_DO6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_D_CY;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_D_XOR;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_A;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_A1;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_A2;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_A3;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_A4;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_A5;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_A6;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_AO5;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_AO6;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_A_CY;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_A_XOR;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_B;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_B1;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_B2;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_B3;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_B4;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_B5;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_B6;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_BMUX;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_BO5;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_BO6;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_B_CY;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_B_XOR;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_C;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_C1;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_C2;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_C3;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_C4;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_C5;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_C6;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_CO5;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_CO6;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_C_CY;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_C_XOR;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_D;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_D1;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_D2;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_D3;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_D4;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_D5;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_D6;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_DO5;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_DO6;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_D_CY;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_D_XOR;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_A;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_A1;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_A2;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_A3;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_A4;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_A5;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_A6;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_AMUX;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_AO5;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_AO6;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_A_CY;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_A_XOR;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_B;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_B1;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_B2;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_B3;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_B4;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_B5;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_B6;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_BO5;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_BO6;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_B_CY;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_B_XOR;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_C;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_C1;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_C2;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_C3;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_C4;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_C5;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_C6;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_CO5;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_CO6;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_C_CY;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_C_XOR;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_D;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_D1;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_D2;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_D3;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_D4;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_D5;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_D6;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_DMUX;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_DO5;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_DO6;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_D_CY;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_D_XOR;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_A;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_A1;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_A2;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_A3;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_A4;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_A5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_A6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_AMUX;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_AO5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_AO6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_A_CY;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_A_XOR;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_B;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_B1;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_B2;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_B3;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_B4;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_B5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_B6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_BO5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_BO6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_B_CY;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_B_XOR;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_C;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_C1;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_C2;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_C3;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_C4;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_C5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_C6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_CO5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_CO6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_C_CY;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_C_XOR;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_D;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_D1;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_D2;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_D3;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_D4;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_D5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_D6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_DO5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_DO6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_D_CY;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_D_XOR;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_A;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_A1;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_A2;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_A3;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_A4;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_A5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_A6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_AMUX;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_AO5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_AO6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_A_CY;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_A_XOR;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_B;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_B1;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_B2;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_B3;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_B4;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_B5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_B6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_BO5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_BO6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_B_CY;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_B_XOR;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_C;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_C1;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_C2;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_C3;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_C4;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_C5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_C6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_CO5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_CO6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_C_CY;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_C_XOR;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_D;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_D1;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_D2;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_D3;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_D4;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_D5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_D6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_DO5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_DO6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_D_CY;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_D_XOR;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_A;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_A1;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_A2;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_A3;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_A4;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_A5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_A6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_AMUX;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_AO5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_AO6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_A_CY;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_A_XOR;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_B;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_B1;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_B2;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_B3;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_B4;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_B5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_B6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_BMUX;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_BO5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_BO6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_B_CY;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_B_XOR;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_C;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_C1;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_C2;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_C3;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_C4;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_C5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_C6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_CO5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_CO6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_C_CY;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_C_XOR;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_D;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_D1;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_D2;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_D3;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_D4;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_D5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_D6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_DO5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_DO6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_D_CY;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_D_XOR;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_A;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_A1;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_A2;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_A3;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_A4;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_A5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_A6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_AMUX;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_AO5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_AO6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_A_CY;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_A_XOR;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_B;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_B1;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_B2;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_B3;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_B4;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_B5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_B6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_BO5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_BO6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_B_CY;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_B_XOR;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_C;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_C1;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_C2;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_C3;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_C4;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_C5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_C6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_CO5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_CO6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_C_CY;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_C_XOR;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_D;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_D1;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_D2;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_D3;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_D4;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_D5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_D6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_DO5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_DO6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_D_CY;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_D_XOR;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_A;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_A1;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_A2;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_A3;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_A4;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_A5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_A6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_AMUX;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_AO5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_AO6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_A_CY;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_A_XOR;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_B;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_B1;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_B2;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_B3;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_B4;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_B5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_B6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_BO5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_BO6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_B_CY;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_B_XOR;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_C;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_C1;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_C2;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_C3;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_C4;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_C5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_C6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_CMUX;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_CO5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_CO6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_C_CY;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_C_XOR;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_D;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_D1;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_D2;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_D3;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_D4;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_D5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_D6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_DO5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_DO6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_D_CY;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_D_XOR;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_A;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_A1;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_A2;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_A3;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_A4;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_A5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_A6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_AMUX;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_AO5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_AO6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_A_CY;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_A_XOR;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_B;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_B1;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_B2;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_B3;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_B4;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_B5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_B6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_BO5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_BO6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_B_CY;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_B_XOR;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_C;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_C1;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_C2;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_C3;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_C4;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_C5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_C6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_CMUX;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_CO5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_CO6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_C_CY;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_C_XOR;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_D;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_D1;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_D2;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_D3;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_D4;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_D5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_D6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_DO5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_DO6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_D_CY;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_D_XOR;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_A;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_A1;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_A2;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_A3;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_A4;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_A5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_A6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_AMUX;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_AO5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_AO6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_A_CY;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_A_XOR;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_B;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_B1;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_B2;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_B3;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_B4;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_B5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_B6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_BO5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_BO6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_B_CY;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_B_XOR;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_C;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_C1;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_C2;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_C3;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_C4;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_C5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_C6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_CMUX;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_CO5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_CO6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_C_CY;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_C_XOR;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_D;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_D1;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_D2;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_D3;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_D4;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_D5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_D6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_DO5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_DO6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_D_CY;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_D_XOR;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_A;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_A1;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_A2;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_A3;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_A4;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_A5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_A6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_AMUX;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_AO5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_AO6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_A_CY;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_A_XOR;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_B;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_B1;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_B2;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_B3;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_B4;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_B5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_B6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_BO5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_BO6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_B_CY;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_B_XOR;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_C;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_C1;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_C2;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_C3;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_C4;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_C5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_C6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_CO5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_CO6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_C_CY;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_C_XOR;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_D;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_D1;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_D2;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_D3;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_D4;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_D5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_D6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_DO5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_DO6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_D_CY;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_D_XOR;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_A;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_A1;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_A2;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_A3;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_A4;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_A5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_A6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_AMUX;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_AO5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_AO6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_A_CY;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_A_XOR;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_B;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_B1;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_B2;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_B3;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_B4;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_B5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_B6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_BMUX;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_BO5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_BO6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_B_CY;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_B_XOR;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_C;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_C1;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_C2;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_C3;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_C4;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_C5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_C6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_CO5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_CO6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_C_CY;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_C_XOR;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_D;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_D1;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_D2;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_D3;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_D4;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_D5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_D6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_DO5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_DO6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_D_CY;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_D_XOR;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_A;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_A1;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_A2;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_A3;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_A4;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_A5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_A6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_AO5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_AO6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_A_CY;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_A_XOR;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_B;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_B1;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_B2;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_B3;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_B4;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_B5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_B6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_BMUX;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_BO5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_BO6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_B_CY;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_B_XOR;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_C;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_C1;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_C2;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_C3;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_C4;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_C5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_C6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_CO5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_CO6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_C_CY;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_C_XOR;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_D;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_D1;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_D2;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_D3;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_D4;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_D5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_D6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_DO5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_DO6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_D_CY;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_D_XOR;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_A;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_A1;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_A2;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_A3;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_A4;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_A5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_A6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_AMUX;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_AO5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_AO6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_A_CY;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_A_XOR;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_B;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_B1;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_B2;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_B3;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_B4;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_B5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_B6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_BO5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_BO6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_B_CY;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_B_XOR;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_C;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_C1;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_C2;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_C3;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_C4;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_C5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_C6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_CO5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_CO6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_C_CY;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_C_XOR;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_D;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_D1;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_D2;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_D3;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_D4;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_D5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_D6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_DO5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_DO6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_D_CY;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_D_XOR;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_A;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_A1;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_A2;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_A3;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_A4;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_A5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_A6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_AO5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_AO6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_A_CY;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_A_XOR;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_B;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_B1;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_B2;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_B3;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_B4;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_B5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_B6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_BO5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_BO6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_B_CY;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_B_XOR;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_C;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_C1;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_C2;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_C3;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_C4;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_C5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_C6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_CO5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_CO6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_C_CY;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_C_XOR;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_D;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_D1;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_D2;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_D3;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_D4;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_D5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_D6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_DO5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_DO6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_D_CY;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_D_XOR;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_A;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_A1;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_A2;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_A3;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_A4;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_A5;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_A6;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_AO5;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_AO6;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_A_CY;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_A_XOR;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_B;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_B1;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_B2;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_B3;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_B4;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_B5;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_B6;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_BO5;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_BO6;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_B_CY;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_B_XOR;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_C;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_C1;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_C2;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_C3;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_C4;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_C5;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_C6;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_CO5;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_CO6;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_C_CY;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_C_XOR;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_D;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_D1;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_D2;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_D3;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_D4;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_D5;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_D6;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_DO5;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_DO6;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_D_CY;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_D_XOR;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_A;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_A1;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_A2;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_A3;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_A4;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_A5;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_A6;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_AMUX;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_AO5;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_AO6;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_A_CY;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_A_XOR;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_B;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_B1;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_B2;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_B3;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_B4;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_B5;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_B6;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_BO5;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_BO6;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_B_CY;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_B_XOR;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_C;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_C1;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_C2;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_C3;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_C4;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_C5;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_C6;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_CO5;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_CO6;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_C_CY;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_C_XOR;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_D;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_D1;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_D2;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_D3;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_D4;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_D5;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_D6;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_DO5;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_DO6;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_D_CY;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_D_XOR;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_A;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_A1;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_A2;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_A3;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_A4;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_A5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_A6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_AO5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_AO6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_A_CY;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_A_XOR;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_B;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_B1;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_B2;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_B3;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_B4;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_B5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_B6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_BMUX;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_BO5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_BO6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_B_CY;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_B_XOR;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_C;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_C1;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_C2;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_C3;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_C4;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_C5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_C6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_CO5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_CO6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_C_CY;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_C_XOR;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_D;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_D1;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_D2;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_D3;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_D4;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_D5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_D6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_DO5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_D_CY;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_D_XOR;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_A;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_A1;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_A2;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_A3;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_A4;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_A5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_A6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_AMUX;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_AO5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_AO6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_A_CY;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_A_XOR;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_B;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_B1;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_B2;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_B3;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_B4;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_B5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_B6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_BO5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_BO6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_B_CY;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_B_XOR;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_C;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_C1;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_C2;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_C3;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_C4;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_C5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_C6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_CO5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_CO6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_C_CY;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_C_XOR;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_D;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_D1;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_D2;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_D3;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_D4;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_D5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_D6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_DO5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_DO6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_D_CY;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_D_XOR;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_A;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_A1;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_A2;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_A3;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_A4;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_A5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_A6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_AO5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_AO6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_A_CY;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_A_XOR;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_B;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_B1;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_B2;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_B3;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_B4;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_B5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_B6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_BO5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_BO6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_B_CY;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_B_XOR;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_C;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_C1;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_C2;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_C3;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_C4;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_C5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_C6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_CO5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_CO6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_C_CY;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_C_XOR;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_D;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_D1;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_D2;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_D3;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_D4;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_D5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_D6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_DO5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_DO6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_D_CY;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_D_XOR;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_A;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_A1;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_A2;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_A3;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_A4;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_A5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_A6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_AO5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_AO6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_A_CY;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_A_XOR;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_B;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_B1;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_B2;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_B3;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_B4;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_B5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_B6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_BO5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_BO6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_B_CY;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_B_XOR;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_C;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_C1;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_C2;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_C3;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_C4;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_C5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_C6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_CO5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_CO6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_C_CY;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_C_XOR;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_D;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_D1;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_D2;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_D3;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_D4;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_D5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_D6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_DO5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_DO6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_D_CY;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_D_XOR;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_A;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_A1;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_A2;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_A3;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_A4;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_A5;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_A6;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_AO5;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_AO6;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_A_CY;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_A_XOR;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_B;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_B1;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_B2;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_B3;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_B4;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_B5;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_B6;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_BO5;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_BO6;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_B_CY;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_B_XOR;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_C;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_C1;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_C2;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_C3;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_C4;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_C5;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_C6;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_CO5;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_CO6;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_C_CY;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_C_XOR;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_D;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_D1;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_D2;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_D3;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_D4;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_D5;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_D6;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_DO5;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_DO6;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_D_CY;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_D_XOR;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_A;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_A1;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_A2;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_A3;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_A4;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_A5;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_A6;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_AMUX;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_AO5;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_AO6;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_A_CY;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_A_XOR;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_B;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_B1;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_B2;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_B3;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_B4;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_B5;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_B6;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_BO5;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_BO6;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_B_CY;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_B_XOR;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_C;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_C1;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_C2;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_C3;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_C4;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_C5;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_C6;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_CO5;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_CO6;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_C_CY;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_C_XOR;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_D;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_D1;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_D2;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_D3;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_D4;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_D5;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_D6;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_DO5;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_DO6;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_D_CY;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_D_XOR;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_A;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_A1;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_A2;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_A3;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_A4;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_A5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_A6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_AO5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_AO6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_A_CY;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_A_XOR;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_B;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_B1;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_B2;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_B3;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_B4;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_B5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_B6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_BO5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_BO6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_B_CY;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_B_XOR;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_C;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_C1;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_C2;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_C3;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_C4;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_C5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_C6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_CO5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_CO6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_C_CY;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_C_XOR;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_D;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_D1;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_D2;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_D3;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_D4;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_D5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_D6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_DO5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_DO6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_D_CY;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_D_XOR;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_A;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_A1;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_A2;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_A3;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_A4;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_A5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_A6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_AMUX;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_AO5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_AO6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_A_CY;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_A_XOR;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_B;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_B1;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_B2;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_B3;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_B4;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_B5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_B6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_BO5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_BO6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_B_CY;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_B_XOR;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_C;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_C1;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_C2;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_C3;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_C4;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_C5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_C6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_CO5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_CO6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_C_CY;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_C_XOR;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_D;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_D1;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_D2;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_D3;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_D4;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_D5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_D6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_DO5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_DO6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_D_CY;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_D_XOR;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_A;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_A1;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_A2;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_A3;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_A4;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_A5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_A6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_AO5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_AO6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_A_CY;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_A_XOR;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_B;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_B1;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_B2;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_B3;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_B4;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_B5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_B6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_BO5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_BO6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_B_CY;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_B_XOR;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_C;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_C1;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_C2;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_C3;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_C4;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_C5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_C6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_CO5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_CO6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_C_CY;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_C_XOR;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_D;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_D1;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_D2;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_D3;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_D4;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_D5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_D6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_DO5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_DO6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_D_CY;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_D_XOR;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_A;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_A1;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_A2;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_A3;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_A4;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_A5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_A6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_AMUX;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_AO5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_AO6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_A_CY;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_A_XOR;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_B;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_B1;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_B2;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_B3;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_B4;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_B5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_B6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_BMUX;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_BO5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_BO6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_B_CY;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_B_XOR;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_C;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_C1;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_C2;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_C3;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_C4;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_C5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_C6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_CO5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_CO6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_C_CY;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_C_XOR;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_D;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_D1;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_D2;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_D3;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_D4;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_D5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_D6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_DO5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_DO6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_D_CY;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_D_XOR;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_A;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_A1;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_A2;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_A3;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_A4;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_A5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_A6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_AMUX;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_AO5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_AO6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_A_CY;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_A_XOR;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_B;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_B1;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_B2;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_B3;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_B4;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_B5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_B6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_BO5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_BO6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_B_CY;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_B_XOR;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_C;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_C1;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_C2;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_C3;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_C4;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_C5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_C6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_CO5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_CO6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_C_CY;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_C_XOR;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_D;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_D1;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_D2;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_D3;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_D4;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_D5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_D6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_DO5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_DO6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_D_CY;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_D_XOR;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_A;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_A1;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_A2;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_A3;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_A4;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_A5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_A6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_AO5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_AO6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_A_CY;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_A_XOR;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_B;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_B1;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_B2;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_B3;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_B4;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_B5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_B6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_BO5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_BO6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_B_CY;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_B_XOR;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_C;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_C1;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_C2;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_C3;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_C4;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_C5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_C6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_CO5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_CO6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_C_CY;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_C_XOR;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_D;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_D1;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_D2;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_D3;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_D4;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_D5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_D6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_DO5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_DO6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_D_CY;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_D_XOR;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_A;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_A1;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_A2;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_A3;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_A4;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_A5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_A6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_AMUX;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_AO5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_AO6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_A_CY;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_A_XOR;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_B;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_B1;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_B2;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_B3;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_B4;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_B5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_B6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_BO5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_BO6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_B_CY;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_B_XOR;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_C;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_C1;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_C2;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_C3;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_C4;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_C5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_C6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_CMUX;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_CO5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_CO6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_C_CY;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_C_XOR;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_D;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_D1;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_D2;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_D3;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_D4;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_D5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_D6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_DO5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_DO6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_D_CY;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_D_XOR;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_A;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_A1;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_A2;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_A3;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_A4;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_A5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_A6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_AO5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_AO6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_A_CY;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_A_XOR;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_B;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_B1;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_B2;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_B3;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_B4;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_B5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_B6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_BO5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_BO6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_B_CY;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_B_XOR;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_C;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_C1;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_C2;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_C3;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_C4;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_C5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_C6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_CO5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_CO6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_C_CY;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_C_XOR;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_D;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_D1;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_D2;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_D3;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_D4;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_D5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_D6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_DO5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_DO6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_D_CY;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_D_XOR;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_A;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_A1;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_A2;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_A3;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_A4;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_A5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_A6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_AO5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_AO6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_A_CY;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_A_XOR;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_B;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_B1;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_B2;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_B3;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_B4;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_B5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_B6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_BO5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_BO6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_B_CY;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_B_XOR;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_C;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_C1;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_C2;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_C3;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_C4;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_C5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_C6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_CO5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_CO6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_C_CY;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_C_XOR;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_D;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_D1;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_D2;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_D3;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_D4;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_D5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_D6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_DO5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_DO6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_D_CY;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_D_XOR;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_A;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_A1;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_A2;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_A3;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_A4;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_A5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_A6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_AO5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_AO6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_A_CY;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_A_XOR;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_B;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_B1;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_B2;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_B3;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_B4;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_B5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_B6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_BO5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_BO6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_B_CY;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_B_XOR;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_C;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_C1;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_C2;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_C3;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_C4;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_C5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_C6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_CO5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_CO6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_C_CY;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_C_XOR;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_D;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_D1;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_D2;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_D3;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_D4;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_D5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_D6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_DO5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_DO6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_D_CY;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_D_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_AO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_AO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_BO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_BO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_CO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_CO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_DO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_DO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_AO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_AO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_BO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_BO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_CO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_CO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_DO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_DO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D_XOR;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A1;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A2;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A3;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A4;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_AO5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_AO6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A_CY;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A_XOR;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B1;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B2;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B3;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B4;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_BO5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_BO6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B_CY;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B_XOR;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C1;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C2;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C3;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C4;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_CO5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_CO6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C_CY;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C_XOR;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D1;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D2;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D3;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D4;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_DO5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_DO6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D_CY;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D_XOR;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A1;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A2;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A3;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A4;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_AMUX;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_AO5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_AO6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A_CY;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A_XOR;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B1;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B2;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B3;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B4;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_BO5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_BO6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B_CY;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B_XOR;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C1;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C2;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C3;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C4;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_CO5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_CO6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C_CY;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C_XOR;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D1;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D2;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D3;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D4;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_DMUX;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_DO5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_DO6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D_CY;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D_XOR;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A1;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A2;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A3;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A4;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_AMUX;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_AO5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_AO6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A_CY;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A_XOR;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B1;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B2;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B3;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B4;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_BO5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_BO6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B_CY;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B_XOR;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C1;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C2;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C3;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C4;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_CO5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_CO6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C_CY;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C_XOR;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D1;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D2;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D3;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D4;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_DO5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_DO6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D_CY;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D_XOR;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A1;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A2;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A3;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A4;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_AMUX;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_AO5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_AO6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A_CY;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A_XOR;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B1;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B2;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B3;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B4;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_BO5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_BO6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B_CY;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B_XOR;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C1;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C2;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C3;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C4;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_CO5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_CO6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C_CY;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C_XOR;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D1;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D2;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D3;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D4;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_DMUX;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_DO5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_DO6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D_CY;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_AMUX;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_AO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_AO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_BO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_BO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_CO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_CO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_DO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_DO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_AO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_AO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_BO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_BO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_CO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_CO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_DO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_DO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D_XOR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A1;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A2;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A3;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A4;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_AO5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_AO6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A_CY;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A_XOR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B1;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B2;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B3;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B4;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_BO5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_BO6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B_CY;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B_XOR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C1;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C2;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C3;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C4;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_CO5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_CO6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C_CY;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C_XOR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D1;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D2;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D3;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D4;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_DO5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_DO6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D_CY;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D_XOR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A1;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A2;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A3;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A4;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_AMUX;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_AO5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_AO6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A_CY;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A_XOR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B1;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B2;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B3;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B4;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_BO5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_BO6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B_CY;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B_XOR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C1;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C2;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C3;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C4;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_CO5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_CO6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C_CY;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C_XOR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D1;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D2;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D3;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D4;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_DO5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_DO6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D_CY;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D_XOR;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A1;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A2;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A3;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A4;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_AO5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_AO6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A_CY;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A_XOR;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B1;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B2;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B3;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B4;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_BO5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_BO6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B_CY;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B_XOR;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C1;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C2;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C3;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C4;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_CO5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_CO6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C_CY;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C_XOR;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D1;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D2;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D3;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D4;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_DO5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_DO6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D_CY;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D_XOR;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A1;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A2;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A3;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A4;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_AMUX;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_AO5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_AO6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A_CY;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A_XOR;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B1;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B2;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B3;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B4;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_BO5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_BO6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B_CY;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B_XOR;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C1;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C2;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C3;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C4;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_CO5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_CO6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C_CY;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C_XOR;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D1;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D2;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D3;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D4;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_DO5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_DO6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D_CY;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D_XOR;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_A;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_A1;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_A2;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_A3;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_A4;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_A5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_A6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_AO5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_AO6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_A_CY;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_A_XOR;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_B;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_B1;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_B2;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_B3;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_B4;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_B5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_B6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_BO5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_BO6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_B_CY;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_B_XOR;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_C;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_C1;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_C2;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_C3;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_C4;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_C5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_C6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_CO5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_CO6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_C_CY;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_C_XOR;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_D;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_D1;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_D2;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_D3;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_D4;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_D5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_D6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_DO5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_DO6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_D_CY;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_D_XOR;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_A;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_A1;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_A2;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_A3;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_A4;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_A5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_A6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_AO5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_AO6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_A_CY;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_A_XOR;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_B;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_B1;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_B2;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_B3;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_B4;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_B5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_B6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_BO5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_BO6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_B_CY;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_B_XOR;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_C;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_C1;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_C2;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_C3;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_C4;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_C5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_C6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_CO5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_CO6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_C_CY;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_C_XOR;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_D;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_D1;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_D2;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_D3;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_D4;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_D5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_D6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_DO5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_DO6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_D_CY;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_D_XOR;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_A;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_A1;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_A2;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_A3;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_A4;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_A5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_A6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_AO5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_AO6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_A_CY;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_A_XOR;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_B;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_B1;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_B2;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_B3;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_B4;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_B5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_B6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_BO5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_BO6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_B_CY;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_B_XOR;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_C;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_C1;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_C2;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_C3;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_C4;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_C5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_C6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_CO5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_CO6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_C_CY;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_C_XOR;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_D;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_D1;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_D2;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_D3;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_D4;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_D5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_D6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_DO5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_DO6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_D_CY;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_D_XOR;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_A;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_A1;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_A2;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_A3;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_A4;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_A5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_A6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_AO5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_AO6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_A_CY;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_A_XOR;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_B;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_B1;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_B2;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_B3;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_B4;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_B5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_B6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_BO5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_BO6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_B_CY;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_B_XOR;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_C;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_C1;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_C2;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_C3;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_C4;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_C5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_C6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_CMUX;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_CO5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_CO6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_C_CY;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_C_XOR;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_D;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_D1;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_D2;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_D3;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_D4;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_D5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_D6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_DO5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_DO6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_D_CY;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_D_XOR;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_A;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_A1;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_A2;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_A3;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_A4;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_A5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_A6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_AMUX;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_AO5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_AO6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_A_CY;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_A_XOR;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_B;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_B1;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_B2;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_B3;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_B4;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_B5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_B6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_BMUX;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_BO5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_BO6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_B_CY;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_B_XOR;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_C;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_C1;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_C2;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_C3;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_C4;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_C5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_C6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_CMUX;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_CO5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_CO6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_C_CY;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_C_XOR;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_D;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_D1;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_D2;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_D3;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_D4;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_D5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_D6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_DMUX;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_DO5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_DO6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_D_CY;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_D_XOR;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_A;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_A1;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_A2;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_A3;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_A4;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_A5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_A6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_AMUX;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_AO5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_AO6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_A_CY;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_A_XOR;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_B;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_B1;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_B2;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_B3;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_B4;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_B5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_B6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_BO5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_BO6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_B_CY;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_B_XOR;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_C;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_C1;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_C2;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_C3;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_C4;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_C5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_C6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_CO5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_CO6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_C_CY;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_C_XOR;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_D;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_D1;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_D2;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_D3;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_D4;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_D5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_D6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_DO5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_DO6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_D_CY;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_D_XOR;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_A;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_A1;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_A2;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_A3;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_A4;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_A5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_A6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_AO5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_AO6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_A_CY;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_A_XOR;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_B;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_B1;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_B2;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_B3;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_B4;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_B5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_B6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_BO5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_BO6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_B_CY;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_B_XOR;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_C;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_C1;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_C2;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_C3;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_C4;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_C5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_C6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_CO5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_CO6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_C_CY;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_C_XOR;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_D;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_D1;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_D2;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_D3;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_D4;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_D5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_D6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_DO5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_DO6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_D_CY;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_D_XOR;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_A;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_A1;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_A2;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_A3;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_A4;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_A5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_A6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_AMUX;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_AO5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_AO6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_A_CY;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_A_XOR;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_B;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_B1;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_B2;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_B3;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_B4;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_B5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_B6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_BO5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_BO6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_B_CY;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_B_XOR;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_C;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_C1;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_C2;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_C3;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_C4;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_C5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_C6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_CO5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_CO6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_C_CY;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_C_XOR;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_D;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_D1;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_D2;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_D3;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_D4;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_D5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_D6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_DO5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_DO6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_D_CY;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_D_XOR;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_A;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_A1;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_A2;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_A3;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_A4;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_A5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_A6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_AO5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_AO6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_A_CY;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_A_XOR;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_B;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_B1;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_B2;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_B3;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_B4;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_B5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_B6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_BO5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_BO6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_B_CY;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_B_XOR;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_C;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_C1;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_C2;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_C3;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_C4;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_C5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_C6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_CO5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_CO6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_C_CY;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_C_XOR;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_D;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_D1;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_D2;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_D3;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_D4;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_D5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_D6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_DO5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_DO6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_D_CY;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_D_XOR;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_A;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_A1;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_A2;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_A3;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_A4;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_A5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_A6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_AO5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_AO6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_A_CY;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_A_XOR;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_B;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_B1;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_B2;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_B3;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_B4;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_B5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_B6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_BO5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_BO6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_B_CY;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_B_XOR;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_C;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_C1;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_C2;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_C3;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_C4;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_C5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_C6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_CO5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_CO6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_C_CY;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_C_XOR;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_D;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_D1;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_D2;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_D3;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_D4;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_D5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_D6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_DO5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_DO6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_D_CY;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_D_XOR;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A1;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A2;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A3;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A4;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_AMUX;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_AO5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_AO6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A_CY;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A_XOR;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B1;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B2;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B3;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B4;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_BO5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_BO6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B_CY;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B_XOR;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C1;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C2;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C3;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C4;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_CO5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_CO6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C_CY;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C_XOR;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D1;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D2;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D3;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D4;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_DO5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_DO6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D_CY;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D_XOR;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A1;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A2;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A3;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A4;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_AMUX;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_AO5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_AO6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A_CY;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A_XOR;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B1;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B2;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B3;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B4;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_BO5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_BO6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B_CY;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B_XOR;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C1;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C2;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C3;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C4;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_CO5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_CO6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C_CY;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C_XOR;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D1;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D2;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D3;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D4;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_DO5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_DO6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D_CY;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D_XOR;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A1;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A2;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A3;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A4;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_AO5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_AO6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A_CY;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A_XOR;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B1;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B2;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B3;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B4;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_BO5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_BO6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B_CY;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B_XOR;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C1;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C2;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C3;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C4;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_CO5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_CO6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C_CY;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C_XOR;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D1;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D2;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D3;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D4;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_DO5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_DO6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D_CY;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D_XOR;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A1;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A2;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A3;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A4;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_AMUX;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_AO5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_AO6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A_CY;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A_XOR;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B1;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B2;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B3;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B4;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_BMUX;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_BO5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_BO6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B_CY;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B_XOR;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C1;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C2;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C3;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C4;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_CO5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_CO6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C_CY;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C_XOR;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D1;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D2;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D3;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D4;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_DO5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_DO6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D_CY;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D_XOR;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A1;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A2;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A3;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A4;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_AMUX;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_AO5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_AO6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A_CY;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A_XOR;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B1;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B2;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B3;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B4;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_BO5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_BO6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B_CY;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B_XOR;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C1;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C2;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C3;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C4;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_CO5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_CO6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C_CY;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C_XOR;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D1;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D2;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D3;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D4;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_DO5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_DO6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D_CY;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D_XOR;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A1;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A2;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A3;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A4;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_AO5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_AO6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A_CY;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A_XOR;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B1;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B2;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B3;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B4;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_BMUX;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_BO5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_BO6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B_CY;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B_XOR;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C1;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C2;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C3;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C4;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_CO5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_CO6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C_CY;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C_XOR;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D1;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D2;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D3;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D4;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_DO5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_DO6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D_CY;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D_XOR;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A1;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A2;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A3;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A4;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_AMUX;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_AO5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_AO6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A_CY;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A_XOR;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B1;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B2;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B3;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B4;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_BO5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_BO6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B_CY;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B_XOR;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C1;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C2;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C3;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C4;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_CMUX;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_CO5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_CO6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C_CY;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C_XOR;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D1;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D2;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D3;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D4;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_DO5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_DO6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D_CY;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D_XOR;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A1;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A2;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A3;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A4;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_AMUX;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_AO5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_AO6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A_CY;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A_XOR;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B1;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B2;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B3;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B4;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_BO5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_BO6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B_CY;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B_XOR;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C1;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C2;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C3;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C4;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_CO5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_CO6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C_CY;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C_XOR;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D1;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D2;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D3;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D4;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_DO5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_DO6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D_CY;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D_XOR;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A1;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A2;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A3;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A4;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_AO5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_AO6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A_CY;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A_XOR;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B1;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B2;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B3;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B4;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_BO5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_BO6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B_CY;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B_XOR;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C1;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C2;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C3;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C4;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_CO5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_CO6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C_CY;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C_XOR;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D1;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D2;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D3;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D4;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_DO5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_DO6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D_CY;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D_XOR;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A1;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A2;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A3;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A4;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_AO5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_AO6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A_CY;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A_XOR;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B1;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B2;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B3;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B4;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_BO5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_BO6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B_CY;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B_XOR;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C1;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C2;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C3;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C4;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_CO5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_CO6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C_CY;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C_XOR;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D1;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D2;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D3;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D4;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_DO5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_DO6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D_CY;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D_XOR;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_A;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_A1;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_A2;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_A3;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_A4;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_A5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_A6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_AMUX;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_AO5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_AO6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_A_CY;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_A_XOR;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_B;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_B1;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_B2;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_B3;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_B4;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_B5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_B6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_BO5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_BO6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_B_CY;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_B_XOR;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_C;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_C1;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_C2;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_C3;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_C4;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_C5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_C6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_CO5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_CO6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_C_CY;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_C_XOR;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_D;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_D1;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_D2;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_D3;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_D4;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_D5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_D6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_DO5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_DO6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_D_CY;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_D_XOR;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_A;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_A1;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_A2;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_A3;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_A4;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_A5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_A6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_AO5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_AO6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_A_CY;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_A_XOR;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_B;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_B1;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_B2;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_B3;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_B4;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_B5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_B6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_BO5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_BO6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_B_CY;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_B_XOR;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_C;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_C1;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_C2;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_C3;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_C4;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_C5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_C6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_CO5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_CO6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_C_CY;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_C_XOR;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_D;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_D1;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_D2;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_D3;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_D4;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_D5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_D6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_DO5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_DO6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_D_CY;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_D_XOR;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A1;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A2;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A3;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A4;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_AMUX;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_AO5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_AO6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A_CY;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A_XOR;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B1;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B2;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B3;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B4;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_BO5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_BO6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B_CY;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B_XOR;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C1;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C2;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C3;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C4;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_CO5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_CO6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C_CY;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C_XOR;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D1;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D2;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D3;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D4;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_DO5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_DO6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D_CY;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D_XOR;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A1;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A2;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A3;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A4;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_AMUX;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_AO5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_AO6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A_CY;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A_XOR;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B1;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B2;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B3;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B4;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_BO5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_BO6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B_CY;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B_XOR;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C1;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C2;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C3;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C4;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_CO5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_CO6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C_CY;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C_XOR;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D1;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D2;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D3;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D4;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_DO5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_DO6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D_CY;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D_XOR;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A1;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A2;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A3;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A4;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_AMUX;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_AO5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_AO6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A_CY;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A_XOR;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B1;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B2;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B3;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B4;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_BO5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_BO6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B_CY;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B_XOR;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C1;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C2;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C3;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C4;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_CO5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_CO6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C_CY;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C_XOR;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D1;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D2;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D3;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D4;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_DO5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_DO6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D_CY;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D_XOR;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A1;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A2;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A3;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A4;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_AMUX;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_AO5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_AO6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A_CY;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A_XOR;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B1;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B2;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B3;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B4;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_BMUX;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_BO5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_BO6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B_CY;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B_XOR;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C1;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C2;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C3;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C4;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_CO5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_CO6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C_CY;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C_XOR;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D1;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D2;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D3;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D4;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_DO5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D_CY;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D_XOR;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_A;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_A1;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_A2;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_A3;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_A4;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_A5;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_A6;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_AO5;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_AO6;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_A_CY;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_A_XOR;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_B;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_B1;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_B2;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_B3;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_B4;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_B5;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_B6;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_BO5;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_BO6;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_B_CY;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_B_XOR;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_C;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_C1;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_C2;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_C3;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_C4;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_C5;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_C6;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_CO5;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_CO6;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_C_CY;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_C_XOR;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_D;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_D1;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_D2;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_D3;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_D4;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_D5;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_D6;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_DO5;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_DO6;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_D_CY;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_D_XOR;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_A;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_A1;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_A2;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_A3;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_A4;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_A5;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_A6;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_AMUX;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_AO5;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_AO6;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_A_CY;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_A_XOR;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_B;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_B1;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_B2;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_B3;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_B4;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_B5;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_B6;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_BO5;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_BO6;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_B_CY;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_B_XOR;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_C;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_C1;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_C2;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_C3;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_C4;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_C5;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_C6;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_CMUX;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_CO5;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_CO6;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_C_CY;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_C_XOR;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_D;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_D1;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_D2;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_D3;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_D4;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_D5;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_D6;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_DO5;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_DO6;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_D_CY;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_D_XOR;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_A;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_A1;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_A2;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_A3;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_A4;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_A5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_A6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_AMUX;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_AO5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_AO6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_A_CY;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_A_XOR;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_B;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_B1;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_B2;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_B3;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_B4;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_B5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_B6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_BMUX;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_BO5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_BO6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_B_CY;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_B_XOR;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_C;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_C1;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_C2;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_C3;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_C4;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_C5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_C6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_CO5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_CO6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_C_CY;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_C_XOR;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_D;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_D1;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_D2;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_D3;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_D4;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_D5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_D6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_DO5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_DO6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_D_CY;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_D_XOR;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_A;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_A1;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_A2;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_A3;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_A4;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_A5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_A6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_AO5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_AO6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_A_CY;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_A_XOR;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_B;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_B1;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_B2;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_B3;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_B4;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_B5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_B6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_BO5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_BO6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_B_CY;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_B_XOR;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_C;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_C1;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_C2;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_C3;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_C4;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_C5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_C6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_CO5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_CO6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_C_CY;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_C_XOR;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_D;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_D1;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_D2;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_D3;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_D4;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_D5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_D6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_DO5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_DO6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_D_CY;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_D_XOR;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_A;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_A1;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_A2;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_A3;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_A4;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_A5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_A6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_AMUX;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_AO5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_AO6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_A_CY;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_A_XOR;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_B;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_B1;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_B2;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_B3;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_B4;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_B5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_B6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_BMUX;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_BO5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_BO6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_B_CY;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_B_XOR;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_C;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_C1;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_C2;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_C3;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_C4;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_C5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_C6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_CMUX;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_CO5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_CO6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_C_CY;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_C_XOR;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_D;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_D1;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_D2;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_D3;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_D4;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_D5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_D6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_DO5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_DO6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_D_CY;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_D_XOR;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_A;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_A1;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_A2;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_A3;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_A4;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_A5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_A6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_AMUX;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_AO5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_AO6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_A_CY;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_A_XOR;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_B;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_B1;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_B2;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_B3;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_B4;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_B5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_B6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_BO5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_BO6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_B_CY;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_B_XOR;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_C;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_C1;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_C2;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_C3;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_C4;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_C5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_C6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_CO5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_CO6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_C_CY;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_C_XOR;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_D;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_D1;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_D2;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_D3;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_D4;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_D5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_D6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_DO5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_DO6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_D_CY;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_D_XOR;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_A;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_A1;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_A2;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_A3;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_A4;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_A5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_A6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_AO5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_AO6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_A_CY;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_A_XOR;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_B;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_B1;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_B2;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_B3;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_B4;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_B5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_B6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_BO5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_BO6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_B_CY;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_B_XOR;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_C;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_C1;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_C2;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_C3;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_C4;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_C5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_C6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_CO5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_CO6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_C_CY;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_C_XOR;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_D;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_D1;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_D2;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_D3;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_D4;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_D5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_D6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_DO5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_DO6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_D_CY;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_D_XOR;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_A;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_A1;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_A2;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_A3;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_A4;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_A5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_A6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_AO5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_AO6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_A_CY;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_A_XOR;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_B;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_B1;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_B2;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_B3;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_B4;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_B5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_B6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_BO5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_BO6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_B_CY;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_B_XOR;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_C;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_C1;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_C2;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_C3;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_C4;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_C5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_C6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_CO5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_CO6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_C_CY;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_C_XOR;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_D;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_D1;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_D2;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_D3;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_D4;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_D5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_D6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_DO5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_DO6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_D_CY;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_D_XOR;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_A;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_A1;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_A2;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_A3;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_A4;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_A5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_A6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_AMUX;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_AO5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_AO6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_A_CY;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_A_XOR;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_B;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_B1;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_B2;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_B3;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_B4;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_B5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_B6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_BO5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_BO6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_B_CY;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_B_XOR;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_C;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_C1;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_C2;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_C3;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_C4;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_C5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_C6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_CO5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_CO6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_C_CY;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_C_XOR;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_D;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_D1;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_D2;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_D3;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_D4;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_D5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_D6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_DO5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_DO6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_D_CY;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_D_XOR;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_A;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_A1;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_A2;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_A3;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_A4;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_A5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_A6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_AMUX;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_AO5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_AO6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_A_CY;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_A_XOR;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_B;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_B1;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_B2;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_B3;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_B4;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_B5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_B6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_BO5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_BO6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_B_CY;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_B_XOR;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_C;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_C1;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_C2;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_C3;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_C4;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_C5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_C6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_CO5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_CO6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_C_CY;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_C_XOR;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_D;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_D1;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_D2;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_D3;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_D4;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_D5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_D6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_DO5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_DO6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_D_CY;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_D_XOR;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A1;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A2;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A3;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A4;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_AMUX;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_AO5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_AO6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A_CY;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A_XOR;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B1;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B2;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B3;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B4;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_BO5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_BO6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B_CY;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B_XOR;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C1;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C2;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C3;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C4;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_CO5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_CO6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C_CY;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C_XOR;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D1;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D2;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D3;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D4;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_DO5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_DO6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D_CY;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D_XOR;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A1;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A2;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A3;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A4;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_AMUX;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_AO5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_AO6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A_CY;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A_XOR;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B1;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B2;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B3;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B4;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_BMUX;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_BO5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_BO6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B_CY;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B_XOR;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C1;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C2;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C3;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C4;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_CO5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_CO6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C_CY;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C_XOR;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D1;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D2;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D3;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D4;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_DO5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_DO6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D_CY;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D_XOR;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A1;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A2;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A3;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A4;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_AO5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_AO6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A_CY;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A_XOR;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B1;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B2;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B3;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B4;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_BO5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_BO6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B_CY;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B_XOR;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C1;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C2;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C3;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C4;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_CO5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_CO6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C_CY;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C_XOR;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D1;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D2;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D3;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D4;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_DO5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_DO6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D_CY;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D_XOR;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A1;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A2;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A3;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A4;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_AMUX;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_AO5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_AO6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A_CY;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A_XOR;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B1;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B2;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B3;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B4;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_BMUX;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_BO5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_BO6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B_CY;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B_XOR;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C1;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C2;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C3;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C4;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_CO5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_CO6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C_CY;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C_XOR;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D1;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D2;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D3;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D4;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_DO5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_DO6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D_CY;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D_XOR;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A1;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A2;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A3;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A4;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_AMUX;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_AO5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_AO6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A_CY;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A_XOR;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B1;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B2;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B3;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B4;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_BO5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_BO6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B_CY;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B_XOR;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C1;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C2;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C3;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C4;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_CO5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_CO6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C_CY;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C_XOR;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D1;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D2;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D3;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D4;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_DO5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_DO6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D_CY;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D_XOR;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A1;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A2;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A3;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A4;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_AO5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_AO6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A_CY;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A_XOR;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B1;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B2;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B3;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B4;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_BO5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_BO6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B_CY;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B_XOR;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C1;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C2;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C3;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C4;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_CO5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_CO6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C_CY;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C_XOR;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D1;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D2;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D3;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D4;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_DO5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_DO6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D_CY;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D_XOR;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A1;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A2;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A3;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A4;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_AO5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_AO6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A_CY;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A_XOR;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B1;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B2;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B3;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B4;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_BO5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_BO6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B_CY;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B_XOR;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C1;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C2;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C3;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C4;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_CO5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_CO6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C_CY;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C_XOR;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D1;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D2;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D3;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D4;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_DO5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_DO6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D_CY;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D_XOR;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A1;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A2;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A3;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A4;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_AMUX;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_AO5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_AO6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A_CY;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A_XOR;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B1;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B2;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B3;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B4;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_BMUX;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_BO5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_BO6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B_CY;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B_XOR;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C1;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C2;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C3;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C4;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_CO5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_CO6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C_CY;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C_XOR;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D1;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D2;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D3;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D4;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_DO5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_DO6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D_CY;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D_XOR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A1;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A2;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A3;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A4;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_AO5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_AO6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A_CY;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A_XOR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B1;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B2;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B3;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B4;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_BO5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_BO6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B_CY;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B_XOR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C1;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C2;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C3;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C4;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_CO5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_CO6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C_CY;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C_XOR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D1;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D2;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D3;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D4;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_DO5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_DO6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D_CY;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D_XOR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A1;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A2;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A3;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A4;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_AO5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_AO6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A_CY;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A_XOR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B1;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B2;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B3;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B4;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_BO5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_BO6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B_CY;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B_XOR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C1;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C2;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C3;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C4;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_CO5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_CO6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C_CY;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C_XOR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D1;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D2;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D3;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D4;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_DO5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_DO6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D_CY;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D_XOR;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A1;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A2;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A3;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A4;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_AMUX;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_AO5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_AO6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A_CY;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A_XOR;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B1;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B2;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B3;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B4;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_BO5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_BO6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B_CY;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B_XOR;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C1;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C2;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C3;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C4;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_CO5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_CO6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C_CY;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C_XOR;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D1;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D2;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D3;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D4;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_DO5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_DO6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D_CY;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D_XOR;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A1;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A2;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A3;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A4;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_AMUX;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_AO5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_AO6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A_CY;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A_XOR;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B1;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B2;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B3;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B4;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_BO5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_BO6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B_CY;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B_XOR;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C1;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C2;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C3;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C4;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_CO5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_CO6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C_CY;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C_XOR;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D1;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D2;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D3;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D4;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_DO5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_DO6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D_CY;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D_XOR;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A1;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A2;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A3;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A4;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_AO5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_AO6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A_CY;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A_XOR;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B1;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B2;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B3;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B4;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_BO5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_BO6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B_CY;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B_XOR;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C1;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C2;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C3;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C4;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_CO5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_CO6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C_CY;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C_XOR;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D1;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D2;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D3;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D4;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_DO5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_DO6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D_CY;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D_XOR;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A1;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A2;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A3;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A4;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_AO5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_AO6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A_CY;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A_XOR;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B1;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B2;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B3;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B4;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_BO5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_BO6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B_CY;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B_XOR;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C1;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C2;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C3;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C4;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_CO5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_CO6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C_CY;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C_XOR;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D1;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D2;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D3;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D4;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_DO5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_DO6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D_CY;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D_XOR;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_A;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_A1;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_A2;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_A3;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_A4;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_A5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_A6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_AO5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_AO6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_A_CY;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_A_XOR;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_B;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_B1;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_B2;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_B3;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_B4;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_B5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_B6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_BO5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_BO6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_B_CY;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_B_XOR;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_C;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_C1;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_C2;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_C3;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_C4;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_C5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_C6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_CO5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_CO6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_C_CY;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_C_XOR;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_D;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_D1;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_D2;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_D3;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_D4;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_D5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_D6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_DO5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_DO6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_D_CY;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_D_XOR;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_A;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_A1;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_A2;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_A3;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_A4;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_A5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_A6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_AO5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_AO6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_A_CY;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_A_XOR;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_B;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_B1;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_B2;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_B3;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_B4;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_B5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_B6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_BO5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_BO6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_B_CY;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_B_XOR;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_C;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_C1;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_C2;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_C3;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_C4;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_C5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_C6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_CO5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_CO6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_C_CY;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_C_XOR;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_D;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_D1;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_D2;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_D3;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_D4;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_D5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_D6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_DO5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_DO6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_D_CY;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_D_XOR;
  wire [0:0] LIOB33_SING_X0Y100_IOB_X0Y100_I;
  wire [0:0] LIOB33_SING_X0Y149_IOB_X0Y149_O;
  wire [0:0] LIOB33_X0Y101_IOB_X0Y101_I;
  wire [0:0] LIOB33_X0Y101_IOB_X0Y102_I;
  wire [0:0] LIOB33_X0Y103_IOB_X0Y103_I;
  wire [0:0] LIOB33_X0Y103_IOB_X0Y104_I;
  wire [0:0] LIOB33_X0Y105_IOB_X0Y105_I;
  wire [0:0] LIOB33_X0Y105_IOB_X0Y106_I;
  wire [0:0] LIOB33_X0Y107_IOB_X0Y107_I;
  wire [0:0] LIOB33_X0Y107_IOB_X0Y108_I;
  wire [0:0] LIOB33_X0Y109_IOB_X0Y109_I;
  wire [0:0] LIOB33_X0Y109_IOB_X0Y110_I;
  wire [0:0] LIOB33_X0Y111_IOB_X0Y111_I;
  wire [0:0] LIOB33_X0Y111_IOB_X0Y112_I;
  wire [0:0] LIOB33_X0Y113_IOB_X0Y113_I;
  wire [0:0] LIOB33_X0Y113_IOB_X0Y114_I;
  wire [0:0] LIOB33_X0Y115_IOB_X0Y115_I;
  wire [0:0] LIOB33_X0Y115_IOB_X0Y116_I;
  wire [0:0] LIOB33_X0Y117_IOB_X0Y117_I;
  wire [0:0] LIOB33_X0Y117_IOB_X0Y118_O;
  wire [0:0] LIOB33_X0Y119_IOB_X0Y119_O;
  wire [0:0] LIOB33_X0Y119_IOB_X0Y120_O;
  wire [0:0] LIOB33_X0Y121_IOB_X0Y121_O;
  wire [0:0] LIOB33_X0Y121_IOB_X0Y122_O;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y123_O;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y124_O;
  wire [0:0] LIOB33_X0Y125_IOB_X0Y125_O;
  wire [0:0] LIOB33_X0Y125_IOB_X0Y126_O;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y127_O;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y128_O;
  wire [0:0] LIOB33_X0Y129_IOB_X0Y129_O;
  wire [0:0] LIOB33_X0Y129_IOB_X0Y130_O;
  wire [0:0] LIOB33_X0Y131_IOB_X0Y131_O;
  wire [0:0] LIOB33_X0Y131_IOB_X0Y132_O;
  wire [0:0] LIOB33_X0Y133_IOB_X0Y133_O;
  wire [0:0] LIOB33_X0Y133_IOB_X0Y134_O;
  wire [0:0] LIOB33_X0Y135_IOB_X0Y135_O;
  wire [0:0] LIOB33_X0Y135_IOB_X0Y136_O;
  wire [0:0] LIOB33_X0Y137_IOB_X0Y137_O;
  wire [0:0] LIOB33_X0Y137_IOB_X0Y138_O;
  wire [0:0] LIOB33_X0Y139_IOB_X0Y139_O;
  wire [0:0] LIOB33_X0Y139_IOB_X0Y140_O;
  wire [0:0] LIOB33_X0Y141_IOB_X0Y141_O;
  wire [0:0] LIOB33_X0Y141_IOB_X0Y142_O;
  wire [0:0] LIOB33_X0Y143_IOB_X0Y143_O;
  wire [0:0] LIOB33_X0Y145_IOB_X0Y145_O;
  wire [0:0] LIOB33_X0Y145_IOB_X0Y146_O;
  wire [0:0] LIOB33_X0Y147_IOB_X0Y147_O;
  wire [0:0] LIOB33_X0Y147_IOB_X0Y148_O;
  wire [0:0] LIOI3_SING_X0Y100_ILOGIC_X0Y100_D;
  wire [0:0] LIOI3_SING_X0Y100_ILOGIC_X0Y100_O;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_D1;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_OQ;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_T1;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y107_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y107_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y108_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y108_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y113_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y113_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y114_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y114_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_TQ;
  wire [0:0] LIOI3_X0Y101_ILOGIC_X0Y101_D;
  wire [0:0] LIOI3_X0Y101_ILOGIC_X0Y101_O;
  wire [0:0] LIOI3_X0Y101_ILOGIC_X0Y102_D;
  wire [0:0] LIOI3_X0Y101_ILOGIC_X0Y102_O;
  wire [0:0] LIOI3_X0Y103_ILOGIC_X0Y103_D;
  wire [0:0] LIOI3_X0Y103_ILOGIC_X0Y103_O;
  wire [0:0] LIOI3_X0Y103_ILOGIC_X0Y104_D;
  wire [0:0] LIOI3_X0Y103_ILOGIC_X0Y104_O;
  wire [0:0] LIOI3_X0Y105_ILOGIC_X0Y105_D;
  wire [0:0] LIOI3_X0Y105_ILOGIC_X0Y105_O;
  wire [0:0] LIOI3_X0Y105_ILOGIC_X0Y106_D;
  wire [0:0] LIOI3_X0Y105_ILOGIC_X0Y106_O;
  wire [0:0] LIOI3_X0Y109_ILOGIC_X0Y109_D;
  wire [0:0] LIOI3_X0Y109_ILOGIC_X0Y109_O;
  wire [0:0] LIOI3_X0Y109_ILOGIC_X0Y110_D;
  wire [0:0] LIOI3_X0Y109_ILOGIC_X0Y110_O;
  wire [0:0] LIOI3_X0Y111_ILOGIC_X0Y111_D;
  wire [0:0] LIOI3_X0Y111_ILOGIC_X0Y111_O;
  wire [0:0] LIOI3_X0Y111_ILOGIC_X0Y112_D;
  wire [0:0] LIOI3_X0Y111_ILOGIC_X0Y112_O;
  wire [0:0] LIOI3_X0Y115_ILOGIC_X0Y115_D;
  wire [0:0] LIOI3_X0Y115_ILOGIC_X0Y115_O;
  wire [0:0] LIOI3_X0Y115_ILOGIC_X0Y116_D;
  wire [0:0] LIOI3_X0Y115_ILOGIC_X0Y116_O;
  wire [0:0] LIOI3_X0Y117_ILOGIC_X0Y117_D;
  wire [0:0] LIOI3_X0Y117_ILOGIC_X0Y117_O;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_D1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_OQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_T1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_TQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_D1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_OQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_T1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_TQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_D1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_OQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_T1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_TQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_D1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_OQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_T1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_TQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_D1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_OQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_T1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_TQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_D1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_OQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_T1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_TQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_D1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_OQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_T1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_TQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_D1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_OQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_T1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_TQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_D1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_OQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_T1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_TQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_D1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_OQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_T1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_TQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_D1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_OQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_T1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_TQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_D1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_OQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_T1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_TQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_D1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_OQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_T1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_TQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_D1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_OQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_T1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_TQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_D1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_OQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_T1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_TQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_D1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_OQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_T1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_TQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_D1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_OQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_T1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_TQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_D1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_OQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_T1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_TQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_D1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_OQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_T1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_TQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_D1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_OQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_T1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_TQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_D1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_OQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_T1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_TQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_D1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_OQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_T1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_TQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_D1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_OQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_T1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_TQ;
  wire [0:0] RIOB33_SING_X105Y100_IOB_X1Y100_I;
  wire [0:0] RIOB33_X105Y101_IOB_X1Y101_I;
  wire [0:0] RIOB33_X105Y101_IOB_X1Y102_I;
  wire [0:0] RIOB33_X105Y103_IOB_X1Y103_I;
  wire [0:0] RIOB33_X105Y103_IOB_X1Y104_I;
  wire [0:0] RIOB33_X105Y105_IOB_X1Y105_I;
  wire [0:0] RIOB33_X105Y105_IOB_X1Y106_I;
  wire [0:0] RIOB33_X105Y107_IOB_X1Y107_I;
  wire [0:0] RIOB33_X105Y107_IOB_X1Y108_I;
  wire [0:0] RIOB33_X105Y109_IOB_X1Y109_I;
  wire [0:0] RIOB33_X105Y109_IOB_X1Y110_I;
  wire [0:0] RIOB33_X105Y111_IOB_X1Y111_I;
  wire [0:0] RIOB33_X105Y111_IOB_X1Y112_I;
  wire [0:0] RIOB33_X105Y113_IOB_X1Y113_I;
  wire [0:0] RIOI3_SING_X105Y100_ILOGIC_X1Y100_D;
  wire [0:0] RIOI3_SING_X105Y100_ILOGIC_X1Y100_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_O;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y101_D;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y101_O;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y102_D;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y102_O;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y103_D;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y103_O;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y104_D;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y104_O;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y105_D;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y105_O;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y106_D;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y106_O;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y109_D;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y109_O;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y110_D;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y110_O;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y111_D;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y111_O;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y112_D;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y112_O;


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h4b5ab4a5b4a54b5a)
  ) CLBLL_L_X2Y106_SLICE_X0Y106_DLUT (
.I0(CLBLL_L_X2Y106_SLICE_X1Y106_CO6),
.I1(CLBLL_L_X2Y106_SLICE_X1Y106_AO6),
.I2(CLBLM_R_X3Y105_SLICE_X2Y105_AO6),
.I3(CLBLL_L_X2Y107_SLICE_X0Y107_AO6),
.I4(CLBLL_L_X2Y106_SLICE_X0Y106_BO5),
.I5(CLBLM_R_X3Y104_SLICE_X3Y104_AO5),
.O5(CLBLL_L_X2Y106_SLICE_X0Y106_DO5),
.O6(CLBLL_L_X2Y106_SLICE_X0Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbbfb00bfaafa00a)
  ) CLBLL_L_X2Y106_SLICE_X0Y106_CLUT (
.I0(CLBLL_L_X2Y106_SLICE_X1Y106_CO6),
.I1(CLBLL_L_X2Y106_SLICE_X1Y106_AO6),
.I2(CLBLM_R_X3Y105_SLICE_X2Y105_AO6),
.I3(CLBLM_R_X3Y104_SLICE_X3Y104_AO5),
.I4(CLBLL_L_X2Y106_SLICE_X0Y106_BO5),
.I5(CLBLL_L_X2Y107_SLICE_X0Y107_AO6),
.O5(CLBLL_L_X2Y106_SLICE_X0Y106_CO5),
.O6(CLBLL_L_X2Y106_SLICE_X0Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h777777773f3f3f3f)
  ) CLBLL_L_X2Y106_SLICE_X0Y106_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y106_I),
.I1(LIOB33_X0Y101_IOB_X0Y102_I),
.I2(LIOB33_X0Y103_IOB_X0Y103_I),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y106_SLICE_X0Y106_BO5),
.O6(CLBLL_L_X2Y106_SLICE_X0Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc3c30f0fababafaf)
  ) CLBLL_L_X2Y106_SLICE_X0Y106_ALUT (
.I0(CLBLL_L_X2Y106_SLICE_X1Y106_CO6),
.I1(LIOB33_X0Y101_IOB_X0Y101_I),
.I2(CLBLL_L_X2Y106_SLICE_X1Y106_AO6),
.I3(1'b1),
.I4(LIOB33_X0Y103_IOB_X0Y103_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y106_SLICE_X0Y106_AO5),
.O6(CLBLL_L_X2Y106_SLICE_X0Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6696969999696966)
  ) CLBLL_L_X2Y106_SLICE_X1Y106_DLUT (
.I0(CLBLM_R_X3Y104_SLICE_X3Y104_DO6),
.I1(CLBLL_L_X2Y106_SLICE_X0Y106_CO6),
.I2(CLBLL_L_X2Y106_SLICE_X0Y106_DO6),
.I3(CLBLL_L_X2Y108_SLICE_X1Y108_AO5),
.I4(CLBLL_L_X2Y107_SLICE_X0Y107_DO6),
.I5(CLBLM_R_X3Y105_SLICE_X3Y105_BO6),
.O5(CLBLL_L_X2Y106_SLICE_X1Y106_DO5),
.O6(CLBLL_L_X2Y106_SLICE_X1Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3444550033440000)
  ) CLBLL_L_X2Y106_SLICE_X1Y106_CLUT (
.I0(LIOB33_X0Y103_IOB_X0Y103_I),
.I1(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I2(RIOB33_X105Y111_IOB_X1Y112_I),
.I3(RIOB33_X105Y113_IOB_X1Y113_I),
.I4(LIOB33_X0Y113_IOB_X0Y114_I),
.I5(LIOB33_X0Y115_IOB_X0Y116_I),
.O5(CLBLL_L_X2Y106_SLICE_X1Y106_CO5),
.O6(CLBLL_L_X2Y106_SLICE_X1Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5aaa5aaaa5559a6a)
  ) CLBLL_L_X2Y106_SLICE_X1Y106_BLUT (
.I0(CLBLM_R_X3Y105_SLICE_X2Y105_AO6),
.I1(LIOB33_X0Y103_IOB_X0Y103_I),
.I2(LIOB33_X0Y101_IOB_X0Y101_I),
.I3(LIOB33_X0Y113_IOB_X0Y114_I),
.I4(CLBLL_L_X2Y106_SLICE_X1Y106_AO6),
.I5(CLBLL_L_X2Y106_SLICE_X1Y106_CO6),
.O5(CLBLL_L_X2Y106_SLICE_X1Y106_BO5),
.O6(CLBLL_L_X2Y106_SLICE_X1Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h074388cc3cf00cc0)
  ) CLBLL_L_X2Y106_SLICE_X1Y106_ALUT (
.I0(RIOB33_X105Y111_IOB_X1Y112_I),
.I1(RIOB33_X105Y113_IOB_X1Y113_I),
.I2(LIOB33_X0Y103_IOB_X0Y103_I),
.I3(LIOB33_X0Y115_IOB_X0Y116_I),
.I4(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I5(LIOB33_X0Y113_IOB_X0Y114_I),
.O5(CLBLL_L_X2Y106_SLICE_X1Y106_AO5),
.O6(CLBLL_L_X2Y106_SLICE_X1Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf9f9f9f990f99090)
  ) CLBLL_L_X2Y107_SLICE_X0Y107_DLUT (
.I0(CLBLL_L_X2Y107_SLICE_X0Y107_AO6),
.I1(CLBLL_L_X2Y106_SLICE_X1Y106_AO6),
.I2(CLBLL_L_X2Y106_SLICE_X0Y106_BO6),
.I3(CLBLL_L_X2Y110_SLICE_X0Y110_AO6),
.I4(CLBLL_L_X2Y107_SLICE_X0Y107_AO5),
.I5(CLBLL_L_X2Y107_SLICE_X0Y107_BO6),
.O5(CLBLL_L_X2Y107_SLICE_X0Y107_DO5),
.O6(CLBLL_L_X2Y107_SLICE_X0Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hda705df7258fa208)
  ) CLBLL_L_X2Y107_SLICE_X0Y107_CLUT (
.I0(LIOB33_X0Y101_IOB_X0Y102_I),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(CLBLL_L_X2Y108_SLICE_X1Y108_BO5),
.I3(LIOB33_X0Y103_IOB_X0Y103_I),
.I4(CLBLL_L_X2Y106_SLICE_X0Y106_AO6),
.I5(CLBLL_L_X2Y106_SLICE_X1Y106_BO6),
.O5(CLBLL_L_X2Y107_SLICE_X0Y107_CO5),
.O6(CLBLL_L_X2Y107_SLICE_X0Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h087800cc0c3c0000)
  ) CLBLL_L_X2Y107_SLICE_X0Y107_BLUT (
.I0(RIOB33_X105Y111_IOB_X1Y112_I),
.I1(RIOB33_X105Y113_IOB_X1Y113_I),
.I2(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I3(RIOB33_X105Y105_IOB_X1Y106_I),
.I4(LIOB33_X0Y103_IOB_X0Y103_I),
.I5(LIOB33_X0Y113_IOB_X0Y114_I),
.O5(CLBLL_L_X2Y107_SLICE_X0Y107_BO5),
.O6(CLBLL_L_X2Y107_SLICE_X0Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333ffff00ffffff)
  ) CLBLL_L_X2Y107_SLICE_X0Y107_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y103_IOB_X0Y103_I),
.I2(1'b1),
.I3(RIOB33_X105Y105_IOB_X1Y106_I),
.I4(LIOB33_X0Y101_IOB_X0Y101_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y107_SLICE_X0Y107_AO5),
.O6(CLBLL_L_X2Y107_SLICE_X0Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y107_SLICE_X1Y107_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y107_SLICE_X1Y107_DO5),
.O6(CLBLL_L_X2Y107_SLICE_X1Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h71d4f3fcd4d4fcfc)
  ) CLBLL_L_X2Y107_SLICE_X1Y107_CLUT (
.I0(LIOB33_X0Y105_IOB_X0Y105_I),
.I1(CLBLL_L_X2Y107_SLICE_X0Y107_CO6),
.I2(CLBLL_L_X2Y108_SLICE_X1Y108_DO6),
.I3(RIOB33_X105Y105_IOB_X1Y106_I),
.I4(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I5(LIOB33_X0Y103_IOB_X0Y104_I),
.O5(CLBLL_L_X2Y107_SLICE_X1Y107_CO5),
.O6(CLBLL_L_X2Y107_SLICE_X1Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3ccc2fdfc333d020)
  ) CLBLL_L_X2Y107_SLICE_X1Y107_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y106_I),
.I1(CLBLL_L_X2Y107_SLICE_X0Y107_BO6),
.I2(LIOB33_X0Y101_IOB_X0Y101_I),
.I3(LIOB33_X0Y103_IOB_X0Y103_I),
.I4(CLBLL_L_X2Y110_SLICE_X0Y110_AO6),
.I5(CLBLL_L_X2Y106_SLICE_X1Y106_AO6),
.O5(CLBLL_L_X2Y107_SLICE_X1Y107_BO5),
.O6(CLBLL_L_X2Y107_SLICE_X1Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h33ff33ff66aa9955)
  ) CLBLL_L_X2Y107_SLICE_X1Y107_ALUT (
.I0(CLBLM_R_X3Y107_SLICE_X2Y107_BO6),
.I1(LIOB33_X0Y105_IOB_X0Y106_I),
.I2(1'b1),
.I3(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I4(CLBLL_L_X2Y107_SLICE_X1Y107_CO6),
.I5(1'b1),
.O5(CLBLL_L_X2Y107_SLICE_X1Y107_AO5),
.O6(CLBLL_L_X2Y107_SLICE_X1Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfaf5a050faf5e8d4)
  ) CLBLL_L_X2Y108_SLICE_X0Y108_DLUT (
.I0(CLBLL_L_X2Y110_SLICE_X0Y110_AO6),
.I1(CLBLL_L_X2Y109_SLICE_X0Y109_BO6),
.I2(CLBLL_L_X2Y108_SLICE_X0Y108_AO6),
.I3(CLBLL_L_X2Y107_SLICE_X0Y107_AO5),
.I4(CLBLL_L_X2Y109_SLICE_X0Y109_DO6),
.I5(CLBLL_L_X2Y109_SLICE_X0Y109_CO6),
.O5(CLBLL_L_X2Y108_SLICE_X0Y108_DO5),
.O6(CLBLL_L_X2Y108_SLICE_X0Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996c33ca55a0ff0)
  ) CLBLL_L_X2Y108_SLICE_X0Y108_CLUT (
.I0(LIOB33_X0Y105_IOB_X0Y105_I),
.I1(LIOB33_X0Y103_IOB_X0Y104_I),
.I2(CLBLL_L_X2Y108_SLICE_X1Y108_DO6),
.I3(CLBLL_L_X2Y107_SLICE_X0Y107_CO6),
.I4(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I5(RIOB33_X105Y105_IOB_X1Y106_I),
.O5(CLBLL_L_X2Y108_SLICE_X0Y108_CO5),
.O6(CLBLL_L_X2Y108_SLICE_X0Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6978a5b4693ca5f0)
  ) CLBLL_L_X2Y108_SLICE_X0Y108_BLUT (
.I0(CLBLL_L_X2Y109_SLICE_X0Y109_DO6),
.I1(LIOB33_X0Y101_IOB_X0Y101_I),
.I2(CLBLL_L_X2Y110_SLICE_X0Y110_AO6),
.I3(CLBLL_L_X2Y109_SLICE_X0Y109_CO6),
.I4(RIOB33_X105Y105_IOB_X1Y106_I),
.I5(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.O5(CLBLL_L_X2Y108_SLICE_X0Y108_BO5),
.O6(CLBLL_L_X2Y108_SLICE_X0Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h7777777788778877)
  ) CLBLL_L_X2Y108_SLICE_X0Y108_ALUT (
.I0(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I1(LIOB33_X0Y101_IOB_X0Y102_I),
.I2(1'b1),
.I3(CLBLL_L_X2Y108_SLICE_X0Y108_BO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y108_SLICE_X0Y108_AO5),
.O6(CLBLL_L_X2Y108_SLICE_X0Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h71f5b2faf3ff30f0)
  ) CLBLL_L_X2Y108_SLICE_X1Y108_DLUT (
.I0(LIOB33_X0Y101_IOB_X0Y102_I),
.I1(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I2(CLBLL_L_X2Y108_SLICE_X0Y108_DO6),
.I3(LIOB33_X0Y103_IOB_X0Y104_I),
.I4(CLBLL_L_X2Y107_SLICE_X1Y107_BO6),
.I5(RIOB33_X105Y105_IOB_X1Y106_I),
.O5(CLBLL_L_X2Y108_SLICE_X1Y108_DO5),
.O6(CLBLL_L_X2Y108_SLICE_X1Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hc639aa55639cff00)
  ) CLBLL_L_X2Y108_SLICE_X1Y108_CLUT (
.I0(CLBLL_L_X2Y109_SLICE_X0Y109_AO6),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I3(CLBLL_L_X2Y107_SLICE_X1Y107_BO6),
.I4(LIOB33_X0Y101_IOB_X0Y102_I),
.I5(CLBLL_L_X2Y108_SLICE_X1Y108_BO6),
.O5(CLBLL_L_X2Y108_SLICE_X1Y108_CO5),
.O6(CLBLL_L_X2Y108_SLICE_X1Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc0033fff0f0f3ff)
  ) CLBLL_L_X2Y108_SLICE_X1Y108_BLUT (
.I0(1'b1),
.I1(LIOB33_X0Y101_IOB_X0Y101_I),
.I2(CLBLL_L_X2Y107_SLICE_X0Y107_BO6),
.I3(RIOB33_X105Y105_IOB_X1Y106_I),
.I4(CLBLL_L_X2Y110_SLICE_X0Y110_AO6),
.I5(1'b1),
.O5(CLBLL_L_X2Y108_SLICE_X1Y108_BO5),
.O6(CLBLL_L_X2Y108_SLICE_X1Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a05f5f55ff55ff)
  ) CLBLL_L_X2Y108_SLICE_X1Y108_ALUT (
.I0(LIOB33_X0Y103_IOB_X0Y104_I),
.I1(1'b1),
.I2(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I3(RIOB33_X105Y105_IOB_X1Y106_I),
.I4(CLBLL_L_X2Y108_SLICE_X1Y108_CO6),
.I5(1'b1),
.O5(CLBLL_L_X2Y108_SLICE_X1Y108_AO5),
.O6(CLBLL_L_X2Y108_SLICE_X1Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h404400006a66cc00)
  ) CLBLL_L_X2Y109_SLICE_X0Y109_DLUT (
.I0(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I1(RIOB33_X105Y113_IOB_X1Y113_I),
.I2(RIOB33_X105Y111_IOB_X1Y112_I),
.I3(LIOB33_X0Y103_IOB_X0Y103_I),
.I4(RIOB33_X105Y105_IOB_X1Y106_I),
.I5(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.O5(CLBLL_L_X2Y109_SLICE_X0Y109_DO5),
.O6(CLBLL_L_X2Y109_SLICE_X0Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h404c22ee6a66cc00)
  ) CLBLL_L_X2Y109_SLICE_X0Y109_CLUT (
.I0(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I1(RIOB33_X105Y113_IOB_X1Y113_I),
.I2(RIOB33_X105Y111_IOB_X1Y112_I),
.I3(LIOB33_X0Y103_IOB_X0Y103_I),
.I4(RIOB33_X105Y105_IOB_X1Y106_I),
.I5(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.O5(CLBLL_L_X2Y109_SLICE_X0Y109_CO5),
.O6(CLBLL_L_X2Y109_SLICE_X0Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0ffffff000f000)
  ) CLBLL_L_X2Y109_SLICE_X0Y109_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I3(RIOB33_X105Y111_IOB_X1Y112_I),
.I4(LIOB33_X0Y101_IOB_X0Y101_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y109_SLICE_X0Y109_BO5),
.O6(CLBLL_L_X2Y109_SLICE_X0Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaabbffcc0033ff)
  ) CLBLL_L_X2Y109_SLICE_X0Y109_ALUT (
.I0(CLBLL_L_X2Y109_SLICE_X0Y109_DO6),
.I1(LIOB33_X0Y101_IOB_X0Y101_I),
.I2(1'b1),
.I3(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I4(CLBLL_L_X2Y109_SLICE_X0Y109_CO6),
.I5(1'b1),
.O5(CLBLL_L_X2Y109_SLICE_X0Y109_AO5),
.O6(CLBLL_L_X2Y109_SLICE_X0Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y109_SLICE_X1Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y109_SLICE_X1Y109_DO5),
.O6(CLBLL_L_X2Y109_SLICE_X1Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y109_SLICE_X1Y109_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y109_SLICE_X1Y109_CO5),
.O6(CLBLL_L_X2Y109_SLICE_X1Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y109_SLICE_X1Y109_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y109_SLICE_X1Y109_BO5),
.O6(CLBLL_L_X2Y109_SLICE_X1Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y109_SLICE_X1Y109_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y109_SLICE_X1Y109_AO5),
.O6(CLBLL_L_X2Y109_SLICE_X1Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y110_SLICE_X0Y110_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y110_SLICE_X0Y110_DO5),
.O6(CLBLL_L_X2Y110_SLICE_X0Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y110_SLICE_X0Y110_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y110_SLICE_X0Y110_CO5),
.O6(CLBLL_L_X2Y110_SLICE_X0Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y110_SLICE_X0Y110_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y110_SLICE_X0Y110_BO5),
.O6(CLBLL_L_X2Y110_SLICE_X0Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h07708bfc3c3c0000)
  ) CLBLL_L_X2Y110_SLICE_X0Y110_ALUT (
.I0(RIOB33_X105Y111_IOB_X1Y112_I),
.I1(LIOB33_X0Y103_IOB_X0Y103_I),
.I2(RIOB33_X105Y105_IOB_X1Y106_I),
.I3(LIOB33_X0Y113_IOB_X0Y114_I),
.I4(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I5(RIOB33_X105Y113_IOB_X1Y113_I),
.O5(CLBLL_L_X2Y110_SLICE_X0Y110_AO5),
.O6(CLBLL_L_X2Y110_SLICE_X0Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y110_SLICE_X1Y110_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y110_SLICE_X1Y110_DO5),
.O6(CLBLL_L_X2Y110_SLICE_X1Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y110_SLICE_X1Y110_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y110_SLICE_X1Y110_CO5),
.O6(CLBLL_L_X2Y110_SLICE_X1Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y110_SLICE_X1Y110_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y110_SLICE_X1Y110_BO5),
.O6(CLBLL_L_X2Y110_SLICE_X1Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y110_SLICE_X1Y110_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y110_SLICE_X1Y110_AO5),
.O6(CLBLL_L_X2Y110_SLICE_X1Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y111_SLICE_X0Y111_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y111_SLICE_X0Y111_DO5),
.O6(CLBLL_L_X2Y111_SLICE_X0Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y111_SLICE_X0Y111_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y111_SLICE_X0Y111_CO5),
.O6(CLBLL_L_X2Y111_SLICE_X0Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y111_SLICE_X0Y111_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y111_SLICE_X0Y111_BO5),
.O6(CLBLL_L_X2Y111_SLICE_X0Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y111_SLICE_X0Y111_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y111_SLICE_X0Y111_AO5),
.O6(CLBLL_L_X2Y111_SLICE_X0Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y111_SLICE_X1Y111_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y111_SLICE_X1Y111_DO5),
.O6(CLBLL_L_X2Y111_SLICE_X1Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y111_SLICE_X1Y111_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y111_SLICE_X1Y111_CO5),
.O6(CLBLL_L_X2Y111_SLICE_X1Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y111_SLICE_X1Y111_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y111_SLICE_X1Y111_BO5),
.O6(CLBLL_L_X2Y111_SLICE_X1Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'he7889ccc2b445000)
  ) CLBLL_L_X2Y111_SLICE_X1Y111_ALUT (
.I0(CLBLL_L_X4Y111_SLICE_X4Y111_DO6),
.I1(RIOB33_X105Y109_IOB_X1Y110_I),
.I2(LIOB33_X0Y109_IOB_X0Y110_I),
.I3(RIOB33_X105Y111_IOB_X1Y111_I),
.I4(LIOB33_X0Y111_IOB_X0Y111_I),
.I5(LIOB33_X0Y111_IOB_X0Y112_I),
.O5(CLBLL_L_X2Y111_SLICE_X1Y111_AO5),
.O6(CLBLL_L_X2Y111_SLICE_X1Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y112_SLICE_X0Y112_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y112_SLICE_X0Y112_DO5),
.O6(CLBLL_L_X2Y112_SLICE_X0Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y112_SLICE_X0Y112_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y112_SLICE_X0Y112_CO5),
.O6(CLBLL_L_X2Y112_SLICE_X0Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y112_SLICE_X0Y112_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y112_SLICE_X0Y112_BO5),
.O6(CLBLL_L_X2Y112_SLICE_X0Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h9d1d37b777777777)
  ) CLBLL_L_X2Y112_SLICE_X0Y112_ALUT (
.I0(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I1(RIOB33_X105Y113_IOB_X1Y113_I),
.I2(RIOB33_X105Y105_IOB_X1Y106_I),
.I3(RIOB33_X105Y111_IOB_X1Y112_I),
.I4(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y112_SLICE_X0Y112_AO5),
.O6(CLBLL_L_X2Y112_SLICE_X0Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y112_SLICE_X1Y112_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y112_SLICE_X1Y112_DO5),
.O6(CLBLL_L_X2Y112_SLICE_X1Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y112_SLICE_X1Y112_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y112_SLICE_X1Y112_CO5),
.O6(CLBLL_L_X2Y112_SLICE_X1Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y112_SLICE_X1Y112_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y112_SLICE_X1Y112_BO5),
.O6(CLBLL_L_X2Y112_SLICE_X1Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y112_SLICE_X1Y112_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y112_SLICE_X1Y112_AO5),
.O6(CLBLL_L_X2Y112_SLICE_X1Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff0f220ff0f2f02)
  ) CLBLL_L_X4Y105_SLICE_X4Y105_DLUT (
.I0(CLBLL_L_X4Y105_SLICE_X4Y105_AO6),
.I1(CLBLM_R_X5Y104_SLICE_X6Y104_AO6),
.I2(CLBLM_R_X7Y106_SLICE_X8Y106_CO6),
.I3(CLBLL_L_X4Y105_SLICE_X4Y105_AO5),
.I4(CLBLM_R_X5Y106_SLICE_X6Y106_CO6),
.I5(CLBLM_R_X7Y106_SLICE_X8Y106_AO6),
.O5(CLBLL_L_X4Y105_SLICE_X4Y105_DO5),
.O6(CLBLL_L_X4Y105_SLICE_X4Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h33ccc936cccc6666)
  ) CLBLL_L_X4Y105_SLICE_X4Y105_CLUT (
.I0(CLBLM_R_X5Y104_SLICE_X6Y104_AO6),
.I1(CLBLM_R_X7Y106_SLICE_X8Y106_CO6),
.I2(LIOB33_X0Y115_IOB_X0Y116_I),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(CLBLM_R_X5Y106_SLICE_X6Y106_CO6),
.I5(LIOB33_X0Y101_IOB_X0Y101_I),
.O5(CLBLL_L_X4Y105_SLICE_X4Y105_CO5),
.O6(CLBLL_L_X4Y105_SLICE_X4Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5aa51ee1a55ae11e)
  ) CLBLL_L_X4Y105_SLICE_X4Y105_BLUT (
.I0(CLBLM_R_X5Y106_SLICE_X6Y106_CO6),
.I1(CLBLL_L_X4Y105_SLICE_X4Y105_AO6),
.I2(CLBLM_R_X7Y106_SLICE_X8Y106_CO6),
.I3(CLBLM_R_X7Y106_SLICE_X8Y106_AO6),
.I4(CLBLM_R_X5Y104_SLICE_X6Y104_AO6),
.I5(CLBLL_L_X4Y105_SLICE_X4Y105_AO5),
.O5(CLBLL_L_X4Y105_SLICE_X4Y105_BO5),
.O6(CLBLL_L_X4Y105_SLICE_X4Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h777777775f5f5f5f)
  ) CLBLL_L_X4Y105_SLICE_X4Y105_ALUT (
.I0(LIOB33_X0Y115_IOB_X0Y116_I),
.I1(LIOB33_X0Y101_IOB_X0Y101_I),
.I2(LIOB33_X0Y101_IOB_X0Y102_I),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y105_SLICE_X4Y105_AO5),
.O6(CLBLL_L_X4Y105_SLICE_X4Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y105_SLICE_X5Y105_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y105_SLICE_X5Y105_DO5),
.O6(CLBLL_L_X4Y105_SLICE_X5Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y105_SLICE_X5Y105_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y105_SLICE_X5Y105_CO5),
.O6(CLBLL_L_X4Y105_SLICE_X5Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y105_SLICE_X5Y105_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y105_SLICE_X5Y105_BO5),
.O6(CLBLL_L_X4Y105_SLICE_X5Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h59a6a6599a65659a)
  ) CLBLL_L_X4Y105_SLICE_X5Y105_ALUT (
.I0(CLBLM_R_X7Y105_SLICE_X8Y105_BO6),
.I1(CLBLL_L_X4Y105_SLICE_X4Y105_BO6),
.I2(CLBLM_R_X3Y104_SLICE_X3Y104_CO6),
.I3(CLBLL_L_X4Y105_SLICE_X4Y105_DO6),
.I4(CLBLM_R_X7Y105_SLICE_X8Y105_AO6),
.I5(CLBLM_R_X3Y105_SLICE_X3Y105_BO5),
.O5(CLBLL_L_X4Y105_SLICE_X5Y105_AO5),
.O6(CLBLL_L_X4Y105_SLICE_X5Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefbc832ecb38020)
  ) CLBLL_L_X4Y106_SLICE_X4Y106_DLUT (
.I0(CLBLM_R_X3Y106_SLICE_X2Y106_BO6),
.I1(CLBLM_R_X3Y105_SLICE_X3Y105_DO6),
.I2(CLBLM_R_X3Y106_SLICE_X2Y106_AO6),
.I3(CLBLM_R_X5Y106_SLICE_X6Y106_BO6),
.I4(CLBLL_L_X4Y106_SLICE_X4Y106_AO6),
.I5(CLBLM_R_X3Y106_SLICE_X3Y106_AO6),
.O5(CLBLL_L_X4Y106_SLICE_X4Y106_DO5),
.O6(CLBLL_L_X4Y106_SLICE_X4Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h96cc66cc993396cc)
  ) CLBLL_L_X4Y106_SLICE_X4Y106_CLUT (
.I0(LIOB33_X0Y115_IOB_X0Y116_I),
.I1(CLBLL_L_X4Y105_SLICE_X4Y105_CO6),
.I2(LIOB33_X0Y113_IOB_X0Y114_I),
.I3(LIOB33_X0Y101_IOB_X0Y102_I),
.I4(CLBLM_R_X5Y106_SLICE_X6Y106_AO6),
.I5(CLBLM_R_X3Y105_SLICE_X3Y105_AO5),
.O5(CLBLL_L_X4Y106_SLICE_X4Y106_CO5),
.O6(CLBLL_L_X4Y106_SLICE_X4Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h59aaa6aa9aa565a5)
  ) CLBLL_L_X4Y106_SLICE_X4Y106_BLUT (
.I0(CLBLM_R_X3Y105_SLICE_X3Y105_DO6),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(CLBLM_R_X3Y106_SLICE_X2Y106_BO6),
.I3(LIOB33_X0Y105_IOB_X0Y105_I),
.I4(LIOB33_X0Y103_IOB_X0Y103_I),
.I5(CLBLM_R_X3Y106_SLICE_X3Y106_AO6),
.O5(CLBLL_L_X4Y106_SLICE_X4Y106_BO5),
.O6(CLBLL_L_X4Y106_SLICE_X4Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h55ff55ff5f5f5f5f)
  ) CLBLL_L_X4Y106_SLICE_X4Y106_ALUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(1'b1),
.I2(LIOB33_X0Y103_IOB_X0Y103_I),
.I3(RIOB33_X105Y105_IOB_X1Y106_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y106_SLICE_X4Y106_AO5),
.O6(CLBLL_L_X4Y106_SLICE_X4Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcd4d4c0cf4d4d0c)
  ) CLBLL_L_X4Y106_SLICE_X5Y106_DLUT (
.I0(CLBLL_L_X4Y106_SLICE_X5Y106_AO6),
.I1(CLBLL_L_X4Y106_SLICE_X4Y106_AO5),
.I2(CLBLM_R_X5Y106_SLICE_X6Y106_BO5),
.I3(CLBLM_R_X3Y106_SLICE_X3Y106_BO6),
.I4(CLBLM_R_X5Y106_SLICE_X6Y106_BO6),
.I5(CLBLL_L_X4Y105_SLICE_X5Y105_AO6),
.O5(CLBLL_L_X4Y106_SLICE_X5Y106_DO5),
.O6(CLBLL_L_X4Y106_SLICE_X5Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h2abfbfbf80eaeaea)
  ) CLBLL_L_X4Y106_SLICE_X5Y106_CLUT (
.I0(CLBLM_R_X3Y104_SLICE_X3Y104_CO6),
.I1(LIOB33_X0Y101_IOB_X0Y102_I),
.I2(LIOB33_X0Y115_IOB_X0Y116_I),
.I3(LIOB33_X0Y113_IOB_X0Y114_I),
.I4(LIOB33_X0Y103_IOB_X0Y104_I),
.I5(CLBLL_L_X4Y105_SLICE_X4Y105_CO6),
.O5(CLBLL_L_X4Y106_SLICE_X5Y106_CO5),
.O6(CLBLL_L_X4Y106_SLICE_X5Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hd2a54bf02da5b4f0)
  ) CLBLL_L_X4Y106_SLICE_X5Y106_BLUT (
.I0(CLBLM_R_X3Y106_SLICE_X3Y106_BO6),
.I1(LIOB33_X0Y103_IOB_X0Y103_I),
.I2(CLBLL_L_X4Y105_SLICE_X5Y105_AO6),
.I3(LIOB33_X0Y105_IOB_X0Y105_I),
.I4(CLBLL_L_X4Y106_SLICE_X5Y106_AO6),
.I5(LIOB33_X0Y113_IOB_X0Y114_I),
.O5(CLBLL_L_X4Y106_SLICE_X5Y106_BO5),
.O6(CLBLL_L_X4Y106_SLICE_X5Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6c93936c93936c6c)
  ) CLBLL_L_X4Y106_SLICE_X5Y106_ALUT (
.I0(LIOB33_X0Y113_IOB_X0Y114_I),
.I1(CLBLM_R_X3Y104_SLICE_X3Y104_CO6),
.I2(LIOB33_X0Y103_IOB_X0Y104_I),
.I3(LIOB33_X0Y115_IOB_X0Y116_I),
.I4(CLBLL_L_X4Y105_SLICE_X4Y105_CO6),
.I5(LIOB33_X0Y101_IOB_X0Y102_I),
.O5(CLBLL_L_X4Y106_SLICE_X5Y106_AO5),
.O6(CLBLL_L_X4Y106_SLICE_X5Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y107_SLICE_X4Y107_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y107_SLICE_X4Y107_DO5),
.O6(CLBLL_L_X4Y107_SLICE_X4Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h4dd4cffcd4d4fcfc)
  ) CLBLL_L_X4Y107_SLICE_X4Y107_CLUT (
.I0(LIOB33_X0Y103_IOB_X0Y103_I),
.I1(CLBLM_R_X3Y106_SLICE_X3Y106_BO6),
.I2(CLBLL_L_X4Y106_SLICE_X4Y106_CO6),
.I3(LIOB33_X0Y103_IOB_X0Y104_I),
.I4(LIOB33_X0Y105_IOB_X0Y105_I),
.I5(LIOB33_X0Y113_IOB_X0Y114_I),
.O5(CLBLL_L_X4Y107_SLICE_X4Y107_CO5),
.O6(CLBLL_L_X4Y107_SLICE_X4Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h2b8e8e8ebbeeeeee)
  ) CLBLL_L_X4Y107_SLICE_X4Y107_BLUT (
.I0(CLBLL_L_X4Y106_SLICE_X4Y106_DO6),
.I1(CLBLL_L_X4Y106_SLICE_X5Y106_BO6),
.I2(RIOB33_X105Y105_IOB_X1Y106_I),
.I3(LIOB33_X0Y105_IOB_X0Y106_I),
.I4(LIOB33_X0Y103_IOB_X0Y103_I),
.I5(LIOB33_X0Y107_IOB_X0Y107_I),
.O5(CLBLL_L_X4Y107_SLICE_X4Y107_BO5),
.O6(CLBLL_L_X4Y107_SLICE_X4Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6c939393936c6c6c)
  ) CLBLL_L_X4Y107_SLICE_X4Y107_ALUT (
.I0(LIOB33_X0Y105_IOB_X0Y105_I),
.I1(CLBLL_L_X4Y106_SLICE_X4Y106_CO6),
.I2(LIOB33_X0Y103_IOB_X0Y103_I),
.I3(LIOB33_X0Y113_IOB_X0Y114_I),
.I4(LIOB33_X0Y103_IOB_X0Y104_I),
.I5(CLBLM_R_X3Y106_SLICE_X3Y106_BO6),
.O5(CLBLL_L_X4Y107_SLICE_X4Y107_AO5),
.O6(CLBLL_L_X4Y107_SLICE_X4Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y107_SLICE_X5Y107_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y107_SLICE_X5Y107_DO5),
.O6(CLBLL_L_X4Y107_SLICE_X5Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y107_SLICE_X5Y107_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y107_SLICE_X5Y107_CO5),
.O6(CLBLL_L_X4Y107_SLICE_X5Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y107_SLICE_X5Y107_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y107_SLICE_X5Y107_BO5),
.O6(CLBLL_L_X4Y107_SLICE_X5Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y107_SLICE_X5Y107_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y107_SLICE_X5Y107_AO5),
.O6(CLBLL_L_X4Y107_SLICE_X5Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y108_SLICE_X4Y108_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y108_SLICE_X4Y108_DO5),
.O6(CLBLL_L_X4Y108_SLICE_X4Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7dddffff14443ccc)
  ) CLBLL_L_X4Y108_SLICE_X4Y108_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y106_I),
.I1(CLBLL_L_X4Y108_SLICE_X5Y108_AO6),
.I2(LIOB33_X0Y103_IOB_X0Y103_I),
.I3(LIOB33_X0Y107_IOB_X0Y107_I),
.I4(LIOB33_X0Y107_IOB_X0Y108_I),
.I5(CLBLL_L_X4Y107_SLICE_X4Y107_BO6),
.O5(CLBLL_L_X4Y108_SLICE_X4Y108_CO5),
.O6(CLBLL_L_X4Y108_SLICE_X4Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h96a55a96aa66aa66)
  ) CLBLL_L_X4Y108_SLICE_X4Y108_BLUT (
.I0(CLBLM_R_X5Y107_SLICE_X7Y107_AO6),
.I1(CLBLL_L_X4Y108_SLICE_X5Y108_BO6),
.I2(LIOB33_X0Y103_IOB_X0Y103_I),
.I3(CLBLL_L_X4Y107_SLICE_X4Y107_BO6),
.I4(RIOB33_X105Y105_IOB_X1Y106_I),
.I5(LIOB33_X0Y107_IOB_X0Y108_I),
.O5(CLBLL_L_X4Y108_SLICE_X4Y108_BO5),
.O6(CLBLL_L_X4Y108_SLICE_X4Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996c33ca55a0ff0)
  ) CLBLL_L_X4Y108_SLICE_X4Y108_ALUT (
.I0(LIOB33_X0Y107_IOB_X0Y108_I),
.I1(LIOB33_X0Y103_IOB_X0Y103_I),
.I2(CLBLL_L_X4Y108_SLICE_X5Y108_AO6),
.I3(CLBLL_L_X4Y107_SLICE_X4Y107_BO6),
.I4(RIOB33_X105Y105_IOB_X1Y106_I),
.I5(LIOB33_X0Y107_IOB_X0Y107_I),
.O5(CLBLL_L_X4Y108_SLICE_X4Y108_AO5),
.O6(CLBLL_L_X4Y108_SLICE_X4Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y108_SLICE_X5Y108_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y108_SLICE_X5Y108_DO5),
.O6(CLBLL_L_X4Y108_SLICE_X5Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'he68acc6c2a4600a0)
  ) CLBLL_L_X4Y108_SLICE_X5Y108_CLUT (
.I0(RIOB33_X105Y111_IOB_X1Y111_I),
.I1(RIOB33_X105Y109_IOB_X1Y110_I),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(CLBLM_R_X5Y108_SLICE_X6Y108_DO6),
.I4(LIOB33_X0Y107_IOB_X0Y107_I),
.I5(LIOB33_X0Y107_IOB_X0Y108_I),
.O5(CLBLL_L_X4Y108_SLICE_X5Y108_CO5),
.O6(CLBLL_L_X4Y108_SLICE_X5Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996c33ca55a0ff0)
  ) CLBLL_L_X4Y108_SLICE_X5Y108_BLUT (
.I0(LIOB33_X0Y107_IOB_X0Y107_I),
.I1(LIOB33_X0Y113_IOB_X0Y114_I),
.I2(CLBLM_R_X5Y106_SLICE_X7Y106_BO6),
.I3(CLBLL_L_X4Y106_SLICE_X5Y106_DO6),
.I4(LIOB33_X0Y103_IOB_X0Y103_I),
.I5(LIOB33_X0Y105_IOB_X0Y106_I),
.O5(CLBLL_L_X4Y108_SLICE_X5Y108_BO5),
.O6(CLBLL_L_X4Y108_SLICE_X5Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h96c33c96f05af05a)
  ) CLBLL_L_X4Y108_SLICE_X5Y108_ALUT (
.I0(CLBLM_R_X5Y107_SLICE_X6Y107_AO6),
.I1(LIOB33_X0Y113_IOB_X0Y114_I),
.I2(CLBLM_R_X5Y106_SLICE_X7Y106_BO6),
.I3(CLBLL_L_X4Y107_SLICE_X4Y107_CO6),
.I4(LIOB33_X0Y103_IOB_X0Y103_I),
.I5(LIOB33_X0Y105_IOB_X0Y106_I),
.O5(CLBLL_L_X4Y108_SLICE_X5Y108_AO5),
.O6(CLBLL_L_X4Y108_SLICE_X5Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffc3d741d741c300)
  ) CLBLL_L_X4Y109_SLICE_X4Y109_DLUT (
.I0(CLBLL_L_X4Y108_SLICE_X5Y108_BO6),
.I1(CLBLL_L_X4Y110_SLICE_X4Y110_AO6),
.I2(CLBLM_R_X5Y107_SLICE_X7Y107_AO6),
.I3(CLBLL_L_X4Y109_SLICE_X4Y109_AO5),
.I4(CLBLL_L_X4Y110_SLICE_X4Y110_AO5),
.I5(CLBLL_L_X4Y107_SLICE_X4Y107_BO6),
.O5(CLBLL_L_X4Y109_SLICE_X4Y109_DO5),
.O6(CLBLL_L_X4Y109_SLICE_X4Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h2dd2b44bd22d4bb4)
  ) CLBLL_L_X4Y109_SLICE_X4Y109_CLUT (
.I0(CLBLL_L_X4Y108_SLICE_X5Y108_BO6),
.I1(CLBLL_L_X4Y107_SLICE_X4Y107_BO6),
.I2(CLBLM_R_X5Y107_SLICE_X7Y107_AO6),
.I3(CLBLL_L_X4Y109_SLICE_X4Y109_AO5),
.I4(CLBLL_L_X4Y110_SLICE_X4Y110_AO5),
.I5(CLBLL_L_X4Y110_SLICE_X4Y110_AO6),
.O5(CLBLL_L_X4Y109_SLICE_X4Y109_CO5),
.O6(CLBLL_L_X4Y109_SLICE_X4Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h444c5d5f5fdfdfff)
  ) CLBLL_L_X4Y109_SLICE_X4Y109_BLUT (
.I0(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I1(CLBLM_R_X3Y108_SLICE_X3Y108_BO6),
.I2(LIOB33_X0Y109_IOB_X0Y110_I),
.I3(LIOB33_X0Y109_IOB_X0Y109_I),
.I4(CLBLL_L_X4Y108_SLICE_X4Y108_AO6),
.I5(CLBLL_L_X4Y109_SLICE_X4Y109_CO6),
.O5(CLBLL_L_X4Y109_SLICE_X4Y109_BO5),
.O6(CLBLL_L_X4Y109_SLICE_X4Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5fa0a05f3f3f3f3f)
  ) CLBLL_L_X4Y109_SLICE_X4Y109_ALUT (
.I0(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(LIOB33_X0Y109_IOB_X0Y109_I),
.I3(CLBLM_R_X3Y108_SLICE_X3Y108_BO6),
.I4(CLBLL_L_X4Y108_SLICE_X4Y108_AO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y109_SLICE_X4Y109_AO5),
.O6(CLBLL_L_X4Y109_SLICE_X4Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y109_SLICE_X5Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y109_SLICE_X5Y109_DO5),
.O6(CLBLL_L_X4Y109_SLICE_X5Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hb43c78f0d2961e5a)
  ) CLBLL_L_X4Y109_SLICE_X5Y109_CLUT (
.I0(CLBLM_R_X5Y108_SLICE_X6Y108_BO6),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(CLBLM_R_X5Y109_SLICE_X6Y109_CO6),
.I3(LIOB33_X0Y109_IOB_X0Y109_I),
.I4(LIOB33_X0Y109_IOB_X0Y110_I),
.I5(CLBLL_L_X4Y108_SLICE_X4Y108_CO6),
.O5(CLBLL_L_X4Y109_SLICE_X5Y109_CO5),
.O6(CLBLL_L_X4Y109_SLICE_X5Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h1f055f1f7f55ff7f)
  ) CLBLL_L_X4Y109_SLICE_X5Y109_BLUT (
.I0(CLBLM_R_X5Y109_SLICE_X6Y109_CO6),
.I1(LIOB33_X0Y109_IOB_X0Y109_I),
.I2(RIOB33_X105Y105_IOB_X1Y106_I),
.I3(CLBLL_L_X4Y108_SLICE_X4Y108_CO6),
.I4(CLBLM_R_X5Y108_SLICE_X6Y108_BO6),
.I5(LIOB33_X0Y109_IOB_X0Y110_I),
.O5(CLBLL_L_X4Y109_SLICE_X5Y109_BO5),
.O6(CLBLL_L_X4Y109_SLICE_X5Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hd78877d728778828)
  ) CLBLL_L_X4Y109_SLICE_X5Y109_ALUT (
.I0(LIOB33_X0Y109_IOB_X0Y109_I),
.I1(LIOB33_X0Y103_IOB_X0Y103_I),
.I2(RIOB33_X105Y105_IOB_X1Y106_I),
.I3(CLBLL_L_X4Y108_SLICE_X4Y108_CO6),
.I4(CLBLM_R_X5Y108_SLICE_X6Y108_BO6),
.I5(CLBLM_R_X5Y109_SLICE_X6Y109_BO6),
.O5(CLBLL_L_X4Y109_SLICE_X5Y109_AO5),
.O6(CLBLL_L_X4Y109_SLICE_X5Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf9ff909999f90090)
  ) CLBLL_L_X4Y110_SLICE_X4Y110_DLUT (
.I0(CLBLM_R_X5Y110_SLICE_X6Y110_BO6),
.I1(CLBLM_R_X3Y111_SLICE_X2Y111_AO6),
.I2(CLBLL_L_X4Y109_SLICE_X4Y109_BO6),
.I3(CLBLL_L_X4Y109_SLICE_X5Y109_CO6),
.I4(CLBLL_L_X4Y111_SLICE_X4Y111_AO5),
.I5(CLBLL_L_X4Y110_SLICE_X4Y110_BO6),
.O5(CLBLL_L_X4Y110_SLICE_X4Y110_DO5),
.O6(CLBLL_L_X4Y110_SLICE_X4Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6fffafff06660aaa)
  ) CLBLL_L_X4Y110_SLICE_X4Y110_CLUT (
.I0(CLBLL_L_X4Y109_SLICE_X5Y109_AO6),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I3(LIOB33_X0Y111_IOB_X0Y111_I),
.I4(LIOB33_X0Y109_IOB_X0Y110_I),
.I5(CLBLL_L_X4Y109_SLICE_X4Y109_BO6),
.O5(CLBLL_L_X4Y110_SLICE_X4Y110_CO5),
.O6(CLBLL_L_X4Y110_SLICE_X4Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f3f3f3f66aa9955)
  ) CLBLL_L_X4Y110_SLICE_X4Y110_BLUT (
.I0(CLBLM_R_X7Y110_SLICE_X9Y110_BO5),
.I1(LIOB33_X0Y111_IOB_X0Y111_I),
.I2(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I3(RIOB33_X105Y107_IOB_X1Y107_I),
.I4(CLBLM_R_X5Y109_SLICE_X7Y109_DO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y110_SLICE_X4Y110_BO5),
.O6(CLBLL_L_X4Y110_SLICE_X4Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h33ff33ff55ff55ff)
  ) CLBLL_L_X4Y110_SLICE_X4Y110_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y106_I),
.I1(LIOB33_X0Y103_IOB_X0Y103_I),
.I2(1'b1),
.I3(LIOB33_X0Y107_IOB_X0Y108_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y110_SLICE_X4Y110_AO5),
.O6(CLBLL_L_X4Y110_SLICE_X4Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hd4af2baf2b50d450)
  ) CLBLL_L_X4Y110_SLICE_X5Y110_DLUT (
.I0(CLBLM_R_X5Y109_SLICE_X7Y109_CO6),
.I1(LIOB33_X0Y111_IOB_X0Y111_I),
.I2(CLBLM_R_X5Y110_SLICE_X6Y110_AO6),
.I3(RIOB33_X105Y107_IOB_X1Y108_I),
.I4(LIOB33_X0Y111_IOB_X0Y112_I),
.I5(CLBLL_L_X4Y110_SLICE_X5Y110_BO6),
.O5(CLBLL_L_X4Y110_SLICE_X5Y110_DO5),
.O6(CLBLL_L_X4Y110_SLICE_X5Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7177f7f775f7ffff)
  ) CLBLL_L_X4Y110_SLICE_X5Y110_CLUT (
.I0(LIOB33_X0Y107_IOB_X0Y107_I),
.I1(RIOB33_X105Y109_IOB_X1Y110_I),
.I2(CLBLM_R_X5Y108_SLICE_X6Y108_DO6),
.I3(LIOB33_X0Y105_IOB_X0Y106_I),
.I4(RIOB33_X105Y111_IOB_X1Y111_I),
.I5(LIOB33_X0Y107_IOB_X0Y108_I),
.O5(CLBLL_L_X4Y110_SLICE_X5Y110_CO5),
.O6(CLBLL_L_X4Y110_SLICE_X5Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h9a5aa6966aaa5666)
  ) CLBLL_L_X4Y110_SLICE_X5Y110_BLUT (
.I0(CLBLM_R_X3Y110_SLICE_X3Y110_DO6),
.I1(CLBLM_R_X5Y109_SLICE_X7Y109_AO5),
.I2(RIOB33_X105Y109_IOB_X1Y109_I),
.I3(LIOB33_X0Y109_IOB_X0Y110_I),
.I4(CLBLM_R_X5Y108_SLICE_X7Y108_AO6),
.I5(LIOB33_X0Y111_IOB_X0Y111_I),
.O5(CLBLL_L_X4Y110_SLICE_X5Y110_BO5),
.O6(CLBLL_L_X4Y110_SLICE_X5Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h1f075f177f57ff77)
  ) CLBLL_L_X4Y110_SLICE_X5Y110_ALUT (
.I0(CLBLM_R_X3Y110_SLICE_X3Y110_DO6),
.I1(CLBLM_R_X5Y109_SLICE_X7Y109_AO5),
.I2(RIOB33_X105Y109_IOB_X1Y109_I),
.I3(CLBLM_R_X5Y108_SLICE_X7Y108_AO6),
.I4(LIOB33_X0Y109_IOB_X0Y110_I),
.I5(LIOB33_X0Y111_IOB_X0Y111_I),
.O5(CLBLL_L_X4Y110_SLICE_X5Y110_AO5),
.O6(CLBLL_L_X4Y110_SLICE_X5Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3713ff77ff3fffff)
  ) CLBLL_L_X4Y111_SLICE_X4Y111_DLUT (
.I0(LIOB33_X0Y109_IOB_X0Y110_I),
.I1(LIOB33_X0Y109_IOB_X0Y109_I),
.I2(LIOB33_X0Y107_IOB_X0Y108_I),
.I3(CLBLL_L_X4Y110_SLICE_X5Y110_CO6),
.I4(RIOB33_X105Y111_IOB_X1Y111_I),
.I5(RIOB33_X105Y109_IOB_X1Y110_I),
.O5(CLBLL_L_X4Y111_SLICE_X4Y111_DO5),
.O6(CLBLL_L_X4Y111_SLICE_X4Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h507075ff55f7f7ff)
  ) CLBLL_L_X4Y111_SLICE_X4Y111_CLUT (
.I0(RIOB33_X105Y107_IOB_X1Y107_I),
.I1(LIOB33_X0Y111_IOB_X0Y111_I),
.I2(CLBLM_R_X7Y110_SLICE_X9Y110_BO5),
.I3(LIOB33_X0Y111_IOB_X0Y112_I),
.I4(CLBLM_R_X3Y111_SLICE_X3Y111_AO5),
.I5(CLBLM_R_X5Y109_SLICE_X7Y109_DO6),
.O5(CLBLL_L_X4Y111_SLICE_X4Y111_CO5),
.O6(CLBLL_L_X4Y111_SLICE_X4Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha95969996a9a5aaa)
  ) CLBLL_L_X4Y111_SLICE_X4Y111_BLUT (
.I0(CLBLM_R_X3Y111_SLICE_X3Y111_AO5),
.I1(CLBLM_R_X7Y110_SLICE_X9Y110_BO5),
.I2(RIOB33_X105Y107_IOB_X1Y107_I),
.I3(LIOB33_X0Y111_IOB_X0Y112_I),
.I4(LIOB33_X0Y111_IOB_X0Y111_I),
.I5(CLBLM_R_X5Y109_SLICE_X7Y109_DO6),
.O5(CLBLL_L_X4Y111_SLICE_X4Y111_BO5),
.O6(CLBLL_L_X4Y111_SLICE_X4Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h7887788777777777)
  ) CLBLL_L_X4Y111_SLICE_X4Y111_ALUT (
.I0(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I1(LIOB33_X0Y111_IOB_X0Y112_I),
.I2(CLBLL_L_X4Y111_SLICE_X5Y111_AO6),
.I3(CLBLL_L_X4Y110_SLICE_X4Y110_CO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y111_SLICE_X4Y111_AO5),
.O6(CLBLL_L_X4Y111_SLICE_X4Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h45455ddf4dcfffff)
  ) CLBLL_L_X4Y111_SLICE_X5Y111_DLUT (
.I0(RIOB33_X105Y107_IOB_X1Y108_I),
.I1(CLBLM_R_X5Y109_SLICE_X7Y109_CO6),
.I2(CLBLM_R_X5Y110_SLICE_X6Y110_AO6),
.I3(LIOB33_X0Y111_IOB_X0Y111_I),
.I4(CLBLL_L_X4Y110_SLICE_X5Y110_BO6),
.I5(LIOB33_X0Y111_IOB_X0Y112_I),
.O5(CLBLL_L_X4Y111_SLICE_X5Y111_DO5),
.O6(CLBLL_L_X4Y111_SLICE_X5Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fbf152aff3f3f00)
  ) CLBLL_L_X4Y111_SLICE_X5Y111_CLUT (
.I0(LIOB33_X0Y113_IOB_X0Y114_I),
.I1(LIOB33_X0Y111_IOB_X0Y111_I),
.I2(LIOB33_X0Y103_IOB_X0Y103_I),
.I3(CLBLM_R_X7Y110_SLICE_X9Y110_DO6),
.I4(CLBLM_R_X5Y110_SLICE_X7Y110_DO6),
.I5(LIOB33_X0Y109_IOB_X0Y110_I),
.O5(CLBLL_L_X4Y111_SLICE_X5Y111_CO5),
.O6(CLBLL_L_X4Y111_SLICE_X5Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6a959595956a6a6a)
  ) CLBLL_L_X4Y111_SLICE_X5Y111_BLUT (
.I0(CLBLM_R_X7Y110_SLICE_X9Y110_DO6),
.I1(LIOB33_X0Y103_IOB_X0Y103_I),
.I2(LIOB33_X0Y111_IOB_X0Y111_I),
.I3(LIOB33_X0Y109_IOB_X0Y110_I),
.I4(LIOB33_X0Y113_IOB_X0Y114_I),
.I5(CLBLM_R_X5Y110_SLICE_X7Y110_DO6),
.O5(CLBLL_L_X4Y111_SLICE_X5Y111_BO5),
.O6(CLBLL_L_X4Y111_SLICE_X5Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6a95956ac03f3fc0)
  ) CLBLL_L_X4Y111_SLICE_X5Y111_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y106_I),
.I1(LIOB33_X0Y103_IOB_X0Y103_I),
.I2(LIOB33_X0Y109_IOB_X0Y110_I),
.I3(CLBLL_L_X4Y109_SLICE_X5Y109_BO6),
.I4(CLBLM_R_X5Y109_SLICE_X7Y109_BO6),
.I5(LIOB33_X0Y111_IOB_X0Y111_I),
.O5(CLBLL_L_X4Y111_SLICE_X5Y111_AO5),
.O6(CLBLL_L_X4Y111_SLICE_X5Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y112_SLICE_X4Y112_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y112_SLICE_X4Y112_DO5),
.O6(CLBLL_L_X4Y112_SLICE_X4Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hd57fbd77d5ff957f)
  ) CLBLL_L_X4Y112_SLICE_X4Y112_CLUT (
.I0(RIOB33_X105Y111_IOB_X1Y111_I),
.I1(LIOB33_X0Y111_IOB_X0Y111_I),
.I2(RIOB33_X105Y109_IOB_X1Y110_I),
.I3(LIOB33_X0Y111_IOB_X0Y112_I),
.I4(CLBLL_L_X4Y111_SLICE_X4Y111_DO6),
.I5(LIOB33_X0Y109_IOB_X0Y110_I),
.O5(CLBLL_L_X4Y112_SLICE_X4Y112_CO5),
.O6(CLBLL_L_X4Y112_SLICE_X4Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6999a55596665aaa)
  ) CLBLL_L_X4Y112_SLICE_X4Y112_BLUT (
.I0(CLBLM_R_X3Y111_SLICE_X2Y111_DO6),
.I1(LIOB33_X0Y115_IOB_X0Y115_I),
.I2(RIOB33_X105Y109_IOB_X1Y110_I),
.I3(LIOB33_X0Y113_IOB_X0Y113_I),
.I4(RIOB33_X105Y109_IOB_X1Y109_I),
.I5(CLBLL_L_X4Y112_SLICE_X4Y112_CO6),
.O5(CLBLL_L_X4Y112_SLICE_X4Y112_BO5),
.O6(CLBLL_L_X4Y112_SLICE_X4Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h7887878787787878)
  ) CLBLL_L_X4Y112_SLICE_X4Y112_ALUT (
.I0(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I1(LIOB33_X0Y115_IOB_X0Y115_I),
.I2(CLBLM_R_X5Y111_SLICE_X6Y111_BO6),
.I3(LIOB33_X0Y113_IOB_X0Y113_I),
.I4(RIOB33_X105Y105_IOB_X1Y106_I),
.I5(CLBLM_R_X3Y111_SLICE_X3Y111_CO6),
.O5(CLBLL_L_X4Y112_SLICE_X4Y112_AO5),
.O6(CLBLL_L_X4Y112_SLICE_X4Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f3f3f3f3f3f3f3f)
  ) CLBLL_L_X4Y112_SLICE_X5Y112_DLUT (
.I0(1'b1),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(LIOB33_X0Y113_IOB_X0Y113_I),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y112_SLICE_X5Y112_DO5),
.O6(CLBLL_L_X4Y112_SLICE_X5Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h4bd2b42db42d4bd2)
  ) CLBLL_L_X4Y112_SLICE_X5Y112_CLUT (
.I0(CLBLL_L_X4Y112_SLICE_X5Y112_AO6),
.I1(CLBLM_R_X5Y111_SLICE_X7Y111_CO6),
.I2(CLBLL_L_X4Y111_SLICE_X4Y111_BO6),
.I3(CLBLM_R_X7Y111_SLICE_X8Y111_DO6),
.I4(CLBLM_R_X5Y111_SLICE_X7Y111_DO6),
.I5(CLBLL_L_X4Y112_SLICE_X5Y112_DO6),
.O5(CLBLL_L_X4Y112_SLICE_X5Y112_CO5),
.O6(CLBLL_L_X4Y112_SLICE_X5Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h2abf2abf6a956a95)
  ) CLBLL_L_X4Y112_SLICE_X5Y112_BLUT (
.I0(CLBLM_R_X5Y111_SLICE_X7Y111_DO6),
.I1(LIOB33_X0Y113_IOB_X0Y113_I),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLL_L_X4Y111_SLICE_X4Y111_BO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y112_SLICE_X5Y112_BO5),
.O6(CLBLL_L_X4Y112_SLICE_X5Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333ffff5aa5aa55)
  ) CLBLL_L_X4Y112_SLICE_X5Y112_ALUT (
.I0(CLBLL_L_X4Y111_SLICE_X5Y111_DO6),
.I1(RIOB33_X105Y103_IOB_X1Y104_I),
.I2(RIOB33_X105Y107_IOB_X1Y108_I),
.I3(CLBLM_R_X3Y111_SLICE_X2Y111_BO6),
.I4(LIOB33_X0Y113_IOB_X0Y113_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y112_SLICE_X5Y112_AO5),
.O6(CLBLL_L_X4Y112_SLICE_X5Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y113_SLICE_X4Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y113_SLICE_X4Y113_DO5),
.O6(CLBLL_L_X4Y113_SLICE_X4Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hd4d4d444ddddddd4)
  ) CLBLL_L_X4Y113_SLICE_X4Y113_CLUT (
.I0(CLBLL_L_X4Y112_SLICE_X4Y112_BO6),
.I1(CLBLM_R_X3Y112_SLICE_X2Y112_BO6),
.I2(CLBLL_L_X4Y113_SLICE_X5Y113_DO6),
.I3(CLBLL_L_X4Y113_SLICE_X5Y113_BO6),
.I4(CLBLL_L_X4Y115_SLICE_X4Y115_CO6),
.I5(CLBLM_R_X3Y112_SLICE_X2Y112_AO6),
.O5(CLBLL_L_X4Y113_SLICE_X4Y113_CO5),
.O6(CLBLL_L_X4Y113_SLICE_X4Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'he1f01e0f0fe1f01e)
  ) CLBLL_L_X4Y113_SLICE_X4Y113_BLUT (
.I0(CLBLL_L_X4Y115_SLICE_X4Y115_CO6),
.I1(CLBLL_L_X4Y113_SLICE_X5Y113_BO6),
.I2(CLBLM_R_X3Y112_SLICE_X2Y112_BO6),
.I3(CLBLM_R_X3Y112_SLICE_X2Y112_AO6),
.I4(CLBLL_L_X4Y112_SLICE_X4Y112_BO6),
.I5(CLBLL_L_X4Y113_SLICE_X5Y113_DO6),
.O5(CLBLL_L_X4Y113_SLICE_X4Y113_BO5),
.O6(CLBLL_L_X4Y113_SLICE_X4Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0fffff69996999)
  ) CLBLL_L_X4Y113_SLICE_X4Y113_ALUT (
.I0(CLBLL_L_X4Y110_SLICE_X5Y110_DO6),
.I1(CLBLL_L_X4Y111_SLICE_X4Y111_CO6),
.I2(LIOB33_X0Y113_IOB_X0Y113_I),
.I3(RIOB33_X105Y107_IOB_X1Y107_I),
.I4(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y113_SLICE_X4Y113_AO5),
.O6(CLBLL_L_X4Y113_SLICE_X4Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h577f77ff0077577f)
  ) CLBLL_L_X4Y113_SLICE_X5Y113_DLUT (
.I0(RIOB33_X105Y107_IOB_X1Y107_I),
.I1(LIOB33_X0Y115_IOB_X0Y115_I),
.I2(LIOB33_X0Y113_IOB_X0Y113_I),
.I3(CLBLL_L_X4Y112_SLICE_X5Y112_AO5),
.I4(CLBLL_L_X4Y110_SLICE_X5Y110_DO6),
.I5(CLBLL_L_X4Y111_SLICE_X4Y111_CO6),
.O5(CLBLL_L_X4Y113_SLICE_X5Y113_DO5),
.O6(CLBLL_L_X4Y113_SLICE_X5Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h9f603fc0c03f9f60)
  ) CLBLL_L_X4Y113_SLICE_X5Y113_CLUT (
.I0(LIOB33_X0Y113_IOB_X0Y113_I),
.I1(LIOB33_X0Y115_IOB_X0Y115_I),
.I2(RIOB33_X105Y107_IOB_X1Y107_I),
.I3(CLBLL_L_X4Y112_SLICE_X5Y112_AO5),
.I4(CLBLL_L_X4Y110_SLICE_X5Y110_DO6),
.I5(CLBLL_L_X4Y111_SLICE_X4Y111_CO6),
.O5(CLBLL_L_X4Y113_SLICE_X5Y113_CO5),
.O6(CLBLL_L_X4Y113_SLICE_X5Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00007f1580ea7f15)
  ) CLBLL_L_X4Y113_SLICE_X5Y113_BLUT (
.I0(CLBLL_L_X4Y113_SLICE_X4Y113_AO5),
.I1(LIOB33_X0Y115_IOB_X0Y115_I),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLL_L_X4Y112_SLICE_X5Y112_BO6),
.I4(CLBLL_L_X4Y113_SLICE_X5Y113_CO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y113_SLICE_X5Y113_BO5),
.O6(CLBLL_L_X4Y113_SLICE_X5Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f3f3f3f6699aa55)
  ) CLBLL_L_X4Y113_SLICE_X5Y113_ALUT (
.I0(CLBLL_L_X4Y113_SLICE_X4Y113_AO5),
.I1(LIOB33_X0Y115_IOB_X0Y115_I),
.I2(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I3(CLBLL_L_X4Y112_SLICE_X5Y112_BO6),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y113_SLICE_X5Y113_AO5),
.O6(CLBLL_L_X4Y113_SLICE_X5Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y114_SLICE_X4Y114_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y114_SLICE_X4Y114_DO5),
.O6(CLBLL_L_X4Y114_SLICE_X4Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y114_SLICE_X4Y114_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y114_SLICE_X4Y114_CO5),
.O6(CLBLL_L_X4Y114_SLICE_X4Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0fffffffff)
  ) CLBLL_L_X4Y114_SLICE_X4Y114_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(LIOB33_X0Y115_IOB_X0Y115_I),
.I3(1'b1),
.I4(1'b1),
.I5(RIOB33_X105Y103_IOB_X1Y104_I),
.O5(CLBLL_L_X4Y114_SLICE_X4Y114_BO5),
.O6(CLBLL_L_X4Y114_SLICE_X4Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'he11ee11ee11ee11e)
  ) CLBLL_L_X4Y114_SLICE_X4Y114_ALUT (
.I0(CLBLL_L_X4Y115_SLICE_X4Y115_CO6),
.I1(CLBLL_L_X4Y113_SLICE_X5Y113_BO6),
.I2(CLBLM_R_X3Y112_SLICE_X2Y112_AO6),
.I3(CLBLL_L_X4Y113_SLICE_X5Y113_DO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y114_SLICE_X4Y114_AO5),
.O6(CLBLL_L_X4Y114_SLICE_X4Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y114_SLICE_X5Y114_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y114_SLICE_X5Y114_DO5),
.O6(CLBLL_L_X4Y114_SLICE_X5Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y114_SLICE_X5Y114_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y114_SLICE_X5Y114_CO5),
.O6(CLBLL_L_X4Y114_SLICE_X5Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y114_SLICE_X5Y114_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y114_SLICE_X5Y114_BO5),
.O6(CLBLL_L_X4Y114_SLICE_X5Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h699969992bbb2bbb)
  ) CLBLL_L_X4Y114_SLICE_X5Y114_ALUT (
.I0(CLBLM_R_X7Y111_SLICE_X8Y111_DO6),
.I1(CLBLM_R_X5Y111_SLICE_X7Y111_CO6),
.I2(LIOB33_X0Y113_IOB_X0Y113_I),
.I3(RIOB33_X105Y103_IOB_X1Y104_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y114_SLICE_X5Y114_AO5),
.O6(CLBLL_L_X4Y114_SLICE_X5Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h9699969966966696)
  ) CLBLL_L_X4Y115_SLICE_X4Y115_DLUT (
.I0(CLBLL_L_X4Y115_SLICE_X4Y115_AO6),
.I1(CLBLL_L_X4Y113_SLICE_X5Y113_AO5),
.I2(CLBLM_R_X5Y115_SLICE_X7Y115_AO5),
.I3(CLBLL_L_X4Y115_SLICE_X4Y115_AO5),
.I4(1'b1),
.I5(CLBLL_L_X4Y116_SLICE_X5Y116_DO6),
.O5(CLBLL_L_X4Y115_SLICE_X4Y115_DO5),
.O6(CLBLL_L_X4Y115_SLICE_X4Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h080a0e0f00080a0e)
  ) CLBLL_L_X4Y115_SLICE_X4Y115_CLUT (
.I0(CLBLL_L_X4Y115_SLICE_X4Y115_AO6),
.I1(CLBLM_R_X5Y115_SLICE_X7Y115_AO5),
.I2(CLBLL_L_X4Y113_SLICE_X5Y113_BO5),
.I3(CLBLL_L_X4Y115_SLICE_X4Y115_AO5),
.I4(CLBLL_L_X4Y113_SLICE_X5Y113_AO5),
.I5(CLBLL_L_X4Y116_SLICE_X5Y116_DO6),
.O5(CLBLL_L_X4Y115_SLICE_X4Y115_CO5),
.O6(CLBLL_L_X4Y115_SLICE_X4Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8f0eef8f0e088f0e)
  ) CLBLL_L_X4Y115_SLICE_X4Y115_BLUT (
.I0(CLBLM_R_X5Y115_SLICE_X7Y115_AO5),
.I1(CLBLL_L_X4Y116_SLICE_X5Y116_DO6),
.I2(CLBLL_L_X4Y113_SLICE_X5Y113_AO5),
.I3(CLBLL_L_X4Y114_SLICE_X4Y114_BO6),
.I4(CLBLL_L_X4Y112_SLICE_X5Y112_BO5),
.I5(CLBLL_L_X4Y114_SLICE_X5Y114_AO5),
.O5(CLBLL_L_X4Y115_SLICE_X4Y115_BO5),
.O6(CLBLL_L_X4Y115_SLICE_X4Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h2a2abfbfc03fc03f)
  ) CLBLL_L_X4Y115_SLICE_X4Y115_ALUT (
.I0(CLBLL_L_X4Y114_SLICE_X5Y114_AO5),
.I1(RIOB33_X105Y103_IOB_X1Y104_I),
.I2(LIOB33_X0Y115_IOB_X0Y115_I),
.I3(CLBLL_L_X4Y112_SLICE_X5Y112_CO6),
.I4(CLBLL_L_X4Y112_SLICE_X5Y112_BO5),
.I5(1'b1),
.O5(CLBLL_L_X4Y115_SLICE_X4Y115_AO5),
.O6(CLBLL_L_X4Y115_SLICE_X4Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y115_SLICE_X5Y115_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y115_SLICE_X5Y115_DO5),
.O6(CLBLL_L_X4Y115_SLICE_X5Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y115_SLICE_X5Y115_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y115_SLICE_X5Y115_CO5),
.O6(CLBLL_L_X4Y115_SLICE_X5Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y115_SLICE_X5Y115_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y115_SLICE_X5Y115_BO5),
.O6(CLBLL_L_X4Y115_SLICE_X5Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88887777a50fa50f)
  ) CLBLL_L_X4Y115_SLICE_X5Y115_ALUT (
.I0(LIOB33_X0Y113_IOB_X0Y113_I),
.I1(RIOB33_X105Y101_IOB_X1Y102_I),
.I2(CLBLM_R_X7Y114_SLICE_X9Y114_DO6),
.I3(RIOB33_X105Y103_IOB_X1Y103_I),
.I4(CLBLM_R_X7Y114_SLICE_X8Y114_BO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y115_SLICE_X5Y115_AO5),
.O6(CLBLL_L_X4Y115_SLICE_X5Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y116_SLICE_X4Y116_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y116_SLICE_X4Y116_DO5),
.O6(CLBLL_L_X4Y116_SLICE_X4Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h55aa55aa55aa55aa)
  ) CLBLL_L_X4Y116_SLICE_X4Y116_CLUT (
.I0(CLBLL_L_X4Y115_SLICE_X4Y115_BO6),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLL_L_X4Y113_SLICE_X5Y113_BO5),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y116_SLICE_X4Y116_CO5),
.O6(CLBLL_L_X4Y116_SLICE_X4Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3c3c3c3c3c3c3c3c)
  ) CLBLL_L_X4Y116_SLICE_X4Y116_BLUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y116_SLICE_X5Y116_DO6),
.I2(CLBLM_R_X5Y115_SLICE_X7Y115_DO6),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y116_SLICE_X4Y116_BO5),
.O6(CLBLL_L_X4Y116_SLICE_X4Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h33ff33ff55ff55ff)
  ) CLBLL_L_X4Y116_SLICE_X4Y116_ALUT (
.I0(RIOB33_X105Y101_IOB_X1Y102_I),
.I1(LIOB33_X0Y113_IOB_X0Y114_I),
.I2(1'b1),
.I3(LIOB33_X0Y115_IOB_X0Y115_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y116_SLICE_X4Y116_AO5),
.O6(CLBLL_L_X4Y116_SLICE_X4Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h80e80080feffe8fe)
  ) CLBLL_L_X4Y116_SLICE_X5Y116_DLUT (
.I0(CLBLM_R_X7Y114_SLICE_X8Y114_CO6),
.I1(CLBLL_L_X4Y116_SLICE_X4Y116_AO5),
.I2(CLBLM_R_X5Y116_SLICE_X6Y116_DO6),
.I3(CLBLL_L_X4Y115_SLICE_X5Y115_AO5),
.I4(CLBLM_R_X5Y116_SLICE_X7Y116_AO6),
.I5(CLBLM_R_X5Y115_SLICE_X7Y115_AO6),
.O5(CLBLL_L_X4Y116_SLICE_X5Y116_DO5),
.O6(CLBLL_L_X4Y116_SLICE_X5Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6999966696669666)
  ) CLBLL_L_X4Y116_SLICE_X5Y116_CLUT (
.I0(CLBLM_R_X7Y116_SLICE_X9Y116_AO6),
.I1(CLBLM_R_X7Y116_SLICE_X8Y116_AO6),
.I2(LIOB33_X0Y113_IOB_X0Y113_I),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(LIOB33_X0Y115_IOB_X0Y116_I),
.I5(LIOB33_X0Y115_IOB_X0Y115_I),
.O5(CLBLL_L_X4Y116_SLICE_X5Y116_CO5),
.O6(CLBLL_L_X4Y116_SLICE_X5Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h99669966d24b2db4)
  ) CLBLL_L_X4Y116_SLICE_X5Y116_BLUT (
.I0(CLBLM_R_X5Y116_SLICE_X7Y116_BO6),
.I1(CLBLM_R_X5Y116_SLICE_X6Y116_AO6),
.I2(CLBLM_R_X5Y116_SLICE_X7Y116_AO6),
.I3(CLBLM_R_X7Y116_SLICE_X8Y116_CO6),
.I4(CLBLM_R_X5Y115_SLICE_X7Y115_BO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y116_SLICE_X5Y116_BO5),
.O6(CLBLL_L_X4Y116_SLICE_X5Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc3c33c3c956aa956)
  ) CLBLL_L_X4Y116_SLICE_X5Y116_ALUT (
.I0(CLBLM_R_X5Y115_SLICE_X6Y115_DO6),
.I1(CLBLM_R_X5Y114_SLICE_X6Y114_CO6),
.I2(CLBLM_R_X5Y115_SLICE_X6Y115_CO6),
.I3(CLBLM_R_X7Y116_SLICE_X8Y116_BO6),
.I4(CLBLL_L_X4Y116_SLICE_X5Y116_CO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y116_SLICE_X5Y116_AO5),
.O6(CLBLL_L_X4Y116_SLICE_X5Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y104_SLICE_X10Y104_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y104_SLICE_X10Y104_DO5),
.O6(CLBLM_L_X8Y104_SLICE_X10Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y104_SLICE_X10Y104_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y104_SLICE_X10Y104_CO5),
.O6(CLBLM_L_X8Y104_SLICE_X10Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y104_SLICE_X10Y104_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y104_SLICE_X10Y104_BO5),
.O6(CLBLM_L_X8Y104_SLICE_X10Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0a5a728822d27288)
  ) CLBLM_L_X8Y104_SLICE_X10Y104_ALUT (
.I0(RIOB33_X105Y113_IOB_X1Y113_I),
.I1(RIOB33_X105Y103_IOB_X1Y104_I),
.I2(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I3(RIOB33_X105Y101_IOB_X1Y102_I),
.I4(RIOB33_X105Y103_IOB_X1Y103_I),
.I5(RIOB33_X105Y111_IOB_X1Y112_I),
.O5(CLBLM_L_X8Y104_SLICE_X10Y104_AO5),
.O6(CLBLM_L_X8Y104_SLICE_X10Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y104_SLICE_X11Y104_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y104_SLICE_X11Y104_DO5),
.O6(CLBLM_L_X8Y104_SLICE_X11Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y104_SLICE_X11Y104_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y104_SLICE_X11Y104_CO5),
.O6(CLBLM_L_X8Y104_SLICE_X11Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y104_SLICE_X11Y104_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y104_SLICE_X11Y104_BO5),
.O6(CLBLM_L_X8Y104_SLICE_X11Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y104_SLICE_X11Y104_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y104_SLICE_X11Y104_AO5),
.O6(CLBLM_L_X8Y104_SLICE_X11Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5f7fffff171f5fff)
  ) CLBLM_L_X8Y105_SLICE_X10Y105_DLUT (
.I0(RIOB33_X105Y109_IOB_X1Y110_I),
.I1(LIOB33_X0Y101_IOB_X0Y101_I),
.I2(LIOB33_X0Y101_IOB_X0Y102_I),
.I3(LIOB33_X0Y103_IOB_X0Y104_I),
.I4(RIOB33_X105Y111_IOB_X1Y111_I),
.I5(CLBLM_L_X10Y105_SLICE_X12Y105_BO6),
.O5(CLBLM_L_X8Y105_SLICE_X10Y105_DO5),
.O6(CLBLM_L_X8Y105_SLICE_X10Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafaf5f5b2a07150)
  ) CLBLM_L_X8Y105_SLICE_X10Y105_CLUT (
.I0(CLBLM_L_X10Y108_SLICE_X13Y108_AO6),
.I1(CLBLM_L_X8Y104_SLICE_X10Y104_AO6),
.I2(CLBLM_L_X8Y105_SLICE_X10Y105_AO5),
.I3(CLBLM_L_X8Y105_SLICE_X10Y105_AO6),
.I4(CLBLM_L_X10Y107_SLICE_X13Y107_BO6),
.I5(CLBLM_L_X8Y107_SLICE_X10Y107_BO6),
.O5(CLBLM_L_X8Y105_SLICE_X10Y105_CO5),
.O6(CLBLM_L_X8Y105_SLICE_X10Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h55a6aa59aa5955a6)
  ) CLBLM_L_X8Y105_SLICE_X10Y105_BLUT (
.I0(CLBLM_L_X10Y107_SLICE_X13Y107_BO6),
.I1(CLBLM_L_X8Y105_SLICE_X10Y105_AO6),
.I2(CLBLM_L_X8Y104_SLICE_X10Y104_AO6),
.I3(CLBLM_L_X8Y107_SLICE_X10Y107_BO6),
.I4(CLBLM_L_X10Y108_SLICE_X13Y108_AO6),
.I5(CLBLM_L_X8Y105_SLICE_X10Y105_AO5),
.O5(CLBLM_L_X8Y105_SLICE_X10Y105_BO5),
.O6(CLBLM_L_X8Y105_SLICE_X10Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h33ff33ff55ff55ff)
  ) CLBLM_L_X8Y105_SLICE_X10Y105_ALUT (
.I0(LIOB33_X0Y101_IOB_X0Y102_I),
.I1(LIOB33_X0Y101_IOB_X0Y101_I),
.I2(1'b1),
.I3(RIOB33_X105Y101_IOB_X1Y102_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y105_SLICE_X10Y105_AO5),
.O6(CLBLM_L_X8Y105_SLICE_X10Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y105_SLICE_X11Y105_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y105_SLICE_X11Y105_DO5),
.O6(CLBLM_L_X8Y105_SLICE_X11Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y105_SLICE_X11Y105_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y105_SLICE_X11Y105_CO5),
.O6(CLBLM_L_X8Y105_SLICE_X11Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y105_SLICE_X11Y105_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y105_SLICE_X11Y105_BO5),
.O6(CLBLM_L_X8Y105_SLICE_X11Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hb2a0dfdf5ddfffff)
  ) CLBLM_L_X8Y105_SLICE_X11Y105_ALUT (
.I0(LIOB33_X0Y101_IOB_X0Y102_I),
.I1(CLBLM_L_X10Y105_SLICE_X12Y105_BO6),
.I2(RIOB33_X105Y109_IOB_X1Y110_I),
.I3(LIOB33_X0Y101_IOB_X0Y101_I),
.I4(RIOB33_X105Y111_IOB_X1Y111_I),
.I5(LIOB33_X0Y103_IOB_X0Y104_I),
.O5(CLBLM_L_X8Y105_SLICE_X11Y105_AO5),
.O6(CLBLM_L_X8Y105_SLICE_X11Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hd24baaff2db45500)
  ) CLBLM_L_X8Y106_SLICE_X10Y106_DLUT (
.I0(CLBLM_L_X10Y105_SLICE_X12Y105_AO6),
.I1(LIOB33_X0Y105_IOB_X0Y106_I),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(CLBLM_L_X10Y106_SLICE_X12Y106_AO6),
.I4(RIOB33_X105Y109_IOB_X1Y109_I),
.I5(CLBLM_L_X8Y106_SLICE_X10Y106_BO6),
.O5(CLBLM_L_X8Y106_SLICE_X10Y106_DO5),
.O6(CLBLM_L_X8Y106_SLICE_X10Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h020baaff2fbfffff)
  ) CLBLM_L_X8Y106_SLICE_X10Y106_CLUT (
.I0(CLBLM_L_X10Y105_SLICE_X12Y105_AO6),
.I1(LIOB33_X0Y105_IOB_X0Y106_I),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(CLBLM_L_X10Y106_SLICE_X12Y106_AO6),
.I4(RIOB33_X105Y109_IOB_X1Y109_I),
.I5(CLBLM_L_X8Y106_SLICE_X10Y106_BO6),
.O5(CLBLM_L_X8Y106_SLICE_X10Y106_CO5),
.O6(CLBLM_L_X8Y106_SLICE_X10Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'he69eaa224c340088)
  ) CLBLM_L_X8Y106_SLICE_X10Y106_BLUT (
.I0(RIOB33_X105Y109_IOB_X1Y110_I),
.I1(LIOB33_X0Y105_IOB_X0Y105_I),
.I2(LIOB33_X0Y103_IOB_X0Y104_I),
.I3(CLBLM_L_X8Y105_SLICE_X10Y105_DO6),
.I4(RIOB33_X105Y111_IOB_X1Y111_I),
.I5(LIOB33_X0Y105_IOB_X0Y106_I),
.O5(CLBLM_L_X8Y106_SLICE_X10Y106_BO5),
.O6(CLBLM_L_X8Y106_SLICE_X10Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h4ddd8eee8eee8eee)
  ) CLBLM_L_X8Y106_SLICE_X10Y106_ALUT (
.I0(CLBLM_R_X7Y106_SLICE_X9Y106_CO6),
.I1(CLBLM_R_X7Y105_SLICE_X8Y105_DO6),
.I2(LIOB33_X0Y103_IOB_X0Y104_I),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(RIOB33_X105Y101_IOB_X1Y101_I),
.I5(LIOB33_X0Y101_IOB_X0Y102_I),
.O5(CLBLM_L_X8Y106_SLICE_X10Y106_AO5),
.O6(CLBLM_L_X8Y106_SLICE_X10Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y106_SLICE_X11Y106_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y106_SLICE_X11Y106_DO5),
.O6(CLBLM_L_X8Y106_SLICE_X11Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y106_SLICE_X11Y106_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y106_SLICE_X11Y106_CO5),
.O6(CLBLM_L_X8Y106_SLICE_X11Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y106_SLICE_X11Y106_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y106_SLICE_X11Y106_BO5),
.O6(CLBLM_L_X8Y106_SLICE_X11Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996c33ca55a0ff0)
  ) CLBLM_L_X8Y106_SLICE_X11Y106_ALUT (
.I0(RIOB33_X105Y109_IOB_X1Y110_I),
.I1(RIOB33_X105Y109_IOB_X1Y109_I),
.I2(CLBLM_L_X8Y105_SLICE_X11Y105_AO6),
.I3(CLBLM_L_X10Y105_SLICE_X12Y105_AO6),
.I4(LIOB33_X0Y105_IOB_X0Y105_I),
.I5(LIOB33_X0Y105_IOB_X0Y106_I),
.O5(CLBLM_L_X8Y106_SLICE_X11Y106_AO5),
.O6(CLBLM_L_X8Y106_SLICE_X11Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h33ccff00d92615ea)
  ) CLBLM_L_X8Y107_SLICE_X10Y107_DLUT (
.I0(CLBLM_L_X8Y104_SLICE_X10Y104_AO6),
.I1(LIOB33_X0Y101_IOB_X0Y101_I),
.I2(RIOB33_X105Y101_IOB_X1Y102_I),
.I3(CLBLM_L_X10Y107_SLICE_X13Y107_BO6),
.I4(RIOB33_X105Y103_IOB_X1Y103_I),
.I5(CLBLM_L_X8Y107_SLICE_X10Y107_BO6),
.O5(CLBLM_L_X8Y107_SLICE_X10Y107_DO5),
.O6(CLBLM_L_X8Y107_SLICE_X10Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h4bb4d22db44b2dd2)
  ) CLBLM_L_X8Y107_SLICE_X10Y107_CLUT (
.I0(CLBLM_L_X8Y107_SLICE_X10Y107_AO6),
.I1(CLBLM_L_X8Y105_SLICE_X10Y105_BO6),
.I2(CLBLM_L_X10Y108_SLICE_X13Y108_BO6),
.I3(CLBLM_L_X12Y108_SLICE_X16Y108_AO6),
.I4(CLBLM_R_X7Y104_SLICE_X9Y104_DO6),
.I5(CLBLM_L_X8Y105_SLICE_X10Y105_CO6),
.O5(CLBLM_L_X8Y107_SLICE_X10Y107_CO5),
.O6(CLBLM_L_X8Y107_SLICE_X10Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h260c0a0a26260000)
  ) CLBLM_L_X8Y107_SLICE_X10Y107_BLUT (
.I0(RIOB33_X105Y113_IOB_X1Y113_I),
.I1(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I2(RIOB33_X105Y101_IOB_X1Y102_I),
.I3(RIOB33_X105Y111_IOB_X1Y112_I),
.I4(RIOB33_X105Y103_IOB_X1Y103_I),
.I5(RIOB33_X105Y103_IOB_X1Y104_I),
.O5(CLBLM_L_X8Y107_SLICE_X10Y107_BO5),
.O6(CLBLM_L_X8Y107_SLICE_X10Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0fff0fff0f0fffff)
  ) CLBLM_L_X8Y107_SLICE_X10Y107_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(RIOB33_X105Y101_IOB_X1Y101_I),
.I3(LIOB33_X0Y103_IOB_X0Y104_I),
.I4(LIOB33_X0Y105_IOB_X0Y105_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y107_SLICE_X10Y107_AO5),
.O6(CLBLM_L_X8Y107_SLICE_X10Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y107_SLICE_X11Y107_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y107_SLICE_X11Y107_DO5),
.O6(CLBLM_L_X8Y107_SLICE_X11Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0080000000000000)
  ) CLBLM_L_X8Y107_SLICE_X11Y107_CLUT (
.I0(LIOB33_X0Y103_IOB_X0Y104_I),
.I1(CLBLM_L_X10Y107_SLICE_X13Y107_BO6),
.I2(CLBLM_L_X10Y107_SLICE_X12Y107_DO6),
.I3(CLBLL_L_X2Y107_SLICE_X0Y107_CO6),
.I4(RIOB33_X105Y105_IOB_X1Y106_I),
.I5(CLBLM_L_X12Y107_SLICE_X16Y107_AO6),
.O5(CLBLM_L_X8Y107_SLICE_X11Y107_CO5),
.O6(CLBLM_L_X8Y107_SLICE_X11Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hd72877888877d728)
  ) CLBLM_L_X8Y107_SLICE_X11Y107_BLUT (
.I0(LIOB33_X0Y101_IOB_X0Y102_I),
.I1(RIOB33_X105Y101_IOB_X1Y102_I),
.I2(RIOB33_X105Y101_IOB_X1Y101_I),
.I3(CLBLM_L_X8Y107_SLICE_X10Y107_DO6),
.I4(CLBLM_L_X8Y107_SLICE_X11Y107_AO6),
.I5(CLBLM_R_X7Y106_SLICE_X9Y106_AO5),
.O5(CLBLM_L_X8Y107_SLICE_X11Y107_BO5),
.O6(CLBLM_L_X8Y107_SLICE_X11Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa0055ffccccddff)
  ) CLBLM_L_X8Y107_SLICE_X11Y107_ALUT (
.I0(RIOB33_X105Y101_IOB_X1Y102_I),
.I1(CLBLM_L_X8Y107_SLICE_X10Y107_BO6),
.I2(1'b1),
.I3(LIOB33_X0Y101_IOB_X0Y101_I),
.I4(CLBLM_L_X8Y104_SLICE_X10Y104_AO6),
.I5(1'b1),
.O5(CLBLM_L_X8Y107_SLICE_X11Y107_AO5),
.O6(CLBLM_L_X8Y107_SLICE_X11Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'he6192ad5738cbf40)
  ) CLBLM_L_X8Y108_SLICE_X10Y108_DLUT (
.I0(CLBLM_L_X8Y106_SLICE_X10Y106_AO6),
.I1(LIOB33_X0Y105_IOB_X0Y105_I),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(CLBLM_L_X8Y107_SLICE_X10Y107_CO6),
.I4(RIOB33_X105Y101_IOB_X1Y101_I),
.I5(CLBLM_L_X8Y108_SLICE_X10Y108_BO6),
.O5(CLBLM_L_X8Y108_SLICE_X10Y108_DO5),
.O6(CLBLM_L_X8Y108_SLICE_X10Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'he8b2c030fcf3e8b2)
  ) CLBLM_L_X8Y108_SLICE_X10Y108_CLUT (
.I0(CLBLM_L_X8Y106_SLICE_X10Y106_AO6),
.I1(CLBLM_L_X8Y107_SLICE_X10Y107_AO5),
.I2(CLBLM_L_X8Y108_SLICE_X11Y108_AO6),
.I3(CLBLM_L_X8Y107_SLICE_X10Y107_CO6),
.I4(CLBLM_R_X7Y108_SLICE_X9Y108_AO6),
.I5(CLBLM_L_X8Y108_SLICE_X10Y108_BO6),
.O5(CLBLM_L_X8Y108_SLICE_X10Y108_CO5),
.O6(CLBLM_L_X8Y108_SLICE_X10Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996a55a996655aa)
  ) CLBLM_L_X8Y108_SLICE_X10Y108_BLUT (
.I0(CLBLM_R_X7Y104_SLICE_X9Y104_DO6),
.I1(LIOB33_X0Y101_IOB_X0Y102_I),
.I2(RIOB33_X105Y101_IOB_X1Y101_I),
.I3(CLBLM_L_X8Y107_SLICE_X10Y107_DO6),
.I4(RIOB33_X105Y101_IOB_X1Y102_I),
.I5(LIOB33_X0Y103_IOB_X0Y104_I),
.O5(CLBLM_L_X8Y108_SLICE_X10Y108_BO5),
.O6(CLBLM_L_X8Y108_SLICE_X10Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h693cc36996c33c96)
  ) CLBLM_L_X8Y108_SLICE_X10Y108_ALUT (
.I0(CLBLM_R_X7Y108_SLICE_X9Y108_AO6),
.I1(CLBLM_L_X8Y107_SLICE_X10Y107_AO5),
.I2(CLBLM_L_X8Y108_SLICE_X11Y108_AO6),
.I3(CLBLM_L_X8Y108_SLICE_X10Y108_BO6),
.I4(CLBLM_L_X8Y106_SLICE_X10Y106_AO6),
.I5(CLBLM_L_X8Y107_SLICE_X10Y107_CO6),
.O5(CLBLM_L_X8Y108_SLICE_X10Y108_AO5),
.O6(CLBLM_L_X8Y108_SLICE_X10Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7f15ff3fd540ffc0)
  ) CLBLM_L_X8Y108_SLICE_X11Y108_DLUT (
.I0(LIOB33_X0Y105_IOB_X0Y105_I),
.I1(LIOB33_X0Y103_IOB_X0Y104_I),
.I2(RIOB33_X105Y101_IOB_X1Y101_I),
.I3(CLBLM_L_X8Y106_SLICE_X10Y106_AO6),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(CLBLM_L_X8Y107_SLICE_X11Y107_BO6),
.O5(CLBLM_L_X8Y108_SLICE_X11Y108_DO5),
.O6(CLBLM_L_X8Y108_SLICE_X11Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6fff0666cfff0ccc)
  ) CLBLM_L_X8Y108_SLICE_X11Y108_CLUT (
.I0(RIOB33_X105Y101_IOB_X1Y102_I),
.I1(CLBLM_L_X8Y107_SLICE_X10Y107_DO6),
.I2(RIOB33_X105Y101_IOB_X1Y101_I),
.I3(LIOB33_X0Y103_IOB_X0Y104_I),
.I4(CLBLM_R_X7Y104_SLICE_X9Y104_DO6),
.I5(LIOB33_X0Y101_IOB_X0Y102_I),
.O5(CLBLM_L_X8Y108_SLICE_X11Y108_CO5),
.O6(CLBLM_L_X8Y108_SLICE_X11Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996c33c96963c3c)
  ) CLBLM_L_X8Y108_SLICE_X11Y108_BLUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(CLBLM_L_X8Y107_SLICE_X11Y107_BO6),
.I2(CLBLM_L_X8Y106_SLICE_X10Y106_AO6),
.I3(RIOB33_X105Y101_IOB_X1Y101_I),
.I4(LIOB33_X0Y105_IOB_X0Y105_I),
.I5(LIOB33_X0Y103_IOB_X0Y104_I),
.O5(CLBLM_L_X8Y108_SLICE_X11Y108_BO5),
.O6(CLBLM_L_X8Y108_SLICE_X11Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5f5f5f5f0fff0fff)
  ) CLBLM_L_X8Y108_SLICE_X11Y108_ALUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(1'b1),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(RIOB33_X105Y101_IOB_X1Y101_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y108_SLICE_X11Y108_AO5),
.O6(CLBLM_L_X8Y108_SLICE_X11Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y109_SLICE_X10Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y109_SLICE_X10Y109_DO5),
.O6(CLBLM_L_X8Y109_SLICE_X10Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996a55ac33c0ff0)
  ) CLBLM_L_X8Y109_SLICE_X10Y109_CLUT (
.I0(LIOB33_X0Y107_IOB_X0Y107_I),
.I1(LIOB33_X0Y115_IOB_X0Y116_I),
.I2(CLBLM_L_X8Y109_SLICE_X11Y109_DO6),
.I3(CLBLM_R_X7Y109_SLICE_X9Y109_DO6),
.I4(LIOB33_X0Y107_IOB_X0Y108_I),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLM_L_X8Y109_SLICE_X10Y109_CO5),
.O6(CLBLM_L_X8Y109_SLICE_X10Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc639639caf50af50)
  ) CLBLM_L_X8Y109_SLICE_X10Y109_BLUT (
.I0(CLBLM_L_X10Y106_SLICE_X13Y106_CO6),
.I1(LIOB33_X0Y107_IOB_X0Y108_I),
.I2(CLBLM_L_X8Y106_SLICE_X11Y106_AO6),
.I3(CLBLM_L_X8Y106_SLICE_X10Y106_DO6),
.I4(LIOB33_X0Y107_IOB_X0Y107_I),
.I5(RIOB33_X105Y107_IOB_X1Y108_I),
.O5(CLBLM_L_X8Y109_SLICE_X10Y109_BO5),
.O6(CLBLM_L_X8Y109_SLICE_X10Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h02af23af3bffbfff)
  ) CLBLM_L_X8Y109_SLICE_X10Y109_ALUT (
.I0(CLBLM_L_X10Y106_SLICE_X13Y106_CO6),
.I1(LIOB33_X0Y107_IOB_X0Y108_I),
.I2(CLBLM_L_X8Y106_SLICE_X11Y106_AO6),
.I3(RIOB33_X105Y107_IOB_X1Y108_I),
.I4(LIOB33_X0Y107_IOB_X0Y107_I),
.I5(CLBLM_L_X8Y106_SLICE_X10Y106_DO6),
.O5(CLBLM_L_X8Y109_SLICE_X10Y109_AO5),
.O6(CLBLM_L_X8Y109_SLICE_X10Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hd27887877878d278)
  ) CLBLM_L_X8Y109_SLICE_X11Y109_DLUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(RIOB33_X105Y101_IOB_X1Y101_I),
.I2(CLBLM_L_X10Y109_SLICE_X12Y109_DO6),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(CLBLM_L_X8Y108_SLICE_X11Y108_DO6),
.I5(CLBLM_L_X8Y109_SLICE_X11Y109_BO6),
.O5(CLBLM_L_X8Y109_SLICE_X11Y109_DO5),
.O6(CLBLM_L_X8Y109_SLICE_X11Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h4cdfdf4cdfdf4c4c)
  ) CLBLM_L_X8Y109_SLICE_X11Y109_CLUT (
.I0(LIOB33_X0Y115_IOB_X0Y116_I),
.I1(CLBLM_R_X7Y109_SLICE_X9Y109_DO6),
.I2(LIOB33_X0Y107_IOB_X0Y108_I),
.I3(LIOB33_X0Y107_IOB_X0Y107_I),
.I4(CLBLM_L_X8Y109_SLICE_X11Y109_DO6),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLM_L_X8Y109_SLICE_X11Y109_CO5),
.O6(CLBLM_L_X8Y109_SLICE_X11Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h69c3963c993366cc)
  ) CLBLM_L_X8Y109_SLICE_X11Y109_BLUT (
.I0(LIOB33_X0Y105_IOB_X0Y105_I),
.I1(CLBLM_L_X10Y107_SLICE_X12Y107_CO6),
.I2(RIOB33_X105Y101_IOB_X1Y102_I),
.I3(RIOB33_X105Y101_IOB_X1Y101_I),
.I4(CLBLM_L_X8Y108_SLICE_X11Y108_CO6),
.I5(LIOB33_X0Y103_IOB_X0Y104_I),
.O5(CLBLM_L_X8Y109_SLICE_X11Y109_BO5),
.O6(CLBLM_L_X8Y109_SLICE_X11Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5f5f5f5f0fff0fff)
  ) CLBLM_L_X8Y109_SLICE_X11Y109_ALUT (
.I0(LIOB33_X0Y115_IOB_X0Y116_I),
.I1(1'b1),
.I2(LIOB33_X0Y109_IOB_X0Y109_I),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y109_SLICE_X11Y109_AO5),
.O6(CLBLM_L_X8Y109_SLICE_X11Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'he765189a4dcfb230)
  ) CLBLM_L_X8Y110_SLICE_X10Y110_DLUT (
.I0(LIOB33_X0Y107_IOB_X0Y108_I),
.I1(CLBLM_R_X7Y109_SLICE_X9Y109_DO6),
.I2(CLBLM_L_X8Y110_SLICE_X11Y110_BO6),
.I3(LIOB33_X0Y115_IOB_X0Y116_I),
.I4(CLBLM_L_X10Y110_SLICE_X12Y110_DO6),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLM_L_X8Y110_SLICE_X10Y110_DO5),
.O6(CLBLM_L_X8Y110_SLICE_X10Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h10f531f573fff7ff)
  ) CLBLM_L_X8Y110_SLICE_X10Y110_CLUT (
.I0(CLBLM_L_X8Y110_SLICE_X10Y110_AO6),
.I1(LIOB33_X0Y109_IOB_X0Y109_I),
.I2(CLBLM_L_X10Y109_SLICE_X12Y109_BO6),
.I3(RIOB33_X105Y107_IOB_X1Y107_I),
.I4(LIOB33_X0Y107_IOB_X0Y108_I),
.I5(CLBLM_L_X8Y109_SLICE_X10Y109_BO6),
.O5(CLBLM_L_X8Y110_SLICE_X10Y110_CO5),
.O6(CLBLM_L_X8Y110_SLICE_X10Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'he619758a4cb3df20)
  ) CLBLM_L_X8Y110_SLICE_X10Y110_BLUT (
.I0(RIOB33_X105Y107_IOB_X1Y107_I),
.I1(CLBLM_L_X10Y109_SLICE_X12Y109_BO6),
.I2(LIOB33_X0Y107_IOB_X0Y108_I),
.I3(CLBLM_L_X8Y109_SLICE_X10Y109_BO6),
.I4(CLBLM_L_X8Y110_SLICE_X10Y110_AO6),
.I5(LIOB33_X0Y109_IOB_X0Y109_I),
.O5(CLBLM_L_X8Y110_SLICE_X10Y110_BO5),
.O6(CLBLM_L_X8Y110_SLICE_X10Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h7887788777777777)
  ) CLBLM_L_X8Y110_SLICE_X10Y110_ALUT (
.I0(LIOB33_X0Y107_IOB_X0Y107_I),
.I1(RIOB33_X105Y107_IOB_X1Y108_I),
.I2(CLBLM_L_X8Y106_SLICE_X11Y106_AO6),
.I3(CLBLM_L_X10Y106_SLICE_X13Y106_CO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y110_SLICE_X10Y110_AO5),
.O6(CLBLM_L_X8Y110_SLICE_X10Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'he8a08e0afae8af8e)
  ) CLBLM_L_X8Y110_SLICE_X11Y110_DLUT (
.I0(CLBLM_L_X8Y109_SLICE_X11Y109_AO6),
.I1(CLBLM_R_X7Y109_SLICE_X8Y109_AO5),
.I2(CLBLM_L_X10Y110_SLICE_X12Y110_DO6),
.I3(CLBLM_R_X7Y109_SLICE_X9Y109_DO6),
.I4(CLBLM_L_X10Y111_SLICE_X13Y111_AO6),
.I5(CLBLM_L_X8Y110_SLICE_X11Y110_BO6),
.O5(CLBLM_L_X8Y110_SLICE_X11Y110_DO5),
.O6(CLBLM_L_X8Y110_SLICE_X11Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h377f15157f7f377f)
  ) CLBLM_L_X8Y110_SLICE_X11Y110_CLUT (
.I0(CLBLM_L_X10Y108_SLICE_X12Y108_BO6),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(LIOB33_X0Y105_IOB_X0Y106_I),
.I4(CLBLM_L_X8Y108_SLICE_X11Y108_DO6),
.I5(CLBLM_L_X8Y109_SLICE_X11Y109_BO6),
.O5(CLBLM_L_X8Y110_SLICE_X11Y110_CO5),
.O6(CLBLM_L_X8Y110_SLICE_X11Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc6af395063af9c50)
  ) CLBLM_L_X8Y110_SLICE_X11Y110_BLUT (
.I0(CLBLM_L_X8Y108_SLICE_X11Y108_DO6),
.I1(LIOB33_X0Y107_IOB_X0Y107_I),
.I2(CLBLM_L_X8Y109_SLICE_X11Y109_BO6),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(CLBLM_L_X10Y108_SLICE_X12Y108_BO6),
.I5(LIOB33_X0Y105_IOB_X0Y106_I),
.O5(CLBLM_L_X8Y110_SLICE_X11Y110_BO5),
.O6(CLBLM_L_X8Y110_SLICE_X11Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h39c6c6399c63639c)
  ) CLBLM_L_X8Y110_SLICE_X11Y110_ALUT (
.I0(CLBLM_L_X8Y110_SLICE_X11Y110_BO6),
.I1(CLBLM_L_X10Y111_SLICE_X13Y111_AO6),
.I2(CLBLM_R_X7Y109_SLICE_X9Y109_DO6),
.I3(CLBLM_L_X8Y109_SLICE_X11Y109_AO6),
.I4(CLBLM_L_X10Y110_SLICE_X12Y110_DO6),
.I5(CLBLM_R_X7Y109_SLICE_X8Y109_AO5),
.O5(CLBLM_L_X8Y110_SLICE_X11Y110_AO5),
.O6(CLBLM_L_X8Y110_SLICE_X11Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h17ff03773fff1777)
  ) CLBLM_L_X8Y111_SLICE_X10Y111_DLUT (
.I0(CLBLM_L_X8Y111_SLICE_X10Y111_AO6),
.I1(CLBLM_L_X8Y110_SLICE_X10Y110_BO6),
.I2(LIOB33_X0Y109_IOB_X0Y110_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_L_X10Y111_SLICE_X12Y111_AO5),
.I5(LIOB33_X0Y109_IOB_X0Y109_I),
.O5(CLBLM_L_X8Y111_SLICE_X10Y111_DO5),
.O6(CLBLM_L_X8Y111_SLICE_X10Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h69c33c69963cc396)
  ) CLBLM_L_X8Y111_SLICE_X10Y111_CLUT (
.I0(CLBLM_R_X7Y109_SLICE_X8Y109_CO6),
.I1(CLBLM_L_X8Y112_SLICE_X10Y112_AO5),
.I2(CLBLM_L_X8Y110_SLICE_X11Y110_DO6),
.I3(CLBLM_R_X7Y110_SLICE_X9Y110_AO5),
.I4(CLBLM_L_X8Y110_SLICE_X11Y110_AO6),
.I5(CLBLM_L_X10Y110_SLICE_X13Y110_BO6),
.O5(CLBLM_L_X8Y111_SLICE_X10Y111_CO5),
.O6(CLBLM_L_X8Y111_SLICE_X10Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc369693ca5a5f0f0)
  ) CLBLM_L_X8Y111_SLICE_X10Y111_BLUT (
.I0(CLBLM_L_X10Y111_SLICE_X12Y111_AO5),
.I1(LIOB33_X0Y109_IOB_X0Y110_I),
.I2(CLBLM_L_X8Y110_SLICE_X10Y110_BO6),
.I3(LIOB33_X0Y109_IOB_X0Y109_I),
.I4(CLBLM_L_X8Y111_SLICE_X10Y111_AO6),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X8Y111_SLICE_X10Y111_BO5),
.O6(CLBLM_L_X8Y111_SLICE_X10Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3cf0c30f33ff33ff)
  ) CLBLM_L_X8Y111_SLICE_X10Y111_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y107_IOB_X1Y107_I),
.I2(CLBLM_L_X8Y110_SLICE_X10Y110_AO6),
.I3(LIOB33_X0Y107_IOB_X0Y108_I),
.I4(CLBLM_L_X10Y109_SLICE_X12Y109_BO6),
.I5(1'b1),
.O5(CLBLM_L_X8Y111_SLICE_X10Y111_AO5),
.O6(CLBLM_L_X8Y111_SLICE_X10Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y111_SLICE_X11Y111_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y111_SLICE_X11Y111_DO5),
.O6(CLBLM_L_X8Y111_SLICE_X11Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y111_SLICE_X11Y111_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y111_SLICE_X11Y111_CO5),
.O6(CLBLM_L_X8Y111_SLICE_X11Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y111_SLICE_X11Y111_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y111_SLICE_X11Y111_BO5),
.O6(CLBLM_L_X8Y111_SLICE_X11Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y111_SLICE_X11Y111_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y111_SLICE_X11Y111_AO5),
.O6(CLBLM_L_X8Y111_SLICE_X11Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y112_SLICE_X10Y112_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y112_SLICE_X10Y112_DO5),
.O6(CLBLM_L_X8Y112_SLICE_X10Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5a96a56996a5695a)
  ) CLBLM_L_X8Y112_SLICE_X10Y112_CLUT (
.I0(CLBLM_L_X8Y112_SLICE_X10Y112_AO6),
.I1(CLBLM_L_X10Y110_SLICE_X13Y110_BO6),
.I2(CLBLM_R_X11Y112_SLICE_X14Y112_AO6),
.I3(CLBLM_L_X8Y112_SLICE_X10Y112_AO5),
.I4(CLBLM_L_X10Y110_SLICE_X13Y110_DO6),
.I5(CLBLM_L_X8Y110_SLICE_X11Y110_DO6),
.O5(CLBLM_L_X8Y112_SLICE_X10Y112_CO5),
.O6(CLBLM_L_X8Y112_SLICE_X10Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha96a695a599a99aa)
  ) CLBLM_L_X8Y112_SLICE_X10Y112_BLUT (
.I0(CLBLM_L_X10Y110_SLICE_X13Y110_CO6),
.I1(CLBLM_L_X8Y109_SLICE_X11Y109_CO6),
.I2(LIOB33_X0Y109_IOB_X0Y109_I),
.I3(CLBLM_L_X10Y113_SLICE_X12Y113_AO6),
.I4(LIOB33_X0Y115_IOB_X0Y116_I),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLM_L_X8Y112_SLICE_X10Y112_BO5),
.O6(CLBLM_L_X8Y112_SLICE_X10Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ffffff5555ffff)
  ) CLBLM_L_X8Y112_SLICE_X10Y112_ALUT (
.I0(LIOB33_X0Y115_IOB_X0Y116_I),
.I1(1'b1),
.I2(1'b1),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(LIOB33_X0Y109_IOB_X0Y110_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y112_SLICE_X10Y112_AO5),
.O6(CLBLM_L_X8Y112_SLICE_X10Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y112_SLICE_X11Y112_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y112_SLICE_X11Y112_DO5),
.O6(CLBLM_L_X8Y112_SLICE_X11Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y112_SLICE_X11Y112_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y112_SLICE_X11Y112_CO5),
.O6(CLBLM_L_X8Y112_SLICE_X11Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y112_SLICE_X11Y112_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y112_SLICE_X11Y112_BO5),
.O6(CLBLM_L_X8Y112_SLICE_X11Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y112_SLICE_X11Y112_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y112_SLICE_X11Y112_AO5),
.O6(CLBLM_L_X8Y112_SLICE_X11Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h1f7f5fff035f137f)
  ) CLBLM_L_X8Y113_SLICE_X10Y113_DLUT (
.I0(LIOB33_X0Y109_IOB_X0Y110_I),
.I1(CLBLM_L_X10Y113_SLICE_X12Y113_AO6),
.I2(LIOB33_X0Y115_IOB_X0Y116_I),
.I3(CLBLM_L_X10Y110_SLICE_X13Y110_BO6),
.I4(LIOB33_X0Y109_IOB_X0Y109_I),
.I5(CLBLM_L_X8Y109_SLICE_X11Y109_CO6),
.O5(CLBLM_L_X8Y113_SLICE_X10Y113_DO5),
.O6(CLBLM_L_X8Y113_SLICE_X10Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6696969999696966)
  ) CLBLM_L_X8Y113_SLICE_X10Y113_CLUT (
.I0(CLBLM_L_X8Y114_SLICE_X11Y114_AO6),
.I1(CLBLM_L_X8Y113_SLICE_X10Y113_AO6),
.I2(CLBLM_L_X8Y114_SLICE_X11Y114_BO6),
.I3(CLBLM_L_X8Y113_SLICE_X10Y113_AO5),
.I4(CLBLM_L_X8Y113_SLICE_X10Y113_DO6),
.I5(CLBLM_L_X10Y114_SLICE_X12Y114_AO6),
.O5(CLBLM_L_X8Y113_SLICE_X10Y113_CO5),
.O6(CLBLM_L_X8Y113_SLICE_X10Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hd7b15f93284ea06c)
  ) CLBLM_L_X8Y113_SLICE_X10Y113_BLUT (
.I0(LIOB33_X0Y115_IOB_X0Y116_I),
.I1(CLBLM_L_X10Y113_SLICE_X12Y113_AO6),
.I2(LIOB33_X0Y109_IOB_X0Y110_I),
.I3(CLBLM_L_X8Y109_SLICE_X11Y109_CO6),
.I4(LIOB33_X0Y109_IOB_X0Y109_I),
.I5(CLBLM_L_X10Y110_SLICE_X13Y110_BO6),
.O5(CLBLM_L_X8Y113_SLICE_X10Y113_BO5),
.O6(CLBLM_L_X8Y113_SLICE_X10Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f3f3f3f0fff0fff)
  ) CLBLM_L_X8Y113_SLICE_X10Y113_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(LIOB33_X0Y111_IOB_X0Y111_I),
.I3(LIOB33_X0Y115_IOB_X0Y116_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y113_SLICE_X10Y113_AO5),
.O6(CLBLM_L_X8Y113_SLICE_X10Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y113_SLICE_X11Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y113_SLICE_X11Y113_DO5),
.O6(CLBLM_L_X8Y113_SLICE_X11Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y113_SLICE_X11Y113_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y113_SLICE_X11Y113_CO5),
.O6(CLBLM_L_X8Y113_SLICE_X11Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fdfdfdf134c4c4c)
  ) CLBLM_L_X8Y113_SLICE_X11Y113_BLUT (
.I0(RIOB33_X105Y101_IOB_X1Y102_I),
.I1(CLBLM_L_X10Y112_SLICE_X12Y112_CO6),
.I2(LIOB33_X0Y111_IOB_X0Y111_I),
.I3(RIOB33_X105Y103_IOB_X1Y103_I),
.I4(LIOB33_X0Y109_IOB_X0Y110_I),
.I5(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.O5(CLBLM_L_X8Y113_SLICE_X11Y113_BO5),
.O6(CLBLM_L_X8Y113_SLICE_X11Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6999c33396663ccc)
  ) CLBLM_L_X8Y113_SLICE_X11Y113_ALUT (
.I0(RIOB33_X105Y101_IOB_X1Y102_I),
.I1(CLBLM_L_X10Y112_SLICE_X12Y112_CO6),
.I2(LIOB33_X0Y109_IOB_X0Y110_I),
.I3(RIOB33_X105Y103_IOB_X1Y103_I),
.I4(LIOB33_X0Y111_IOB_X0Y111_I),
.I5(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.O5(CLBLM_L_X8Y113_SLICE_X11Y113_AO5),
.O6(CLBLM_L_X8Y113_SLICE_X11Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y114_SLICE_X10Y114_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y114_SLICE_X10Y114_DO5),
.O6(CLBLM_L_X8Y114_SLICE_X10Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y114_SLICE_X10Y114_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y114_SLICE_X10Y114_CO5),
.O6(CLBLM_L_X8Y114_SLICE_X10Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y114_SLICE_X10Y114_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y114_SLICE_X10Y114_BO5),
.O6(CLBLM_L_X8Y114_SLICE_X10Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6c939393936c6c6c)
  ) CLBLM_L_X8Y114_SLICE_X10Y114_ALUT (
.I0(LIOB33_X0Y111_IOB_X0Y112_I),
.I1(CLBLM_L_X8Y113_SLICE_X11Y113_BO6),
.I2(RIOB33_X105Y101_IOB_X1Y102_I),
.I3(LIOB33_X0Y111_IOB_X0Y111_I),
.I4(RIOB33_X105Y103_IOB_X1Y103_I),
.I5(CLBLM_L_X10Y112_SLICE_X12Y112_AO6),
.O5(CLBLM_L_X8Y114_SLICE_X10Y114_AO5),
.O6(CLBLM_L_X8Y114_SLICE_X10Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7bf31230ffff5af0)
  ) CLBLM_L_X8Y114_SLICE_X11Y114_DLUT (
.I0(LIOB33_X0Y109_IOB_X0Y110_I),
.I1(RIOB33_X105Y101_IOB_X1Y101_I),
.I2(CLBLM_R_X11Y114_SLICE_X14Y114_DO6),
.I3(RIOB33_X105Y101_IOB_X1Y102_I),
.I4(CLBLM_L_X10Y114_SLICE_X12Y114_CO6),
.I5(LIOB33_X0Y111_IOB_X0Y111_I),
.O5(CLBLM_L_X8Y114_SLICE_X11Y114_DO5),
.O6(CLBLM_L_X8Y114_SLICE_X11Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996c33ca55a0ff0)
  ) CLBLM_L_X8Y114_SLICE_X11Y114_CLUT (
.I0(LIOB33_X0Y109_IOB_X0Y110_I),
.I1(RIOB33_X105Y101_IOB_X1Y101_I),
.I2(CLBLM_R_X11Y114_SLICE_X14Y114_DO6),
.I3(CLBLM_L_X10Y114_SLICE_X12Y114_CO6),
.I4(RIOB33_X105Y101_IOB_X1Y102_I),
.I5(LIOB33_X0Y111_IOB_X0Y111_I),
.O5(CLBLM_L_X8Y114_SLICE_X11Y114_CO5),
.O6(CLBLM_L_X8Y114_SLICE_X11Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha6956a956aa66a6a)
  ) CLBLM_L_X8Y114_SLICE_X11Y114_BLUT (
.I0(CLBLM_R_X11Y112_SLICE_X14Y112_AO6),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(LIOB33_X0Y109_IOB_X0Y110_I),
.I3(CLBLM_L_X10Y113_SLICE_X12Y113_DO6),
.I4(LIOB33_X0Y109_IOB_X0Y109_I),
.I5(CLBLM_L_X10Y113_SLICE_X12Y113_CO6),
.O5(CLBLM_L_X8Y114_SLICE_X11Y114_BO5),
.O6(CLBLM_L_X8Y114_SLICE_X11Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h37157f157f377f7f)
  ) CLBLM_L_X8Y114_SLICE_X11Y114_ALUT (
.I0(CLBLM_R_X11Y112_SLICE_X14Y112_AO6),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(LIOB33_X0Y109_IOB_X0Y110_I),
.I3(CLBLM_L_X10Y113_SLICE_X12Y113_DO6),
.I4(LIOB33_X0Y109_IOB_X0Y109_I),
.I5(CLBLM_L_X10Y113_SLICE_X12Y113_CO6),
.O5(CLBLM_L_X8Y114_SLICE_X11Y114_AO5),
.O6(CLBLM_L_X8Y114_SLICE_X11Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h695aa56996a55a96)
  ) CLBLM_L_X8Y115_SLICE_X10Y115_DLUT (
.I0(CLBLM_L_X8Y115_SLICE_X10Y115_AO6),
.I1(CLBLM_L_X8Y114_SLICE_X11Y114_AO6),
.I2(CLBLM_L_X10Y112_SLICE_X13Y112_CO6),
.I3(CLBLM_L_X10Y114_SLICE_X12Y114_AO6),
.I4(CLBLM_L_X8Y113_SLICE_X10Y113_AO6),
.I5(CLBLM_L_X8Y116_SLICE_X10Y116_AO6),
.O5(CLBLM_L_X8Y115_SLICE_X10Y115_DO5),
.O6(CLBLM_L_X8Y115_SLICE_X10Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h2888beeebeeebeee)
  ) CLBLM_L_X8Y115_SLICE_X10Y115_CLUT (
.I0(CLBLM_L_X8Y114_SLICE_X11Y114_AO6),
.I1(CLBLM_L_X10Y114_SLICE_X12Y114_DO6),
.I2(RIOB33_X105Y101_IOB_X1Y101_I),
.I3(LIOB33_X0Y109_IOB_X0Y110_I),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(LIOB33_X0Y111_IOB_X0Y111_I),
.O5(CLBLM_L_X8Y115_SLICE_X10Y115_CO5),
.O6(CLBLM_L_X8Y115_SLICE_X10Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h59a69a65a659659a)
  ) CLBLM_L_X8Y115_SLICE_X10Y115_BLUT (
.I0(CLBLM_R_X11Y114_SLICE_X14Y114_BO6),
.I1(CLBLM_L_X10Y114_SLICE_X12Y114_AO6),
.I2(CLBLM_L_X8Y114_SLICE_X11Y114_AO6),
.I3(CLBLM_L_X8Y116_SLICE_X10Y116_AO6),
.I4(CLBLM_L_X8Y113_SLICE_X10Y113_AO6),
.I5(CLBLM_L_X10Y114_SLICE_X12Y114_CO6),
.O5(CLBLM_L_X8Y115_SLICE_X10Y115_BO5),
.O6(CLBLM_L_X8Y115_SLICE_X10Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h55ff55ff77ff1133)
  ) CLBLM_L_X8Y115_SLICE_X10Y115_ALUT (
.I0(LIOB33_X0Y111_IOB_X0Y112_I),
.I1(CLBLM_L_X8Y114_SLICE_X11Y114_CO6),
.I2(1'b1),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(CLBLM_L_X8Y115_SLICE_X10Y115_CO6),
.I5(1'b1),
.O5(CLBLM_L_X8Y115_SLICE_X10Y115_AO5),
.O6(CLBLM_L_X8Y115_SLICE_X10Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y115_SLICE_X11Y115_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y115_SLICE_X11Y115_DO5),
.O6(CLBLM_L_X8Y115_SLICE_X11Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y115_SLICE_X11Y115_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y115_SLICE_X11Y115_CO5),
.O6(CLBLM_L_X8Y115_SLICE_X11Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y115_SLICE_X11Y115_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y115_SLICE_X11Y115_BO5),
.O6(CLBLM_L_X8Y115_SLICE_X11Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y115_SLICE_X11Y115_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y115_SLICE_X11Y115_AO5),
.O6(CLBLM_L_X8Y115_SLICE_X11Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y116_SLICE_X10Y116_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y116_SLICE_X10Y116_DO5),
.O6(CLBLM_L_X8Y116_SLICE_X10Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h2bd4d42bd42b2bd4)
  ) CLBLM_L_X8Y116_SLICE_X10Y116_CLUT (
.I0(CLBLM_R_X11Y114_SLICE_X14Y114_BO6),
.I1(CLBLM_L_X8Y116_SLICE_X10Y116_AO6),
.I2(CLBLM_L_X10Y114_SLICE_X12Y114_CO6),
.I3(CLBLM_L_X8Y116_SLICE_X10Y116_AO5),
.I4(CLBLM_L_X10Y112_SLICE_X13Y112_BO6),
.I5(CLBLM_R_X7Y114_SLICE_X9Y114_AO6),
.O5(CLBLM_L_X8Y116_SLICE_X10Y116_CO5),
.O6(CLBLM_L_X8Y116_SLICE_X10Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha9696a6665a5a6aa)
  ) CLBLM_L_X8Y116_SLICE_X10Y116_BLUT (
.I0(CLBLM_L_X10Y112_SLICE_X13Y112_BO6),
.I1(LIOB33_X0Y111_IOB_X0Y111_I),
.I2(CLBLM_L_X10Y114_SLICE_X12Y114_CO6),
.I3(RIOB33_X105Y101_IOB_X1Y101_I),
.I4(CLBLM_R_X11Y114_SLICE_X14Y114_BO6),
.I5(RIOB33_X105Y101_IOB_X1Y102_I),
.O5(CLBLM_L_X8Y116_SLICE_X10Y116_BO5),
.O6(CLBLM_L_X8Y116_SLICE_X10Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h33ff33ff77777777)
  ) CLBLM_L_X8Y116_SLICE_X10Y116_ALUT (
.I0(RIOB33_X105Y101_IOB_X1Y102_I),
.I1(LIOB33_X0Y111_IOB_X0Y111_I),
.I2(1'b1),
.I3(RIOB33_X105Y101_IOB_X1Y101_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y116_SLICE_X10Y116_AO5),
.O6(CLBLM_L_X8Y116_SLICE_X10Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y116_SLICE_X11Y116_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y116_SLICE_X11Y116_DO5),
.O6(CLBLM_L_X8Y116_SLICE_X11Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y116_SLICE_X11Y116_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y116_SLICE_X11Y116_CO5),
.O6(CLBLM_L_X8Y116_SLICE_X11Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y116_SLICE_X11Y116_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y116_SLICE_X11Y116_BO5),
.O6(CLBLM_L_X8Y116_SLICE_X11Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y116_SLICE_X11Y116_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y116_SLICE_X11Y116_AO5),
.O6(CLBLM_L_X8Y116_SLICE_X11Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y105_SLICE_X12Y105_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y105_SLICE_X12Y105_DO5),
.O6(CLBLM_L_X10Y105_SLICE_X12Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hbc70cc00d61a0cc0)
  ) CLBLM_L_X10Y105_SLICE_X12Y105_CLUT (
.I0(LIOB33_X0Y101_IOB_X0Y101_I),
.I1(RIOB33_X105Y109_IOB_X1Y110_I),
.I2(LIOB33_X0Y101_IOB_X0Y102_I),
.I3(LIOB33_X0Y103_IOB_X0Y104_I),
.I4(RIOB33_X105Y111_IOB_X1Y111_I),
.I5(CLBLM_L_X10Y105_SLICE_X12Y105_BO6),
.O5(CLBLM_L_X10Y105_SLICE_X12Y105_CO5),
.O6(CLBLM_L_X10Y105_SLICE_X12Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5f577f7f7f7fffff)
  ) CLBLM_L_X10Y105_SLICE_X12Y105_BLUT (
.I0(RIOB33_X105Y109_IOB_X1Y110_I),
.I1(LIOB33_X0Y101_IOB_X0Y101_I),
.I2(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I3(RIOB33_X105Y111_IOB_X1Y112_I),
.I4(RIOB33_X105Y111_IOB_X1Y111_I),
.I5(RIOB33_X105Y113_IOB_X1Y113_I),
.O5(CLBLM_L_X10Y105_SLICE_X12Y105_BO5),
.O6(CLBLM_L_X10Y105_SLICE_X12Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h1f007f5f5f1fff7f)
  ) CLBLM_L_X10Y105_SLICE_X12Y105_ALUT (
.I0(LIOB33_X0Y105_IOB_X0Y105_I),
.I1(LIOB33_X0Y103_IOB_X0Y104_I),
.I2(RIOB33_X105Y109_IOB_X1Y109_I),
.I3(CLBLM_R_X11Y105_SLICE_X14Y105_AO6),
.I4(CLBLM_L_X10Y105_SLICE_X12Y105_CO6),
.I5(CLBLM_L_X10Y106_SLICE_X12Y106_AO5),
.O5(CLBLM_L_X10Y105_SLICE_X12Y105_AO5),
.O6(CLBLM_L_X10Y105_SLICE_X12Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'he55fa0a01aa0a0a0)
  ) CLBLM_L_X10Y105_SLICE_X13Y105_DLUT (
.I0(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I1(RIOB33_X105Y111_IOB_X1Y112_I),
.I2(RIOB33_X105Y111_IOB_X1Y111_I),
.I3(RIOB33_X105Y113_IOB_X1Y113_I),
.I4(RIOB33_X105Y109_IOB_X1Y110_I),
.I5(LIOB33_X0Y101_IOB_X0Y101_I),
.O5(CLBLM_L_X10Y105_SLICE_X13Y105_DO5),
.O6(CLBLM_L_X10Y105_SLICE_X13Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6696969999696966)
  ) CLBLM_L_X10Y105_SLICE_X13Y105_CLUT (
.I0(CLBLM_L_X10Y105_SLICE_X13Y105_AO6),
.I1(CLBLM_L_X10Y106_SLICE_X12Y106_AO5),
.I2(CLBLM_R_X11Y105_SLICE_X14Y105_BO6),
.I3(CLBLM_L_X10Y105_SLICE_X13Y105_AO5),
.I4(CLBLM_R_X11Y105_SLICE_X14Y105_CO6),
.I5(CLBLM_R_X11Y105_SLICE_X14Y105_AO6),
.O5(CLBLM_L_X10Y105_SLICE_X13Y105_CO5),
.O6(CLBLM_L_X10Y105_SLICE_X13Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha569c3c3695af0f0)
  ) CLBLM_L_X10Y105_SLICE_X13Y105_BLUT (
.I0(LIOB33_X0Y105_IOB_X0Y105_I),
.I1(CLBLM_R_X11Y105_SLICE_X14Y105_AO6),
.I2(CLBLM_L_X10Y105_SLICE_X12Y105_CO6),
.I3(LIOB33_X0Y103_IOB_X0Y104_I),
.I4(RIOB33_X105Y109_IOB_X1Y109_I),
.I5(CLBLM_L_X10Y106_SLICE_X12Y106_AO5),
.O5(CLBLM_L_X10Y105_SLICE_X13Y105_BO5),
.O6(CLBLM_L_X10Y105_SLICE_X13Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h55ff55ff77777777)
  ) CLBLM_L_X10Y105_SLICE_X13Y105_ALUT (
.I0(LIOB33_X0Y103_IOB_X0Y104_I),
.I1(RIOB33_X105Y107_IOB_X1Y108_I),
.I2(1'b1),
.I3(RIOB33_X105Y109_IOB_X1Y109_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y105_SLICE_X13Y105_AO5),
.O6(CLBLM_L_X10Y105_SLICE_X13Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y106_SLICE_X12Y106_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y106_SLICE_X12Y106_DO5),
.O6(CLBLM_L_X10Y106_SLICE_X12Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y106_SLICE_X12Y106_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y106_SLICE_X12Y106_CO5),
.O6(CLBLM_L_X10Y106_SLICE_X12Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf43f3fff00ffffff)
  ) CLBLM_L_X10Y106_SLICE_X12Y106_BLUT (
.I0(RIOB33_X105Y111_IOB_X1Y112_I),
.I1(RIOB33_X105Y113_IOB_X1Y113_I),
.I2(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I3(LIOB33_X0Y101_IOB_X0Y101_I),
.I4(RIOB33_X105Y111_IOB_X1Y111_I),
.I5(RIOB33_X105Y109_IOB_X1Y110_I),
.O5(CLBLM_L_X10Y106_SLICE_X12Y106_BO5),
.O6(CLBLM_L_X10Y106_SLICE_X12Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c03f3fa05fa05f)
  ) CLBLM_L_X10Y106_SLICE_X12Y106_ALUT (
.I0(LIOB33_X0Y101_IOB_X0Y102_I),
.I1(LIOB33_X0Y105_IOB_X0Y105_I),
.I2(RIOB33_X105Y109_IOB_X1Y110_I),
.I3(CLBLM_L_X10Y106_SLICE_X12Y106_BO6),
.I4(CLBLM_L_X8Y105_SLICE_X11Y105_AO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y106_SLICE_X12Y106_AO5),
.O6(CLBLM_L_X10Y106_SLICE_X12Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hc6aa395563ff9c00)
  ) CLBLM_L_X10Y106_SLICE_X13Y106_DLUT (
.I0(CLBLM_R_X11Y105_SLICE_X15Y105_BO6),
.I1(LIOB33_X0Y105_IOB_X0Y106_I),
.I2(LIOB33_X0Y105_IOB_X0Y105_I),
.I3(RIOB33_X105Y107_IOB_X1Y108_I),
.I4(CLBLM_L_X10Y105_SLICE_X13Y105_BO6),
.I5(CLBLM_L_X10Y106_SLICE_X13Y106_BO6),
.O5(CLBLM_L_X10Y106_SLICE_X13Y106_DO5),
.O6(CLBLM_L_X10Y106_SLICE_X13Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h02aa3bff23ffbfff)
  ) CLBLM_L_X10Y106_SLICE_X13Y106_CLUT (
.I0(CLBLM_R_X11Y105_SLICE_X15Y105_BO6),
.I1(LIOB33_X0Y105_IOB_X0Y106_I),
.I2(LIOB33_X0Y105_IOB_X0Y105_I),
.I3(RIOB33_X105Y107_IOB_X1Y108_I),
.I4(CLBLM_L_X10Y105_SLICE_X13Y105_BO6),
.I5(CLBLM_L_X10Y106_SLICE_X13Y106_BO6),
.O5(CLBLM_L_X10Y106_SLICE_X13Y106_CO5),
.O6(CLBLM_L_X10Y106_SLICE_X13Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996c33c96963c3c)
  ) CLBLM_L_X10Y106_SLICE_X13Y106_BLUT (
.I0(LIOB33_X0Y101_IOB_X0Y102_I),
.I1(CLBLM_L_X10Y106_SLICE_X12Y106_BO6),
.I2(CLBLM_R_X11Y105_SLICE_X14Y105_AO6),
.I3(RIOB33_X105Y109_IOB_X1Y109_I),
.I4(RIOB33_X105Y109_IOB_X1Y110_I),
.I5(LIOB33_X0Y103_IOB_X0Y104_I),
.O5(CLBLM_L_X10Y106_SLICE_X13Y106_BO5),
.O6(CLBLM_L_X10Y106_SLICE_X13Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h7788887777777777)
  ) CLBLM_L_X10Y106_SLICE_X13Y106_ALUT (
.I0(LIOB33_X0Y105_IOB_X0Y105_I),
.I1(RIOB33_X105Y107_IOB_X1Y108_I),
.I2(1'b1),
.I3(CLBLM_L_X10Y106_SLICE_X13Y106_BO6),
.I4(CLBLM_R_X11Y105_SLICE_X15Y105_BO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y106_SLICE_X13Y106_AO5),
.O6(CLBLM_L_X10Y106_SLICE_X13Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h4488458a8a8a8a8a)
  ) CLBLM_L_X10Y107_SLICE_X12Y107_DLUT (
.I0(CLBLM_L_X10Y108_SLICE_X12Y108_DO6),
.I1(CLBLM_L_X10Y107_SLICE_X13Y107_CO6),
.I2(CLBLM_L_X10Y107_SLICE_X13Y107_BO6),
.I3(RIOB33_X105Y103_IOB_X1Y104_I),
.I4(RIOB33_X105Y103_IOB_X1Y103_I),
.I5(LIOB33_X0Y101_IOB_X0Y101_I),
.O5(CLBLM_L_X10Y107_SLICE_X12Y107_DO5),
.O6(CLBLM_L_X10Y107_SLICE_X12Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hbd2d4ddd42d2b222)
  ) CLBLM_L_X10Y107_SLICE_X12Y107_CLUT (
.I0(CLBLM_L_X10Y108_SLICE_X12Y108_AO6),
.I1(CLBLM_L_X8Y107_SLICE_X11Y107_AO5),
.I2(LIOB33_X0Y101_IOB_X0Y102_I),
.I3(RIOB33_X105Y101_IOB_X1Y102_I),
.I4(RIOB33_X105Y103_IOB_X1Y103_I),
.I5(CLBLM_L_X10Y107_SLICE_X12Y107_BO6),
.O5(CLBLM_L_X10Y107_SLICE_X12Y107_CO5),
.O6(CLBLM_L_X10Y107_SLICE_X12Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0ef3f10cf1f30e0c)
  ) CLBLM_L_X10Y107_SLICE_X12Y107_BLUT (
.I0(RIOB33_X105Y103_IOB_X1Y103_I),
.I1(CLBLM_L_X10Y107_SLICE_X13Y107_BO6),
.I2(CLBLM_L_X10Y107_SLICE_X13Y107_CO6),
.I3(LIOB33_X0Y101_IOB_X0Y101_I),
.I4(CLBLM_L_X10Y108_SLICE_X12Y108_DO6),
.I5(RIOB33_X105Y103_IOB_X1Y104_I),
.O5(CLBLM_L_X10Y107_SLICE_X12Y107_BO5),
.O6(CLBLM_L_X10Y107_SLICE_X12Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h7887877887788778)
  ) CLBLM_L_X10Y107_SLICE_X12Y107_ALUT (
.I0(LIOB33_X0Y101_IOB_X0Y102_I),
.I1(RIOB33_X105Y103_IOB_X1Y103_I),
.I2(CLBLM_L_X8Y105_SLICE_X10Y105_CO6),
.I3(CLBLM_L_X10Y107_SLICE_X12Y107_BO6),
.I4(LIOB33_X0Y103_IOB_X0Y104_I),
.I5(RIOB33_X105Y101_IOB_X1Y102_I),
.O5(CLBLM_L_X10Y107_SLICE_X12Y107_AO5),
.O6(CLBLM_L_X10Y107_SLICE_X12Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y107_SLICE_X13Y107_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y107_SLICE_X13Y107_DO5),
.O6(CLBLM_L_X10Y107_SLICE_X13Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h46550f000a0a0000)
  ) CLBLM_L_X10Y107_SLICE_X13Y107_CLUT (
.I0(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I1(RIOB33_X105Y111_IOB_X1Y112_I),
.I2(RIOB33_X105Y103_IOB_X1Y103_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(RIOB33_X105Y103_IOB_X1Y104_I),
.I5(RIOB33_X105Y113_IOB_X1Y113_I),
.O5(CLBLM_L_X10Y107_SLICE_X13Y107_CO5),
.O6(CLBLM_L_X10Y107_SLICE_X13Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h1d302ec05530a6c0)
  ) CLBLM_L_X10Y107_SLICE_X13Y107_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(RIOB33_X105Y103_IOB_X1Y104_I),
.I2(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I3(RIOB33_X105Y113_IOB_X1Y113_I),
.I4(RIOB33_X105Y103_IOB_X1Y103_I),
.I5(RIOB33_X105Y111_IOB_X1Y112_I),
.O5(CLBLM_L_X10Y107_SLICE_X13Y107_BO5),
.O6(CLBLM_L_X10Y107_SLICE_X13Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h60c0f6fcf6fcf6fc)
  ) CLBLM_L_X10Y107_SLICE_X13Y107_ALUT (
.I0(LIOB33_X0Y101_IOB_X0Y102_I),
.I1(CLBLM_L_X10Y107_SLICE_X12Y107_BO6),
.I2(CLBLM_L_X8Y105_SLICE_X10Y105_CO6),
.I3(RIOB33_X105Y103_IOB_X1Y103_I),
.I4(LIOB33_X0Y103_IOB_X0Y104_I),
.I5(RIOB33_X105Y101_IOB_X1Y102_I),
.O5(CLBLM_L_X10Y107_SLICE_X13Y107_AO5),
.O6(CLBLM_L_X10Y107_SLICE_X13Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h15255aaac0f050a0)
  ) CLBLM_L_X10Y108_SLICE_X12Y108_DLUT (
.I0(RIOB33_X105Y103_IOB_X1Y104_I),
.I1(RIOB33_X105Y111_IOB_X1Y112_I),
.I2(RIOB33_X105Y113_IOB_X1Y113_I),
.I3(RIOB33_X105Y107_IOB_X1Y107_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.O5(CLBLM_L_X10Y108_SLICE_X12Y108_DO5),
.O6(CLBLM_L_X10Y108_SLICE_X12Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffc3d741d741c300)
  ) CLBLM_L_X10Y108_SLICE_X12Y108_CLUT (
.I0(CLBLM_L_X10Y107_SLICE_X12Y107_AO6),
.I1(CLBLM_L_X10Y108_SLICE_X13Y108_CO6),
.I2(CLBLM_L_X12Y108_SLICE_X16Y108_AO5),
.I3(CLBLM_L_X8Y108_SLICE_X11Y108_AO5),
.I4(CLBLM_L_X8Y107_SLICE_X10Y107_AO5),
.I5(CLBLM_L_X8Y108_SLICE_X11Y108_CO6),
.O5(CLBLM_L_X10Y108_SLICE_X12Y108_CO5),
.O6(CLBLM_L_X10Y108_SLICE_X12Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h69a55a69965aa596)
  ) CLBLM_L_X10Y108_SLICE_X12Y108_BLUT (
.I0(CLBLM_L_X12Y108_SLICE_X16Y108_AO5),
.I1(CLBLM_L_X8Y107_SLICE_X10Y107_AO5),
.I2(CLBLM_L_X10Y108_SLICE_X13Y108_CO6),
.I3(CLBLM_L_X8Y108_SLICE_X11Y108_CO6),
.I4(CLBLM_L_X10Y107_SLICE_X12Y107_AO6),
.I5(CLBLM_L_X8Y108_SLICE_X11Y108_AO5),
.O5(CLBLM_L_X10Y108_SLICE_X12Y108_BO5),
.O6(CLBLM_L_X10Y108_SLICE_X12Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf00f00ffcccfccff)
  ) CLBLM_L_X10Y108_SLICE_X12Y108_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y107_SLICE_X13Y107_CO6),
.I2(LIOB33_X0Y101_IOB_X0Y101_I),
.I3(CLBLM_L_X10Y107_SLICE_X13Y107_BO6),
.I4(RIOB33_X105Y103_IOB_X1Y103_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y108_SLICE_X12Y108_AO5),
.O6(CLBLM_L_X10Y108_SLICE_X12Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff0ff0ff2202f02)
  ) CLBLM_L_X10Y108_SLICE_X13Y108_DLUT (
.I0(CLBLM_L_X10Y108_SLICE_X13Y108_AO6),
.I1(CLBLM_L_X10Y107_SLICE_X13Y107_BO6),
.I2(CLBLM_L_X10Y108_SLICE_X12Y108_DO6),
.I3(CLBLM_L_X10Y108_SLICE_X13Y108_AO5),
.I4(CLBLM_R_X11Y107_SLICE_X14Y107_AO6),
.I5(CLBLM_L_X10Y107_SLICE_X13Y107_CO6),
.O5(CLBLM_L_X10Y108_SLICE_X13Y108_DO5),
.O6(CLBLM_L_X10Y108_SLICE_X13Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6c93936c36c9c936)
  ) CLBLM_L_X10Y108_SLICE_X13Y108_CLUT (
.I0(CLBLM_L_X12Y108_SLICE_X16Y108_AO6),
.I1(CLBLM_R_X11Y108_SLICE_X15Y108_AO6),
.I2(CLBLM_L_X8Y105_SLICE_X10Y105_CO6),
.I3(CLBLM_R_X11Y107_SLICE_X14Y107_BO6),
.I4(CLBLM_L_X10Y108_SLICE_X13Y108_DO6),
.I5(CLBLM_L_X10Y108_SLICE_X13Y108_BO6),
.O5(CLBLM_L_X10Y108_SLICE_X13Y108_CO5),
.O6(CLBLM_L_X10Y108_SLICE_X13Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5a965aa5a569a55a)
  ) CLBLM_L_X10Y108_SLICE_X13Y108_BLUT (
.I0(CLBLM_L_X10Y108_SLICE_X12Y108_DO6),
.I1(CLBLM_L_X10Y107_SLICE_X13Y107_BO6),
.I2(CLBLM_R_X11Y107_SLICE_X14Y107_AO6),
.I3(CLBLM_L_X10Y107_SLICE_X13Y107_CO6),
.I4(CLBLM_L_X10Y108_SLICE_X13Y108_AO6),
.I5(CLBLM_L_X10Y108_SLICE_X13Y108_AO5),
.O5(CLBLM_L_X10Y108_SLICE_X13Y108_BO5),
.O6(CLBLM_L_X10Y108_SLICE_X13Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0fffff3f3f3f3f)
  ) CLBLM_L_X10Y108_SLICE_X13Y108_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y101_IOB_X0Y102_I),
.I2(RIOB33_X105Y103_IOB_X1Y103_I),
.I3(1'b1),
.I4(LIOB33_X0Y101_IOB_X0Y101_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y108_SLICE_X13Y108_AO5),
.O6(CLBLM_L_X10Y108_SLICE_X13Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h9f3f60c0c5953a6a)
  ) CLBLM_L_X10Y109_SLICE_X12Y109_DLUT (
.I0(CLBLM_L_X10Y107_SLICE_X12Y107_AO6),
.I1(RIOB33_X105Y101_IOB_X1Y102_I),
.I2(LIOB33_X0Y105_IOB_X0Y105_I),
.I3(RIOB33_X105Y101_IOB_X1Y101_I),
.I4(CLBLM_L_X10Y108_SLICE_X13Y108_CO6),
.I5(CLBLM_L_X8Y108_SLICE_X11Y108_CO6),
.O5(CLBLM_L_X10Y109_SLICE_X12Y109_DO5),
.O6(CLBLM_L_X10Y109_SLICE_X12Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fdfff5f134c5f00)
  ) CLBLM_L_X10Y109_SLICE_X12Y109_CLUT (
.I0(RIOB33_X105Y101_IOB_X1Y101_I),
.I1(LIOB33_X0Y103_IOB_X0Y104_I),
.I2(LIOB33_X0Y105_IOB_X0Y105_I),
.I3(CLBLM_L_X10Y107_SLICE_X12Y107_CO6),
.I4(RIOB33_X105Y101_IOB_X1Y102_I),
.I5(CLBLM_L_X8Y108_SLICE_X11Y108_CO6),
.O5(CLBLM_L_X10Y109_SLICE_X12Y109_CO5),
.O6(CLBLM_L_X10Y109_SLICE_X12Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h444c5d5f5fdfdfff)
  ) CLBLM_L_X10Y109_SLICE_X12Y109_BLUT (
.I0(RIOB33_X105Y107_IOB_X1Y107_I),
.I1(CLBLM_R_X11Y109_SLICE_X14Y109_AO6),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(LIOB33_X0Y105_IOB_X0Y106_I),
.I4(CLBLM_L_X10Y106_SLICE_X13Y106_AO6),
.I5(CLBLM_L_X10Y106_SLICE_X13Y106_DO6),
.O5(CLBLM_L_X10Y109_SLICE_X12Y109_BO5),
.O6(CLBLM_L_X10Y109_SLICE_X12Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hb78877b748778848)
  ) CLBLM_L_X10Y109_SLICE_X12Y109_ALUT (
.I0(LIOB33_X0Y107_IOB_X0Y107_I),
.I1(RIOB33_X105Y107_IOB_X1Y107_I),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(CLBLM_R_X11Y109_SLICE_X14Y109_AO6),
.I4(CLBLM_L_X10Y106_SLICE_X13Y106_AO6),
.I5(CLBLM_L_X10Y106_SLICE_X13Y106_DO6),
.O5(CLBLM_L_X10Y109_SLICE_X12Y109_AO5),
.O6(CLBLM_L_X10Y109_SLICE_X12Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h373f03377fff0f7f)
  ) CLBLM_L_X10Y109_SLICE_X13Y109_DLUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(RIOB33_X105Y101_IOB_X1Y101_I),
.I2(CLBLM_R_X11Y110_SLICE_X15Y110_AO6),
.I3(CLBLM_L_X10Y109_SLICE_X13Y109_CO6),
.I4(CLBLM_L_X10Y109_SLICE_X12Y109_CO6),
.I5(LIOB33_X0Y107_IOB_X0Y107_I),
.O5(CLBLM_L_X10Y109_SLICE_X13Y109_DO5),
.O6(CLBLM_L_X10Y109_SLICE_X13Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7887877888777788)
  ) CLBLM_L_X10Y109_SLICE_X13Y109_CLUT (
.I0(RIOB33_X105Y103_IOB_X1Y103_I),
.I1(LIOB33_X0Y103_IOB_X0Y104_I),
.I2(LIOB33_X0Y105_IOB_X0Y105_I),
.I3(CLBLM_R_X11Y108_SLICE_X14Y108_DO6),
.I4(CLBLM_L_X10Y107_SLICE_X13Y107_AO6),
.I5(RIOB33_X105Y101_IOB_X1Y102_I),
.O5(CLBLM_L_X10Y109_SLICE_X13Y109_CO5),
.O6(CLBLM_L_X10Y109_SLICE_X13Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'he62a19d573bf8c40)
  ) CLBLM_L_X10Y109_SLICE_X13Y109_BLUT (
.I0(CLBLM_L_X10Y109_SLICE_X12Y109_CO6),
.I1(LIOB33_X0Y105_IOB_X0Y106_I),
.I2(RIOB33_X105Y101_IOB_X1Y101_I),
.I3(RIOB33_X105Y101_IOB_X1Y102_I),
.I4(CLBLM_R_X11Y109_SLICE_X15Y109_BO6),
.I5(CLBLM_L_X10Y109_SLICE_X13Y109_CO6),
.O5(CLBLM_L_X10Y109_SLICE_X13Y109_BO5),
.O6(CLBLM_L_X10Y109_SLICE_X13Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc96939996c3c9ccc)
  ) CLBLM_L_X10Y109_SLICE_X13Y109_ALUT (
.I0(CLBLM_L_X10Y109_SLICE_X12Y109_CO6),
.I1(CLBLM_R_X11Y110_SLICE_X15Y110_AO6),
.I2(RIOB33_X105Y101_IOB_X1Y101_I),
.I3(LIOB33_X0Y105_IOB_X0Y106_I),
.I4(LIOB33_X0Y107_IOB_X0Y107_I),
.I5(CLBLM_L_X10Y109_SLICE_X13Y109_CO6),
.O5(CLBLM_L_X10Y109_SLICE_X13Y109_AO5),
.O6(CLBLM_L_X10Y109_SLICE_X13Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h639c9c63c63939c6)
  ) CLBLM_L_X10Y110_SLICE_X12Y110_DLUT (
.I0(CLBLM_L_X10Y110_SLICE_X12Y110_AO6),
.I1(CLBLM_R_X11Y110_SLICE_X14Y110_AO6),
.I2(CLBLM_L_X10Y108_SLICE_X12Y108_BO6),
.I3(CLBLM_L_X10Y108_SLICE_X12Y108_CO6),
.I4(CLBLM_R_X11Y110_SLICE_X15Y110_AO6),
.I5(CLBLM_L_X8Y108_SLICE_X10Y108_CO6),
.O5(CLBLM_L_X10Y110_SLICE_X12Y110_DO5),
.O6(CLBLM_L_X10Y110_SLICE_X12Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h59a6a6599a65659a)
  ) CLBLM_L_X10Y110_SLICE_X12Y110_CLUT (
.I0(CLBLM_L_X8Y106_SLICE_X11Y106_AO6),
.I1(CLBLM_L_X10Y106_SLICE_X13Y106_DO6),
.I2(CLBLM_L_X10Y110_SLICE_X12Y110_AO5),
.I3(CLBLM_L_X8Y110_SLICE_X10Y110_AO5),
.I4(CLBLM_L_X10Y106_SLICE_X13Y106_CO6),
.I5(CLBLM_R_X11Y109_SLICE_X14Y109_BO6),
.O5(CLBLM_L_X10Y110_SLICE_X12Y110_CO5),
.O6(CLBLM_L_X10Y110_SLICE_X12Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5f5f5f5f77777777)
  ) CLBLM_L_X10Y110_SLICE_X12Y110_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(LIOB33_X0Y109_IOB_X0Y109_I),
.I2(LIOB33_X0Y107_IOB_X0Y108_I),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y110_SLICE_X12Y110_BO5),
.O6(CLBLM_L_X10Y110_SLICE_X12Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h55ff55ff5555ffff)
  ) CLBLM_L_X10Y110_SLICE_X12Y110_ALUT (
.I0(LIOB33_X0Y107_IOB_X0Y107_I),
.I1(1'b1),
.I2(1'b1),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(RIOB33_X105Y107_IOB_X1Y107_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y110_SLICE_X12Y110_AO5),
.O6(CLBLM_L_X10Y110_SLICE_X12Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hea80fea880eaa8fe)
  ) CLBLM_L_X10Y110_SLICE_X13Y110_DLUT (
.I0(CLBLM_L_X8Y109_SLICE_X11Y109_AO5),
.I1(CLBLM_L_X10Y111_SLICE_X13Y111_AO6),
.I2(CLBLM_L_X8Y110_SLICE_X11Y110_CO6),
.I3(CLBLM_L_X10Y111_SLICE_X13Y111_AO5),
.I4(CLBLM_L_X10Y109_SLICE_X13Y109_AO6),
.I5(CLBLM_R_X11Y110_SLICE_X14Y110_CO6),
.O5(CLBLM_L_X10Y110_SLICE_X13Y110_DO5),
.O6(CLBLM_L_X10Y110_SLICE_X13Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h96c3cc663c96cc66)
  ) CLBLM_L_X10Y110_SLICE_X13Y110_CLUT (
.I0(CLBLM_L_X10Y109_SLICE_X13Y109_AO6),
.I1(CLBLM_R_X11Y110_SLICE_X14Y110_CO6),
.I2(RIOB33_X105Y101_IOB_X1Y101_I),
.I3(CLBLM_L_X8Y110_SLICE_X11Y110_CO6),
.I4(LIOB33_X0Y107_IOB_X0Y108_I),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLM_L_X10Y110_SLICE_X13Y110_CO5),
.O6(CLBLM_L_X10Y110_SLICE_X13Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h718e8e718e71718e)
  ) CLBLM_L_X10Y110_SLICE_X13Y110_BLUT (
.I0(CLBLM_L_X8Y110_SLICE_X11Y110_CO6),
.I1(CLBLM_L_X10Y111_SLICE_X13Y111_AO6),
.I2(CLBLM_L_X10Y109_SLICE_X13Y109_AO6),
.I3(CLBLM_R_X11Y110_SLICE_X14Y110_CO6),
.I4(CLBLM_L_X8Y109_SLICE_X11Y109_AO5),
.I5(CLBLM_L_X10Y111_SLICE_X13Y111_AO5),
.O5(CLBLM_L_X10Y110_SLICE_X13Y110_BO5),
.O6(CLBLM_L_X10Y110_SLICE_X13Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h659a9a65a65959a6)
  ) CLBLM_L_X10Y110_SLICE_X13Y110_ALUT (
.I0(CLBLM_L_X10Y110_SLICE_X12Y110_AO5),
.I1(CLBLM_L_X12Y109_SLICE_X16Y109_AO5),
.I2(CLBLM_R_X11Y109_SLICE_X14Y109_DO6),
.I3(CLBLM_R_X11Y109_SLICE_X14Y109_BO6),
.I4(CLBLM_L_X10Y106_SLICE_X13Y106_DO6),
.I5(CLBLM_R_X13Y108_SLICE_X18Y108_CO6),
.O5(CLBLM_L_X10Y110_SLICE_X13Y110_AO5),
.O6(CLBLM_L_X10Y110_SLICE_X13Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h93c9ff556c3600aa)
  ) CLBLM_L_X10Y111_SLICE_X12Y111_DLUT (
.I0(CLBLM_L_X10Y111_SLICE_X12Y111_AO6),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(RIOB33_X105Y103_IOB_X1Y104_I),
.I3(CLBLM_R_X11Y111_SLICE_X15Y111_DO6),
.I4(LIOB33_X0Y109_IOB_X0Y109_I),
.I5(CLBLM_L_X10Y111_SLICE_X12Y111_BO6),
.O5(CLBLM_L_X10Y111_SLICE_X12Y111_DO5),
.O6(CLBLM_L_X10Y111_SLICE_X12Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfddff44fd00d4004)
  ) CLBLM_L_X10Y111_SLICE_X12Y111_CLUT (
.I0(CLBLM_L_X10Y109_SLICE_X12Y109_AO6),
.I1(CLBLM_L_X10Y111_SLICE_X13Y111_CO6),
.I2(CLBLM_L_X10Y110_SLICE_X12Y110_CO6),
.I3(CLBLM_L_X8Y111_SLICE_X10Y111_AO5),
.I4(CLBLM_L_X10Y110_SLICE_X12Y110_BO6),
.I5(CLBLM_L_X10Y110_SLICE_X12Y110_BO5),
.O5(CLBLM_L_X10Y111_SLICE_X12Y111_CO5),
.O6(CLBLM_L_X10Y111_SLICE_X12Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hd78d778728728878)
  ) CLBLM_L_X10Y111_SLICE_X12Y111_BLUT (
.I0(LIOB33_X0Y107_IOB_X0Y108_I),
.I1(RIOB33_X105Y107_IOB_X1Y107_I),
.I2(CLBLM_L_X10Y109_SLICE_X12Y109_AO6),
.I3(CLBLM_L_X10Y111_SLICE_X13Y111_CO6),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_L_X10Y110_SLICE_X12Y110_CO6),
.O5(CLBLM_L_X10Y111_SLICE_X12Y111_BO5),
.O6(CLBLM_L_X10Y111_SLICE_X12Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5aa5f00f5f05ff0f)
  ) CLBLM_L_X10Y111_SLICE_X12Y111_ALUT (
.I0(LIOB33_X0Y107_IOB_X0Y108_I),
.I1(1'b1),
.I2(CLBLM_L_X10Y109_SLICE_X12Y109_AO6),
.I3(CLBLM_L_X10Y111_SLICE_X13Y111_CO6),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y111_SLICE_X12Y111_AO5),
.O6(CLBLM_L_X10Y111_SLICE_X12Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hc69c399c639c9c9c)
  ) CLBLM_L_X10Y111_SLICE_X13Y111_DLUT (
.I0(CLBLM_R_X11Y111_SLICE_X15Y111_AO6),
.I1(CLBLM_L_X10Y110_SLICE_X13Y110_AO6),
.I2(CLBLM_R_X11Y111_SLICE_X14Y111_CO6),
.I3(LIOB33_X0Y107_IOB_X0Y108_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(RIOB33_X105Y103_IOB_X1Y104_I),
.O5(CLBLM_L_X10Y111_SLICE_X13Y111_DO5),
.O6(CLBLM_L_X10Y111_SLICE_X13Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h78ffffff00787878)
  ) CLBLM_L_X10Y111_SLICE_X13Y111_CLUT (
.I0(RIOB33_X105Y107_IOB_X1Y107_I),
.I1(LIOB33_X0Y105_IOB_X0Y106_I),
.I2(CLBLM_R_X11Y109_SLICE_X14Y109_CO6),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(LIOB33_X0Y107_IOB_X0Y107_I),
.I5(CLBLM_R_X13Y108_SLICE_X18Y108_CO6),
.O5(CLBLM_L_X10Y111_SLICE_X13Y111_CO5),
.O6(CLBLM_L_X10Y111_SLICE_X13Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7dff143cddff44cc)
  ) CLBLM_L_X10Y111_SLICE_X13Y111_BLUT (
.I0(RIOB33_X105Y103_IOB_X1Y104_I),
.I1(CLBLM_L_X10Y111_SLICE_X12Y111_BO6),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(LIOB33_X0Y109_IOB_X0Y110_I),
.I4(CLBLM_R_X11Y111_SLICE_X14Y111_BO6),
.I5(LIOB33_X0Y109_IOB_X0Y109_I),
.O5(CLBLM_L_X10Y111_SLICE_X13Y111_BO5),
.O6(CLBLM_L_X10Y111_SLICE_X13Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h777777775f5f5f5f)
  ) CLBLM_L_X10Y111_SLICE_X13Y111_ALUT (
.I0(LIOB33_X0Y107_IOB_X0Y108_I),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(RIOB33_X105Y101_IOB_X1Y101_I),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y111_SLICE_X13Y111_AO5),
.O6(CLBLM_L_X10Y111_SLICE_X13Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0d4d4f5f5ddddfff)
  ) CLBLM_L_X10Y112_SLICE_X12Y112_DLUT (
.I0(CLBLM_R_X11Y111_SLICE_X14Y111_DO6),
.I1(CLBLM_R_X11Y112_SLICE_X14Y112_DO6),
.I2(RIOB33_X105Y103_IOB_X1Y103_I),
.I3(LIOB33_X0Y109_IOB_X0Y109_I),
.I4(CLBLM_R_X11Y112_SLICE_X15Y112_DO6),
.I5(LIOB33_X0Y109_IOB_X0Y110_I),
.O5(CLBLM_L_X10Y112_SLICE_X12Y112_DO5),
.O6(CLBLM_L_X10Y112_SLICE_X12Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h9af059ff650fa600)
  ) CLBLM_L_X10Y112_SLICE_X12Y112_CLUT (
.I0(RIOB33_X105Y103_IOB_X1Y104_I),
.I1(RIOB33_X105Y103_IOB_X1Y103_I),
.I2(CLBLM_R_X11Y112_SLICE_X14Y112_DO6),
.I3(LIOB33_X0Y109_IOB_X0Y109_I),
.I4(CLBLM_R_X11Y112_SLICE_X15Y112_DO6),
.I5(CLBLM_L_X10Y111_SLICE_X13Y111_DO6),
.O5(CLBLM_L_X10Y112_SLICE_X12Y112_CO5),
.O6(CLBLM_L_X10Y112_SLICE_X12Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h4bb4d22db44b2dd2)
  ) CLBLM_L_X10Y112_SLICE_X12Y112_BLUT (
.I0(CLBLM_L_X10Y110_SLICE_X13Y110_DO6),
.I1(CLBLM_R_X11Y112_SLICE_X14Y112_AO6),
.I2(CLBLM_L_X10Y112_SLICE_X13Y112_AO6),
.I3(CLBLM_R_X11Y113_SLICE_X14Y113_AO6),
.I4(CLBLM_L_X8Y112_SLICE_X10Y112_AO6),
.I5(CLBLM_R_X11Y112_SLICE_X14Y112_CO6),
.O5(CLBLM_L_X10Y112_SLICE_X12Y112_BO5),
.O6(CLBLM_L_X10Y112_SLICE_X12Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h66999999aa555555)
  ) CLBLM_L_X10Y112_SLICE_X12Y112_ALUT (
.I0(CLBLM_L_X10Y111_SLICE_X12Y111_DO6),
.I1(CLBLM_L_X10Y112_SLICE_X12Y112_DO6),
.I2(1'b1),
.I3(LIOB33_X0Y109_IOB_X0Y110_I),
.I4(RIOB33_X105Y103_IOB_X1Y104_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y112_SLICE_X12Y112_AO5),
.O6(CLBLM_L_X10Y112_SLICE_X12Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ffffffffffff)
  ) CLBLM_L_X10Y112_SLICE_X13Y112_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(RIOB33_X105Y103_IOB_X1Y103_I),
.I5(LIOB33_X0Y109_IOB_X0Y110_I),
.O5(CLBLM_L_X10Y112_SLICE_X13Y112_DO5),
.O6(CLBLM_L_X10Y112_SLICE_X13Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h69963cc3c33c6996)
  ) CLBLM_L_X10Y112_SLICE_X13Y112_CLUT (
.I0(CLBLM_L_X10Y112_SLICE_X13Y112_AO6),
.I1(CLBLM_R_X11Y112_SLICE_X15Y112_BO6),
.I2(CLBLM_R_X11Y113_SLICE_X14Y113_CO6),
.I3(CLBLM_L_X10Y112_SLICE_X13Y112_AO5),
.I4(CLBLM_R_X11Y113_SLICE_X14Y113_AO6),
.I5(CLBLM_R_X11Y112_SLICE_X14Y112_CO6),
.O5(CLBLM_L_X10Y112_SLICE_X13Y112_CO5),
.O6(CLBLM_L_X10Y112_SLICE_X13Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h69963cc3c33c6996)
  ) CLBLM_L_X10Y112_SLICE_X13Y112_BLUT (
.I0(CLBLM_R_X11Y113_SLICE_X14Y113_CO6),
.I1(CLBLM_R_X11Y111_SLICE_X15Y111_CO6),
.I2(CLBLM_R_X11Y111_SLICE_X14Y111_DO6),
.I3(CLBLM_L_X10Y112_SLICE_X13Y112_DO6),
.I4(CLBLM_R_X11Y112_SLICE_X15Y112_BO6),
.I5(CLBLM_L_X10Y112_SLICE_X13Y112_AO5),
.O5(CLBLM_L_X10Y112_SLICE_X13Y112_BO5),
.O6(CLBLM_L_X10Y112_SLICE_X13Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ffffff55ff55ff)
  ) CLBLM_L_X10Y112_SLICE_X13Y112_ALUT (
.I0(RIOB33_X105Y101_IOB_X1Y102_I),
.I1(1'b1),
.I2(1'b1),
.I3(LIOB33_X0Y109_IOB_X0Y110_I),
.I4(RIOB33_X105Y101_IOB_X1Y101_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y112_SLICE_X13Y112_AO5),
.O6(CLBLM_L_X10Y112_SLICE_X13Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7f07ff778f08ff88)
  ) CLBLM_L_X10Y113_SLICE_X12Y113_DLUT (
.I0(RIOB33_X105Y101_IOB_X1Y101_I),
.I1(LIOB33_X0Y107_IOB_X0Y107_I),
.I2(LIOB33_X0Y107_IOB_X0Y108_I),
.I3(CLBLM_L_X8Y110_SLICE_X11Y110_CO6),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(CLBLM_L_X10Y109_SLICE_X13Y109_BO6),
.O5(CLBLM_L_X10Y113_SLICE_X12Y113_DO5),
.O6(CLBLM_L_X10Y113_SLICE_X12Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996c33c996633cc)
  ) CLBLM_L_X10Y113_SLICE_X12Y113_CLUT (
.I0(RIOB33_X105Y101_IOB_X1Y101_I),
.I1(CLBLM_L_X10Y109_SLICE_X13Y109_DO6),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(CLBLM_L_X12Y111_SLICE_X16Y111_BO6),
.I4(LIOB33_X0Y107_IOB_X0Y108_I),
.I5(RIOB33_X105Y101_IOB_X1Y102_I),
.O5(CLBLM_L_X10Y113_SLICE_X12Y113_CO5),
.O6(CLBLM_L_X10Y113_SLICE_X12Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hd2a52da54bf0b4f0)
  ) CLBLM_L_X10Y113_SLICE_X12Y113_BLUT (
.I0(CLBLM_L_X10Y113_SLICE_X12Y113_DO6),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(CLBLM_R_X11Y112_SLICE_X14Y112_BO6),
.I3(LIOB33_X0Y109_IOB_X0Y109_I),
.I4(RIOB33_X105Y101_IOB_X1Y101_I),
.I5(CLBLM_L_X10Y113_SLICE_X12Y113_CO6),
.O5(CLBLM_L_X10Y113_SLICE_X12Y113_BO5),
.O6(CLBLM_L_X10Y113_SLICE_X12Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6a95c03f956a3fc0)
  ) CLBLM_L_X10Y113_SLICE_X12Y113_ALUT (
.I0(LIOB33_X0Y107_IOB_X0Y107_I),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(LIOB33_X0Y107_IOB_X0Y108_I),
.I3(CLBLM_L_X10Y109_SLICE_X13Y109_BO6),
.I4(RIOB33_X105Y101_IOB_X1Y101_I),
.I5(CLBLM_L_X8Y110_SLICE_X11Y110_CO6),
.O5(CLBLM_L_X10Y113_SLICE_X12Y113_AO5),
.O6(CLBLM_L_X10Y113_SLICE_X12Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y113_SLICE_X13Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y113_SLICE_X13Y113_DO5),
.O6(CLBLM_L_X10Y113_SLICE_X13Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y113_SLICE_X13Y113_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y113_SLICE_X13Y113_CO5),
.O6(CLBLM_L_X10Y113_SLICE_X13Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y113_SLICE_X13Y113_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y113_SLICE_X13Y113_BO5),
.O6(CLBLM_L_X10Y113_SLICE_X13Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333ffff77777777)
  ) CLBLM_L_X10Y113_SLICE_X13Y113_ALUT (
.I0(LIOB33_X0Y107_IOB_X0Y108_I),
.I1(RIOB33_X105Y101_IOB_X1Y102_I),
.I2(1'b1),
.I3(1'b1),
.I4(LIOB33_X0Y109_IOB_X0Y109_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y113_SLICE_X13Y113_AO5),
.O6(CLBLM_L_X10Y113_SLICE_X13Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8778f0f0e11e3c3c)
  ) CLBLM_L_X10Y114_SLICE_X12Y114_DLUT (
.I0(RIOB33_X105Y101_IOB_X1Y101_I),
.I1(CLBLM_R_X11Y114_SLICE_X14Y114_AO6),
.I2(CLBLM_R_X11Y113_SLICE_X14Y113_BO6),
.I3(RIOB33_X105Y101_IOB_X1Y102_I),
.I4(LIOB33_X0Y109_IOB_X0Y109_I),
.I5(CLBLM_L_X10Y114_SLICE_X12Y114_BO6),
.O5(CLBLM_L_X10Y114_SLICE_X12Y114_DO5),
.O6(CLBLM_L_X10Y114_SLICE_X12Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h1f7f5fff07571777)
  ) CLBLM_L_X10Y114_SLICE_X12Y114_CLUT (
.I0(CLBLM_R_X11Y113_SLICE_X14Y113_AO6),
.I1(CLBLM_R_X11Y114_SLICE_X14Y114_AO6),
.I2(RIOB33_X105Y101_IOB_X1Y101_I),
.I3(LIOB33_X0Y109_IOB_X0Y110_I),
.I4(LIOB33_X0Y109_IOB_X0Y109_I),
.I5(CLBLM_L_X10Y114_SLICE_X12Y114_BO6),
.O5(CLBLM_L_X10Y114_SLICE_X12Y114_CO5),
.O6(CLBLM_L_X10Y114_SLICE_X12Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6f06ff66cf0cffcc)
  ) CLBLM_L_X10Y114_SLICE_X12Y114_BLUT (
.I0(LIOB33_X0Y107_IOB_X0Y107_I),
.I1(CLBLM_L_X12Y111_SLICE_X16Y111_BO6),
.I2(LIOB33_X0Y107_IOB_X0Y108_I),
.I3(CLBLM_L_X10Y109_SLICE_X13Y109_DO6),
.I4(RIOB33_X105Y101_IOB_X1Y101_I),
.I5(RIOB33_X105Y101_IOB_X1Y102_I),
.O5(CLBLM_L_X10Y114_SLICE_X12Y114_BO5),
.O6(CLBLM_L_X10Y114_SLICE_X12Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8fe3701c7f1380ec)
  ) CLBLM_L_X10Y114_SLICE_X12Y114_ALUT (
.I0(LIOB33_X0Y109_IOB_X0Y109_I),
.I1(CLBLM_R_X11Y114_SLICE_X14Y114_AO6),
.I2(RIOB33_X105Y101_IOB_X1Y101_I),
.I3(CLBLM_L_X10Y114_SLICE_X12Y114_BO6),
.I4(CLBLM_R_X11Y113_SLICE_X14Y113_AO6),
.I5(LIOB33_X0Y109_IOB_X0Y110_I),
.O5(CLBLM_L_X10Y114_SLICE_X12Y114_AO5),
.O6(CLBLM_L_X10Y114_SLICE_X12Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y114_SLICE_X13Y114_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y114_SLICE_X13Y114_DO5),
.O6(CLBLM_L_X10Y114_SLICE_X13Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y114_SLICE_X13Y114_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y114_SLICE_X13Y114_CO5),
.O6(CLBLM_L_X10Y114_SLICE_X13Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y114_SLICE_X13Y114_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y114_SLICE_X13Y114_BO5),
.O6(CLBLM_L_X10Y114_SLICE_X13Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y114_SLICE_X13Y114_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y114_SLICE_X13Y114_AO5),
.O6(CLBLM_L_X10Y114_SLICE_X13Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h220266c60000a0a0)
  ) CLBLM_L_X12Y105_SLICE_X16Y105_DLUT (
.I0(RIOB33_X105Y113_IOB_X1Y113_I),
.I1(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I2(RIOB33_X105Y109_IOB_X1Y110_I),
.I3(RIOB33_X105Y111_IOB_X1Y112_I),
.I4(RIOB33_X105Y107_IOB_X1Y108_I),
.I5(RIOB33_X105Y109_IOB_X1Y109_I),
.O5(CLBLM_L_X12Y105_SLICE_X16Y105_DO5),
.O6(CLBLM_L_X12Y105_SLICE_X16Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'he7efc545951db7b7)
  ) CLBLM_L_X12Y105_SLICE_X16Y105_CLUT (
.I0(RIOB33_X105Y113_IOB_X1Y113_I),
.I1(RIOB33_X105Y109_IOB_X1Y110_I),
.I2(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I3(RIOB33_X105Y111_IOB_X1Y112_I),
.I4(RIOB33_X105Y111_IOB_X1Y111_I),
.I5(RIOB33_X105Y109_IOB_X1Y109_I),
.O5(CLBLM_L_X12Y105_SLICE_X16Y105_CO5),
.O6(CLBLM_L_X12Y105_SLICE_X16Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h66aa63ff99559c00)
  ) CLBLM_L_X12Y105_SLICE_X16Y105_BLUT (
.I0(CLBLM_L_X12Y105_SLICE_X16Y105_DO6),
.I1(RIOB33_X105Y109_IOB_X1Y109_I),
.I2(RIOB33_X105Y107_IOB_X1Y108_I),
.I3(LIOB33_X0Y101_IOB_X0Y101_I),
.I4(CLBLM_R_X11Y107_SLICE_X14Y107_DO6),
.I5(CLBLM_L_X12Y105_SLICE_X16Y105_CO6),
.O5(CLBLM_L_X12Y105_SLICE_X16Y105_BO5),
.O6(CLBLM_L_X12Y105_SLICE_X16Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc333c333abbbabbb)
  ) CLBLM_L_X12Y105_SLICE_X16Y105_ALUT (
.I0(CLBLM_L_X12Y105_SLICE_X16Y105_DO6),
.I1(CLBLM_R_X11Y107_SLICE_X14Y107_DO6),
.I2(RIOB33_X105Y107_IOB_X1Y108_I),
.I3(LIOB33_X0Y101_IOB_X0Y101_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y105_SLICE_X16Y105_AO5),
.O6(CLBLM_L_X12Y105_SLICE_X16Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y105_SLICE_X17Y105_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y105_SLICE_X17Y105_DO5),
.O6(CLBLM_L_X12Y105_SLICE_X17Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y105_SLICE_X17Y105_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y105_SLICE_X17Y105_CO5),
.O6(CLBLM_L_X12Y105_SLICE_X17Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y105_SLICE_X17Y105_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y105_SLICE_X17Y105_BO5),
.O6(CLBLM_L_X12Y105_SLICE_X17Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y105_SLICE_X17Y105_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y105_SLICE_X17Y105_AO5),
.O6(CLBLM_L_X12Y105_SLICE_X17Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y106_SLICE_X16Y106_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y106_SLICE_X16Y106_DO5),
.O6(CLBLM_L_X12Y106_SLICE_X16Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h96996696aa55aaaa)
  ) CLBLM_L_X12Y106_SLICE_X16Y106_CLUT (
.I0(CLBLM_L_X12Y105_SLICE_X16Y105_BO6),
.I1(RIOB33_X105Y107_IOB_X1Y108_I),
.I2(RIOB33_X105Y107_IOB_X1Y107_I),
.I3(CLBLM_L_X12Y106_SLICE_X16Y106_AO5),
.I4(CLBLM_L_X12Y105_SLICE_X16Y105_AO6),
.I5(LIOB33_X0Y101_IOB_X0Y102_I),
.O5(CLBLM_L_X12Y106_SLICE_X16Y106_CO5),
.O6(CLBLM_L_X12Y106_SLICE_X16Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h004c00f0b0bc0000)
  ) CLBLM_L_X12Y106_SLICE_X16Y106_BLUT (
.I0(RIOB33_X105Y111_IOB_X1Y112_I),
.I1(RIOB33_X105Y109_IOB_X1Y109_I),
.I2(RIOB33_X105Y107_IOB_X1Y108_I),
.I3(RIOB33_X105Y107_IOB_X1Y107_I),
.I4(RIOB33_X105Y113_IOB_X1Y113_I),
.I5(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.O5(CLBLM_L_X12Y106_SLICE_X16Y106_BO5),
.O6(CLBLM_L_X12Y106_SLICE_X16Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c03f3fff00ff3f)
  ) CLBLM_L_X12Y106_SLICE_X16Y106_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y101_IOB_X0Y101_I),
.I2(RIOB33_X105Y107_IOB_X1Y107_I),
.I3(CLBLM_L_X12Y106_SLICE_X16Y106_BO6),
.I4(CLBLM_L_X12Y107_SLICE_X17Y107_AO6),
.I5(1'b1),
.O5(CLBLM_L_X12Y106_SLICE_X16Y106_AO5),
.O6(CLBLM_L_X12Y106_SLICE_X16Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y106_SLICE_X17Y106_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y106_SLICE_X17Y106_DO5),
.O6(CLBLM_L_X12Y106_SLICE_X17Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y106_SLICE_X17Y106_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y106_SLICE_X17Y106_CO5),
.O6(CLBLM_L_X12Y106_SLICE_X17Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y106_SLICE_X17Y106_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y106_SLICE_X17Y106_BO5),
.O6(CLBLM_L_X12Y106_SLICE_X17Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y106_SLICE_X17Y106_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y106_SLICE_X17Y106_AO5),
.O6(CLBLM_L_X12Y106_SLICE_X17Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h87e1ff55781e00aa)
  ) CLBLM_L_X12Y107_SLICE_X16Y107_DLUT (
.I0(CLBLM_L_X12Y106_SLICE_X16Y106_AO6),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(RIOB33_X105Y107_IOB_X1Y107_I),
.I3(CLBLM_L_X12Y107_SLICE_X16Y107_AO5),
.I4(LIOB33_X0Y101_IOB_X0Y102_I),
.I5(CLBLM_L_X12Y107_SLICE_X16Y107_BO6),
.O5(CLBLM_L_X12Y107_SLICE_X16Y107_DO5),
.O6(CLBLM_L_X12Y107_SLICE_X16Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h202200007d228888)
  ) CLBLM_L_X12Y107_SLICE_X16Y107_CLUT (
.I0(RIOB33_X105Y107_IOB_X1Y107_I),
.I1(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I2(RIOB33_X105Y111_IOB_X1Y112_I),
.I3(RIOB33_X105Y107_IOB_X1Y108_I),
.I4(RIOB33_X105Y113_IOB_X1Y113_I),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X12Y107_SLICE_X16Y107_CO5),
.O6(CLBLM_L_X12Y107_SLICE_X16Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h55ffad07aa0052f8)
  ) CLBLM_L_X12Y107_SLICE_X16Y107_BLUT (
.I0(LIOB33_X0Y101_IOB_X0Y101_I),
.I1(RIOB33_X105Y107_IOB_X1Y107_I),
.I2(CLBLM_L_X12Y107_SLICE_X17Y107_AO6),
.I3(RIOB33_X105Y107_IOB_X1Y108_I),
.I4(CLBLM_L_X12Y106_SLICE_X16Y106_BO6),
.I5(CLBLM_R_X11Y107_SLICE_X14Y107_DO6),
.O5(CLBLM_L_X12Y107_SLICE_X16Y107_BO5),
.O6(CLBLM_L_X12Y107_SLICE_X16Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc333c333ffff0333)
  ) CLBLM_L_X12Y107_SLICE_X16Y107_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X12Y107_SLICE_X17Y107_BO6),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(LIOB33_X0Y101_IOB_X0Y101_I),
.I4(CLBLM_L_X12Y107_SLICE_X16Y107_CO6),
.I5(1'b1),
.O5(CLBLM_L_X12Y107_SLICE_X16Y107_AO5),
.O6(CLBLM_L_X12Y107_SLICE_X16Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y107_SLICE_X17Y107_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y107_SLICE_X17Y107_DO5),
.O6(CLBLM_L_X12Y107_SLICE_X17Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y107_SLICE_X17Y107_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y107_SLICE_X17Y107_CO5),
.O6(CLBLM_L_X12Y107_SLICE_X17Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h073c880c43f0ccc0)
  ) CLBLM_L_X12Y107_SLICE_X17Y107_BLUT (
.I0(RIOB33_X105Y111_IOB_X1Y112_I),
.I1(RIOB33_X105Y113_IOB_X1Y113_I),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(RIOB33_X105Y107_IOB_X1Y107_I),
.I4(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I5(RIOB33_X105Y107_IOB_X1Y108_I),
.O5(CLBLM_L_X12Y107_SLICE_X17Y107_BO5),
.O6(CLBLM_L_X12Y107_SLICE_X17Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h074388cc3cf00cc0)
  ) CLBLM_L_X12Y107_SLICE_X17Y107_ALUT (
.I0(RIOB33_X105Y111_IOB_X1Y112_I),
.I1(RIOB33_X105Y113_IOB_X1Y113_I),
.I2(RIOB33_X105Y107_IOB_X1Y107_I),
.I3(RIOB33_X105Y109_IOB_X1Y109_I),
.I4(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I5(RIOB33_X105Y107_IOB_X1Y108_I),
.O5(CLBLM_L_X12Y107_SLICE_X17Y107_AO5),
.O6(CLBLM_L_X12Y107_SLICE_X17Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6a95956a956a956a)
  ) CLBLM_L_X12Y108_SLICE_X16Y108_DLUT (
.I0(CLBLM_R_X13Y108_SLICE_X19Y108_BO6),
.I1(LIOB33_X0Y103_IOB_X0Y104_I),
.I2(RIOB33_X105Y103_IOB_X1Y104_I),
.I3(CLBLM_R_X11Y108_SLICE_X15Y108_DO6),
.I4(RIOB33_X105Y103_IOB_X1Y103_I),
.I5(LIOB33_X0Y105_IOB_X0Y105_I),
.O5(CLBLM_L_X12Y108_SLICE_X16Y108_DO5),
.O6(CLBLM_L_X12Y108_SLICE_X16Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h2a80bfeabfeabfea)
  ) CLBLM_L_X12Y108_SLICE_X16Y108_CLUT (
.I0(CLBLM_R_X13Y108_SLICE_X19Y108_BO6),
.I1(RIOB33_X105Y103_IOB_X1Y104_I),
.I2(LIOB33_X0Y103_IOB_X0Y104_I),
.I3(CLBLM_R_X11Y108_SLICE_X15Y108_DO6),
.I4(RIOB33_X105Y103_IOB_X1Y103_I),
.I5(LIOB33_X0Y105_IOB_X0Y105_I),
.O5(CLBLM_L_X12Y108_SLICE_X16Y108_CO5),
.O6(CLBLM_L_X12Y108_SLICE_X16Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0fff0fff3f3f3f3f)
  ) CLBLM_L_X12Y108_SLICE_X16Y108_BLUT (
.I0(1'b1),
.I1(LIOB33_X0Y103_IOB_X0Y104_I),
.I2(RIOB33_X105Y103_IOB_X1Y104_I),
.I3(LIOB33_X0Y105_IOB_X0Y105_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y108_SLICE_X16Y108_BO5),
.O6(CLBLM_L_X12Y108_SLICE_X16Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f3f3f3f0fff0fff)
  ) CLBLM_L_X12Y108_SLICE_X16Y108_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y103_IOB_X0Y104_I),
.I2(RIOB33_X105Y101_IOB_X1Y102_I),
.I3(LIOB33_X0Y105_IOB_X0Y105_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y108_SLICE_X16Y108_AO5),
.O6(CLBLM_L_X12Y108_SLICE_X16Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6999966696669666)
  ) CLBLM_L_X12Y108_SLICE_X17Y108_DLUT (
.I0(CLBLM_R_X11Y107_SLICE_X14Y107_CO6),
.I1(CLBLM_R_X11Y107_SLICE_X15Y107_CO6),
.I2(RIOB33_X105Y103_IOB_X1Y104_I),
.I3(LIOB33_X0Y103_IOB_X0Y104_I),
.I4(LIOB33_X0Y101_IOB_X0Y102_I),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X12Y108_SLICE_X17Y108_DO5),
.O6(CLBLM_L_X12Y108_SLICE_X17Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hb37fd9154c8026ea)
  ) CLBLM_L_X12Y108_SLICE_X17Y108_CLUT (
.I0(CLBLM_R_X11Y106_SLICE_X15Y106_CO6),
.I1(LIOB33_X0Y105_IOB_X0Y105_I),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(RIOB33_X105Y107_IOB_X1Y107_I),
.I4(CLBLM_R_X13Y108_SLICE_X18Y108_AO6),
.I5(CLBLM_R_X11Y106_SLICE_X14Y106_BO6),
.O5(CLBLM_L_X12Y108_SLICE_X17Y108_CO5),
.O6(CLBLM_L_X12Y108_SLICE_X17Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h4d8ecf0cddeeffcc)
  ) CLBLM_L_X12Y108_SLICE_X17Y108_BLUT (
.I0(LIOB33_X0Y101_IOB_X0Y102_I),
.I1(CLBLM_R_X11Y107_SLICE_X14Y107_CO6),
.I2(RIOB33_X105Y103_IOB_X1Y104_I),
.I3(CLBLM_R_X11Y107_SLICE_X15Y107_CO6),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(LIOB33_X0Y103_IOB_X0Y104_I),
.O5(CLBLM_L_X12Y108_SLICE_X17Y108_BO5),
.O6(CLBLM_L_X12Y108_SLICE_X17Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h33ff33ff55ff55ff)
  ) CLBLM_L_X12Y108_SLICE_X17Y108_ALUT (
.I0(LIOB33_X0Y103_IOB_X0Y104_I),
.I1(LIOB33_X0Y105_IOB_X0Y105_I),
.I2(1'b1),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y108_SLICE_X17Y108_AO5),
.O6(CLBLM_L_X12Y108_SLICE_X17Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha659659a9a9a9a9a)
  ) CLBLM_L_X12Y109_SLICE_X16Y109_DLUT (
.I0(CLBLM_R_X11Y108_SLICE_X15Y108_CO6),
.I1(CLBLM_R_X13Y108_SLICE_X19Y108_BO6),
.I2(CLBLM_L_X12Y108_SLICE_X17Y108_DO6),
.I3(RIOB33_X105Y103_IOB_X1Y104_I),
.I4(RIOB33_X105Y103_IOB_X1Y103_I),
.I5(LIOB33_X0Y105_IOB_X0Y105_I),
.O5(CLBLM_L_X12Y109_SLICE_X16Y109_DO5),
.O6(CLBLM_L_X12Y109_SLICE_X16Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hefdfae5d8a450804)
  ) CLBLM_L_X12Y109_SLICE_X16Y109_CLUT (
.I0(CLBLM_R_X11Y108_SLICE_X15Y108_CO6),
.I1(CLBLM_R_X13Y108_SLICE_X19Y108_BO6),
.I2(CLBLM_L_X12Y108_SLICE_X17Y108_DO6),
.I3(CLBLM_L_X12Y108_SLICE_X16Y108_BO6),
.I4(CLBLM_R_X11Y108_SLICE_X15Y108_AO5),
.I5(CLBLM_L_X12Y110_SLICE_X16Y110_AO6),
.O5(CLBLM_L_X12Y109_SLICE_X16Y109_CO5),
.O6(CLBLM_L_X12Y109_SLICE_X16Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h2dd2d22db44b4bb4)
  ) CLBLM_L_X12Y109_SLICE_X16Y109_BLUT (
.I0(CLBLM_L_X12Y108_SLICE_X17Y108_DO6),
.I1(CLBLM_R_X13Y108_SLICE_X19Y108_BO6),
.I2(CLBLM_R_X11Y108_SLICE_X15Y108_CO6),
.I3(CLBLM_L_X12Y110_SLICE_X16Y110_AO6),
.I4(CLBLM_L_X12Y108_SLICE_X16Y108_BO6),
.I5(CLBLM_R_X11Y108_SLICE_X15Y108_AO5),
.O5(CLBLM_L_X12Y109_SLICE_X16Y109_BO5),
.O6(CLBLM_L_X12Y109_SLICE_X16Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0fffff5555ffff)
  ) CLBLM_L_X12Y109_SLICE_X16Y109_ALUT (
.I0(LIOB33_X0Y107_IOB_X0Y107_I),
.I1(1'b1),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(1'b1),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_L_X12Y109_SLICE_X16Y109_AO5),
.O6(CLBLM_L_X12Y109_SLICE_X16Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h60c0f6fcf6fcf6fc)
  ) CLBLM_L_X12Y109_SLICE_X17Y109_DLUT (
.I0(RIOB33_X105Y107_IOB_X1Y107_I),
.I1(CLBLM_L_X12Y106_SLICE_X16Y106_CO6),
.I2(CLBLM_R_X13Y108_SLICE_X18Y108_AO6),
.I3(LIOB33_X0Y103_IOB_X0Y104_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(LIOB33_X0Y105_IOB_X0Y105_I),
.O5(CLBLM_L_X12Y109_SLICE_X17Y109_DO5),
.O6(CLBLM_L_X12Y109_SLICE_X17Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h695a96a5a5695a96)
  ) CLBLM_L_X12Y109_SLICE_X17Y109_CLUT (
.I0(CLBLM_L_X12Y109_SLICE_X17Y109_AO6),
.I1(CLBLM_L_X12Y108_SLICE_X16Y108_BO6),
.I2(CLBLM_R_X11Y106_SLICE_X15Y106_DO6),
.I3(CLBLM_R_X13Y108_SLICE_X18Y108_BO6),
.I4(CLBLM_L_X12Y108_SLICE_X17Y108_AO6),
.I5(CLBLM_L_X12Y108_SLICE_X17Y108_BO6),
.O5(CLBLM_L_X12Y109_SLICE_X17Y109_CO5),
.O6(CLBLM_L_X12Y109_SLICE_X17Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'head58040fefda854)
  ) CLBLM_L_X12Y109_SLICE_X17Y109_BLUT (
.I0(CLBLM_R_X11Y106_SLICE_X15Y106_DO6),
.I1(CLBLM_L_X12Y108_SLICE_X17Y108_BO6),
.I2(CLBLM_L_X12Y108_SLICE_X16Y108_BO6),
.I3(CLBLM_L_X12Y108_SLICE_X17Y108_AO6),
.I4(CLBLM_L_X12Y109_SLICE_X17Y109_AO6),
.I5(CLBLM_R_X13Y108_SLICE_X18Y108_BO6),
.O5(CLBLM_L_X12Y109_SLICE_X17Y109_BO5),
.O6(CLBLM_L_X12Y109_SLICE_X17Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f3f3f3f77777777)
  ) CLBLM_L_X12Y109_SLICE_X17Y109_ALUT (
.I0(LIOB33_X0Y107_IOB_X0Y107_I),
.I1(RIOB33_X105Y103_IOB_X1Y104_I),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y109_SLICE_X17Y109_AO5),
.O6(CLBLM_L_X12Y109_SLICE_X17Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h9f5f60a0a3935c6c)
  ) CLBLM_L_X12Y110_SLICE_X16Y110_DLUT (
.I0(RIOB33_X105Y107_IOB_X1Y107_I),
.I1(CLBLM_R_X11Y109_SLICE_X14Y109_AO5),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X11Y109_SLICE_X14Y109_CO6),
.I5(CLBLM_L_X12Y109_SLICE_X17Y109_DO6),
.O5(CLBLM_L_X12Y110_SLICE_X16Y110_DO5),
.O6(CLBLM_L_X12Y110_SLICE_X16Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7df5ffff14503cf0)
  ) CLBLM_L_X12Y110_SLICE_X16Y110_CLUT (
.I0(RIOB33_X105Y103_IOB_X1Y104_I),
.I1(LIOB33_X0Y103_IOB_X0Y104_I),
.I2(CLBLM_L_X12Y107_SLICE_X16Y107_DO6),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(LIOB33_X0Y105_IOB_X0Y105_I),
.I5(CLBLM_L_X12Y108_SLICE_X17Y108_BO6),
.O5(CLBLM_L_X12Y110_SLICE_X16Y110_CO5),
.O6(CLBLM_L_X12Y110_SLICE_X16Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h4ddd8eeecfff0ccc)
  ) CLBLM_L_X12Y110_SLICE_X16Y110_BLUT (
.I0(RIOB33_X105Y103_IOB_X1Y103_I),
.I1(CLBLM_L_X10Y107_SLICE_X13Y107_AO6),
.I2(RIOB33_X105Y101_IOB_X1Y102_I),
.I3(LIOB33_X0Y105_IOB_X0Y105_I),
.I4(CLBLM_R_X11Y108_SLICE_X14Y108_DO6),
.I5(LIOB33_X0Y103_IOB_X0Y104_I),
.O5(CLBLM_L_X12Y110_SLICE_X16Y110_BO5),
.O6(CLBLM_L_X12Y110_SLICE_X16Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h55ff55ff5f5f5f5f)
  ) CLBLM_L_X12Y110_SLICE_X16Y110_ALUT (
.I0(RIOB33_X105Y103_IOB_X1Y103_I),
.I1(1'b1),
.I2(LIOB33_X0Y107_IOB_X0Y108_I),
.I3(LIOB33_X0Y105_IOB_X0Y106_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y110_SLICE_X16Y110_AO5),
.O6(CLBLM_L_X12Y110_SLICE_X16Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6ac0953f953f6ac0)
  ) CLBLM_L_X12Y110_SLICE_X17Y110_DLUT (
.I0(RIOB33_X105Y107_IOB_X1Y107_I),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(LIOB33_X0Y105_IOB_X0Y105_I),
.I3(LIOB33_X0Y103_IOB_X0Y104_I),
.I4(CLBLM_R_X13Y108_SLICE_X18Y108_AO6),
.I5(CLBLM_L_X12Y106_SLICE_X16Y106_CO6),
.O5(CLBLM_L_X12Y110_SLICE_X17Y110_DO5),
.O6(CLBLM_L_X12Y110_SLICE_X17Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hb4783cf0d21e965a)
  ) CLBLM_L_X12Y110_SLICE_X17Y110_CLUT (
.I0(CLBLM_R_X13Y108_SLICE_X18Y108_BO6),
.I1(LIOB33_X0Y105_IOB_X0Y105_I),
.I2(CLBLM_R_X11Y106_SLICE_X15Y106_DO6),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(RIOB33_X105Y103_IOB_X1Y104_I),
.I5(CLBLM_L_X12Y108_SLICE_X17Y108_BO6),
.O5(CLBLM_L_X12Y110_SLICE_X17Y110_CO5),
.O6(CLBLM_L_X12Y110_SLICE_X17Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6999966696669666)
  ) CLBLM_L_X12Y110_SLICE_X17Y110_BLUT (
.I0(CLBLM_L_X12Y107_SLICE_X16Y107_DO6),
.I1(CLBLM_L_X12Y108_SLICE_X17Y108_BO6),
.I2(RIOB33_X105Y103_IOB_X1Y104_I),
.I3(LIOB33_X0Y105_IOB_X0Y105_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(LIOB33_X0Y103_IOB_X0Y104_I),
.O5(CLBLM_L_X12Y110_SLICE_X17Y110_BO5),
.O6(CLBLM_L_X12Y110_SLICE_X17Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hd75f28a0a0d75f28)
  ) CLBLM_L_X12Y110_SLICE_X17Y110_ALUT (
.I0(RIOB33_X105Y103_IOB_X1Y103_I),
.I1(LIOB33_X0Y105_IOB_X0Y106_I),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(CLBLM_L_X12Y110_SLICE_X17Y110_BO6),
.I4(CLBLM_L_X12Y109_SLICE_X17Y109_CO6),
.I5(CLBLM_L_X12Y108_SLICE_X16Y108_CO6),
.O5(CLBLM_L_X12Y110_SLICE_X17Y110_AO5),
.O6(CLBLM_L_X12Y110_SLICE_X17Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'he14b78d269c35af0)
  ) CLBLM_L_X12Y111_SLICE_X16Y111_DLUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(CLBLM_L_X12Y110_SLICE_X16Y110_CO6),
.I2(CLBLM_L_X12Y108_SLICE_X17Y108_CO6),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_L_X12Y110_SLICE_X17Y110_DO6),
.I5(RIOB33_X105Y103_IOB_X1Y104_I),
.O5(CLBLM_L_X12Y111_SLICE_X16Y111_DO5),
.O6(CLBLM_L_X12Y111_SLICE_X16Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h87f078f0e13c1e3c)
  ) CLBLM_L_X12Y111_SLICE_X16Y111_CLUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(CLBLM_L_X12Y108_SLICE_X16Y108_DO6),
.I2(CLBLM_L_X12Y109_SLICE_X16Y109_BO6),
.I3(RIOB33_X105Y101_IOB_X1Y102_I),
.I4(LIOB33_X0Y107_IOB_X0Y107_I),
.I5(CLBLM_L_X12Y110_SLICE_X16Y110_BO6),
.O5(CLBLM_L_X12Y111_SLICE_X16Y111_CO5),
.O6(CLBLM_L_X12Y111_SLICE_X16Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hb48778b478877878)
  ) CLBLM_L_X12Y111_SLICE_X16Y111_BLUT (
.I0(RIOB33_X105Y103_IOB_X1Y103_I),
.I1(LIOB33_X0Y105_IOB_X0Y106_I),
.I2(CLBLM_L_X12Y109_SLICE_X16Y109_DO6),
.I3(CLBLM_L_X12Y110_SLICE_X16Y110_BO6),
.I4(CLBLM_L_X12Y108_SLICE_X16Y108_DO6),
.I5(RIOB33_X105Y101_IOB_X1Y102_I),
.O5(CLBLM_L_X12Y111_SLICE_X16Y111_BO5),
.O6(CLBLM_L_X12Y111_SLICE_X16Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h032b2b3fbbbbffff)
  ) CLBLM_L_X12Y111_SLICE_X16Y111_ALUT (
.I0(CLBLM_L_X12Y110_SLICE_X16Y110_BO6),
.I1(CLBLM_L_X12Y109_SLICE_X16Y109_BO6),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(LIOB33_X0Y105_IOB_X0Y106_I),
.I4(CLBLM_L_X12Y108_SLICE_X16Y108_DO6),
.I5(RIOB33_X105Y101_IOB_X1Y102_I),
.O5(CLBLM_L_X12Y111_SLICE_X16Y111_AO5),
.O6(CLBLM_L_X12Y111_SLICE_X16Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y111_SLICE_X17Y111_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y111_SLICE_X17Y111_DO5),
.O6(CLBLM_L_X12Y111_SLICE_X17Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y111_SLICE_X17Y111_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y111_SLICE_X17Y111_CO5),
.O6(CLBLM_L_X12Y111_SLICE_X17Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y111_SLICE_X17Y111_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y111_SLICE_X17Y111_BO5),
.O6(CLBLM_L_X12Y111_SLICE_X17Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y111_SLICE_X17Y111_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y111_SLICE_X17Y111_AO5),
.O6(CLBLM_L_X12Y111_SLICE_X17Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y104_SLICE_X2Y104_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y104_SLICE_X2Y104_DO5),
.O6(CLBLM_R_X3Y104_SLICE_X2Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y104_SLICE_X2Y104_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y104_SLICE_X2Y104_CO5),
.O6(CLBLM_R_X3Y104_SLICE_X2Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y104_SLICE_X2Y104_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y104_SLICE_X2Y104_BO5),
.O6(CLBLM_R_X3Y104_SLICE_X2Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y104_SLICE_X2Y104_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y104_SLICE_X2Y104_AO5),
.O6(CLBLM_R_X3Y104_SLICE_X2Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5a5aa5a596a5695a)
  ) CLBLM_R_X3Y104_SLICE_X3Y104_DLUT (
.I0(CLBLM_R_X3Y104_SLICE_X3Y104_AO6),
.I1(CLBLM_R_X3Y105_SLICE_X2Y105_AO6),
.I2(CLBLM_R_X5Y104_SLICE_X6Y104_AO6),
.I3(CLBLM_R_X3Y104_SLICE_X3Y104_AO5),
.I4(CLBLL_L_X4Y105_SLICE_X4Y105_AO6),
.I5(CLBLM_R_X3Y104_SLICE_X3Y104_BO6),
.O5(CLBLM_R_X3Y104_SLICE_X3Y104_DO5),
.O6(CLBLM_R_X3Y104_SLICE_X3Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafaafafb2a02b0a)
  ) CLBLM_R_X3Y104_SLICE_X3Y104_CLUT (
.I0(CLBLM_R_X3Y104_SLICE_X3Y104_AO6),
.I1(CLBLM_R_X3Y105_SLICE_X2Y105_AO6),
.I2(CLBLM_R_X5Y104_SLICE_X6Y104_AO6),
.I3(CLBLM_R_X3Y104_SLICE_X3Y104_AO5),
.I4(CLBLL_L_X4Y105_SLICE_X4Y105_AO6),
.I5(CLBLM_R_X3Y104_SLICE_X3Y104_BO6),
.O5(CLBLM_R_X3Y104_SLICE_X3Y104_CO5),
.O6(CLBLM_R_X3Y104_SLICE_X3Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h550a0c00190a0c00)
  ) CLBLM_R_X3Y104_SLICE_X3Y104_BLUT (
.I0(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(LIOB33_X0Y113_IOB_X0Y114_I),
.I3(RIOB33_X105Y113_IOB_X1Y113_I),
.I4(LIOB33_X0Y115_IOB_X0Y116_I),
.I5(RIOB33_X105Y111_IOB_X1Y112_I),
.O5(CLBLM_R_X3Y104_SLICE_X3Y104_BO5),
.O6(CLBLM_R_X3Y104_SLICE_X3Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0fff0fff55ff55ff)
  ) CLBLM_R_X3Y104_SLICE_X3Y104_ALUT (
.I0(LIOB33_X0Y101_IOB_X0Y101_I),
.I1(1'b1),
.I2(LIOB33_X0Y101_IOB_X0Y102_I),
.I3(LIOB33_X0Y113_IOB_X0Y114_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y104_SLICE_X3Y104_AO5),
.O6(CLBLM_R_X3Y104_SLICE_X3Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y105_SLICE_X2Y105_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y105_SLICE_X2Y105_DO5),
.O6(CLBLM_R_X3Y105_SLICE_X2Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y105_SLICE_X2Y105_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y105_SLICE_X2Y105_CO5),
.O6(CLBLM_R_X3Y105_SLICE_X2Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hd42baf502bd4af50)
  ) CLBLM_R_X3Y105_SLICE_X2Y105_BLUT (
.I0(CLBLL_L_X2Y106_SLICE_X0Y106_AO5),
.I1(LIOB33_X0Y103_IOB_X0Y103_I),
.I2(CLBLM_R_X3Y105_SLICE_X3Y105_AO6),
.I3(CLBLM_R_X3Y105_SLICE_X3Y105_CO6),
.I4(LIOB33_X0Y101_IOB_X0Y102_I),
.I5(LIOB33_X0Y113_IOB_X0Y114_I),
.O5(CLBLM_R_X3Y105_SLICE_X2Y105_BO5),
.O6(CLBLM_R_X3Y105_SLICE_X2Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h424e02ce6c60ac60)
  ) CLBLM_R_X3Y105_SLICE_X2Y105_ALUT (
.I0(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I1(RIOB33_X105Y113_IOB_X1Y113_I),
.I2(LIOB33_X0Y115_IOB_X0Y116_I),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(RIOB33_X105Y111_IOB_X1Y112_I),
.I5(LIOB33_X0Y113_IOB_X0Y114_I),
.O5(CLBLM_R_X3Y105_SLICE_X2Y105_AO5),
.O6(CLBLM_R_X3Y105_SLICE_X2Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6696996996996966)
  ) CLBLM_R_X3Y105_SLICE_X3Y105_DLUT (
.I0(CLBLM_R_X3Y104_SLICE_X3Y104_CO6),
.I1(CLBLL_L_X4Y105_SLICE_X4Y105_BO6),
.I2(CLBLM_R_X3Y104_SLICE_X3Y104_DO6),
.I3(CLBLL_L_X2Y106_SLICE_X0Y106_CO6),
.I4(CLBLM_R_X3Y105_SLICE_X3Y105_BO5),
.I5(CLBLM_R_X3Y105_SLICE_X3Y105_BO6),
.O5(CLBLM_R_X3Y105_SLICE_X3Y105_DO5),
.O6(CLBLM_R_X3Y105_SLICE_X3Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6c6c6c6c939c936c)
  ) CLBLM_R_X3Y105_SLICE_X3Y105_CLUT (
.I0(LIOB33_X0Y115_IOB_X0Y116_I),
.I1(CLBLM_R_X5Y104_SLICE_X6Y104_AO6),
.I2(LIOB33_X0Y101_IOB_X0Y101_I),
.I3(CLBLM_R_X3Y105_SLICE_X2Y105_AO6),
.I4(LIOB33_X0Y113_IOB_X0Y114_I),
.I5(CLBLM_R_X3Y104_SLICE_X3Y104_BO6),
.O5(CLBLM_R_X3Y105_SLICE_X3Y105_CO5),
.O6(CLBLM_R_X3Y105_SLICE_X3Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f3f3f3f5f5f5f5f)
  ) CLBLM_R_X3Y105_SLICE_X3Y105_BLUT (
.I0(LIOB33_X0Y113_IOB_X0Y114_I),
.I1(LIOB33_X0Y103_IOB_X0Y103_I),
.I2(LIOB33_X0Y103_IOB_X0Y104_I),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y105_SLICE_X3Y105_BO5),
.O6(CLBLM_R_X3Y105_SLICE_X3Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h87878787ff07ff07)
  ) CLBLM_R_X3Y105_SLICE_X3Y105_ALUT (
.I0(LIOB33_X0Y113_IOB_X0Y114_I),
.I1(LIOB33_X0Y101_IOB_X0Y101_I),
.I2(CLBLM_R_X3Y105_SLICE_X2Y105_AO6),
.I3(CLBLM_R_X3Y104_SLICE_X3Y104_BO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y105_SLICE_X3Y105_AO5),
.O6(CLBLM_R_X3Y105_SLICE_X3Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hee8e8e88dd4d4d44)
  ) CLBLM_R_X3Y106_SLICE_X2Y106_DLUT (
.I0(CLBLM_R_X3Y106_SLICE_X2Y106_AO6),
.I1(CLBLL_L_X2Y107_SLICE_X1Y107_AO6),
.I2(CLBLM_R_X3Y106_SLICE_X2Y106_CO6),
.I3(CLBLM_R_X3Y106_SLICE_X2Y106_AO5),
.I4(CLBLL_L_X2Y108_SLICE_X1Y108_DO6),
.I5(CLBLL_L_X2Y106_SLICE_X1Y106_DO6),
.O5(CLBLM_R_X3Y106_SLICE_X2Y106_DO5),
.O6(CLBLM_R_X3Y106_SLICE_X2Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h69969966a55a55aa)
  ) CLBLM_R_X3Y106_SLICE_X2Y106_CLUT (
.I0(CLBLL_L_X2Y106_SLICE_X1Y106_BO6),
.I1(LIOB33_X0Y101_IOB_X0Y102_I),
.I2(LIOB33_X0Y103_IOB_X0Y104_I),
.I3(CLBLL_L_X2Y107_SLICE_X0Y107_DO6),
.I4(RIOB33_X105Y105_IOB_X1Y106_I),
.I5(LIOB33_X0Y103_IOB_X0Y103_I),
.O5(CLBLM_R_X3Y106_SLICE_X2Y106_CO5),
.O6(CLBLM_R_X3Y106_SLICE_X2Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7ff7f7f707707070)
  ) CLBLM_R_X3Y106_SLICE_X2Y106_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y106_I),
.I1(LIOB33_X0Y103_IOB_X0Y104_I),
.I2(CLBLL_L_X2Y106_SLICE_X1Y106_BO6),
.I3(LIOB33_X0Y103_IOB_X0Y103_I),
.I4(LIOB33_X0Y101_IOB_X0Y102_I),
.I5(CLBLL_L_X2Y107_SLICE_X0Y107_DO6),
.O5(CLBLM_R_X3Y106_SLICE_X2Y106_BO5),
.O6(CLBLM_R_X3Y106_SLICE_X2Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h55ff55ff33ff33ff)
  ) CLBLM_R_X3Y106_SLICE_X2Y106_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y106_I),
.I1(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I2(1'b1),
.I3(LIOB33_X0Y105_IOB_X0Y105_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y106_SLICE_X2Y106_AO5),
.O6(CLBLM_R_X3Y106_SLICE_X2Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h4114c33c14143c3c)
  ) CLBLM_R_X3Y106_SLICE_X3Y106_DLUT (
.I0(LIOB33_X0Y103_IOB_X0Y103_I),
.I1(CLBLM_R_X3Y105_SLICE_X3Y105_CO6),
.I2(CLBLL_L_X2Y106_SLICE_X0Y106_CO6),
.I3(LIOB33_X0Y101_IOB_X0Y102_I),
.I4(LIOB33_X0Y103_IOB_X0Y104_I),
.I5(LIOB33_X0Y113_IOB_X0Y114_I),
.O5(CLBLM_R_X3Y106_SLICE_X3Y106_DO5),
.O6(CLBLM_R_X3Y106_SLICE_X3Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h144150053cc3f00f)
  ) CLBLM_R_X3Y106_SLICE_X3Y106_CLUT (
.I0(LIOB33_X0Y103_IOB_X0Y104_I),
.I1(LIOB33_X0Y113_IOB_X0Y114_I),
.I2(CLBLL_L_X2Y106_SLICE_X0Y106_CO6),
.I3(CLBLM_R_X3Y105_SLICE_X3Y105_CO6),
.I4(LIOB33_X0Y101_IOB_X0Y102_I),
.I5(LIOB33_X0Y103_IOB_X0Y103_I),
.O5(CLBLM_R_X3Y106_SLICE_X3Y106_CO5),
.O6(CLBLM_R_X3Y106_SLICE_X3Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fff0777f7777000)
  ) CLBLM_R_X3Y106_SLICE_X3Y106_BLUT (
.I0(LIOB33_X0Y103_IOB_X0Y104_I),
.I1(LIOB33_X0Y103_IOB_X0Y103_I),
.I2(LIOB33_X0Y101_IOB_X0Y102_I),
.I3(LIOB33_X0Y113_IOB_X0Y114_I),
.I4(CLBLL_L_X2Y106_SLICE_X0Y106_CO6),
.I5(CLBLM_R_X3Y105_SLICE_X3Y105_CO6),
.O5(CLBLM_R_X3Y106_SLICE_X3Y106_BO5),
.O6(CLBLM_R_X3Y106_SLICE_X3Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h936c5fa06c93a05f)
  ) CLBLM_R_X3Y106_SLICE_X3Y106_ALUT (
.I0(LIOB33_X0Y103_IOB_X0Y104_I),
.I1(LIOB33_X0Y113_IOB_X0Y114_I),
.I2(LIOB33_X0Y103_IOB_X0Y103_I),
.I3(CLBLL_L_X2Y106_SLICE_X0Y106_CO6),
.I4(LIOB33_X0Y101_IOB_X0Y102_I),
.I5(CLBLM_R_X3Y105_SLICE_X3Y105_CO6),
.O5(CLBLM_R_X3Y106_SLICE_X3Y106_AO5),
.O6(CLBLM_R_X3Y106_SLICE_X3Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7df51450ffff3cf0)
  ) CLBLM_R_X3Y107_SLICE_X2Y107_DLUT (
.I0(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I1(LIOB33_X0Y105_IOB_X0Y106_I),
.I2(CLBLL_L_X4Y106_SLICE_X4Y106_BO6),
.I3(RIOB33_X105Y105_IOB_X1Y106_I),
.I4(CLBLM_R_X3Y106_SLICE_X2Y106_DO6),
.I5(LIOB33_X0Y107_IOB_X0Y107_I),
.O5(CLBLM_R_X3Y107_SLICE_X2Y107_DO5),
.O6(CLBLM_R_X3Y107_SLICE_X2Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hb748c03f3fc0b748)
  ) CLBLM_R_X3Y107_SLICE_X2Y107_CLUT (
.I0(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I1(LIOB33_X0Y105_IOB_X0Y106_I),
.I2(RIOB33_X105Y105_IOB_X1Y106_I),
.I3(CLBLL_L_X4Y106_SLICE_X4Y106_BO6),
.I4(CLBLL_L_X2Y107_SLICE_X1Y107_CO6),
.I5(CLBLM_R_X3Y107_SLICE_X2Y107_BO6),
.O5(CLBLM_R_X3Y107_SLICE_X2Y107_CO5),
.O6(CLBLM_R_X3Y107_SLICE_X2Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6c93936c93936c6c)
  ) CLBLM_R_X3Y107_SLICE_X2Y107_BLUT (
.I0(LIOB33_X0Y103_IOB_X0Y104_I),
.I1(CLBLM_R_X3Y105_SLICE_X2Y105_BO6),
.I2(LIOB33_X0Y103_IOB_X0Y103_I),
.I3(RIOB33_X105Y105_IOB_X1Y106_I),
.I4(CLBLM_R_X3Y106_SLICE_X2Y106_BO6),
.I5(LIOB33_X0Y105_IOB_X0Y105_I),
.O5(CLBLM_R_X3Y107_SLICE_X2Y107_BO5),
.O6(CLBLM_R_X3Y107_SLICE_X2Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0000fff33ff33ff)
  ) CLBLM_R_X3Y107_SLICE_X2Y107_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y103_IOB_X0Y103_I),
.I2(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I3(LIOB33_X0Y107_IOB_X0Y107_I),
.I4(CLBLM_R_X3Y107_SLICE_X2Y107_CO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y107_SLICE_X2Y107_AO5),
.O6(CLBLM_R_X3Y107_SLICE_X2Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000200000202)
  ) CLBLM_R_X3Y107_SLICE_X3Y107_DLUT (
.I0(CLBLM_L_X8Y107_SLICE_X11Y107_CO6),
.I1(CLBLM_R_X3Y106_SLICE_X3Y106_DO6),
.I2(CLBLL_L_X4Y106_SLICE_X4Y106_AO6),
.I3(LIOB33_X0Y103_IOB_X0Y104_I),
.I4(CLBLL_L_X4Y106_SLICE_X4Y106_BO6),
.I5(LIOB33_X0Y103_IOB_X0Y103_I),
.O5(CLBLM_R_X3Y107_SLICE_X3Y107_DO5),
.O6(CLBLM_R_X3Y107_SLICE_X3Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h2000000000000000)
  ) CLBLM_R_X3Y107_SLICE_X3Y107_CLUT (
.I0(CLBLM_L_X8Y107_SLICE_X11Y107_CO6),
.I1(CLBLL_L_X4Y106_SLICE_X4Y106_BO6),
.I2(CLBLM_R_X3Y108_SLICE_X3Y108_CO6),
.I3(RIOB33_X105Y105_IOB_X1Y106_I),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(CLBLM_R_X3Y106_SLICE_X3Y106_CO6),
.O5(CLBLM_R_X3Y107_SLICE_X3Y107_CO5),
.O6(CLBLM_R_X3Y107_SLICE_X3Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h71f3b230f5fffaf0)
  ) CLBLM_R_X3Y107_SLICE_X3Y107_BLUT (
.I0(LIOB33_X0Y103_IOB_X0Y104_I),
.I1(LIOB33_X0Y105_IOB_X0Y105_I),
.I2(CLBLM_R_X3Y106_SLICE_X2Y106_BO6),
.I3(LIOB33_X0Y103_IOB_X0Y103_I),
.I4(CLBLM_R_X3Y105_SLICE_X2Y105_BO6),
.I5(RIOB33_X105Y105_IOB_X1Y106_I),
.O5(CLBLM_R_X3Y107_SLICE_X3Y107_BO5),
.O6(CLBLM_R_X3Y107_SLICE_X3Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8fe37f13701c80ec)
  ) CLBLM_R_X3Y107_SLICE_X3Y107_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y106_I),
.I1(CLBLL_L_X4Y107_SLICE_X4Y107_AO6),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(CLBLM_R_X3Y107_SLICE_X3Y107_BO6),
.I4(LIOB33_X0Y103_IOB_X0Y103_I),
.I5(CLBLL_L_X4Y106_SLICE_X5Y106_BO6),
.O5(CLBLM_R_X3Y107_SLICE_X3Y107_AO5),
.O6(CLBLM_R_X3Y107_SLICE_X3Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y108_SLICE_X2Y108_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y108_SLICE_X2Y108_DO5),
.O6(CLBLM_R_X3Y108_SLICE_X2Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y108_SLICE_X2Y108_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y108_SLICE_X2Y108_CO5),
.O6(CLBLM_R_X3Y108_SLICE_X2Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y108_SLICE_X2Y108_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y108_SLICE_X2Y108_BO5),
.O6(CLBLM_R_X3Y108_SLICE_X2Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y108_SLICE_X2Y108_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y108_SLICE_X2Y108_AO5),
.O6(CLBLM_R_X3Y108_SLICE_X2Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y108_SLICE_X3Y108_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y108_SLICE_X3Y108_DO5),
.O6(CLBLM_R_X3Y108_SLICE_X3Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h122121215aa5a5a5)
  ) CLBLM_R_X3Y108_SLICE_X3Y108_CLUT (
.I0(CLBLM_R_X3Y107_SLICE_X3Y107_AO6),
.I1(LIOB33_X0Y107_IOB_X0Y108_I),
.I2(CLBLM_R_X3Y107_SLICE_X2Y107_DO6),
.I3(LIOB33_X0Y107_IOB_X0Y107_I),
.I4(RIOB33_X105Y105_IOB_X1Y106_I),
.I5(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.O5(CLBLM_R_X3Y108_SLICE_X3Y108_CO5),
.O6(CLBLM_R_X3Y108_SLICE_X3Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h2bafb2fab2fab2fa)
  ) CLBLM_R_X3Y108_SLICE_X3Y108_BLUT (
.I0(CLBLM_R_X3Y107_SLICE_X2Y107_DO6),
.I1(LIOB33_X0Y107_IOB_X0Y108_I),
.I2(CLBLM_R_X3Y107_SLICE_X3Y107_AO6),
.I3(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I4(RIOB33_X105Y105_IOB_X1Y106_I),
.I5(LIOB33_X0Y107_IOB_X0Y107_I),
.O5(CLBLM_R_X3Y108_SLICE_X3Y108_BO5),
.O6(CLBLM_R_X3Y108_SLICE_X3Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996a55a96965a5a)
  ) CLBLM_R_X3Y108_SLICE_X3Y108_ALUT (
.I0(CLBLM_R_X3Y107_SLICE_X2Y107_DO6),
.I1(LIOB33_X0Y107_IOB_X0Y108_I),
.I2(CLBLM_R_X3Y107_SLICE_X3Y107_AO6),
.I3(RIOB33_X105Y105_IOB_X1Y106_I),
.I4(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I5(LIOB33_X0Y107_IOB_X0Y107_I),
.O5(CLBLM_R_X3Y108_SLICE_X3Y108_AO5),
.O6(CLBLM_R_X3Y108_SLICE_X3Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y109_SLICE_X2Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y109_SLICE_X2Y109_DO5),
.O6(CLBLM_R_X3Y109_SLICE_X2Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y109_SLICE_X2Y109_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y109_SLICE_X2Y109_CO5),
.O6(CLBLM_R_X3Y109_SLICE_X2Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y109_SLICE_X2Y109_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y109_SLICE_X2Y109_BO5),
.O6(CLBLM_R_X3Y109_SLICE_X2Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y109_SLICE_X2Y109_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y109_SLICE_X2Y109_AO5),
.O6(CLBLM_R_X3Y109_SLICE_X2Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y109_SLICE_X3Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y109_SLICE_X3Y109_DO5),
.O6(CLBLM_R_X3Y109_SLICE_X3Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y109_SLICE_X3Y109_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y109_SLICE_X3Y109_CO5),
.O6(CLBLM_R_X3Y109_SLICE_X3Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y109_SLICE_X3Y109_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y109_SLICE_X3Y109_BO5),
.O6(CLBLM_R_X3Y109_SLICE_X3Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hb777488888b77748)
  ) CLBLM_R_X3Y109_SLICE_X3Y109_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y106_I),
.I1(LIOB33_X0Y109_IOB_X0Y109_I),
.I2(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I3(CLBLL_L_X4Y108_SLICE_X4Y108_AO6),
.I4(CLBLL_L_X4Y108_SLICE_X4Y108_BO6),
.I5(CLBLM_R_X3Y108_SLICE_X3Y108_BO6),
.O5(CLBLM_R_X3Y109_SLICE_X3Y109_AO5),
.O6(CLBLM_R_X3Y109_SLICE_X3Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y110_SLICE_X2Y110_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y110_SLICE_X2Y110_DO5),
.O6(CLBLM_R_X3Y110_SLICE_X2Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y110_SLICE_X2Y110_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y110_SLICE_X2Y110_CO5),
.O6(CLBLM_R_X3Y110_SLICE_X2Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y110_SLICE_X2Y110_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y110_SLICE_X2Y110_BO5),
.O6(CLBLM_R_X3Y110_SLICE_X2Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y110_SLICE_X2Y110_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y110_SLICE_X2Y110_AO5),
.O6(CLBLM_R_X3Y110_SLICE_X2Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hbcd0cc6c701c00a0)
  ) CLBLM_R_X3Y110_SLICE_X3Y110_DLUT (
.I0(LIOB33_X0Y107_IOB_X0Y108_I),
.I1(RIOB33_X105Y109_IOB_X1Y110_I),
.I2(RIOB33_X105Y111_IOB_X1Y111_I),
.I3(CLBLL_L_X4Y110_SLICE_X5Y110_CO6),
.I4(LIOB33_X0Y109_IOB_X0Y109_I),
.I5(LIOB33_X0Y109_IOB_X0Y110_I),
.O5(CLBLM_R_X3Y110_SLICE_X3Y110_DO5),
.O6(CLBLM_R_X3Y110_SLICE_X3Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0200220008008800)
  ) CLBLM_R_X3Y110_SLICE_X3Y110_CLUT (
.I0(CLBLM_R_X3Y108_SLICE_X3Y108_CO6),
.I1(CLBLM_R_X5Y109_SLICE_X7Y109_CO6),
.I2(LIOB33_X0Y111_IOB_X0Y111_I),
.I3(CLBLM_R_X3Y107_SLICE_X3Y107_DO6),
.I4(RIOB33_X105Y107_IOB_X1Y108_I),
.I5(CLBLM_R_X5Y110_SLICE_X6Y110_AO6),
.O5(CLBLM_R_X3Y110_SLICE_X3Y110_CO5),
.O6(CLBLM_R_X3Y110_SLICE_X3Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7887877888777788)
  ) CLBLM_R_X3Y110_SLICE_X3Y110_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y106_I),
.I1(LIOB33_X0Y109_IOB_X0Y110_I),
.I2(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I3(CLBLL_L_X4Y109_SLICE_X5Y109_AO6),
.I4(CLBLL_L_X4Y109_SLICE_X4Y109_BO6),
.I5(LIOB33_X0Y111_IOB_X0Y111_I),
.O5(CLBLM_R_X3Y110_SLICE_X3Y110_BO5),
.O6(CLBLM_R_X3Y110_SLICE_X3Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c03f3f77777777)
  ) CLBLM_R_X3Y110_SLICE_X3Y110_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y106_I),
.I1(LIOB33_X0Y109_IOB_X0Y110_I),
.I2(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I3(1'b1),
.I4(CLBLM_R_X3Y109_SLICE_X3Y109_AO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y110_SLICE_X3Y110_AO5),
.O6(CLBLM_R_X3Y110_SLICE_X3Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h223b2a3f3fbfbfff)
  ) CLBLM_R_X3Y111_SLICE_X2Y111_DLUT (
.I0(CLBLL_L_X4Y110_SLICE_X5Y110_AO6),
.I1(RIOB33_X105Y109_IOB_X1Y109_I),
.I2(LIOB33_X0Y113_IOB_X0Y113_I),
.I3(CLBLM_R_X3Y111_SLICE_X2Y111_AO5),
.I4(LIOB33_X0Y111_IOB_X0Y112_I),
.I5(CLBLL_L_X2Y111_SLICE_X1Y111_AO6),
.O5(CLBLM_R_X3Y111_SLICE_X2Y111_DO5),
.O6(CLBLM_R_X3Y111_SLICE_X2Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hca6f6a3f359095c0)
  ) CLBLM_R_X3Y111_SLICE_X2Y111_CLUT (
.I0(CLBLL_L_X4Y110_SLICE_X5Y110_AO6),
.I1(LIOB33_X0Y113_IOB_X0Y113_I),
.I2(RIOB33_X105Y109_IOB_X1Y109_I),
.I3(CLBLM_R_X3Y111_SLICE_X2Y111_AO5),
.I4(LIOB33_X0Y111_IOB_X0Y112_I),
.I5(CLBLL_L_X2Y111_SLICE_X1Y111_AO6),
.O5(CLBLM_R_X3Y111_SLICE_X2Y111_CO5),
.O6(CLBLM_R_X3Y111_SLICE_X2Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6c93936c93936c6c)
  ) CLBLM_R_X3Y111_SLICE_X2Y111_BLUT (
.I0(RIOB33_X105Y109_IOB_X1Y109_I),
.I1(CLBLM_R_X3Y111_SLICE_X3Y111_DO6),
.I2(LIOB33_X0Y111_IOB_X0Y112_I),
.I3(LIOB33_X0Y111_IOB_X0Y111_I),
.I4(CLBLL_L_X4Y110_SLICE_X5Y110_AO6),
.I5(RIOB33_X105Y109_IOB_X1Y110_I),
.O5(CLBLM_R_X3Y111_SLICE_X2Y111_BO5),
.O6(CLBLM_R_X3Y111_SLICE_X2Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h55ff55ffc333c333)
  ) CLBLM_R_X3Y111_SLICE_X2Y111_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y106_I),
.I1(CLBLM_R_X3Y111_SLICE_X3Y111_DO6),
.I2(RIOB33_X105Y109_IOB_X1Y110_I),
.I3(LIOB33_X0Y111_IOB_X0Y111_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y111_SLICE_X2Y111_AO5),
.O6(CLBLM_R_X3Y111_SLICE_X2Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h88ffe8777fff57ff)
  ) CLBLM_R_X3Y111_SLICE_X3Y111_DLUT (
.I0(LIOB33_X0Y109_IOB_X0Y109_I),
.I1(RIOB33_X105Y109_IOB_X1Y110_I),
.I2(LIOB33_X0Y107_IOB_X0Y108_I),
.I3(RIOB33_X105Y111_IOB_X1Y111_I),
.I4(CLBLL_L_X4Y110_SLICE_X5Y110_CO6),
.I5(LIOB33_X0Y109_IOB_X0Y110_I),
.O5(CLBLM_R_X3Y111_SLICE_X3Y111_DO5),
.O6(CLBLM_R_X3Y111_SLICE_X3Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'heaaac000bfffeaaa)
  ) CLBLM_R_X3Y111_SLICE_X3Y111_CLUT (
.I0(CLBLL_L_X4Y113_SLICE_X4Y113_AO6),
.I1(CLBLM_R_X3Y112_SLICE_X3Y112_AO6),
.I2(CLBLM_R_X7Y111_SLICE_X8Y111_BO6),
.I3(CLBLM_R_X3Y110_SLICE_X3Y110_CO6),
.I4(CLBLL_L_X4Y110_SLICE_X4Y110_DO6),
.I5(CLBLM_R_X5Y110_SLICE_X6Y110_DO6),
.O5(CLBLM_R_X3Y111_SLICE_X3Y111_CO5),
.O6(CLBLM_R_X3Y111_SLICE_X3Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8f780ff00ff00ff0)
  ) CLBLM_R_X3Y111_SLICE_X3Y111_BLUT (
.I0(CLBLM_R_X7Y111_SLICE_X8Y111_BO6),
.I1(CLBLM_R_X3Y112_SLICE_X3Y112_AO6),
.I2(CLBLL_L_X4Y110_SLICE_X4Y110_DO6),
.I3(CLBLM_R_X5Y110_SLICE_X6Y110_DO6),
.I4(CLBLM_R_X3Y111_SLICE_X3Y111_AO6),
.I5(CLBLM_R_X3Y107_SLICE_X3Y107_CO6),
.O5(CLBLM_R_X3Y111_SLICE_X3Y111_BO5),
.O6(CLBLM_R_X3Y111_SLICE_X3Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h050f50f05af0a50f)
  ) CLBLM_R_X3Y111_SLICE_X3Y111_ALUT (
.I0(RIOB33_X105Y107_IOB_X1Y108_I),
.I1(1'b1),
.I2(CLBLM_R_X5Y110_SLICE_X6Y110_AO6),
.I3(LIOB33_X0Y111_IOB_X0Y111_I),
.I4(CLBLM_R_X5Y109_SLICE_X7Y109_CO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y111_SLICE_X3Y111_AO5),
.O6(CLBLM_R_X3Y111_SLICE_X3Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y112_SLICE_X2Y112_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y112_SLICE_X2Y112_DO5),
.O6(CLBLM_R_X3Y112_SLICE_X2Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y112_SLICE_X2Y112_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y112_SLICE_X2Y112_CO5),
.O6(CLBLM_R_X3Y112_SLICE_X2Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h507055f775fff7ff)
  ) CLBLM_R_X3Y112_SLICE_X2Y112_BLUT (
.I0(RIOB33_X105Y107_IOB_X1Y108_I),
.I1(LIOB33_X0Y113_IOB_X0Y113_I),
.I2(CLBLL_L_X4Y111_SLICE_X5Y111_DO6),
.I3(LIOB33_X0Y115_IOB_X0Y115_I),
.I4(CLBLM_R_X3Y111_SLICE_X2Y111_BO6),
.I5(CLBLM_R_X3Y111_SLICE_X2Y111_CO6),
.O5(CLBLM_R_X3Y112_SLICE_X2Y112_BO5),
.O6(CLBLM_R_X3Y112_SLICE_X2Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hda705df7258fa208)
  ) CLBLM_R_X3Y112_SLICE_X2Y112_ALUT (
.I0(RIOB33_X105Y107_IOB_X1Y108_I),
.I1(LIOB33_X0Y113_IOB_X0Y113_I),
.I2(CLBLL_L_X4Y111_SLICE_X5Y111_DO6),
.I3(LIOB33_X0Y115_IOB_X0Y115_I),
.I4(CLBLM_R_X3Y111_SLICE_X2Y111_BO6),
.I5(CLBLM_R_X3Y111_SLICE_X2Y111_CO6),
.O5(CLBLM_R_X3Y112_SLICE_X2Y112_AO5),
.O6(CLBLM_R_X3Y112_SLICE_X2Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h9fc7bf973fbf3f3f)
  ) CLBLM_R_X3Y112_SLICE_X3Y112_DLUT (
.I0(RIOB33_X105Y109_IOB_X1Y110_I),
.I1(LIOB33_X0Y115_IOB_X0Y115_I),
.I2(RIOB33_X105Y111_IOB_X1Y111_I),
.I3(CLBLM_R_X3Y112_SLICE_X3Y112_CO6),
.I4(LIOB33_X0Y111_IOB_X0Y112_I),
.I5(LIOB33_X0Y113_IOB_X0Y113_I),
.O5(CLBLM_R_X3Y112_SLICE_X3Y112_DO5),
.O6(CLBLM_R_X3Y112_SLICE_X3Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f13ff7f7f1fffff)
  ) CLBLM_R_X3Y112_SLICE_X3Y112_CLUT (
.I0(LIOB33_X0Y109_IOB_X0Y110_I),
.I1(RIOB33_X105Y109_IOB_X1Y110_I),
.I2(RIOB33_X105Y111_IOB_X1Y111_I),
.I3(CLBLL_L_X4Y111_SLICE_X4Y111_DO6),
.I4(LIOB33_X0Y111_IOB_X0Y111_I),
.I5(LIOB33_X0Y111_IOB_X0Y112_I),
.O5(CLBLM_R_X3Y112_SLICE_X3Y112_CO5),
.O6(CLBLM_R_X3Y112_SLICE_X3Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h4dd4cffcdd44ffcc)
  ) CLBLM_R_X3Y112_SLICE_X3Y112_BLUT (
.I0(LIOB33_X0Y115_IOB_X0Y115_I),
.I1(CLBLM_R_X3Y111_SLICE_X2Y111_DO6),
.I2(LIOB33_X0Y113_IOB_X0Y113_I),
.I3(CLBLL_L_X4Y112_SLICE_X4Y112_CO6),
.I4(RIOB33_X105Y109_IOB_X1Y109_I),
.I5(RIOB33_X105Y109_IOB_X1Y110_I),
.O5(CLBLM_R_X3Y112_SLICE_X3Y112_BO5),
.O6(CLBLM_R_X3Y112_SLICE_X3Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h4114c33c14143c3c)
  ) CLBLM_R_X3Y112_SLICE_X3Y112_ALUT (
.I0(LIOB33_X0Y115_IOB_X0Y115_I),
.I1(CLBLM_R_X3Y111_SLICE_X2Y111_DO6),
.I2(CLBLL_L_X4Y112_SLICE_X4Y112_CO6),
.I3(LIOB33_X0Y113_IOB_X0Y113_I),
.I4(RIOB33_X105Y109_IOB_X1Y109_I),
.I5(RIOB33_X105Y109_IOB_X1Y110_I),
.O5(CLBLM_R_X3Y112_SLICE_X3Y112_AO5),
.O6(CLBLM_R_X3Y112_SLICE_X3Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y113_SLICE_X2Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y113_SLICE_X2Y113_DO5),
.O6(CLBLM_R_X3Y113_SLICE_X2Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y113_SLICE_X2Y113_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y113_SLICE_X2Y113_CO5),
.O6(CLBLM_R_X3Y113_SLICE_X2Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y113_SLICE_X2Y113_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y113_SLICE_X2Y113_BO5),
.O6(CLBLM_R_X3Y113_SLICE_X2Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y113_SLICE_X2Y113_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y113_SLICE_X2Y113_AO5),
.O6(CLBLM_R_X3Y113_SLICE_X2Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0dcf4fffdfffdfff)
  ) CLBLM_R_X3Y113_SLICE_X3Y113_DLUT (
.I0(LIOB33_X0Y115_IOB_X0Y115_I),
.I1(CLBLM_R_X3Y112_SLICE_X3Y112_CO6),
.I2(LIOB33_X0Y113_IOB_X0Y113_I),
.I3(RIOB33_X105Y109_IOB_X1Y110_I),
.I4(LIOB33_X0Y111_IOB_X0Y112_I),
.I5(RIOB33_X105Y111_IOB_X1Y111_I),
.O5(CLBLM_R_X3Y113_SLICE_X3Y113_DO5),
.O6(CLBLM_R_X3Y113_SLICE_X3Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h20a0b3ff0020a0b3)
  ) CLBLM_R_X3Y113_SLICE_X3Y113_CLUT (
.I0(RIOB33_X105Y111_IOB_X1Y111_I),
.I1(CLBLL_L_X4Y113_SLICE_X4Y113_CO6),
.I2(LIOB33_X0Y115_IOB_X0Y115_I),
.I3(CLBLM_R_X3Y112_SLICE_X3Y112_BO6),
.I4(CLBLM_R_X3Y113_SLICE_X3Y113_DO6),
.I5(CLBLM_R_X3Y113_SLICE_X3Y113_BO6),
.O5(CLBLM_R_X3Y113_SLICE_X3Y113_CO5),
.O6(CLBLM_R_X3Y113_SLICE_X3Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hbccc7000d60c1ac0)
  ) CLBLM_R_X3Y113_SLICE_X3Y113_BLUT (
.I0(LIOB33_X0Y111_IOB_X0Y112_I),
.I1(RIOB33_X105Y109_IOB_X1Y110_I),
.I2(LIOB33_X0Y113_IOB_X0Y113_I),
.I3(RIOB33_X105Y111_IOB_X1Y111_I),
.I4(LIOB33_X0Y115_IOB_X0Y115_I),
.I5(CLBLM_R_X3Y112_SLICE_X3Y112_CO6),
.O5(CLBLM_R_X3Y113_SLICE_X3Y113_BO5),
.O6(CLBLM_R_X3Y113_SLICE_X3Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc33cc33c6a566a56)
  ) CLBLM_R_X3Y113_SLICE_X3Y113_ALUT (
.I0(CLBLM_R_X3Y112_SLICE_X3Y112_DO6),
.I1(CLBLL_L_X4Y113_SLICE_X4Y113_CO6),
.I2(CLBLM_R_X3Y112_SLICE_X3Y112_BO6),
.I3(CLBLM_R_X3Y113_SLICE_X3Y113_BO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y113_SLICE_X3Y113_AO5),
.O6(CLBLM_R_X3Y113_SLICE_X3Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y114_SLICE_X2Y114_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y114_SLICE_X2Y114_DO5),
.O6(CLBLM_R_X3Y114_SLICE_X2Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y114_SLICE_X2Y114_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y114_SLICE_X2Y114_CO5),
.O6(CLBLM_R_X3Y114_SLICE_X2Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y114_SLICE_X2Y114_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y114_SLICE_X2Y114_BO5),
.O6(CLBLM_R_X3Y114_SLICE_X2Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y114_SLICE_X2Y114_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y114_SLICE_X2Y114_AO5),
.O6(CLBLM_R_X3Y114_SLICE_X2Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y114_SLICE_X3Y114_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y114_SLICE_X3Y114_DO5),
.O6(CLBLM_R_X3Y114_SLICE_X3Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y114_SLICE_X3Y114_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y114_SLICE_X3Y114_CO5),
.O6(CLBLM_R_X3Y114_SLICE_X3Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y114_SLICE_X3Y114_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y114_SLICE_X3Y114_BO5),
.O6(CLBLM_R_X3Y114_SLICE_X3Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h99559955f00f0f0f)
  ) CLBLM_R_X3Y114_SLICE_X3Y114_ALUT (
.I0(CLBLM_R_X7Y113_SLICE_X9Y113_BO6),
.I1(LIOB33_X0Y113_IOB_X0Y114_I),
.I2(CLBLM_R_X3Y111_SLICE_X3Y111_BO6),
.I3(LIOB33_X0Y113_IOB_X0Y113_I),
.I4(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y114_SLICE_X3Y114_AO5),
.O6(CLBLM_R_X3Y114_SLICE_X3Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y104_SLICE_X6Y104_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y104_SLICE_X6Y104_DO5),
.O6(CLBLM_R_X5Y104_SLICE_X6Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y104_SLICE_X6Y104_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y104_SLICE_X6Y104_CO5),
.O6(CLBLM_R_X5Y104_SLICE_X6Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y104_SLICE_X6Y104_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y104_SLICE_X6Y104_BO5),
.O6(CLBLM_R_X5Y104_SLICE_X6Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h503a5ac0303a9ac0)
  ) CLBLM_R_X5Y104_SLICE_X6Y104_ALUT (
.I0(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I1(RIOB33_X105Y101_IOB_X1Y101_I),
.I2(RIOB33_X105Y113_IOB_X1Y113_I),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(LIOB33_X0Y115_IOB_X0Y116_I),
.I5(RIOB33_X105Y111_IOB_X1Y112_I),
.O5(CLBLM_R_X5Y104_SLICE_X6Y104_AO5),
.O6(CLBLM_R_X5Y104_SLICE_X6Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y104_SLICE_X7Y104_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y104_SLICE_X7Y104_DO5),
.O6(CLBLM_R_X5Y104_SLICE_X7Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y104_SLICE_X7Y104_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y104_SLICE_X7Y104_CO5),
.O6(CLBLM_R_X5Y104_SLICE_X7Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y104_SLICE_X7Y104_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y104_SLICE_X7Y104_BO5),
.O6(CLBLM_R_X5Y104_SLICE_X7Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y104_SLICE_X7Y104_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y104_SLICE_X7Y104_AO5),
.O6(CLBLM_R_X5Y104_SLICE_X7Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y105_SLICE_X6Y105_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y105_SLICE_X6Y105_DO5),
.O6(CLBLM_R_X5Y105_SLICE_X6Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y105_SLICE_X6Y105_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y105_SLICE_X6Y105_CO5),
.O6(CLBLM_R_X5Y105_SLICE_X6Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y105_SLICE_X6Y105_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y105_SLICE_X6Y105_BO5),
.O6(CLBLM_R_X5Y105_SLICE_X6Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h7ff7f7f707707070)
  ) CLBLM_R_X5Y105_SLICE_X6Y105_ALUT (
.I0(LIOB33_X0Y115_IOB_X0Y116_I),
.I1(LIOB33_X0Y103_IOB_X0Y104_I),
.I2(CLBLM_R_X5Y105_SLICE_X7Y105_CO6),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(LIOB33_X0Y101_IOB_X0Y102_I),
.I5(CLBLL_L_X4Y105_SLICE_X4Y105_DO6),
.O5(CLBLM_R_X5Y105_SLICE_X6Y105_AO5),
.O6(CLBLM_R_X5Y105_SLICE_X6Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y105_SLICE_X7Y105_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y105_SLICE_X7Y105_DO5),
.O6(CLBLM_R_X5Y105_SLICE_X7Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h54abab54bb44bb44)
  ) CLBLM_R_X5Y105_SLICE_X7Y105_CLUT (
.I0(CLBLM_R_X5Y105_SLICE_X7Y105_AO6),
.I1(CLBLM_R_X7Y106_SLICE_X8Y106_CO6),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(CLBLM_R_X7Y104_SLICE_X8Y104_AO6),
.I4(RIOB33_X105Y101_IOB_X1Y101_I),
.I5(LIOB33_X0Y101_IOB_X0Y101_I),
.O5(CLBLM_R_X5Y105_SLICE_X7Y105_CO5),
.O6(CLBLM_R_X5Y105_SLICE_X7Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6ac0953f953f6ac0)
  ) CLBLM_R_X5Y105_SLICE_X7Y105_BLUT (
.I0(LIOB33_X0Y103_IOB_X0Y104_I),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(LIOB33_X0Y101_IOB_X0Y102_I),
.I3(LIOB33_X0Y115_IOB_X0Y116_I),
.I4(CLBLM_R_X5Y105_SLICE_X7Y105_CO6),
.I5(CLBLL_L_X4Y105_SLICE_X4Y105_DO6),
.O5(CLBLM_R_X5Y105_SLICE_X7Y105_BO5),
.O6(CLBLM_R_X5Y105_SLICE_X7Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5350202023502020)
  ) CLBLM_R_X5Y105_SLICE_X7Y105_ALUT (
.I0(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(RIOB33_X105Y101_IOB_X1Y101_I),
.I3(RIOB33_X105Y101_IOB_X1Y102_I),
.I4(RIOB33_X105Y113_IOB_X1Y113_I),
.I5(RIOB33_X105Y111_IOB_X1Y112_I),
.O5(CLBLM_R_X5Y105_SLICE_X7Y105_AO5),
.O6(CLBLM_R_X5Y105_SLICE_X7Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hc6936c936cc66c6c)
  ) CLBLM_R_X5Y106_SLICE_X6Y106_DLUT (
.I0(LIOB33_X0Y101_IOB_X0Y102_I),
.I1(CLBLM_R_X5Y105_SLICE_X7Y105_CO6),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(CLBLM_R_X5Y106_SLICE_X6Y106_AO5),
.I4(LIOB33_X0Y115_IOB_X0Y116_I),
.I5(CLBLM_R_X7Y106_SLICE_X8Y106_BO6),
.O5(CLBLM_R_X5Y106_SLICE_X6Y106_DO5),
.O6(CLBLM_R_X5Y106_SLICE_X6Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h1d5140400c0c4040)
  ) CLBLM_R_X5Y106_SLICE_X6Y106_CLUT (
.I0(LIOB33_X0Y115_IOB_X0Y116_I),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I3(RIOB33_X105Y111_IOB_X1Y112_I),
.I4(RIOB33_X105Y113_IOB_X1Y113_I),
.I5(RIOB33_X105Y101_IOB_X1Y101_I),
.O5(CLBLM_R_X5Y106_SLICE_X6Y106_CO5),
.O6(CLBLM_R_X5Y106_SLICE_X6Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h33ff33ff77777777)
  ) CLBLM_R_X5Y106_SLICE_X6Y106_BLUT (
.I0(LIOB33_X0Y113_IOB_X0Y114_I),
.I1(LIOB33_X0Y105_IOB_X0Y105_I),
.I2(1'b1),
.I3(LIOB33_X0Y103_IOB_X0Y103_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y106_SLICE_X6Y106_BO5),
.O6(CLBLM_R_X5Y106_SLICE_X6Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc30fc30fffff030f)
  ) CLBLM_R_X5Y106_SLICE_X6Y106_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y101_IOB_X0Y101_I),
.I2(CLBLM_R_X5Y104_SLICE_X6Y104_AO6),
.I3(LIOB33_X0Y115_IOB_X0Y116_I),
.I4(CLBLM_R_X5Y106_SLICE_X6Y106_CO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y106_SLICE_X6Y106_AO5),
.O6(CLBLM_R_X5Y106_SLICE_X6Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdc4dc40f7317310)
  ) CLBLM_R_X5Y106_SLICE_X7Y106_DLUT (
.I0(CLBLM_R_X5Y105_SLICE_X7Y105_BO6),
.I1(CLBLM_R_X7Y105_SLICE_X8Y105_CO6),
.I2(CLBLM_R_X5Y106_SLICE_X6Y106_BO5),
.I3(CLBLM_R_X5Y106_SLICE_X7Y106_AO5),
.I4(CLBLL_L_X4Y106_SLICE_X5Y106_CO6),
.I5(CLBLM_R_X7Y108_SLICE_X9Y108_AO5),
.O5(CLBLM_R_X5Y106_SLICE_X7Y106_DO5),
.O6(CLBLM_R_X5Y106_SLICE_X7Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h39c69c63c639639c)
  ) CLBLM_R_X5Y106_SLICE_X7Y106_CLUT (
.I0(CLBLM_R_X5Y105_SLICE_X7Y105_BO6),
.I1(CLBLM_R_X7Y105_SLICE_X8Y105_CO6),
.I2(CLBLM_R_X5Y106_SLICE_X6Y106_BO5),
.I3(CLBLM_R_X5Y106_SLICE_X7Y106_AO5),
.I4(CLBLL_L_X4Y106_SLICE_X5Y106_CO6),
.I5(CLBLM_R_X7Y108_SLICE_X9Y108_AO5),
.O5(CLBLM_R_X5Y106_SLICE_X7Y106_CO5),
.O6(CLBLM_R_X5Y106_SLICE_X7Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h96669996cccc3c3c)
  ) CLBLM_R_X5Y106_SLICE_X7Y106_BLUT (
.I0(LIOB33_X0Y115_IOB_X0Y116_I),
.I1(CLBLM_R_X7Y105_SLICE_X8Y105_CO6),
.I2(CLBLM_R_X5Y105_SLICE_X7Y105_BO6),
.I3(LIOB33_X0Y113_IOB_X0Y114_I),
.I4(CLBLL_L_X4Y106_SLICE_X5Y106_CO6),
.I5(LIOB33_X0Y105_IOB_X0Y105_I),
.O5(CLBLM_R_X5Y106_SLICE_X7Y106_BO5),
.O6(CLBLM_R_X5Y106_SLICE_X7Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5f5f5f5f55ff55ff)
  ) CLBLM_R_X5Y106_SLICE_X7Y106_ALUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(1'b1),
.I2(LIOB33_X0Y115_IOB_X0Y116_I),
.I3(LIOB33_X0Y113_IOB_X0Y114_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y106_SLICE_X7Y106_AO5),
.O6(CLBLM_R_X5Y106_SLICE_X7Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h60f6a0faf6f6fafa)
  ) CLBLM_R_X5Y107_SLICE_X6Y107_DLUT (
.I0(CLBLM_R_X5Y106_SLICE_X6Y106_DO6),
.I1(LIOB33_X0Y103_IOB_X0Y104_I),
.I2(CLBLL_L_X4Y106_SLICE_X5Y106_CO6),
.I3(LIOB33_X0Y113_IOB_X0Y114_I),
.I4(LIOB33_X0Y115_IOB_X0Y116_I),
.I5(LIOB33_X0Y105_IOB_X0Y105_I),
.O5(CLBLM_R_X5Y107_SLICE_X6Y107_DO5),
.O6(CLBLM_R_X5Y107_SLICE_X6Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h69a5965a965a965a)
  ) CLBLM_R_X5Y107_SLICE_X6Y107_CLUT (
.I0(CLBLM_R_X5Y105_SLICE_X6Y105_AO6),
.I1(LIOB33_X0Y103_IOB_X0Y104_I),
.I2(CLBLM_R_X7Y106_SLICE_X9Y106_DO6),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(LIOB33_X0Y115_IOB_X0Y116_I),
.I5(LIOB33_X0Y105_IOB_X0Y105_I),
.O5(CLBLM_R_X5Y107_SLICE_X6Y107_CO5),
.O6(CLBLM_R_X5Y107_SLICE_X6Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'he21d6a957b843fc0)
  ) CLBLM_R_X5Y107_SLICE_X6Y107_BLUT (
.I0(CLBLM_R_X5Y107_SLICE_X6Y107_DO6),
.I1(LIOB33_X0Y105_IOB_X0Y106_I),
.I2(LIOB33_X0Y115_IOB_X0Y116_I),
.I3(CLBLM_R_X7Y107_SLICE_X9Y107_CO6),
.I4(LIOB33_X0Y113_IOB_X0Y114_I),
.I5(CLBLM_R_X5Y107_SLICE_X6Y107_CO6),
.O5(CLBLM_R_X5Y107_SLICE_X6Y107_BO5),
.O6(CLBLM_R_X5Y107_SLICE_X6Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6a95956a95956a6a)
  ) CLBLM_R_X5Y107_SLICE_X6Y107_ALUT (
.I0(CLBLL_L_X4Y106_SLICE_X5Y106_CO6),
.I1(LIOB33_X0Y115_IOB_X0Y116_I),
.I2(LIOB33_X0Y103_IOB_X0Y104_I),
.I3(LIOB33_X0Y105_IOB_X0Y105_I),
.I4(CLBLM_R_X5Y106_SLICE_X6Y106_DO6),
.I5(LIOB33_X0Y113_IOB_X0Y114_I),
.O5(CLBLM_R_X5Y107_SLICE_X6Y107_AO5),
.O6(CLBLM_R_X5Y107_SLICE_X6Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y107_SLICE_X7Y107_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y107_SLICE_X7Y107_DO5),
.O6(CLBLM_R_X5Y107_SLICE_X7Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y107_SLICE_X7Y107_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y107_SLICE_X7Y107_CO5),
.O6(CLBLM_R_X5Y107_SLICE_X7Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996969699666666)
  ) CLBLM_R_X5Y107_SLICE_X7Y107_BLUT (
.I0(CLBLM_R_X7Y107_SLICE_X9Y107_CO6),
.I1(CLBLM_R_X5Y106_SLICE_X7Y106_DO6),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(LIOB33_X0Y115_IOB_X0Y116_I),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(LIOB33_X0Y113_IOB_X0Y114_I),
.O5(CLBLM_R_X5Y107_SLICE_X7Y107_BO5),
.O6(CLBLM_R_X5Y107_SLICE_X7Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996996666996996)
  ) CLBLM_R_X5Y107_SLICE_X7Y107_ALUT (
.I0(CLBLM_R_X5Y106_SLICE_X7Y106_DO6),
.I1(CLBLM_R_X7Y108_SLICE_X8Y108_AO6),
.I2(CLBLM_R_X3Y107_SLICE_X2Y107_AO5),
.I3(CLBLM_R_X7Y107_SLICE_X9Y107_AO6),
.I4(CLBLL_L_X4Y106_SLICE_X5Y106_DO6),
.I5(CLBLM_R_X5Y106_SLICE_X7Y106_CO6),
.O5(CLBLM_R_X5Y107_SLICE_X7Y107_AO5),
.O6(CLBLM_R_X5Y107_SLICE_X7Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h4ddf5dff4fffdfff)
  ) CLBLM_R_X5Y108_SLICE_X6Y108_DLUT (
.I0(RIOB33_X105Y109_IOB_X1Y110_I),
.I1(CLBLM_L_X8Y105_SLICE_X10Y105_DO6),
.I2(RIOB33_X105Y111_IOB_X1Y111_I),
.I3(LIOB33_X0Y105_IOB_X0Y105_I),
.I4(LIOB33_X0Y103_IOB_X0Y104_I),
.I5(LIOB33_X0Y105_IOB_X0Y106_I),
.O5(CLBLM_R_X5Y108_SLICE_X6Y108_DO5),
.O6(CLBLM_R_X5Y108_SLICE_X6Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h4d8e8e8eddeeeeee)
  ) CLBLM_R_X5Y108_SLICE_X6Y108_CLUT (
.I0(CLBLM_R_X5Y107_SLICE_X6Y107_BO6),
.I1(CLBLM_R_X5Y108_SLICE_X6Y108_AO6),
.I2(LIOB33_X0Y107_IOB_X0Y108_I),
.I3(LIOB33_X0Y107_IOB_X0Y107_I),
.I4(LIOB33_X0Y113_IOB_X0Y114_I),
.I5(LIOB33_X0Y103_IOB_X0Y103_I),
.O5(CLBLM_R_X5Y108_SLICE_X6Y108_CO5),
.O6(CLBLM_R_X5Y108_SLICE_X6Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6c93936ca05f5fa0)
  ) CLBLM_R_X5Y108_SLICE_X6Y108_BLUT (
.I0(LIOB33_X0Y113_IOB_X0Y114_I),
.I1(LIOB33_X0Y103_IOB_X0Y103_I),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(CLBLM_R_X5Y108_SLICE_X6Y108_AO6),
.I4(CLBLM_R_X5Y107_SLICE_X6Y107_BO6),
.I5(LIOB33_X0Y107_IOB_X0Y108_I),
.O5(CLBLM_R_X5Y108_SLICE_X6Y108_BO5),
.O6(CLBLM_R_X5Y108_SLICE_X6Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h7080f7f8f7f8f7f8)
  ) CLBLM_R_X5Y108_SLICE_X6Y108_ALUT (
.I0(LIOB33_X0Y113_IOB_X0Y114_I),
.I1(LIOB33_X0Y105_IOB_X0Y106_I),
.I2(CLBLL_L_X4Y106_SLICE_X5Y106_DO6),
.I3(CLBLM_R_X5Y106_SLICE_X7Y106_BO6),
.I4(LIOB33_X0Y107_IOB_X0Y107_I),
.I5(LIOB33_X0Y103_IOB_X0Y103_I),
.O5(CLBLM_R_X5Y108_SLICE_X6Y108_AO5),
.O6(CLBLM_R_X5Y108_SLICE_X6Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8fe78f877f3fff7f)
  ) CLBLM_R_X5Y108_SLICE_X7Y108_DLUT (
.I0(RIOB33_X105Y109_IOB_X1Y110_I),
.I1(LIOB33_X0Y105_IOB_X0Y105_I),
.I2(RIOB33_X105Y111_IOB_X1Y111_I),
.I3(CLBLM_L_X8Y105_SLICE_X10Y105_DO6),
.I4(LIOB33_X0Y103_IOB_X0Y104_I),
.I5(LIOB33_X0Y105_IOB_X0Y106_I),
.O5(CLBLM_R_X5Y108_SLICE_X7Y108_DO5),
.O6(CLBLM_R_X5Y108_SLICE_X7Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h87f0e15a78f01e5a)
  ) CLBLM_R_X5Y108_SLICE_X7Y108_CLUT (
.I0(CLBLM_R_X5Y109_SLICE_X7Y109_AO6),
.I1(LIOB33_X0Y107_IOB_X0Y108_I),
.I2(CLBLL_L_X4Y108_SLICE_X5Y108_CO6),
.I3(RIOB33_X105Y109_IOB_X1Y109_I),
.I4(CLBLM_L_X8Y106_SLICE_X10Y106_CO6),
.I5(LIOB33_X0Y109_IOB_X0Y109_I),
.O5(CLBLM_R_X5Y108_SLICE_X7Y108_CO5),
.O6(CLBLM_R_X5Y108_SLICE_X7Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h69999666a5555aaa)
  ) CLBLM_R_X5Y108_SLICE_X7Y108_BLUT (
.I0(CLBLM_R_X5Y108_SLICE_X7Y108_DO6),
.I1(LIOB33_X0Y107_IOB_X0Y108_I),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(RIOB33_X105Y109_IOB_X1Y110_I),
.I4(CLBLM_L_X8Y106_SLICE_X10Y106_CO6),
.I5(RIOB33_X105Y109_IOB_X1Y109_I),
.O5(CLBLM_R_X5Y108_SLICE_X7Y108_BO5),
.O6(CLBLM_R_X5Y108_SLICE_X7Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h137f0137ffff0fff)
  ) CLBLM_R_X5Y108_SLICE_X7Y108_ALUT (
.I0(LIOB33_X0Y107_IOB_X0Y108_I),
.I1(LIOB33_X0Y109_IOB_X0Y109_I),
.I2(CLBLM_R_X5Y109_SLICE_X7Y109_AO6),
.I3(CLBLL_L_X4Y108_SLICE_X5Y108_CO6),
.I4(CLBLM_L_X8Y106_SLICE_X10Y106_CO6),
.I5(RIOB33_X105Y109_IOB_X1Y109_I),
.O5(CLBLM_R_X5Y108_SLICE_X7Y108_AO5),
.O6(CLBLM_R_X5Y108_SLICE_X7Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'he88ea00afaafe88e)
  ) CLBLM_R_X5Y109_SLICE_X6Y109_DLUT (
.I0(CLBLM_R_X5Y109_SLICE_X6Y109_AO6),
.I1(CLBLL_L_X4Y110_SLICE_X4Y110_AO6),
.I2(CLBLM_R_X7Y108_SLICE_X8Y108_BO6),
.I3(CLBLM_R_X7Y109_SLICE_X8Y109_AO6),
.I4(CLBLM_R_X5Y108_SLICE_X6Y108_AO6),
.I5(CLBLM_R_X5Y107_SLICE_X7Y107_BO6),
.O5(CLBLM_R_X5Y109_SLICE_X6Y109_DO5),
.O6(CLBLM_R_X5Y109_SLICE_X6Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996969669696996)
  ) CLBLM_R_X5Y109_SLICE_X6Y109_CLUT (
.I0(CLBLM_R_X5Y109_SLICE_X6Y109_AO6),
.I1(CLBLM_R_X7Y109_SLICE_X8Y109_AO6),
.I2(CLBLM_R_X7Y108_SLICE_X8Y108_BO6),
.I3(CLBLL_L_X4Y110_SLICE_X4Y110_AO6),
.I4(CLBLM_R_X5Y108_SLICE_X6Y108_AO6),
.I5(CLBLM_R_X5Y107_SLICE_X7Y107_BO6),
.O5(CLBLM_R_X5Y109_SLICE_X6Y109_CO5),
.O6(CLBLM_R_X5Y109_SLICE_X6Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hd25ab49678f01e3c)
  ) CLBLM_R_X5Y109_SLICE_X6Y109_BLUT (
.I0(LIOB33_X0Y107_IOB_X0Y108_I),
.I1(CLBLM_R_X5Y107_SLICE_X7Y107_BO6),
.I2(CLBLM_R_X7Y108_SLICE_X8Y108_BO6),
.I3(LIOB33_X0Y103_IOB_X0Y103_I),
.I4(CLBLM_R_X5Y108_SLICE_X6Y108_AO6),
.I5(LIOB33_X0Y113_IOB_X0Y114_I),
.O5(CLBLM_R_X5Y109_SLICE_X6Y109_BO5),
.O6(CLBLM_R_X5Y109_SLICE_X6Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h7777777755ff55ff)
  ) CLBLM_R_X5Y109_SLICE_X6Y109_ALUT (
.I0(LIOB33_X0Y109_IOB_X0Y109_I),
.I1(LIOB33_X0Y103_IOB_X0Y103_I),
.I2(1'b1),
.I3(LIOB33_X0Y113_IOB_X0Y114_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y109_SLICE_X6Y109_AO5),
.O6(CLBLM_R_X5Y109_SLICE_X6Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h9aa565a559aaa6aa)
  ) CLBLM_R_X5Y109_SLICE_X7Y109_DLUT (
.I0(CLBLM_R_X5Y108_SLICE_X7Y108_CO6),
.I1(LIOB33_X0Y109_IOB_X0Y109_I),
.I2(CLBLM_L_X8Y109_SLICE_X10Y109_AO6),
.I3(RIOB33_X105Y107_IOB_X1Y108_I),
.I4(LIOB33_X0Y109_IOB_X0Y110_I),
.I5(CLBLM_R_X5Y108_SLICE_X7Y108_BO6),
.O5(CLBLM_R_X5Y109_SLICE_X7Y109_DO5),
.O6(CLBLM_R_X5Y109_SLICE_X7Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h1171f5f57177ffff)
  ) CLBLM_R_X5Y109_SLICE_X7Y109_CLUT (
.I0(CLBLM_R_X5Y108_SLICE_X7Y108_CO6),
.I1(LIOB33_X0Y109_IOB_X0Y110_I),
.I2(CLBLM_L_X8Y109_SLICE_X10Y109_AO6),
.I3(LIOB33_X0Y109_IOB_X0Y109_I),
.I4(RIOB33_X105Y107_IOB_X1Y108_I),
.I5(CLBLM_R_X5Y108_SLICE_X7Y108_BO6),
.O5(CLBLM_R_X5Y109_SLICE_X7Y109_CO5),
.O6(CLBLM_R_X5Y109_SLICE_X7Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h9c3c6cccc6963666)
  ) CLBLM_R_X5Y109_SLICE_X7Y109_BLUT (
.I0(CLBLM_R_X7Y109_SLICE_X9Y109_CO6),
.I1(CLBLM_R_X7Y109_SLICE_X8Y109_BO6),
.I2(LIOB33_X0Y109_IOB_X0Y109_I),
.I3(LIOB33_X0Y103_IOB_X0Y103_I),
.I4(LIOB33_X0Y113_IOB_X0Y114_I),
.I5(CLBLM_R_X5Y108_SLICE_X6Y108_CO6),
.O5(CLBLM_R_X5Y109_SLICE_X7Y109_BO5),
.O6(CLBLM_R_X5Y109_SLICE_X7Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha555a555c0c03f3f)
  ) CLBLM_R_X5Y109_SLICE_X7Y109_ALUT (
.I0(CLBLM_R_X5Y108_SLICE_X7Y108_DO6),
.I1(LIOB33_X0Y109_IOB_X0Y109_I),
.I2(RIOB33_X105Y109_IOB_X1Y110_I),
.I3(LIOB33_X0Y107_IOB_X0Y107_I),
.I4(CLBLM_R_X5Y110_SLICE_X6Y110_CO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y109_SLICE_X7Y109_AO5),
.O6(CLBLM_R_X5Y109_SLICE_X7Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h4bb4d22db44b2dd2)
  ) CLBLM_R_X5Y110_SLICE_X6Y110_DLUT (
.I0(CLBLM_R_X3Y111_SLICE_X2Y111_AO6),
.I1(CLBLM_R_X5Y110_SLICE_X7Y110_CO6),
.I2(CLBLM_R_X5Y110_SLICE_X7Y110_AO6),
.I3(CLBLM_R_X5Y111_SLICE_X6Y111_AO6),
.I4(CLBLL_L_X4Y109_SLICE_X5Y109_BO6),
.I5(CLBLM_R_X7Y110_SLICE_X8Y110_AO6),
.O5(CLBLM_R_X5Y110_SLICE_X6Y110_DO5),
.O6(CLBLM_R_X5Y110_SLICE_X6Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha7e5ff5f0f87ffff)
  ) CLBLM_R_X5Y110_SLICE_X6Y110_CLUT (
.I0(LIOB33_X0Y107_IOB_X0Y107_I),
.I1(LIOB33_X0Y105_IOB_X0Y106_I),
.I2(LIOB33_X0Y107_IOB_X0Y108_I),
.I3(CLBLM_R_X5Y108_SLICE_X6Y108_DO6),
.I4(RIOB33_X105Y111_IOB_X1Y111_I),
.I5(RIOB33_X105Y109_IOB_X1Y110_I),
.O5(CLBLM_R_X5Y110_SLICE_X6Y110_CO5),
.O6(CLBLM_R_X5Y110_SLICE_X6Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6699966996699966)
  ) CLBLM_R_X5Y110_SLICE_X6Y110_BLUT (
.I0(CLBLM_R_X5Y109_SLICE_X6Y109_DO6),
.I1(CLBLM_R_X5Y110_SLICE_X7Y110_BO5),
.I2(CLBLM_R_X5Y109_SLICE_X6Y109_CO6),
.I3(CLBLM_R_X7Y109_SLICE_X8Y109_DO6),
.I4(CLBLL_L_X4Y109_SLICE_X4Y109_DO6),
.I5(CLBLM_R_X3Y110_SLICE_X3Y110_AO5),
.O5(CLBLM_R_X5Y110_SLICE_X6Y110_BO5),
.O6(CLBLM_R_X5Y110_SLICE_X6Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h7887878787787878)
  ) CLBLM_R_X5Y110_SLICE_X6Y110_ALUT (
.I0(LIOB33_X0Y109_IOB_X0Y110_I),
.I1(RIOB33_X105Y109_IOB_X1Y109_I),
.I2(CLBLM_R_X5Y108_SLICE_X7Y108_AO6),
.I3(RIOB33_X105Y109_IOB_X1Y110_I),
.I4(LIOB33_X0Y109_IOB_X0Y109_I),
.I5(CLBLM_R_X5Y110_SLICE_X6Y110_CO6),
.O5(CLBLM_R_X5Y110_SLICE_X6Y110_AO5),
.O6(CLBLM_R_X5Y110_SLICE_X6Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0701ff337f1fffff)
  ) CLBLM_R_X5Y110_SLICE_X7Y110_DLUT (
.I0(LIOB33_X0Y109_IOB_X0Y109_I),
.I1(CLBLM_R_X7Y109_SLICE_X9Y109_CO6),
.I2(LIOB33_X0Y109_IOB_X0Y110_I),
.I3(CLBLM_R_X5Y108_SLICE_X6Y108_CO6),
.I4(LIOB33_X0Y103_IOB_X0Y103_I),
.I5(CLBLM_R_X7Y109_SLICE_X8Y109_DO6),
.O5(CLBLM_R_X5Y110_SLICE_X7Y110_DO5),
.O6(CLBLM_R_X5Y110_SLICE_X7Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h87e1ff33781e00cc)
  ) CLBLM_R_X5Y110_SLICE_X7Y110_CLUT (
.I0(LIOB33_X0Y109_IOB_X0Y109_I),
.I1(CLBLM_R_X7Y109_SLICE_X9Y109_CO6),
.I2(LIOB33_X0Y109_IOB_X0Y110_I),
.I3(CLBLM_R_X5Y108_SLICE_X6Y108_CO6),
.I4(LIOB33_X0Y103_IOB_X0Y103_I),
.I5(CLBLM_R_X7Y109_SLICE_X8Y109_DO6),
.O5(CLBLM_R_X5Y110_SLICE_X7Y110_CO5),
.O6(CLBLM_R_X5Y110_SLICE_X7Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333ffff77777777)
  ) CLBLM_R_X5Y110_SLICE_X7Y110_BLUT (
.I0(LIOB33_X0Y103_IOB_X0Y103_I),
.I1(LIOB33_X0Y109_IOB_X0Y110_I),
.I2(1'b1),
.I3(1'b1),
.I4(RIOB33_X105Y107_IOB_X1Y107_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y110_SLICE_X7Y110_BO5),
.O6(CLBLM_R_X5Y110_SLICE_X7Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h777777773333ffff)
  ) CLBLM_R_X5Y110_SLICE_X7Y110_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y106_I),
.I1(LIOB33_X0Y111_IOB_X0Y112_I),
.I2(1'b1),
.I3(1'b1),
.I4(RIOB33_X105Y103_IOB_X1Y104_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y110_SLICE_X7Y110_AO5),
.O6(CLBLM_R_X5Y110_SLICE_X7Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h07017f1fff3fff3f)
  ) CLBLM_R_X5Y111_SLICE_X6Y111_DLUT (
.I0(LIOB33_X0Y111_IOB_X0Y112_I),
.I1(CLBLL_L_X4Y111_SLICE_X5Y111_BO6),
.I2(CLBLM_R_X5Y111_SLICE_X7Y111_BO6),
.I3(CLBLM_R_X5Y111_SLICE_X6Y111_CO6),
.I4(LIOB33_X0Y113_IOB_X0Y113_I),
.I5(RIOB33_X105Y105_IOB_X1Y106_I),
.O5(CLBLM_R_X5Y111_SLICE_X6Y111_DO5),
.O6(CLBLM_R_X5Y111_SLICE_X6Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h28bebebea0fafafa)
  ) CLBLM_R_X5Y111_SLICE_X6Y111_CLUT (
.I0(CLBLL_L_X4Y109_SLICE_X5Y109_BO6),
.I1(LIOB33_X0Y103_IOB_X0Y103_I),
.I2(CLBLM_R_X5Y109_SLICE_X7Y109_BO6),
.I3(RIOB33_X105Y105_IOB_X1Y106_I),
.I4(LIOB33_X0Y111_IOB_X0Y111_I),
.I5(LIOB33_X0Y109_IOB_X0Y110_I),
.O5(CLBLM_R_X5Y111_SLICE_X6Y111_CO5),
.O6(CLBLM_R_X5Y111_SLICE_X6Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hd27878788787d278)
  ) CLBLM_R_X5Y111_SLICE_X6Y111_BLUT (
.I0(LIOB33_X0Y111_IOB_X0Y112_I),
.I1(LIOB33_X0Y103_IOB_X0Y103_I),
.I2(CLBLM_R_X5Y111_SLICE_X7Y111_AO6),
.I3(RIOB33_X105Y105_IOB_X1Y106_I),
.I4(CLBLL_L_X4Y111_SLICE_X5Y111_BO6),
.I5(CLBLM_R_X5Y111_SLICE_X6Y111_CO6),
.O5(CLBLM_R_X5Y111_SLICE_X6Y111_BO5),
.O6(CLBLM_R_X5Y111_SLICE_X6Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h55ff55ff33ff33ff)
  ) CLBLM_R_X5Y111_SLICE_X6Y111_ALUT (
.I0(LIOB33_X0Y103_IOB_X0Y103_I),
.I1(LIOB33_X0Y113_IOB_X0Y114_I),
.I2(1'b1),
.I3(LIOB33_X0Y111_IOB_X0Y111_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y111_SLICE_X6Y111_AO5),
.O6(CLBLM_R_X5Y111_SLICE_X6Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h007171fff3fff3ff)
  ) CLBLM_R_X5Y111_SLICE_X7Y111_DLUT (
.I0(LIOB33_X0Y111_IOB_X0Y111_I),
.I1(CLBLM_R_X7Y110_SLICE_X9Y110_BO6),
.I2(CLBLM_L_X8Y111_SLICE_X10Y111_DO6),
.I3(CLBLL_L_X4Y110_SLICE_X4Y110_BO5),
.I4(LIOB33_X0Y111_IOB_X0Y112_I),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X5Y111_SLICE_X7Y111_DO5),
.O6(CLBLM_R_X5Y111_SLICE_X7Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8e71718ef3f30c0c)
  ) CLBLM_R_X5Y111_SLICE_X7Y111_CLUT (
.I0(LIOB33_X0Y111_IOB_X0Y111_I),
.I1(CLBLM_R_X7Y110_SLICE_X9Y110_BO6),
.I2(CLBLM_L_X8Y111_SLICE_X10Y111_DO6),
.I3(LIOB33_X0Y111_IOB_X0Y112_I),
.I4(CLBLL_L_X4Y110_SLICE_X4Y110_BO5),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X5Y111_SLICE_X7Y111_CO5),
.O6(CLBLM_R_X5Y111_SLICE_X7Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6a9556a9956aa956)
  ) CLBLM_R_X5Y111_SLICE_X7Y111_BLUT (
.I0(CLBLM_R_X5Y111_SLICE_X6Y111_AO5),
.I1(CLBLM_R_X5Y110_SLICE_X7Y110_DO6),
.I2(CLBLM_R_X5Y111_SLICE_X6Y111_AO6),
.I3(CLBLM_R_X5Y112_SLICE_X7Y112_AO5),
.I4(CLBLM_R_X7Y110_SLICE_X8Y110_CO6),
.I5(CLBLM_L_X8Y111_SLICE_X10Y111_CO6),
.O5(CLBLM_R_X5Y111_SLICE_X7Y111_BO5),
.O6(CLBLM_R_X5Y111_SLICE_X7Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6a9556a9956aa956)
  ) CLBLM_R_X5Y111_SLICE_X7Y111_ALUT (
.I0(CLBLM_R_X5Y111_SLICE_X6Y111_AO5),
.I1(CLBLM_R_X5Y110_SLICE_X7Y110_DO6),
.I2(CLBLM_R_X5Y111_SLICE_X6Y111_AO6),
.I3(CLBLM_R_X7Y110_SLICE_X8Y110_BO6),
.I4(CLBLM_R_X7Y110_SLICE_X8Y110_CO6),
.I5(CLBLM_L_X8Y113_SLICE_X10Y113_BO6),
.O5(CLBLM_R_X5Y111_SLICE_X7Y111_AO5),
.O6(CLBLM_R_X5Y111_SLICE_X7Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hb7d13f95482ec06a)
  ) CLBLM_R_X5Y112_SLICE_X6Y112_DLUT (
.I0(CLBLL_L_X4Y111_SLICE_X5Y111_BO6),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(LIOB33_X0Y113_IOB_X0Y113_I),
.I3(CLBLM_R_X5Y111_SLICE_X6Y111_CO6),
.I4(LIOB33_X0Y111_IOB_X0Y112_I),
.I5(CLBLM_R_X5Y111_SLICE_X7Y111_BO6),
.O5(CLBLM_R_X5Y112_SLICE_X6Y112_DO5),
.O6(CLBLM_R_X5Y112_SLICE_X6Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h956aa9566a9556a9)
  ) CLBLM_R_X5Y112_SLICE_X6Y112_CLUT (
.I0(CLBLM_R_X5Y112_SLICE_X6Y112_AO6),
.I1(CLBLL_L_X4Y113_SLICE_X5Y113_AO6),
.I2(CLBLM_R_X3Y111_SLICE_X3Y111_CO6),
.I3(CLBLM_R_X5Y111_SLICE_X6Y111_DO6),
.I4(CLBLM_R_X5Y112_SLICE_X6Y112_DO6),
.I5(CLBLM_R_X5Y112_SLICE_X6Y112_BO6),
.O5(CLBLM_R_X5Y112_SLICE_X6Y112_CO5),
.O6(CLBLM_R_X5Y112_SLICE_X6Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h965af0f0a5960ff0)
  ) CLBLM_R_X5Y112_SLICE_X6Y112_BLUT (
.I0(LIOB33_X0Y113_IOB_X0Y113_I),
.I1(LIOB33_X0Y111_IOB_X0Y112_I),
.I2(CLBLM_R_X7Y112_SLICE_X8Y112_AO6),
.I3(CLBLM_R_X7Y112_SLICE_X8Y112_BO6),
.I4(LIOB33_X0Y103_IOB_X0Y103_I),
.I5(CLBLL_L_X4Y111_SLICE_X5Y111_CO6),
.O5(CLBLM_R_X5Y112_SLICE_X6Y112_BO5),
.O6(CLBLM_R_X5Y112_SLICE_X6Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h55ff55ff0fff0fff)
  ) CLBLM_R_X5Y112_SLICE_X6Y112_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y106_I),
.I1(1'b1),
.I2(LIOB33_X0Y103_IOB_X0Y103_I),
.I3(LIOB33_X0Y115_IOB_X0Y115_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y112_SLICE_X6Y112_AO5),
.O6(CLBLM_R_X5Y112_SLICE_X6Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y112_SLICE_X7Y112_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y112_SLICE_X7Y112_DO5),
.O6(CLBLM_R_X5Y112_SLICE_X7Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y112_SLICE_X7Y112_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y112_SLICE_X7Y112_CO5),
.O6(CLBLM_R_X5Y112_SLICE_X7Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y112_SLICE_X7Y112_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y112_SLICE_X7Y112_BO5),
.O6(CLBLM_R_X5Y112_SLICE_X7Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h33ff33ff00ffffff)
  ) CLBLM_R_X5Y112_SLICE_X7Y112_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y113_IOB_X0Y114_I),
.I2(1'b1),
.I3(LIOB33_X0Y111_IOB_X0Y112_I),
.I4(LIOB33_X0Y103_IOB_X0Y103_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y112_SLICE_X7Y112_AO5),
.O6(CLBLM_R_X5Y112_SLICE_X7Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fd5ffff15403fc0)
  ) CLBLM_R_X5Y113_SLICE_X6Y113_DLUT (
.I0(LIOB33_X0Y103_IOB_X0Y103_I),
.I1(LIOB33_X0Y113_IOB_X0Y114_I),
.I2(LIOB33_X0Y113_IOB_X0Y113_I),
.I3(CLBLM_R_X7Y113_SLICE_X9Y113_BO6),
.I4(LIOB33_X0Y115_IOB_X0Y115_I),
.I5(CLBLM_R_X5Y113_SLICE_X6Y113_BO6),
.O5(CLBLM_R_X5Y113_SLICE_X6Y113_DO5),
.O6(CLBLM_R_X5Y113_SLICE_X6Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hb42dd2d24bd2d2d2)
  ) CLBLM_R_X5Y113_SLICE_X6Y113_CLUT (
.I0(CLBLM_R_X7Y112_SLICE_X8Y112_BO6),
.I1(CLBLL_L_X4Y111_SLICE_X5Y111_CO6),
.I2(CLBLM_R_X7Y113_SLICE_X8Y113_AO6),
.I3(LIOB33_X0Y103_IOB_X0Y103_I),
.I4(LIOB33_X0Y111_IOB_X0Y112_I),
.I5(LIOB33_X0Y113_IOB_X0Y114_I),
.O5(CLBLM_R_X5Y113_SLICE_X6Y113_CO5),
.O6(CLBLM_R_X5Y113_SLICE_X6Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h15ff7fff010f57ff)
  ) CLBLM_R_X5Y113_SLICE_X6Y113_BLUT (
.I0(LIOB33_X0Y113_IOB_X0Y113_I),
.I1(LIOB33_X0Y111_IOB_X0Y112_I),
.I2(CLBLM_R_X7Y112_SLICE_X8Y112_BO6),
.I3(LIOB33_X0Y103_IOB_X0Y103_I),
.I4(CLBLM_R_X7Y112_SLICE_X8Y112_AO6),
.I5(CLBLL_L_X4Y111_SLICE_X5Y111_CO6),
.O5(CLBLM_R_X5Y113_SLICE_X6Y113_BO5),
.O6(CLBLM_R_X5Y113_SLICE_X6Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h7f13ff5fdf4c5f00)
  ) CLBLM_R_X5Y113_SLICE_X6Y113_ALUT (
.I0(LIOB33_X0Y115_IOB_X0Y115_I),
.I1(LIOB33_X0Y103_IOB_X0Y103_I),
.I2(RIOB33_X105Y105_IOB_X1Y106_I),
.I3(CLBLM_R_X5Y111_SLICE_X6Y111_DO6),
.I4(LIOB33_X0Y113_IOB_X0Y113_I),
.I5(CLBLM_R_X5Y113_SLICE_X6Y113_CO6),
.O5(CLBLM_R_X5Y113_SLICE_X6Y113_AO5),
.O6(CLBLM_R_X5Y113_SLICE_X6Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y113_SLICE_X7Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y113_SLICE_X7Y113_DO5),
.O6(CLBLM_R_X5Y113_SLICE_X7Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y113_SLICE_X7Y113_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y113_SLICE_X7Y113_CO5),
.O6(CLBLM_R_X5Y113_SLICE_X7Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y113_SLICE_X7Y113_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y113_SLICE_X7Y113_BO5),
.O6(CLBLM_R_X5Y113_SLICE_X7Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y113_SLICE_X7Y113_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y113_SLICE_X7Y113_AO5),
.O6(CLBLM_R_X5Y113_SLICE_X7Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffd0fffdff40fff4)
  ) CLBLM_R_X5Y114_SLICE_X6Y114_DLUT (
.I0(CLBLM_R_X5Y113_SLICE_X6Y113_AO6),
.I1(CLBLM_R_X5Y112_SLICE_X6Y112_CO6),
.I2(CLBLM_R_X5Y115_SLICE_X6Y115_BO6),
.I3(CLBLM_R_X5Y116_SLICE_X6Y116_CO6),
.I4(CLBLM_R_X5Y113_SLICE_X6Y113_DO6),
.I5(CLBLM_R_X5Y114_SLICE_X6Y114_BO6),
.O5(CLBLM_R_X5Y114_SLICE_X6Y114_DO5),
.O6(CLBLM_R_X5Y114_SLICE_X6Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h2f0bbf2f0b022f0b)
  ) CLBLM_R_X5Y114_SLICE_X6Y114_CLUT (
.I0(CLBLM_R_X5Y113_SLICE_X6Y113_AO6),
.I1(CLBLM_R_X5Y112_SLICE_X6Y112_CO6),
.I2(CLBLM_R_X5Y115_SLICE_X6Y115_BO6),
.I3(CLBLM_R_X5Y112_SLICE_X6Y112_AO5),
.I4(CLBLM_R_X3Y114_SLICE_X3Y114_AO6),
.I5(CLBLM_R_X5Y113_SLICE_X6Y113_BO6),
.O5(CLBLM_R_X5Y114_SLICE_X6Y114_CO5),
.O6(CLBLM_R_X5Y114_SLICE_X6Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h69969696c33c3c3c)
  ) CLBLM_R_X5Y114_SLICE_X6Y114_BLUT (
.I0(LIOB33_X0Y115_IOB_X0Y115_I),
.I1(CLBLM_R_X5Y113_SLICE_X6Y113_BO6),
.I2(CLBLM_R_X7Y113_SLICE_X9Y113_BO6),
.I3(LIOB33_X0Y113_IOB_X0Y114_I),
.I4(LIOB33_X0Y113_IOB_X0Y113_I),
.I5(LIOB33_X0Y103_IOB_X0Y103_I),
.O5(CLBLM_R_X5Y114_SLICE_X6Y114_BO5),
.O6(CLBLM_R_X5Y114_SLICE_X6Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h699966690ff0f00f)
  ) CLBLM_R_X5Y114_SLICE_X6Y114_ALUT (
.I0(CLBLM_R_X5Y113_SLICE_X6Y113_DO6),
.I1(CLBLM_R_X5Y115_SLICE_X6Y115_BO6),
.I2(CLBLM_R_X5Y112_SLICE_X6Y112_CO6),
.I3(CLBLM_R_X5Y114_SLICE_X6Y114_BO6),
.I4(CLBLM_R_X5Y113_SLICE_X6Y113_AO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y114_SLICE_X6Y114_AO5),
.O6(CLBLM_R_X5Y114_SLICE_X6Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y114_SLICE_X7Y114_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y114_SLICE_X7Y114_DO5),
.O6(CLBLM_R_X5Y114_SLICE_X7Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y114_SLICE_X7Y114_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y114_SLICE_X7Y114_CO5),
.O6(CLBLM_R_X5Y114_SLICE_X7Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y114_SLICE_X7Y114_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y114_SLICE_X7Y114_BO5),
.O6(CLBLM_R_X5Y114_SLICE_X7Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y114_SLICE_X7Y114_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y114_SLICE_X7Y114_AO5),
.O6(CLBLM_R_X5Y114_SLICE_X7Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7f13b320ff5fffa0)
  ) CLBLM_R_X5Y115_SLICE_X6Y115_DLUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(LIOB33_X0Y115_IOB_X0Y116_I),
.I2(LIOB33_X0Y113_IOB_X0Y113_I),
.I3(CLBLM_R_X7Y116_SLICE_X8Y116_AO6),
.I4(CLBLM_R_X7Y116_SLICE_X9Y116_AO6),
.I5(LIOB33_X0Y115_IOB_X0Y115_I),
.O5(CLBLM_R_X5Y115_SLICE_X6Y115_DO5),
.O6(CLBLM_R_X5Y115_SLICE_X6Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6f06af0aff66ffaa)
  ) CLBLM_R_X5Y115_SLICE_X6Y115_CLUT (
.I0(CLBLM_R_X7Y115_SLICE_X8Y115_AO6),
.I1(LIOB33_X0Y115_IOB_X0Y116_I),
.I2(LIOB33_X0Y113_IOB_X0Y114_I),
.I3(CLBLM_R_X7Y113_SLICE_X9Y113_CO6),
.I4(LIOB33_X0Y113_IOB_X0Y113_I),
.I5(LIOB33_X0Y115_IOB_X0Y115_I),
.O5(CLBLM_R_X5Y115_SLICE_X6Y115_CO5),
.O6(CLBLM_R_X5Y115_SLICE_X6Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996a55ac33c0ff0)
  ) CLBLM_R_X5Y115_SLICE_X6Y115_BLUT (
.I0(LIOB33_X0Y113_IOB_X0Y113_I),
.I1(LIOB33_X0Y113_IOB_X0Y114_I),
.I2(CLBLM_R_X7Y115_SLICE_X8Y115_AO6),
.I3(CLBLM_R_X7Y113_SLICE_X9Y113_CO6),
.I4(LIOB33_X0Y115_IOB_X0Y115_I),
.I5(LIOB33_X0Y115_IOB_X0Y116_I),
.O5(CLBLM_R_X5Y115_SLICE_X6Y115_BO5),
.O6(CLBLM_R_X5Y115_SLICE_X6Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h7777777733ff33ff)
  ) CLBLM_R_X5Y115_SLICE_X6Y115_ALUT (
.I0(LIOB33_X0Y111_IOB_X0Y112_I),
.I1(LIOB33_X0Y115_IOB_X0Y116_I),
.I2(1'b1),
.I3(LIOB33_X0Y115_IOB_X0Y115_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y115_SLICE_X6Y115_AO5),
.O6(CLBLM_R_X5Y115_SLICE_X6Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hc369693ca5a5f0f0)
  ) CLBLM_R_X5Y115_SLICE_X7Y115_DLUT (
.I0(CLBLM_R_X7Y114_SLICE_X9Y114_CO6),
.I1(RIOB33_X105Y103_IOB_X1Y104_I),
.I2(CLBLL_L_X4Y112_SLICE_X5Y112_CO6),
.I3(RIOB33_X105Y103_IOB_X1Y103_I),
.I4(CLBLL_L_X4Y114_SLICE_X5Y114_AO6),
.I5(LIOB33_X0Y115_IOB_X0Y115_I),
.O5(CLBLM_R_X5Y115_SLICE_X7Y115_DO5),
.O6(CLBLM_R_X5Y115_SLICE_X7Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h48de88eededeeeee)
  ) CLBLM_R_X5Y115_SLICE_X7Y115_CLUT (
.I0(CLBLM_R_X7Y114_SLICE_X9Y114_DO6),
.I1(CLBLM_R_X7Y114_SLICE_X8Y114_CO6),
.I2(LIOB33_X0Y113_IOB_X0Y113_I),
.I3(RIOB33_X105Y101_IOB_X1Y102_I),
.I4(RIOB33_X105Y103_IOB_X1Y103_I),
.I5(LIOB33_X0Y115_IOB_X0Y115_I),
.O5(CLBLM_R_X5Y115_SLICE_X7Y115_CO5),
.O6(CLBLM_R_X5Y115_SLICE_X7Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6c93936c93936c6c)
  ) CLBLM_R_X5Y115_SLICE_X7Y115_BLUT (
.I0(LIOB33_X0Y113_IOB_X0Y113_I),
.I1(CLBLM_R_X7Y114_SLICE_X8Y114_CO6),
.I2(RIOB33_X105Y103_IOB_X1Y103_I),
.I3(LIOB33_X0Y115_IOB_X0Y115_I),
.I4(CLBLM_R_X7Y114_SLICE_X9Y114_DO6),
.I5(RIOB33_X105Y101_IOB_X1Y102_I),
.O5(CLBLM_R_X5Y115_SLICE_X7Y115_BO5),
.O6(CLBLM_R_X5Y115_SLICE_X7Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6a6a95957f7f1515)
  ) CLBLM_R_X5Y115_SLICE_X7Y115_ALUT (
.I0(CLBLL_L_X4Y114_SLICE_X5Y114_AO6),
.I1(LIOB33_X0Y115_IOB_X0Y115_I),
.I2(RIOB33_X105Y103_IOB_X1Y103_I),
.I3(1'b1),
.I4(CLBLM_R_X7Y114_SLICE_X9Y114_CO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y115_SLICE_X7Y115_AO5),
.O6(CLBLM_R_X5Y115_SLICE_X7Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff5f0f057f1f0701)
  ) CLBLM_R_X5Y116_SLICE_X6Y116_DLUT (
.I0(CLBLM_R_X7Y116_SLICE_X8Y116_BO6),
.I1(CLBLM_R_X5Y114_SLICE_X6Y114_DO6),
.I2(CLBLM_R_X5Y116_SLICE_X7Y116_BO6),
.I3(CLBLM_R_X5Y115_SLICE_X6Y115_DO6),
.I4(CLBLM_R_X7Y116_SLICE_X8Y116_CO6),
.I5(CLBLM_R_X5Y116_SLICE_X6Y116_BO6),
.O5(CLBLM_R_X5Y116_SLICE_X6Y116_DO5),
.O6(CLBLM_R_X5Y116_SLICE_X6Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h69965aa5a55a6996)
  ) CLBLM_R_X5Y116_SLICE_X6Y116_CLUT (
.I0(CLBLM_R_X7Y116_SLICE_X9Y116_CO6),
.I1(CLBLM_R_X7Y113_SLICE_X9Y113_CO6),
.I2(CLBLM_R_X7Y116_SLICE_X8Y116_AO6),
.I3(CLBLM_R_X5Y115_SLICE_X6Y115_AO5),
.I4(CLBLM_R_X7Y116_SLICE_X8Y116_DO6),
.I5(CLBLL_L_X4Y116_SLICE_X4Y116_AO6),
.O5(CLBLM_R_X5Y116_SLICE_X6Y116_CO5),
.O6(CLBLM_R_X5Y116_SLICE_X6Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3110c440c4403110)
  ) CLBLM_R_X5Y116_SLICE_X6Y116_BLUT (
.I0(CLBLM_R_X7Y116_SLICE_X8Y116_DO6),
.I1(CLBLM_R_X7Y116_SLICE_X8Y116_AO6),
.I2(CLBLM_R_X7Y113_SLICE_X9Y113_CO6),
.I3(CLBLL_L_X4Y116_SLICE_X4Y116_AO6),
.I4(CLBLM_R_X7Y116_SLICE_X9Y116_CO6),
.I5(CLBLM_R_X5Y115_SLICE_X6Y115_AO5),
.O5(CLBLM_R_X5Y116_SLICE_X6Y116_BO5),
.O6(CLBLM_R_X5Y116_SLICE_X6Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8eff08ef08ef008e)
  ) CLBLM_R_X5Y116_SLICE_X6Y116_ALUT (
.I0(CLBLM_R_X5Y115_SLICE_X6Y115_CO6),
.I1(CLBLM_R_X7Y116_SLICE_X8Y116_AO6),
.I2(CLBLM_R_X7Y116_SLICE_X9Y116_CO6),
.I3(CLBLM_R_X7Y116_SLICE_X8Y116_BO6),
.I4(CLBLM_R_X5Y114_SLICE_X6Y114_CO6),
.I5(CLBLM_R_X5Y115_SLICE_X6Y115_AO5),
.O5(CLBLM_R_X5Y116_SLICE_X6Y116_AO5),
.O6(CLBLM_R_X5Y116_SLICE_X6Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haa55aa5555aa55aa)
  ) CLBLM_R_X5Y116_SLICE_X7Y116_DLUT (
.I0(CLBLM_R_X5Y115_SLICE_X7Y115_AO6),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X5Y116_SLICE_X7Y116_CO6),
.I4(1'b1),
.I5(CLBLM_R_X5Y115_SLICE_X7Y115_CO6),
.O5(CLBLM_R_X5Y116_SLICE_X7Y116_DO5),
.O6(CLBLM_R_X5Y116_SLICE_X7Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000e880fee8fffe)
  ) CLBLM_R_X5Y116_SLICE_X7Y116_CLUT (
.I0(CLBLM_R_X7Y114_SLICE_X9Y114_BO6),
.I1(CLBLM_R_X5Y116_SLICE_X6Y116_AO6),
.I2(CLBLM_R_X7Y116_SLICE_X8Y116_CO6),
.I3(CLBLM_R_X5Y116_SLICE_X7Y116_AO5),
.I4(CLBLL_L_X4Y115_SLICE_X5Y115_AO6),
.I5(CLBLM_R_X5Y115_SLICE_X7Y115_BO6),
.O5(CLBLM_R_X5Y116_SLICE_X7Y116_CO5),
.O6(CLBLM_R_X5Y116_SLICE_X7Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7888877787777888)
  ) CLBLM_R_X5Y116_SLICE_X7Y116_BLUT (
.I0(LIOB33_X0Y113_IOB_X0Y113_I),
.I1(RIOB33_X105Y101_IOB_X1Y102_I),
.I2(LIOB33_X0Y115_IOB_X0Y115_I),
.I3(RIOB33_X105Y101_IOB_X1Y101_I),
.I4(CLBLM_R_X7Y114_SLICE_X8Y114_BO6),
.I5(CLBLM_R_X7Y114_SLICE_X9Y114_BO6),
.O5(CLBLM_R_X5Y116_SLICE_X7Y116_BO5),
.O6(CLBLM_R_X5Y116_SLICE_X7Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0ccfcfcf00ffffff)
  ) CLBLM_R_X5Y116_SLICE_X7Y116_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y114_SLICE_X9Y114_BO6),
.I2(CLBLL_L_X4Y115_SLICE_X5Y115_AO6),
.I3(RIOB33_X105Y101_IOB_X1Y101_I),
.I4(LIOB33_X0Y115_IOB_X0Y115_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y116_SLICE_X7Y116_AO5),
.O6(CLBLM_R_X5Y116_SLICE_X7Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y104_SLICE_X8Y104_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y104_SLICE_X8Y104_DO5),
.O6(CLBLM_R_X7Y104_SLICE_X8Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y104_SLICE_X8Y104_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y104_SLICE_X8Y104_CO5),
.O6(CLBLM_R_X7Y104_SLICE_X8Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y104_SLICE_X8Y104_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y104_SLICE_X8Y104_BO5),
.O6(CLBLM_R_X7Y104_SLICE_X8Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h53235cdc28282828)
  ) CLBLM_R_X7Y104_SLICE_X8Y104_ALUT (
.I0(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I1(RIOB33_X105Y101_IOB_X1Y101_I),
.I2(RIOB33_X105Y101_IOB_X1Y102_I),
.I3(RIOB33_X105Y111_IOB_X1Y112_I),
.I4(RIOB33_X105Y103_IOB_X1Y103_I),
.I5(RIOB33_X105Y113_IOB_X1Y113_I),
.O5(CLBLM_R_X7Y104_SLICE_X8Y104_AO5),
.O6(CLBLM_R_X7Y104_SLICE_X8Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfaa0fee0af0aef0e)
  ) CLBLM_R_X7Y104_SLICE_X9Y104_DLUT (
.I0(CLBLM_R_X7Y104_SLICE_X9Y104_CO6),
.I1(CLBLM_R_X7Y104_SLICE_X9Y104_AO6),
.I2(CLBLM_L_X8Y105_SLICE_X10Y105_AO6),
.I3(CLBLM_R_X7Y104_SLICE_X9Y104_AO5),
.I4(CLBLM_R_X7Y104_SLICE_X8Y104_AO6),
.I5(CLBLM_L_X8Y104_SLICE_X10Y104_AO6),
.O5(CLBLM_R_X7Y104_SLICE_X9Y104_DO5),
.O6(CLBLM_R_X7Y104_SLICE_X9Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h1c0f505055000000)
  ) CLBLM_R_X7Y104_SLICE_X9Y104_CLUT (
.I0(RIOB33_X105Y101_IOB_X1Y101_I),
.I1(RIOB33_X105Y111_IOB_X1Y112_I),
.I2(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I3(RIOB33_X105Y103_IOB_X1Y103_I),
.I4(RIOB33_X105Y113_IOB_X1Y113_I),
.I5(RIOB33_X105Y101_IOB_X1Y102_I),
.O5(CLBLM_R_X7Y104_SLICE_X9Y104_CO5),
.O6(CLBLM_R_X7Y104_SLICE_X9Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h55aaa659aa5559a6)
  ) CLBLM_R_X7Y104_SLICE_X9Y104_BLUT (
.I0(CLBLM_L_X8Y105_SLICE_X10Y105_AO6),
.I1(CLBLM_R_X7Y104_SLICE_X9Y104_AO6),
.I2(CLBLM_R_X7Y104_SLICE_X8Y104_AO6),
.I3(CLBLM_L_X8Y104_SLICE_X10Y104_AO6),
.I4(CLBLM_R_X7Y104_SLICE_X9Y104_CO6),
.I5(CLBLM_R_X7Y104_SLICE_X9Y104_AO5),
.O5(CLBLM_R_X7Y104_SLICE_X9Y104_BO5),
.O6(CLBLM_R_X7Y104_SLICE_X9Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333ffff00ffffff)
  ) CLBLM_R_X7Y104_SLICE_X9Y104_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y101_IOB_X0Y101_I),
.I2(1'b1),
.I3(LIOB33_X0Y101_IOB_X0Y102_I),
.I4(RIOB33_X105Y101_IOB_X1Y101_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y104_SLICE_X9Y104_AO5),
.O6(CLBLM_R_X7Y104_SLICE_X9Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hee88fec8bb22fb32)
  ) CLBLM_R_X7Y105_SLICE_X8Y105_DLUT (
.I0(CLBLM_R_X5Y105_SLICE_X7Y105_AO6),
.I1(CLBLM_R_X7Y104_SLICE_X9Y104_AO6),
.I2(CLBLM_R_X7Y106_SLICE_X8Y106_AO6),
.I3(CLBLM_R_X7Y106_SLICE_X8Y106_AO5),
.I4(CLBLM_R_X7Y106_SLICE_X8Y106_CO6),
.I5(CLBLM_R_X7Y104_SLICE_X8Y104_AO6),
.O5(CLBLM_R_X7Y105_SLICE_X8Y105_DO5),
.O6(CLBLM_R_X7Y105_SLICE_X8Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h78871ee18778e11e)
  ) CLBLM_R_X7Y105_SLICE_X8Y105_CLUT (
.I0(CLBLM_R_X7Y105_SLICE_X8Y105_AO6),
.I1(CLBLL_L_X4Y105_SLICE_X4Y105_DO6),
.I2(CLBLM_R_X7Y105_SLICE_X8Y105_DO6),
.I3(CLBLM_R_X7Y105_SLICE_X8Y105_AO5),
.I4(CLBLM_R_X7Y105_SLICE_X8Y105_BO6),
.I5(CLBLM_R_X7Y104_SLICE_X9Y104_BO6),
.O5(CLBLM_R_X7Y105_SLICE_X8Y105_CO5),
.O6(CLBLM_R_X7Y105_SLICE_X8Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h33cc9c63cc33639c)
  ) CLBLM_R_X7Y105_SLICE_X8Y105_BLUT (
.I0(CLBLM_R_X7Y106_SLICE_X8Y106_CO6),
.I1(CLBLM_R_X7Y104_SLICE_X9Y104_AO6),
.I2(CLBLM_R_X7Y106_SLICE_X8Y106_AO6),
.I3(CLBLM_R_X7Y104_SLICE_X8Y104_AO6),
.I4(CLBLM_R_X5Y105_SLICE_X7Y105_AO6),
.I5(CLBLM_R_X7Y106_SLICE_X8Y106_AO5),
.O5(CLBLM_R_X7Y105_SLICE_X8Y105_BO5),
.O6(CLBLM_R_X7Y105_SLICE_X8Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h7777777733ff33ff)
  ) CLBLM_R_X7Y105_SLICE_X8Y105_ALUT (
.I0(LIOB33_X0Y115_IOB_X0Y116_I),
.I1(LIOB33_X0Y103_IOB_X0Y104_I),
.I2(1'b1),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y105_SLICE_X8Y105_AO5),
.O6(CLBLM_R_X7Y105_SLICE_X8Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y105_SLICE_X9Y105_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y105_SLICE_X9Y105_DO5),
.O6(CLBLM_R_X7Y105_SLICE_X9Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y105_SLICE_X9Y105_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y105_SLICE_X9Y105_CO5),
.O6(CLBLM_R_X7Y105_SLICE_X9Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y105_SLICE_X9Y105_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y105_SLICE_X9Y105_BO5),
.O6(CLBLM_R_X7Y105_SLICE_X9Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h599aa665a665599a)
  ) CLBLM_R_X7Y105_SLICE_X9Y105_ALUT (
.I0(CLBLM_R_X7Y104_SLICE_X9Y104_DO6),
.I1(CLBLM_R_X7Y104_SLICE_X9Y104_BO6),
.I2(CLBLM_R_X7Y105_SLICE_X8Y105_AO5),
.I3(CLBLM_R_X7Y105_SLICE_X8Y105_DO6),
.I4(CLBLM_L_X8Y107_SLICE_X10Y107_AO6),
.I5(CLBLM_L_X8Y105_SLICE_X10Y105_BO6),
.O5(CLBLM_R_X7Y105_SLICE_X9Y105_AO5),
.O6(CLBLM_R_X7Y105_SLICE_X9Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y106_SLICE_X8Y106_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y106_SLICE_X8Y106_DO5),
.O6(CLBLM_R_X7Y106_SLICE_X8Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f6630c0656630c0)
  ) CLBLM_R_X7Y106_SLICE_X8Y106_CLUT (
.I0(RIOB33_X105Y101_IOB_X1Y102_I),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I3(RIOB33_X105Y101_IOB_X1Y101_I),
.I4(RIOB33_X105Y113_IOB_X1Y113_I),
.I5(RIOB33_X105Y111_IOB_X1Y112_I),
.O5(CLBLM_R_X7Y106_SLICE_X8Y106_CO5),
.O6(CLBLM_R_X7Y106_SLICE_X8Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa0055ffccccddff)
  ) CLBLM_R_X7Y106_SLICE_X8Y106_BLUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(CLBLM_R_X5Y105_SLICE_X7Y105_AO6),
.I2(1'b1),
.I3(LIOB33_X0Y101_IOB_X0Y101_I),
.I4(CLBLM_R_X7Y106_SLICE_X8Y106_CO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y106_SLICE_X8Y106_BO5),
.O6(CLBLM_R_X7Y106_SLICE_X8Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h33ff33ff0fff0fff)
  ) CLBLM_R_X7Y106_SLICE_X8Y106_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y101_IOB_X0Y101_I),
.I2(LIOB33_X0Y101_IOB_X0Y102_I),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y106_SLICE_X8Y106_AO5),
.O6(CLBLM_R_X7Y106_SLICE_X8Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hbd42718e39c6f50a)
  ) CLBLM_R_X7Y106_SLICE_X9Y106_DLUT (
.I0(CLBLM_R_X7Y106_SLICE_X9Y106_AO6),
.I1(LIOB33_X0Y101_IOB_X0Y102_I),
.I2(CLBLM_R_X7Y106_SLICE_X8Y106_BO5),
.I3(CLBLM_R_X7Y106_SLICE_X9Y106_CO6),
.I4(RIOB33_X105Y101_IOB_X1Y101_I),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLM_R_X7Y106_SLICE_X9Y106_DO5),
.O6(CLBLM_R_X7Y106_SLICE_X9Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6c6f6c5f939093a0)
  ) CLBLM_R_X7Y106_SLICE_X9Y106_CLUT (
.I0(RIOB33_X105Y101_IOB_X1Y102_I),
.I1(CLBLM_R_X7Y104_SLICE_X9Y104_CO6),
.I2(LIOB33_X0Y101_IOB_X0Y101_I),
.I3(CLBLM_R_X7Y104_SLICE_X8Y104_AO6),
.I4(RIOB33_X105Y101_IOB_X1Y101_I),
.I5(CLBLM_L_X8Y104_SLICE_X10Y104_AO6),
.O5(CLBLM_R_X7Y106_SLICE_X9Y106_CO5),
.O6(CLBLM_R_X7Y106_SLICE_X9Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h69c39933963c66cc)
  ) CLBLM_R_X7Y106_SLICE_X9Y106_BLUT (
.I0(LIOB33_X0Y103_IOB_X0Y104_I),
.I1(CLBLM_R_X7Y105_SLICE_X8Y105_DO6),
.I2(LIOB33_X0Y101_IOB_X0Y102_I),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(RIOB33_X105Y101_IOB_X1Y101_I),
.I5(CLBLM_R_X7Y106_SLICE_X9Y106_CO6),
.O5(CLBLM_R_X7Y106_SLICE_X9Y106_BO5),
.O6(CLBLM_R_X7Y106_SLICE_X9Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa555555ccdddddd)
  ) CLBLM_R_X7Y106_SLICE_X9Y106_ALUT (
.I0(CLBLM_R_X7Y104_SLICE_X8Y104_AO6),
.I1(CLBLM_R_X7Y104_SLICE_X9Y104_CO6),
.I2(1'b1),
.I3(LIOB33_X0Y101_IOB_X0Y101_I),
.I4(RIOB33_X105Y101_IOB_X1Y101_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y106_SLICE_X9Y106_AO5),
.O6(CLBLM_R_X7Y106_SLICE_X9Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y107_SLICE_X8Y107_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y107_SLICE_X8Y107_DO5),
.O6(CLBLM_R_X7Y107_SLICE_X8Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y107_SLICE_X8Y107_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y107_SLICE_X8Y107_CO5),
.O6(CLBLM_R_X7Y107_SLICE_X8Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y107_SLICE_X8Y107_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y107_SLICE_X8Y107_BO5),
.O6(CLBLM_R_X7Y107_SLICE_X8Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y107_SLICE_X8Y107_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y107_SLICE_X8Y107_AO5),
.O6(CLBLM_R_X7Y107_SLICE_X8Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h28bebebea0fafafa)
  ) CLBLM_R_X7Y107_SLICE_X9Y107_DLUT (
.I0(CLBLM_R_X5Y105_SLICE_X6Y105_AO6),
.I1(LIOB33_X0Y103_IOB_X0Y104_I),
.I2(CLBLM_R_X7Y106_SLICE_X9Y106_DO6),
.I3(LIOB33_X0Y115_IOB_X0Y116_I),
.I4(LIOB33_X0Y105_IOB_X0Y105_I),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLM_R_X7Y107_SLICE_X9Y107_DO5),
.O6(CLBLM_R_X7Y107_SLICE_X9Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hda2a25d54fbfb040)
  ) CLBLM_R_X7Y107_SLICE_X9Y107_CLUT (
.I0(CLBLM_R_X5Y105_SLICE_X6Y105_AO6),
.I1(LIOB33_X0Y115_IOB_X0Y116_I),
.I2(LIOB33_X0Y105_IOB_X0Y105_I),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(CLBLM_R_X7Y105_SLICE_X9Y105_AO6),
.I5(CLBLM_R_X7Y106_SLICE_X9Y106_BO6),
.O5(CLBLM_R_X7Y107_SLICE_X9Y107_CO5),
.O6(CLBLM_R_X7Y107_SLICE_X9Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf9ff909999f90090)
  ) CLBLM_R_X7Y107_SLICE_X9Y107_BLUT (
.I0(CLBLM_R_X7Y105_SLICE_X9Y105_AO6),
.I1(CLBLM_R_X7Y108_SLICE_X9Y108_AO6),
.I2(CLBLM_R_X5Y105_SLICE_X6Y105_AO6),
.I3(CLBLM_R_X7Y106_SLICE_X9Y106_BO6),
.I4(CLBLM_R_X5Y106_SLICE_X7Y106_AO6),
.I5(CLBLM_R_X7Y108_SLICE_X9Y108_AO5),
.O5(CLBLM_R_X7Y107_SLICE_X9Y107_BO5),
.O6(CLBLM_R_X7Y107_SLICE_X9Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3cc396699669c33c)
  ) CLBLM_R_X7Y107_SLICE_X9Y107_ALUT (
.I0(CLBLM_R_X7Y106_SLICE_X9Y106_BO6),
.I1(CLBLM_R_X7Y108_SLICE_X9Y108_AO6),
.I2(CLBLM_R_X7Y105_SLICE_X9Y105_AO6),
.I3(CLBLM_R_X5Y106_SLICE_X7Y106_AO6),
.I4(CLBLM_R_X5Y105_SLICE_X6Y105_AO6),
.I5(CLBLM_R_X7Y108_SLICE_X9Y108_AO5),
.O5(CLBLM_R_X7Y107_SLICE_X9Y107_AO5),
.O6(CLBLM_R_X7Y107_SLICE_X9Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y108_SLICE_X8Y108_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y108_SLICE_X8Y108_DO5),
.O6(CLBLM_R_X7Y108_SLICE_X8Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h71d4f3fcf550fff0)
  ) CLBLM_R_X7Y108_SLICE_X8Y108_CLUT (
.I0(LIOB33_X0Y107_IOB_X0Y107_I),
.I1(LIOB33_X0Y115_IOB_X0Y116_I),
.I2(CLBLM_R_X5Y106_SLICE_X7Y106_DO6),
.I3(CLBLM_R_X7Y107_SLICE_X9Y107_CO6),
.I4(LIOB33_X0Y113_IOB_X0Y114_I),
.I5(LIOB33_X0Y105_IOB_X0Y106_I),
.O5(CLBLM_R_X7Y108_SLICE_X8Y108_CO5),
.O6(CLBLM_R_X7Y108_SLICE_X8Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h639cc6399c6339c6)
  ) CLBLM_R_X7Y108_SLICE_X8Y108_BLUT (
.I0(CLBLM_R_X5Y106_SLICE_X7Y106_DO6),
.I1(CLBLM_L_X8Y108_SLICE_X10Y108_AO6),
.I2(CLBLM_R_X7Y107_SLICE_X9Y107_AO6),
.I3(CLBLM_R_X7Y107_SLICE_X9Y107_BO6),
.I4(CLBLM_R_X7Y108_SLICE_X8Y108_AO6),
.I5(CLBLM_R_X7Y108_SLICE_X8Y108_AO5),
.O5(CLBLM_R_X7Y108_SLICE_X8Y108_BO5),
.O6(CLBLM_R_X7Y108_SLICE_X8Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0fffff3f3f3f3f)
  ) CLBLM_R_X7Y108_SLICE_X8Y108_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y115_IOB_X0Y116_I),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(1'b1),
.I4(LIOB33_X0Y113_IOB_X0Y114_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y108_SLICE_X8Y108_AO5),
.O6(CLBLM_R_X7Y108_SLICE_X8Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h4d8ecf0cddeeffcc)
  ) CLBLM_R_X7Y108_SLICE_X9Y108_DLUT (
.I0(LIOB33_X0Y107_IOB_X0Y107_I),
.I1(CLBLM_R_X7Y108_SLICE_X8Y108_CO6),
.I2(LIOB33_X0Y107_IOB_X0Y108_I),
.I3(CLBLM_R_X7Y108_SLICE_X9Y108_CO6),
.I4(LIOB33_X0Y115_IOB_X0Y116_I),
.I5(LIOB33_X0Y113_IOB_X0Y114_I),
.O5(CLBLM_R_X7Y108_SLICE_X9Y108_DO5),
.O6(CLBLM_R_X7Y108_SLICE_X9Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hb44b2dd2dd22dd22)
  ) CLBLM_R_X7Y108_SLICE_X9Y108_CLUT (
.I0(CLBLM_L_X8Y108_SLICE_X11Y108_BO6),
.I1(CLBLM_R_X7Y107_SLICE_X9Y107_DO6),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(CLBLM_L_X8Y108_SLICE_X10Y108_DO6),
.I4(LIOB33_X0Y115_IOB_X0Y116_I),
.I5(LIOB33_X0Y105_IOB_X0Y106_I),
.O5(CLBLM_R_X7Y108_SLICE_X9Y108_CO5),
.O6(CLBLM_R_X7Y108_SLICE_X9Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h4db2b24db24d4db2)
  ) CLBLM_R_X7Y108_SLICE_X9Y108_BLUT (
.I0(CLBLM_R_X7Y108_SLICE_X8Y108_AO5),
.I1(CLBLM_L_X8Y108_SLICE_X10Y108_AO6),
.I2(CLBLM_R_X7Y107_SLICE_X9Y107_BO6),
.I3(CLBLM_L_X8Y108_SLICE_X10Y108_CO6),
.I4(CLBLM_L_X10Y110_SLICE_X12Y110_AO6),
.I5(CLBLM_L_X10Y108_SLICE_X12Y108_BO6),
.O5(CLBLM_R_X7Y108_SLICE_X9Y108_BO5),
.O6(CLBLM_R_X7Y108_SLICE_X9Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f3f3f3f0fff0fff)
  ) CLBLM_R_X7Y108_SLICE_X9Y108_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(LIOB33_X0Y105_IOB_X0Y105_I),
.I3(LIOB33_X0Y115_IOB_X0Y116_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y108_SLICE_X9Y108_AO5),
.O6(CLBLM_R_X7Y108_SLICE_X9Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h639cc6399c6339c6)
  ) CLBLM_R_X7Y109_SLICE_X8Y109_DLUT (
.I0(CLBLM_R_X7Y109_SLICE_X8Y109_AO6),
.I1(CLBLM_R_X5Y109_SLICE_X6Y109_AO5),
.I2(CLBLM_R_X7Y109_SLICE_X9Y109_BO6),
.I3(CLBLM_R_X7Y109_SLICE_X8Y109_AO5),
.I4(CLBLM_R_X7Y108_SLICE_X8Y108_CO6),
.I5(CLBLM_R_X7Y108_SLICE_X9Y108_BO6),
.O5(CLBLM_R_X7Y109_SLICE_X8Y109_DO5),
.O6(CLBLM_R_X7Y109_SLICE_X8Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hef8cce088cef08ce)
  ) CLBLM_R_X7Y109_SLICE_X8Y109_CLUT (
.I0(CLBLM_R_X7Y109_SLICE_X8Y109_AO6),
.I1(CLBLM_R_X5Y109_SLICE_X6Y109_AO5),
.I2(CLBLM_R_X7Y109_SLICE_X9Y109_BO6),
.I3(CLBLM_R_X7Y109_SLICE_X8Y109_AO5),
.I4(CLBLM_R_X7Y108_SLICE_X8Y108_CO6),
.I5(CLBLM_R_X7Y108_SLICE_X9Y108_BO6),
.O5(CLBLM_R_X7Y109_SLICE_X8Y109_CO5),
.O6(CLBLM_R_X7Y109_SLICE_X8Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h956aaaaaa9566666)
  ) CLBLM_R_X7Y109_SLICE_X8Y109_BLUT (
.I0(CLBLM_R_X7Y108_SLICE_X9Y108_BO6),
.I1(CLBLM_R_X7Y109_SLICE_X9Y109_BO6),
.I2(LIOB33_X0Y113_IOB_X0Y114_I),
.I3(LIOB33_X0Y115_IOB_X0Y116_I),
.I4(LIOB33_X0Y107_IOB_X0Y108_I),
.I5(CLBLM_R_X7Y108_SLICE_X8Y108_CO6),
.O5(CLBLM_R_X7Y109_SLICE_X8Y109_BO5),
.O6(CLBLM_R_X7Y109_SLICE_X8Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0fffff3333ffff)
  ) CLBLM_R_X7Y109_SLICE_X8Y109_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y115_IOB_X0Y116_I),
.I2(LIOB33_X0Y113_IOB_X0Y114_I),
.I3(1'b1),
.I4(LIOB33_X0Y107_IOB_X0Y108_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y109_SLICE_X8Y109_AO5),
.O6(CLBLM_R_X7Y109_SLICE_X8Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h2888beeebeeebeee)
  ) CLBLM_R_X7Y109_SLICE_X9Y109_DLUT (
.I0(CLBLM_R_X7Y107_SLICE_X9Y107_BO6),
.I1(CLBLM_L_X8Y108_SLICE_X10Y108_DO6),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(LIOB33_X0Y107_IOB_X0Y107_I),
.I5(LIOB33_X0Y115_IOB_X0Y116_I),
.O5(CLBLM_R_X7Y109_SLICE_X9Y109_DO5),
.O6(CLBLM_R_X7Y109_SLICE_X9Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6a95956a956a956a)
  ) CLBLM_R_X7Y109_SLICE_X9Y109_CLUT (
.I0(CLBLM_R_X7Y108_SLICE_X9Y108_CO6),
.I1(LIOB33_X0Y107_IOB_X0Y108_I),
.I2(LIOB33_X0Y113_IOB_X0Y114_I),
.I3(CLBLM_R_X7Y108_SLICE_X8Y108_CO6),
.I4(LIOB33_X0Y107_IOB_X0Y107_I),
.I5(LIOB33_X0Y115_IOB_X0Y116_I),
.O5(CLBLM_R_X7Y109_SLICE_X9Y109_CO5),
.O6(CLBLM_R_X7Y109_SLICE_X9Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h69969696c33c3c3c)
  ) CLBLM_R_X7Y109_SLICE_X9Y109_BLUT (
.I0(LIOB33_X0Y107_IOB_X0Y107_I),
.I1(CLBLM_L_X8Y108_SLICE_X10Y108_DO6),
.I2(CLBLM_R_X7Y107_SLICE_X9Y107_BO6),
.I3(LIOB33_X0Y105_IOB_X0Y106_I),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(LIOB33_X0Y115_IOB_X0Y116_I),
.O5(CLBLM_R_X7Y109_SLICE_X9Y109_BO5),
.O6(CLBLM_R_X7Y109_SLICE_X9Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0fffff6699cc33)
  ) CLBLM_R_X7Y109_SLICE_X9Y109_ALUT (
.I0(LIOB33_X0Y109_IOB_X0Y109_I),
.I1(CLBLM_R_X5Y108_SLICE_X7Y108_BO6),
.I2(LIOB33_X0Y101_IOB_X0Y101_I),
.I3(CLBLM_L_X8Y109_SLICE_X10Y109_AO6),
.I4(RIOB33_X105Y107_IOB_X1Y108_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y109_SLICE_X9Y109_AO5),
.O6(CLBLM_R_X7Y109_SLICE_X9Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y110_SLICE_X8Y110_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y110_SLICE_X8Y110_DO5),
.O6(CLBLM_R_X7Y110_SLICE_X8Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'he178695a4bd2c3f0)
  ) CLBLM_R_X7Y110_SLICE_X8Y110_CLUT (
.I0(LIOB33_X0Y113_IOB_X0Y114_I),
.I1(CLBLM_R_X7Y108_SLICE_X9Y108_DO6),
.I2(CLBLM_L_X8Y110_SLICE_X11Y110_AO6),
.I3(CLBLM_L_X8Y109_SLICE_X10Y109_CO6),
.I4(LIOB33_X0Y109_IOB_X0Y109_I),
.I5(LIOB33_X0Y109_IOB_X0Y110_I),
.O5(CLBLM_R_X7Y110_SLICE_X8Y110_CO5),
.O6(CLBLM_R_X7Y110_SLICE_X8Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0b3b2bbb2fbf3fff)
  ) CLBLM_R_X7Y110_SLICE_X8Y110_BLUT (
.I0(CLBLM_R_X7Y108_SLICE_X9Y108_DO6),
.I1(CLBLM_L_X8Y110_SLICE_X11Y110_AO6),
.I2(LIOB33_X0Y113_IOB_X0Y114_I),
.I3(LIOB33_X0Y109_IOB_X0Y110_I),
.I4(LIOB33_X0Y109_IOB_X0Y109_I),
.I5(CLBLM_L_X8Y109_SLICE_X10Y109_CO6),
.O5(CLBLM_R_X7Y110_SLICE_X8Y110_BO5),
.O6(CLBLM_R_X7Y110_SLICE_X8Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996c33c3cc36996)
  ) CLBLM_R_X7Y110_SLICE_X8Y110_ALUT (
.I0(CLBLM_R_X5Y109_SLICE_X6Y109_DO6),
.I1(CLBLM_L_X8Y110_SLICE_X11Y110_AO6),
.I2(CLBLM_R_X7Y109_SLICE_X8Y109_CO6),
.I3(CLBLM_R_X7Y110_SLICE_X9Y110_AO5),
.I4(CLBLM_R_X5Y110_SLICE_X7Y110_BO5),
.I5(CLBLM_R_X7Y109_SLICE_X8Y109_DO6),
.O5(CLBLM_R_X7Y110_SLICE_X8Y110_AO5),
.O6(CLBLM_R_X7Y110_SLICE_X8Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8f70e31c7f8013ec)
  ) CLBLM_R_X7Y110_SLICE_X9Y110_DLUT (
.I0(LIOB33_X0Y113_IOB_X0Y114_I),
.I1(CLBLM_L_X8Y109_SLICE_X10Y109_CO6),
.I2(LIOB33_X0Y109_IOB_X0Y109_I),
.I3(CLBLM_L_X8Y110_SLICE_X10Y110_DO6),
.I4(CLBLM_R_X7Y108_SLICE_X9Y108_DO6),
.I5(LIOB33_X0Y115_IOB_X0Y116_I),
.O5(CLBLM_R_X7Y110_SLICE_X9Y110_DO5),
.O6(CLBLM_R_X7Y110_SLICE_X9Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h693cc36996c33c96)
  ) CLBLM_R_X7Y110_SLICE_X9Y110_CLUT (
.I0(CLBLM_R_X7Y110_SLICE_X9Y110_AO6),
.I1(CLBLM_R_X7Y109_SLICE_X9Y109_AO5),
.I2(CLBLM_L_X8Y110_SLICE_X10Y110_CO6),
.I3(CLBLM_L_X8Y110_SLICE_X10Y110_BO6),
.I4(CLBLM_L_X10Y111_SLICE_X12Y111_CO6),
.I5(CLBLM_R_X5Y110_SLICE_X7Y110_BO6),
.O5(CLBLM_R_X7Y110_SLICE_X9Y110_CO5),
.O6(CLBLM_R_X7Y110_SLICE_X9Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6969a5a52b2bafaf)
  ) CLBLM_R_X7Y110_SLICE_X9Y110_BLUT (
.I0(CLBLM_L_X8Y110_SLICE_X10Y110_CO6),
.I1(LIOB33_X0Y109_IOB_X0Y110_I),
.I2(CLBLM_R_X7Y109_SLICE_X9Y109_AO5),
.I3(1'b1),
.I4(RIOB33_X105Y107_IOB_X1Y107_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y110_SLICE_X9Y110_BO5),
.O6(CLBLM_R_X7Y110_SLICE_X9Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h777777773f3f3f3f)
  ) CLBLM_R_X7Y110_SLICE_X9Y110_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(LIOB33_X0Y109_IOB_X0Y110_I),
.I2(LIOB33_X0Y113_IOB_X0Y114_I),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y110_SLICE_X9Y110_AO5),
.O6(CLBLM_R_X7Y110_SLICE_X9Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h307370ff33f7f7ff)
  ) CLBLM_R_X7Y111_SLICE_X8Y111_DLUT (
.I0(LIOB33_X0Y111_IOB_X0Y111_I),
.I1(RIOB33_X105Y103_IOB_X1Y104_I),
.I2(CLBLM_L_X10Y111_SLICE_X13Y111_BO6),
.I3(CLBLM_R_X7Y111_SLICE_X8Y111_AO5),
.I4(LIOB33_X0Y111_IOB_X0Y112_I),
.I5(CLBLM_L_X8Y111_SLICE_X10Y111_BO6),
.O5(CLBLM_R_X7Y111_SLICE_X8Y111_DO5),
.O6(CLBLM_R_X7Y111_SLICE_X8Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h9c3963c6c3ccc3cc)
  ) CLBLM_R_X7Y111_SLICE_X8Y111_CLUT (
.I0(RIOB33_X105Y103_IOB_X1Y104_I),
.I1(CLBLM_R_X7Y110_SLICE_X9Y110_CO6),
.I2(CLBLM_L_X10Y111_SLICE_X13Y111_BO6),
.I3(CLBLM_L_X8Y111_SLICE_X10Y111_BO6),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(LIOB33_X0Y111_IOB_X0Y111_I),
.O5(CLBLM_R_X7Y111_SLICE_X8Y111_CO5),
.O6(CLBLM_R_X7Y111_SLICE_X8Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h4c0480c880c84c04)
  ) CLBLM_R_X7Y111_SLICE_X8Y111_BLUT (
.I0(CLBLM_R_X7Y112_SLICE_X9Y112_BO5),
.I1(CLBLM_R_X5Y110_SLICE_X7Y110_AO5),
.I2(CLBLM_L_X10Y111_SLICE_X13Y111_BO6),
.I3(CLBLM_L_X8Y111_SLICE_X10Y111_BO6),
.I4(CLBLM_R_X7Y111_SLICE_X8Y111_AO6),
.I5(CLBLM_R_X7Y110_SLICE_X9Y110_CO6),
.O5(CLBLM_R_X7Y111_SLICE_X8Y111_BO5),
.O6(CLBLM_R_X7Y111_SLICE_X8Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h55ff55ff66cc9933)
  ) CLBLM_R_X7Y111_SLICE_X8Y111_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X8Y111_SLICE_X10Y111_DO6),
.I2(1'b1),
.I3(LIOB33_X0Y111_IOB_X0Y111_I),
.I4(CLBLM_R_X7Y110_SLICE_X9Y110_BO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y111_SLICE_X8Y111_AO5),
.O6(CLBLM_R_X7Y111_SLICE_X8Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y111_SLICE_X9Y111_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y111_SLICE_X9Y111_DO5),
.O6(CLBLM_R_X7Y111_SLICE_X9Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y111_SLICE_X9Y111_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y111_SLICE_X9Y111_CO5),
.O6(CLBLM_R_X7Y111_SLICE_X9Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y111_SLICE_X9Y111_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y111_SLICE_X9Y111_BO5),
.O6(CLBLM_R_X7Y111_SLICE_X9Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00ffff00ff00)
  ) CLBLM_R_X7Y111_SLICE_X9Y111_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_L_X10Y111_SLICE_X13Y111_BO6),
.I4(1'b1),
.I5(CLBLM_L_X8Y111_SLICE_X10Y111_BO6),
.O5(CLBLM_R_X7Y111_SLICE_X9Y111_AO5),
.O6(CLBLM_R_X7Y111_SLICE_X9Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y112_SLICE_X8Y112_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y112_SLICE_X8Y112_DO5),
.O6(CLBLM_R_X7Y112_SLICE_X8Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y112_SLICE_X8Y112_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y112_SLICE_X8Y112_CO5),
.O6(CLBLM_R_X7Y112_SLICE_X8Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h69999666c3333ccc)
  ) CLBLM_R_X7Y112_SLICE_X8Y112_BLUT (
.I0(LIOB33_X0Y109_IOB_X0Y110_I),
.I1(CLBLM_R_X7Y110_SLICE_X8Y110_BO6),
.I2(LIOB33_X0Y113_IOB_X0Y114_I),
.I3(LIOB33_X0Y111_IOB_X0Y111_I),
.I4(CLBLM_L_X8Y112_SLICE_X10Y112_BO6),
.I5(LIOB33_X0Y115_IOB_X0Y116_I),
.O5(CLBLM_R_X7Y112_SLICE_X8Y112_BO5),
.O6(CLBLM_R_X7Y112_SLICE_X8Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6a5695a995a96a56)
  ) CLBLM_R_X7Y112_SLICE_X8Y112_ALUT (
.I0(CLBLM_L_X8Y113_SLICE_X10Y113_AO5),
.I1(CLBLM_R_X7Y110_SLICE_X8Y110_BO6),
.I2(CLBLM_R_X5Y111_SLICE_X6Y111_AO5),
.I3(CLBLM_L_X8Y113_SLICE_X10Y113_BO6),
.I4(CLBLM_R_X5Y112_SLICE_X7Y112_AO6),
.I5(CLBLM_L_X8Y112_SLICE_X10Y112_CO6),
.O5(CLBLM_R_X7Y112_SLICE_X8Y112_AO5),
.O6(CLBLM_R_X7Y112_SLICE_X8Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h95a9aa666a56aa66)
  ) CLBLM_R_X7Y112_SLICE_X9Y112_DLUT (
.I0(CLBLM_R_X7Y111_SLICE_X9Y111_AO6),
.I1(CLBLM_L_X10Y112_SLICE_X12Y112_AO5),
.I2(RIOB33_X105Y103_IOB_X1Y103_I),
.I3(CLBLM_L_X10Y112_SLICE_X12Y112_DO6),
.I4(LIOB33_X0Y111_IOB_X0Y111_I),
.I5(RIOB33_X105Y103_IOB_X1Y104_I),
.O5(CLBLM_R_X7Y112_SLICE_X9Y112_DO5),
.O6(CLBLM_R_X7Y112_SLICE_X9Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6affffff006a6a6a)
  ) CLBLM_R_X7Y112_SLICE_X9Y112_CLUT (
.I0(CLBLM_L_X8Y112_SLICE_X10Y112_BO6),
.I1(LIOB33_X0Y115_IOB_X0Y116_I),
.I2(LIOB33_X0Y109_IOB_X0Y110_I),
.I3(LIOB33_X0Y113_IOB_X0Y114_I),
.I4(LIOB33_X0Y111_IOB_X0Y111_I),
.I5(CLBLM_R_X7Y110_SLICE_X8Y110_BO6),
.O5(CLBLM_R_X7Y112_SLICE_X9Y112_CO5),
.O6(CLBLM_R_X7Y112_SLICE_X9Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc0033ff33ff33ff)
  ) CLBLM_R_X7Y112_SLICE_X9Y112_BLUT (
.I0(1'b1),
.I1(LIOB33_X0Y111_IOB_X0Y111_I),
.I2(1'b1),
.I3(RIOB33_X105Y103_IOB_X1Y104_I),
.I4(CLBLM_R_X7Y111_SLICE_X9Y111_AO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y112_SLICE_X9Y112_BO5),
.O6(CLBLM_R_X7Y112_SLICE_X9Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0000fff4ddd4ddd)
  ) CLBLM_R_X7Y112_SLICE_X9Y112_ALUT (
.I0(CLBLM_L_X10Y112_SLICE_X12Y112_AO5),
.I1(CLBLM_L_X10Y112_SLICE_X12Y112_DO6),
.I2(RIOB33_X105Y103_IOB_X1Y103_I),
.I3(LIOB33_X0Y111_IOB_X0Y111_I),
.I4(CLBLM_L_X10Y112_SLICE_X12Y112_AO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y112_SLICE_X9Y112_AO5),
.O6(CLBLM_R_X7Y112_SLICE_X9Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y113_SLICE_X8Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y113_SLICE_X8Y113_DO5),
.O6(CLBLM_R_X7Y113_SLICE_X8Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y113_SLICE_X8Y113_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y113_SLICE_X8Y113_CO5),
.O6(CLBLM_R_X7Y113_SLICE_X8Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7ff7ff7707707700)
  ) CLBLM_R_X7Y113_SLICE_X8Y113_BLUT (
.I0(LIOB33_X0Y115_IOB_X0Y116_I),
.I1(LIOB33_X0Y111_IOB_X0Y111_I),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(CLBLM_L_X10Y113_SLICE_X12Y113_BO6),
.I4(LIOB33_X0Y109_IOB_X0Y110_I),
.I5(CLBLM_L_X8Y113_SLICE_X10Y113_DO6),
.O5(CLBLM_R_X7Y113_SLICE_X8Y113_BO5),
.O6(CLBLM_R_X7Y113_SLICE_X8Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996996666996996)
  ) CLBLM_R_X7Y113_SLICE_X8Y113_ALUT (
.I0(CLBLM_L_X8Y113_SLICE_X10Y113_AO5),
.I1(CLBLM_L_X8Y113_SLICE_X10Y113_DO6),
.I2(CLBLM_R_X5Y111_SLICE_X6Y111_AO5),
.I3(CLBLM_L_X8Y114_SLICE_X11Y114_BO6),
.I4(CLBLM_R_X7Y110_SLICE_X8Y110_BO6),
.I5(CLBLM_L_X8Y113_SLICE_X10Y113_BO6),
.O5(CLBLM_R_X7Y113_SLICE_X8Y113_AO5),
.O6(CLBLM_R_X7Y113_SLICE_X8Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996969669696996)
  ) CLBLM_R_X7Y113_SLICE_X9Y113_DLUT (
.I0(CLBLM_L_X8Y113_SLICE_X10Y113_AO6),
.I1(CLBLM_L_X10Y112_SLICE_X12Y112_BO6),
.I2(CLBLM_R_X5Y115_SLICE_X6Y115_AO6),
.I3(CLBLM_L_X8Y113_SLICE_X10Y113_DO6),
.I4(CLBLM_L_X8Y113_SLICE_X10Y113_AO5),
.I5(CLBLM_L_X8Y114_SLICE_X11Y114_BO6),
.O5(CLBLM_R_X7Y113_SLICE_X9Y113_DO5),
.O6(CLBLM_R_X7Y113_SLICE_X9Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h373f7fff11153f7f)
  ) CLBLM_R_X7Y113_SLICE_X9Y113_CLUT (
.I0(CLBLM_R_X7Y113_SLICE_X9Y113_AO6),
.I1(LIOB33_X0Y113_IOB_X0Y114_I),
.I2(LIOB33_X0Y113_IOB_X0Y113_I),
.I3(LIOB33_X0Y111_IOB_X0Y112_I),
.I4(CLBLM_R_X7Y113_SLICE_X9Y113_DO6),
.I5(CLBLM_R_X7Y112_SLICE_X9Y112_CO6),
.O5(CLBLM_R_X7Y113_SLICE_X9Y113_CO5),
.O6(CLBLM_R_X7Y113_SLICE_X9Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hd57fb9132a8046ec)
  ) CLBLM_R_X7Y113_SLICE_X9Y113_BLUT (
.I0(LIOB33_X0Y111_IOB_X0Y112_I),
.I1(CLBLM_R_X7Y113_SLICE_X9Y113_AO6),
.I2(LIOB33_X0Y113_IOB_X0Y114_I),
.I3(LIOB33_X0Y115_IOB_X0Y116_I),
.I4(CLBLM_R_X7Y112_SLICE_X9Y112_CO6),
.I5(CLBLM_L_X8Y113_SLICE_X10Y113_CO6),
.O5(CLBLM_R_X7Y113_SLICE_X9Y113_BO5),
.O6(CLBLM_R_X7Y113_SLICE_X9Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h69c39933963c66cc)
  ) CLBLM_R_X7Y113_SLICE_X9Y113_ALUT (
.I0(LIOB33_X0Y115_IOB_X0Y116_I),
.I1(CLBLM_L_X10Y113_SLICE_X12Y113_BO6),
.I2(LIOB33_X0Y109_IOB_X0Y110_I),
.I3(LIOB33_X0Y111_IOB_X0Y111_I),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(CLBLM_L_X8Y113_SLICE_X10Y113_DO6),
.O5(CLBLM_R_X7Y113_SLICE_X9Y113_AO5),
.O6(CLBLM_R_X7Y113_SLICE_X9Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y114_SLICE_X8Y114_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y114_SLICE_X8Y114_DO5),
.O6(CLBLM_R_X7Y114_SLICE_X8Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h1705ff775f17ff77)
  ) CLBLM_R_X7Y114_SLICE_X8Y114_CLUT (
.I0(CLBLM_R_X7Y114_SLICE_X8Y114_AO6),
.I1(CLBLM_R_X7Y112_SLICE_X9Y112_AO6),
.I2(LIOB33_X0Y113_IOB_X0Y113_I),
.I3(CLBLM_L_X8Y113_SLICE_X11Y113_BO6),
.I4(RIOB33_X105Y101_IOB_X1Y102_I),
.I5(LIOB33_X0Y111_IOB_X0Y112_I),
.O5(CLBLM_R_X7Y114_SLICE_X8Y114_CO5),
.O6(CLBLM_R_X7Y114_SLICE_X8Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h9aa559aa65a5a6aa)
  ) CLBLM_R_X7Y114_SLICE_X8Y114_BLUT (
.I0(CLBLM_R_X7Y112_SLICE_X9Y112_DO6),
.I1(RIOB33_X105Y101_IOB_X1Y102_I),
.I2(CLBLM_L_X8Y113_SLICE_X11Y113_BO6),
.I3(LIOB33_X0Y111_IOB_X0Y112_I),
.I4(CLBLM_R_X7Y112_SLICE_X9Y112_AO6),
.I5(RIOB33_X105Y103_IOB_X1Y103_I),
.O5(CLBLM_R_X7Y114_SLICE_X8Y114_BO5),
.O6(CLBLM_R_X7Y114_SLICE_X8Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa555555c3c33333)
  ) CLBLM_R_X7Y114_SLICE_X8Y114_ALUT (
.I0(CLBLM_R_X7Y112_SLICE_X9Y112_DO6),
.I1(CLBLM_R_X7Y111_SLICE_X8Y111_CO6),
.I2(RIOB33_X105Y103_IOB_X1Y104_I),
.I3(RIOB33_X105Y103_IOB_X1Y103_I),
.I4(LIOB33_X0Y111_IOB_X0Y112_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y114_SLICE_X8Y114_AO5),
.O6(CLBLM_R_X7Y114_SLICE_X8Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h93933333c9c99999)
  ) CLBLM_R_X7Y114_SLICE_X9Y114_DLUT (
.I0(CLBLM_R_X7Y112_SLICE_X9Y112_BO6),
.I1(CLBLM_R_X7Y114_SLICE_X8Y114_AO5),
.I2(LIOB33_X0Y111_IOB_X0Y112_I),
.I3(1'b1),
.I4(RIOB33_X105Y103_IOB_X1Y103_I),
.I5(CLBLM_R_X7Y112_SLICE_X9Y112_AO5),
.O5(CLBLM_R_X7Y114_SLICE_X9Y114_DO5),
.O6(CLBLM_R_X7Y114_SLICE_X9Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h17033f17ff77ff77)
  ) CLBLM_R_X7Y114_SLICE_X9Y114_CLUT (
.I0(CLBLM_R_X7Y112_SLICE_X9Y112_BO6),
.I1(CLBLM_R_X7Y114_SLICE_X8Y114_AO5),
.I2(LIOB33_X0Y113_IOB_X0Y113_I),
.I3(CLBLM_R_X7Y112_SLICE_X9Y112_AO5),
.I4(LIOB33_X0Y111_IOB_X0Y112_I),
.I5(RIOB33_X105Y103_IOB_X1Y103_I),
.O5(CLBLM_R_X7Y114_SLICE_X9Y114_CO5),
.O6(CLBLM_R_X7Y114_SLICE_X9Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h157fffff01570fff)
  ) CLBLM_R_X7Y114_SLICE_X9Y114_BLUT (
.I0(LIOB33_X0Y113_IOB_X0Y113_I),
.I1(LIOB33_X0Y111_IOB_X0Y112_I),
.I2(CLBLM_L_X8Y113_SLICE_X11Y113_AO6),
.I3(CLBLM_L_X8Y114_SLICE_X10Y114_AO6),
.I4(RIOB33_X105Y101_IOB_X1Y101_I),
.I5(CLBLM_L_X8Y114_SLICE_X11Y114_DO6),
.O5(CLBLM_R_X7Y114_SLICE_X9Y114_BO5),
.O6(CLBLM_R_X7Y114_SLICE_X9Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333ffffd42b50af)
  ) CLBLM_R_X7Y114_SLICE_X9Y114_ALUT (
.I0(CLBLM_L_X8Y114_SLICE_X11Y114_DO6),
.I1(LIOB33_X0Y111_IOB_X0Y112_I),
.I2(CLBLM_L_X8Y113_SLICE_X11Y113_AO6),
.I3(CLBLM_L_X8Y114_SLICE_X10Y114_AO6),
.I4(RIOB33_X105Y101_IOB_X1Y101_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y114_SLICE_X9Y114_AO5),
.O6(CLBLM_R_X7Y114_SLICE_X9Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y115_SLICE_X8Y115_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y115_SLICE_X8Y115_DO5),
.O6(CLBLM_R_X7Y115_SLICE_X8Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y115_SLICE_X8Y115_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y115_SLICE_X8Y115_CO5),
.O6(CLBLM_R_X7Y115_SLICE_X8Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y115_SLICE_X8Y115_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y115_SLICE_X8Y115_BO5),
.O6(CLBLM_R_X7Y115_SLICE_X8Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc69c6c366696cc3c)
  ) CLBLM_R_X7Y115_SLICE_X8Y115_ALUT (
.I0(LIOB33_X0Y111_IOB_X0Y112_I),
.I1(CLBLM_L_X8Y115_SLICE_X10Y115_BO6),
.I2(CLBLM_R_X7Y115_SLICE_X9Y115_AO6),
.I3(CLBLM_R_X7Y113_SLICE_X8Y113_BO6),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(LIOB33_X0Y115_IOB_X0Y116_I),
.O5(CLBLM_R_X7Y115_SLICE_X8Y115_AO5),
.O6(CLBLM_R_X7Y115_SLICE_X8Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y115_SLICE_X9Y115_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y115_SLICE_X9Y115_DO5),
.O6(CLBLM_R_X7Y115_SLICE_X9Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y115_SLICE_X9Y115_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y115_SLICE_X9Y115_CO5),
.O6(CLBLM_R_X7Y115_SLICE_X9Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y115_SLICE_X9Y115_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y115_SLICE_X9Y115_BO5),
.O6(CLBLM_R_X7Y115_SLICE_X9Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996c33c996633cc)
  ) CLBLM_R_X7Y115_SLICE_X9Y115_ALUT (
.I0(RIOB33_X105Y101_IOB_X1Y101_I),
.I1(CLBLM_L_X10Y114_SLICE_X12Y114_DO6),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(CLBLM_L_X8Y114_SLICE_X11Y114_AO6),
.I4(LIOB33_X0Y109_IOB_X0Y110_I),
.I5(LIOB33_X0Y111_IOB_X0Y111_I),
.O5(CLBLM_R_X7Y115_SLICE_X9Y115_AO5),
.O6(CLBLM_R_X7Y115_SLICE_X9Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h9666aaaa999655aa)
  ) CLBLM_R_X7Y116_SLICE_X8Y116_DLUT (
.I0(CLBLM_L_X8Y115_SLICE_X10Y115_DO6),
.I1(LIOB33_X0Y113_IOB_X0Y113_I),
.I2(LIOB33_X0Y111_IOB_X0Y112_I),
.I3(CLBLM_R_X7Y115_SLICE_X9Y115_AO6),
.I4(LIOB33_X0Y115_IOB_X0Y116_I),
.I5(CLBLM_R_X7Y113_SLICE_X8Y113_BO6),
.O5(CLBLM_R_X7Y116_SLICE_X8Y116_DO5),
.O6(CLBLM_R_X7Y116_SLICE_X8Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7f15ff3fd540ffc0)
  ) CLBLM_R_X7Y116_SLICE_X8Y116_CLUT (
.I0(LIOB33_X0Y115_IOB_X0Y115_I),
.I1(LIOB33_X0Y113_IOB_X0Y113_I),
.I2(RIOB33_X105Y101_IOB_X1Y101_I),
.I3(CLBLM_R_X7Y116_SLICE_X9Y116_BO6),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(CLBLM_R_X7Y114_SLICE_X9Y114_AO5),
.O5(CLBLM_R_X7Y116_SLICE_X8Y116_CO5),
.O6(CLBLM_R_X7Y116_SLICE_X8Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7887887787787788)
  ) CLBLM_R_X7Y116_SLICE_X8Y116_BLUT (
.I0(LIOB33_X0Y113_IOB_X0Y113_I),
.I1(RIOB33_X105Y101_IOB_X1Y101_I),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(CLBLM_R_X7Y114_SLICE_X9Y114_AO5),
.I4(LIOB33_X0Y115_IOB_X0Y115_I),
.I5(CLBLM_R_X7Y116_SLICE_X9Y116_BO6),
.O5(CLBLM_R_X7Y116_SLICE_X8Y116_BO5),
.O6(CLBLM_R_X7Y116_SLICE_X8Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h054d4d5fcfcfffff)
  ) CLBLM_R_X7Y116_SLICE_X8Y116_ALUT (
.I0(LIOB33_X0Y113_IOB_X0Y113_I),
.I1(CLBLM_R_X7Y113_SLICE_X8Y113_BO6),
.I2(CLBLM_L_X8Y115_SLICE_X10Y115_DO6),
.I3(LIOB33_X0Y111_IOB_X0Y112_I),
.I4(CLBLM_R_X7Y115_SLICE_X9Y115_AO6),
.I5(LIOB33_X0Y115_IOB_X0Y116_I),
.O5(CLBLM_R_X7Y116_SLICE_X8Y116_AO5),
.O6(CLBLM_R_X7Y116_SLICE_X8Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y116_SLICE_X9Y116_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y116_SLICE_X9Y116_DO5),
.O6(CLBLM_R_X7Y116_SLICE_X9Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h87e1ff55781e00aa)
  ) CLBLM_R_X7Y116_SLICE_X9Y116_CLUT (
.I0(CLBLM_L_X8Y114_SLICE_X11Y114_CO6),
.I1(LIOB33_X0Y111_IOB_X0Y112_I),
.I2(LIOB33_X0Y113_IOB_X0Y113_I),
.I3(CLBLM_L_X8Y115_SLICE_X10Y115_CO6),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(CLBLM_L_X8Y116_SLICE_X10Y116_CO6),
.O5(CLBLM_R_X7Y116_SLICE_X9Y116_CO5),
.O6(CLBLM_R_X7Y116_SLICE_X9Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h4cdfdf4cdfdf4c4c)
  ) CLBLM_R_X7Y116_SLICE_X9Y116_BLUT (
.I0(LIOB33_X0Y113_IOB_X0Y113_I),
.I1(CLBLM_L_X8Y115_SLICE_X10Y115_AO5),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(RIOB33_X105Y101_IOB_X1Y101_I),
.I4(CLBLM_L_X8Y116_SLICE_X10Y116_BO6),
.I5(LIOB33_X0Y111_IOB_X0Y112_I),
.O5(CLBLM_R_X7Y116_SLICE_X9Y116_BO5),
.O6(CLBLM_R_X7Y116_SLICE_X9Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hb74877888877b748)
  ) CLBLM_R_X7Y116_SLICE_X9Y116_ALUT (
.I0(RIOB33_X105Y101_IOB_X1Y101_I),
.I1(LIOB33_X0Y111_IOB_X0Y112_I),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(CLBLM_L_X8Y116_SLICE_X10Y116_BO6),
.I4(CLBLM_L_X8Y114_SLICE_X11Y114_CO6),
.I5(CLBLM_L_X8Y115_SLICE_X10Y115_CO6),
.O5(CLBLM_R_X7Y116_SLICE_X9Y116_AO5),
.O6(CLBLM_R_X7Y116_SLICE_X9Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h33ccc639cc3339c6)
  ) CLBLM_R_X11Y105_SLICE_X14Y105_DLUT (
.I0(CLBLM_R_X7Y109_SLICE_X9Y109_AO6),
.I1(CLBLM_R_X11Y105_SLICE_X15Y105_AO5),
.I2(CLBLM_R_X11Y107_SLICE_X14Y107_DO6),
.I3(CLBLM_R_X11Y106_SLICE_X14Y106_AO6),
.I4(CLBLM_L_X12Y105_SLICE_X16Y105_DO6),
.I5(CLBLM_L_X12Y105_SLICE_X16Y105_CO6),
.O5(CLBLM_R_X11Y105_SLICE_X14Y105_DO5),
.O6(CLBLM_R_X11Y105_SLICE_X14Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcc0fec8f330fb32)
  ) CLBLM_R_X11Y105_SLICE_X14Y105_CLUT (
.I0(CLBLM_R_X7Y109_SLICE_X9Y109_AO6),
.I1(CLBLM_R_X11Y105_SLICE_X15Y105_AO5),
.I2(CLBLM_L_X12Y105_SLICE_X16Y105_DO6),
.I3(CLBLM_R_X11Y106_SLICE_X14Y106_AO6),
.I4(CLBLM_R_X11Y107_SLICE_X14Y107_DO6),
.I5(CLBLM_L_X12Y105_SLICE_X16Y105_CO6),
.O5(CLBLM_R_X11Y105_SLICE_X14Y105_CO5),
.O6(CLBLM_R_X11Y105_SLICE_X14Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6665ccff999a3300)
  ) CLBLM_R_X11Y105_SLICE_X14Y105_BLUT (
.I0(LIOB33_X0Y101_IOB_X0Y102_I),
.I1(CLBLM_R_X11Y105_SLICE_X15Y105_DO6),
.I2(LIOB33_X0Y101_IOB_X0Y101_I),
.I3(CLBLM_L_X12Y105_SLICE_X16Y105_CO6),
.I4(RIOB33_X105Y109_IOB_X1Y109_I),
.I5(CLBLM_L_X10Y105_SLICE_X13Y105_DO6),
.O5(CLBLM_R_X11Y105_SLICE_X14Y105_BO5),
.O6(CLBLM_R_X11Y105_SLICE_X14Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h4445ccffdddfffff)
  ) CLBLM_R_X11Y105_SLICE_X14Y105_ALUT (
.I0(LIOB33_X0Y101_IOB_X0Y102_I),
.I1(CLBLM_R_X11Y105_SLICE_X15Y105_DO6),
.I2(LIOB33_X0Y101_IOB_X0Y101_I),
.I3(CLBLM_L_X12Y105_SLICE_X16Y105_CO6),
.I4(RIOB33_X105Y109_IOB_X1Y109_I),
.I5(CLBLM_L_X10Y105_SLICE_X13Y105_DO6),
.O5(CLBLM_R_X11Y105_SLICE_X14Y105_AO5),
.O6(CLBLM_R_X11Y105_SLICE_X14Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0110affb31111ff)
  ) CLBLM_R_X11Y105_SLICE_X15Y105_DLUT (
.I0(RIOB33_X105Y109_IOB_X1Y110_I),
.I1(RIOB33_X105Y109_IOB_X1Y109_I),
.I2(RIOB33_X105Y111_IOB_X1Y112_I),
.I3(RIOB33_X105Y113_IOB_X1Y113_I),
.I4(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I5(RIOB33_X105Y111_IOB_X1Y111_I),
.O5(CLBLM_R_X11Y105_SLICE_X15Y105_DO5),
.O6(CLBLM_R_X11Y105_SLICE_X15Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h87f0e15a78f01e5a)
  ) CLBLM_R_X11Y105_SLICE_X15Y105_CLUT (
.I0(CLBLM_R_X11Y105_SLICE_X15Y105_AO6),
.I1(LIOB33_X0Y101_IOB_X0Y102_I),
.I2(CLBLM_R_X11Y105_SLICE_X14Y105_BO6),
.I3(RIOB33_X105Y107_IOB_X1Y108_I),
.I4(CLBLM_L_X12Y105_SLICE_X16Y105_AO5),
.I5(LIOB33_X0Y103_IOB_X0Y104_I),
.O5(CLBLM_R_X11Y105_SLICE_X15Y105_CO5),
.O6(CLBLM_R_X11Y105_SLICE_X15Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h023b23bfbbbbffff)
  ) CLBLM_R_X11Y105_SLICE_X15Y105_BLUT (
.I0(CLBLM_L_X12Y105_SLICE_X16Y105_AO5),
.I1(CLBLM_R_X11Y105_SLICE_X14Y105_BO6),
.I2(LIOB33_X0Y101_IOB_X0Y102_I),
.I3(LIOB33_X0Y103_IOB_X0Y104_I),
.I4(CLBLM_R_X11Y105_SLICE_X15Y105_AO6),
.I5(RIOB33_X105Y107_IOB_X1Y108_I),
.O5(CLBLM_R_X11Y105_SLICE_X15Y105_BO5),
.O6(CLBLM_R_X11Y105_SLICE_X15Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc333c3330fff0fff)
  ) CLBLM_R_X11Y105_SLICE_X15Y105_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X12Y105_SLICE_X16Y105_CO6),
.I2(LIOB33_X0Y101_IOB_X0Y101_I),
.I3(RIOB33_X105Y109_IOB_X1Y109_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y105_SLICE_X15Y105_AO5),
.O6(CLBLM_R_X11Y105_SLICE_X15Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5aa55aa5a55a6996)
  ) CLBLM_R_X11Y106_SLICE_X14Y106_DLUT (
.I0(CLBLM_R_X7Y109_SLICE_X9Y109_AO6),
.I1(CLBLM_R_X11Y106_SLICE_X15Y106_AO5),
.I2(CLBLM_R_X11Y107_SLICE_X14Y107_DO6),
.I3(CLBLM_R_X11Y106_SLICE_X14Y106_AO5),
.I4(CLBLM_L_X12Y107_SLICE_X17Y107_AO6),
.I5(CLBLM_L_X12Y106_SLICE_X16Y106_BO6),
.O5(CLBLM_R_X11Y106_SLICE_X14Y106_DO5),
.O6(CLBLM_R_X11Y106_SLICE_X14Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffa5ffa5a500ed84)
  ) CLBLM_R_X11Y106_SLICE_X14Y106_CLUT (
.I0(CLBLM_R_X7Y109_SLICE_X9Y109_AO6),
.I1(CLBLM_R_X11Y106_SLICE_X15Y106_AO5),
.I2(CLBLM_R_X11Y107_SLICE_X14Y107_DO6),
.I3(CLBLM_R_X11Y106_SLICE_X14Y106_AO5),
.I4(CLBLM_L_X12Y107_SLICE_X17Y107_AO6),
.I5(CLBLM_L_X12Y106_SLICE_X16Y106_BO6),
.O5(CLBLM_R_X11Y106_SLICE_X14Y106_CO5),
.O6(CLBLM_R_X11Y106_SLICE_X14Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h39c6c6399c63639c)
  ) CLBLM_R_X11Y106_SLICE_X14Y106_BLUT (
.I0(CLBLM_R_X11Y105_SLICE_X14Y105_DO6),
.I1(CLBLM_R_X11Y105_SLICE_X14Y105_CO6),
.I2(CLBLM_R_X11Y106_SLICE_X15Y106_AO6),
.I3(CLBLM_L_X10Y105_SLICE_X13Y105_AO5),
.I4(CLBLM_R_X11Y105_SLICE_X14Y105_BO6),
.I5(CLBLM_R_X11Y106_SLICE_X14Y106_CO6),
.O5(CLBLM_R_X11Y106_SLICE_X14Y106_BO5),
.O6(CLBLM_R_X11Y106_SLICE_X14Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333ffff3f3f3f3f)
  ) CLBLM_R_X11Y106_SLICE_X14Y106_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y101_IOB_X0Y102_I),
.I2(RIOB33_X105Y107_IOB_X1Y107_I),
.I3(1'b1),
.I4(RIOB33_X105Y107_IOB_X1Y108_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y106_SLICE_X14Y106_AO5),
.O6(CLBLM_R_X11Y106_SLICE_X14Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6699966996699966)
  ) CLBLM_R_X11Y106_SLICE_X15Y106_DLUT (
.I0(CLBLM_R_X11Y106_SLICE_X15Y106_AO6),
.I1(CLBLM_R_X11Y106_SLICE_X14Y106_CO6),
.I2(CLBLM_R_X11Y106_SLICE_X14Y106_DO6),
.I3(CLBLM_R_X11Y105_SLICE_X14Y105_DO6),
.I4(CLBLM_L_X12Y108_SLICE_X17Y108_AO5),
.I5(CLBLM_R_X11Y107_SLICE_X15Y107_BO6),
.O5(CLBLM_R_X11Y106_SLICE_X15Y106_DO5),
.O6(CLBLM_R_X11Y106_SLICE_X15Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6c939393936c6c6c)
  ) CLBLM_R_X11Y106_SLICE_X15Y106_CLUT (
.I0(RIOB33_X105Y107_IOB_X1Y107_I),
.I1(CLBLM_R_X11Y106_SLICE_X14Y106_CO6),
.I2(LIOB33_X0Y103_IOB_X0Y104_I),
.I3(LIOB33_X0Y101_IOB_X0Y102_I),
.I4(RIOB33_X105Y107_IOB_X1Y108_I),
.I5(CLBLM_L_X12Y105_SLICE_X16Y105_BO6),
.O5(CLBLM_R_X11Y106_SLICE_X15Y106_CO5),
.O6(CLBLM_R_X11Y106_SLICE_X15Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7d14ff3cdd44ffcc)
  ) CLBLM_R_X11Y106_SLICE_X15Y106_BLUT (
.I0(LIOB33_X0Y103_IOB_X0Y104_I),
.I1(CLBLM_L_X12Y105_SLICE_X16Y105_BO6),
.I2(RIOB33_X105Y107_IOB_X1Y108_I),
.I3(CLBLM_R_X11Y106_SLICE_X14Y106_CO6),
.I4(RIOB33_X105Y107_IOB_X1Y107_I),
.I5(LIOB33_X0Y101_IOB_X0Y102_I),
.O5(CLBLM_R_X11Y106_SLICE_X15Y106_BO5),
.O6(CLBLM_R_X11Y106_SLICE_X15Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h55ff55ff0fff0fff)
  ) CLBLM_R_X11Y106_SLICE_X15Y106_ALUT (
.I0(LIOB33_X0Y103_IOB_X0Y104_I),
.I1(1'b1),
.I2(LIOB33_X0Y101_IOB_X0Y101_I),
.I3(RIOB33_X105Y107_IOB_X1Y107_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y106_SLICE_X15Y106_AO5),
.O6(CLBLM_R_X11Y106_SLICE_X15Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h043f73c08c0c8cc0)
  ) CLBLM_R_X11Y107_SLICE_X14Y107_DLUT (
.I0(RIOB33_X105Y111_IOB_X1Y112_I),
.I1(RIOB33_X105Y113_IOB_X1Y113_I),
.I2(RIOB33_X105Y109_IOB_X1Y110_I),
.I3(RIOB33_X105Y109_IOB_X1Y109_I),
.I4(RIOB33_X105Y107_IOB_X1Y108_I),
.I5(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.O5(CLBLM_R_X11Y107_SLICE_X14Y107_DO5),
.O6(CLBLM_R_X11Y107_SLICE_X14Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcc0f330fec8fb32)
  ) CLBLM_R_X11Y107_SLICE_X14Y107_CLUT (
.I0(CLBLM_R_X11Y107_SLICE_X14Y107_AO6),
.I1(CLBLM_R_X11Y107_SLICE_X15Y107_AO6),
.I2(CLBLM_R_X11Y108_SLICE_X14Y108_BO6),
.I3(CLBLM_R_X11Y107_SLICE_X14Y107_AO5),
.I4(CLBLM_L_X12Y107_SLICE_X17Y107_BO6),
.I5(CLBLM_L_X10Y108_SLICE_X12Y108_DO6),
.O5(CLBLM_R_X11Y107_SLICE_X14Y107_CO5),
.O6(CLBLM_R_X11Y107_SLICE_X14Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h693c696996c39696)
  ) CLBLM_R_X11Y107_SLICE_X14Y107_BLUT (
.I0(CLBLM_R_X11Y108_SLICE_X14Y108_BO6),
.I1(CLBLM_L_X12Y107_SLICE_X17Y107_BO6),
.I2(CLBLM_R_X11Y107_SLICE_X15Y107_AO6),
.I3(CLBLM_L_X10Y108_SLICE_X12Y108_DO6),
.I4(CLBLM_R_X11Y107_SLICE_X14Y107_AO6),
.I5(CLBLM_R_X11Y107_SLICE_X14Y107_AO5),
.O5(CLBLM_R_X11Y107_SLICE_X14Y107_BO5),
.O6(CLBLM_R_X11Y107_SLICE_X14Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0fff0fff55ff55ff)
  ) CLBLM_R_X11Y107_SLICE_X14Y107_ALUT (
.I0(LIOB33_X0Y101_IOB_X0Y102_I),
.I1(1'b1),
.I2(LIOB33_X0Y101_IOB_X0Y101_I),
.I3(RIOB33_X105Y103_IOB_X1Y104_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y107_SLICE_X14Y107_AO5),
.O6(CLBLM_R_X11Y107_SLICE_X14Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6699669996699966)
  ) CLBLM_R_X11Y107_SLICE_X15Y107_DLUT (
.I0(CLBLM_L_X12Y107_SLICE_X17Y107_AO6),
.I1(CLBLM_R_X11Y106_SLICE_X15Y106_AO5),
.I2(CLBLM_L_X12Y107_SLICE_X17Y107_BO6),
.I3(CLBLM_R_X11Y107_SLICE_X15Y107_AO5),
.I4(CLBLM_R_X11Y107_SLICE_X15Y107_AO6),
.I5(CLBLM_L_X12Y107_SLICE_X16Y107_CO6),
.O5(CLBLM_R_X11Y107_SLICE_X15Y107_DO5),
.O6(CLBLM_R_X11Y107_SLICE_X15Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h32ddcdddcd223222)
  ) CLBLM_R_X11Y107_SLICE_X15Y107_CLUT (
.I0(CLBLM_L_X12Y107_SLICE_X17Y107_BO6),
.I1(CLBLM_L_X12Y107_SLICE_X16Y107_CO6),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(LIOB33_X0Y101_IOB_X0Y101_I),
.I4(RIOB33_X105Y107_IOB_X1Y107_I),
.I5(CLBLM_L_X12Y107_SLICE_X17Y107_AO6),
.O5(CLBLM_R_X11Y107_SLICE_X15Y107_CO5),
.O6(CLBLM_R_X11Y107_SLICE_X15Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffc3ffebc300c382)
  ) CLBLM_R_X11Y107_SLICE_X15Y107_BLUT (
.I0(CLBLM_R_X11Y107_SLICE_X15Y107_AO6),
.I1(CLBLM_L_X12Y107_SLICE_X17Y107_AO6),
.I2(CLBLM_R_X11Y106_SLICE_X15Y106_AO5),
.I3(CLBLM_L_X12Y107_SLICE_X16Y107_CO6),
.I4(CLBLM_L_X12Y107_SLICE_X17Y107_BO6),
.I5(CLBLM_R_X11Y107_SLICE_X15Y107_AO5),
.O5(CLBLM_R_X11Y107_SLICE_X15Y107_BO5),
.O6(CLBLM_R_X11Y107_SLICE_X15Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0fff0fff55ff55ff)
  ) CLBLM_R_X11Y107_SLICE_X15Y107_ALUT (
.I0(LIOB33_X0Y101_IOB_X0Y102_I),
.I1(1'b1),
.I2(LIOB33_X0Y101_IOB_X0Y101_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y107_SLICE_X15Y107_AO5),
.O6(CLBLM_R_X11Y107_SLICE_X15Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hbd4239c6718ef50a)
  ) CLBLM_R_X11Y108_SLICE_X14Y108_DLUT (
.I0(CLBLM_R_X11Y108_SLICE_X14Y108_AO6),
.I1(LIOB33_X0Y101_IOB_X0Y102_I),
.I2(CLBLM_L_X10Y108_SLICE_X12Y108_AO5),
.I3(CLBLM_R_X11Y108_SLICE_X14Y108_CO6),
.I4(RIOB33_X105Y103_IOB_X1Y103_I),
.I5(RIOB33_X105Y103_IOB_X1Y104_I),
.O5(CLBLM_R_X11Y108_SLICE_X14Y108_DO5),
.O6(CLBLM_R_X11Y108_SLICE_X14Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h66aa66aa995a965a)
  ) CLBLM_R_X11Y108_SLICE_X14Y108_CLUT (
.I0(CLBLM_L_X12Y107_SLICE_X17Y107_BO6),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_L_X10Y108_SLICE_X12Y108_DO6),
.I3(LIOB33_X0Y101_IOB_X0Y101_I),
.I4(RIOB33_X105Y103_IOB_X1Y104_I),
.I5(CLBLM_R_X11Y108_SLICE_X14Y108_BO6),
.O5(CLBLM_R_X11Y108_SLICE_X14Y108_CO5),
.O6(CLBLM_R_X11Y108_SLICE_X14Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f50440043504400)
  ) CLBLM_R_X11Y108_SLICE_X14Y108_BLUT (
.I0(RIOB33_X105Y103_IOB_X1Y104_I),
.I1(RIOB33_X105Y107_IOB_X1Y107_I),
.I2(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I3(RIOB33_X105Y113_IOB_X1Y113_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(RIOB33_X105Y111_IOB_X1Y112_I),
.O5(CLBLM_R_X11Y108_SLICE_X14Y108_BO5),
.O6(CLBLM_R_X11Y108_SLICE_X14Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h95959595ff15ff15)
  ) CLBLM_R_X11Y108_SLICE_X14Y108_ALUT (
.I0(CLBLM_L_X10Y108_SLICE_X12Y108_DO6),
.I1(RIOB33_X105Y103_IOB_X1Y104_I),
.I2(LIOB33_X0Y101_IOB_X0Y101_I),
.I3(CLBLM_R_X11Y108_SLICE_X14Y108_BO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y108_SLICE_X14Y108_AO5),
.O6(CLBLM_R_X11Y108_SLICE_X14Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha59969aa69995aaa)
  ) CLBLM_R_X11Y108_SLICE_X15Y108_DLUT (
.I0(CLBLM_R_X11Y107_SLICE_X15Y107_CO6),
.I1(CLBLM_R_X11Y108_SLICE_X14Y108_AO5),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(LIOB33_X0Y101_IOB_X0Y102_I),
.I4(CLBLM_L_X12Y107_SLICE_X16Y107_AO6),
.I5(RIOB33_X105Y103_IOB_X1Y104_I),
.O5(CLBLM_R_X11Y108_SLICE_X15Y108_DO5),
.O6(CLBLM_R_X11Y108_SLICE_X15Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h78871ee18778e11e)
  ) CLBLM_R_X11Y108_SLICE_X15Y108_CLUT (
.I0(CLBLM_L_X12Y108_SLICE_X16Y108_BO5),
.I1(CLBLM_R_X11Y107_SLICE_X14Y107_CO6),
.I2(CLBLM_R_X11Y106_SLICE_X14Y106_DO6),
.I3(CLBLM_L_X12Y108_SLICE_X17Y108_AO5),
.I4(CLBLM_R_X11Y107_SLICE_X15Y107_DO6),
.I5(CLBLM_R_X11Y107_SLICE_X15Y107_BO6),
.O5(CLBLM_R_X11Y108_SLICE_X15Y108_CO5),
.O6(CLBLM_R_X11Y108_SLICE_X15Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h59a69a65a659659a)
  ) CLBLM_R_X11Y108_SLICE_X15Y108_BLUT (
.I0(CLBLM_R_X11Y107_SLICE_X15Y107_DO6),
.I1(CLBLM_R_X11Y107_SLICE_X14Y107_BO6),
.I2(CLBLM_L_X10Y108_SLICE_X13Y108_DO6),
.I3(CLBLM_L_X12Y108_SLICE_X16Y108_BO5),
.I4(CLBLM_R_X11Y108_SLICE_X15Y108_AO6),
.I5(CLBLM_R_X11Y107_SLICE_X14Y107_CO6),
.O5(CLBLM_R_X11Y108_SLICE_X15Y108_BO5),
.O6(CLBLM_R_X11Y108_SLICE_X15Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h33ff33ff0fff0fff)
  ) CLBLM_R_X11Y108_SLICE_X15Y108_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y103_IOB_X0Y104_I),
.I2(LIOB33_X0Y105_IOB_X0Y105_I),
.I3(RIOB33_X105Y103_IOB_X1Y103_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y108_SLICE_X15Y108_AO5),
.O6(CLBLM_R_X11Y108_SLICE_X15Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h788787781ee1e11e)
  ) CLBLM_R_X11Y109_SLICE_X14Y109_DLUT (
.I0(CLBLM_R_X11Y106_SLICE_X15Y106_BO6),
.I1(CLBLM_R_X11Y109_SLICE_X15Y109_AO5),
.I2(CLBLM_R_X11Y109_SLICE_X15Y109_AO6),
.I3(CLBLM_L_X10Y106_SLICE_X13Y106_AO5),
.I4(CLBLM_L_X10Y105_SLICE_X13Y105_CO6),
.I5(CLBLM_R_X11Y105_SLICE_X15Y105_CO6),
.O5(CLBLM_R_X11Y109_SLICE_X14Y109_DO5),
.O6(CLBLM_R_X11Y109_SLICE_X14Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'he27b6a3f1d8495c0)
  ) CLBLM_R_X11Y109_SLICE_X14Y109_CLUT (
.I0(CLBLM_R_X11Y106_SLICE_X15Y106_BO6),
.I1(LIOB33_X0Y105_IOB_X0Y105_I),
.I2(RIOB33_X105Y107_IOB_X1Y108_I),
.I3(CLBLM_R_X11Y105_SLICE_X15Y105_CO6),
.I4(RIOB33_X105Y107_IOB_X1Y107_I),
.I5(CLBLM_L_X10Y105_SLICE_X13Y105_CO6),
.O5(CLBLM_R_X11Y109_SLICE_X14Y109_CO5),
.O6(CLBLM_R_X11Y109_SLICE_X14Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbb0f220b0fb20f2)
  ) CLBLM_R_X11Y109_SLICE_X14Y109_BLUT (
.I0(CLBLM_R_X11Y109_SLICE_X15Y109_AO5),
.I1(CLBLM_R_X11Y105_SLICE_X15Y105_CO6),
.I2(CLBLM_R_X11Y109_SLICE_X15Y109_AO6),
.I3(CLBLM_L_X10Y106_SLICE_X13Y106_AO5),
.I4(CLBLM_R_X11Y106_SLICE_X15Y106_BO6),
.I5(CLBLM_L_X10Y105_SLICE_X13Y105_CO6),
.O5(CLBLM_R_X11Y109_SLICE_X14Y109_BO5),
.O6(CLBLM_R_X11Y109_SLICE_X14Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h7171f3f36969c3c3)
  ) CLBLM_R_X11Y109_SLICE_X14Y109_ALUT (
.I0(RIOB33_X105Y107_IOB_X1Y107_I),
.I1(CLBLM_R_X11Y105_SLICE_X15Y105_CO6),
.I2(CLBLM_R_X11Y106_SLICE_X15Y106_BO6),
.I3(1'b1),
.I4(LIOB33_X0Y105_IOB_X0Y105_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y109_SLICE_X14Y109_AO5),
.O6(CLBLM_R_X11Y109_SLICE_X14Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h2dd2b44bd22d4bb4)
  ) CLBLM_R_X11Y109_SLICE_X15Y109_DLUT (
.I0(CLBLM_R_X13Y108_SLICE_X18Y108_DO6),
.I1(CLBLM_L_X12Y109_SLICE_X17Y109_BO6),
.I2(CLBLM_R_X11Y109_SLICE_X14Y109_DO6),
.I3(CLBLM_R_X13Y108_SLICE_X18Y108_CO6),
.I4(CLBLM_L_X12Y109_SLICE_X17Y109_AO5),
.I5(CLBLM_L_X12Y109_SLICE_X16Y109_AO5),
.O5(CLBLM_R_X11Y109_SLICE_X15Y109_DO5),
.O6(CLBLM_R_X11Y109_SLICE_X15Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996969669696996)
  ) CLBLM_R_X11Y109_SLICE_X15Y109_CLUT (
.I0(CLBLM_R_X13Y108_SLICE_X18Y108_DO6),
.I1(CLBLM_L_X12Y109_SLICE_X17Y109_BO6),
.I2(CLBLM_L_X12Y109_SLICE_X17Y109_AO5),
.I3(CLBLM_R_X11Y110_SLICE_X14Y110_AO5),
.I4(CLBLM_L_X12Y109_SLICE_X16Y109_CO6),
.I5(CLBLM_L_X12Y109_SLICE_X17Y109_CO6),
.O5(CLBLM_R_X11Y109_SLICE_X15Y109_CO5),
.O6(CLBLM_R_X11Y109_SLICE_X15Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h9f605fa0a35c936c)
  ) CLBLM_R_X11Y109_SLICE_X15Y109_BLUT (
.I0(RIOB33_X105Y103_IOB_X1Y103_I),
.I1(CLBLM_R_X13Y108_SLICE_X19Y108_AO6),
.I2(LIOB33_X0Y105_IOB_X0Y105_I),
.I3(CLBLM_R_X11Y108_SLICE_X15Y108_BO6),
.I4(RIOB33_X105Y101_IOB_X1Y102_I),
.I5(CLBLM_L_X10Y107_SLICE_X13Y107_AO6),
.O5(CLBLM_R_X11Y109_SLICE_X15Y109_BO5),
.O6(CLBLM_R_X11Y109_SLICE_X15Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h33ff33ff0fff0fff)
  ) CLBLM_R_X11Y109_SLICE_X15Y109_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y105_IOB_X0Y106_I),
.I2(LIOB33_X0Y105_IOB_X0Y105_I),
.I3(RIOB33_X105Y107_IOB_X1Y107_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y109_SLICE_X15Y109_AO5),
.O6(CLBLM_R_X11Y109_SLICE_X15Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h39c69c63c639639c)
  ) CLBLM_R_X11Y110_SLICE_X14Y110_DLUT (
.I0(CLBLM_L_X12Y109_SLICE_X16Y109_BO6),
.I1(CLBLM_L_X12Y109_SLICE_X17Y109_CO6),
.I2(CLBLM_R_X11Y110_SLICE_X15Y110_BO6),
.I3(CLBLM_R_X11Y110_SLICE_X14Y110_AO5),
.I4(CLBLM_R_X11Y110_SLICE_X14Y110_BO5),
.I5(CLBLM_L_X12Y109_SLICE_X16Y109_CO6),
.O5(CLBLM_R_X11Y110_SLICE_X14Y110_DO5),
.O6(CLBLM_R_X11Y110_SLICE_X14Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5a96a56996a5695a)
  ) CLBLM_R_X11Y110_SLICE_X14Y110_CLUT (
.I0(CLBLM_L_X12Y109_SLICE_X16Y109_BO6),
.I1(CLBLM_R_X11Y110_SLICE_X15Y110_AO6),
.I2(CLBLM_R_X11Y110_SLICE_X15Y110_BO6),
.I3(CLBLM_R_X11Y110_SLICE_X14Y110_AO6),
.I4(CLBLM_R_X11Y110_SLICE_X14Y110_BO5),
.I5(CLBLM_L_X10Y108_SLICE_X12Y108_CO6),
.O5(CLBLM_R_X11Y110_SLICE_X14Y110_CO5),
.O6(CLBLM_R_X11Y110_SLICE_X14Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h33ff33ff0fff0fff)
  ) CLBLM_R_X11Y110_SLICE_X14Y110_BLUT (
.I0(1'b1),
.I1(LIOB33_X0Y105_IOB_X0Y106_I),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(RIOB33_X105Y101_IOB_X1Y102_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y110_SLICE_X14Y110_BO5),
.O6(CLBLM_R_X11Y110_SLICE_X14Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0fffff5f5f5f5f)
  ) CLBLM_R_X11Y110_SLICE_X14Y110_ALUT (
.I0(RIOB33_X105Y103_IOB_X1Y103_I),
.I1(1'b1),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(1'b1),
.I4(RIOB33_X105Y101_IOB_X1Y101_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y110_SLICE_X14Y110_AO5),
.O6(CLBLM_R_X11Y110_SLICE_X14Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h1f057f3f3f15ff7f)
  ) CLBLM_R_X11Y110_SLICE_X15Y110_DLUT (
.I0(CLBLM_L_X12Y110_SLICE_X17Y110_BO6),
.I1(LIOB33_X0Y107_IOB_X0Y107_I),
.I2(RIOB33_X105Y103_IOB_X1Y103_I),
.I3(CLBLM_L_X12Y108_SLICE_X16Y108_CO6),
.I4(CLBLM_L_X12Y109_SLICE_X17Y109_CO6),
.I5(LIOB33_X0Y105_IOB_X0Y106_I),
.O5(CLBLM_R_X11Y110_SLICE_X15Y110_DO5),
.O6(CLBLM_R_X11Y110_SLICE_X15Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h96c33c96cc66cc66)
  ) CLBLM_R_X11Y110_SLICE_X15Y110_CLUT (
.I0(CLBLM_L_X12Y110_SLICE_X17Y110_BO6),
.I1(CLBLM_L_X12Y110_SLICE_X17Y110_CO6),
.I2(RIOB33_X105Y103_IOB_X1Y104_I),
.I3(CLBLM_L_X12Y108_SLICE_X16Y108_CO6),
.I4(RIOB33_X105Y103_IOB_X1Y103_I),
.I5(LIOB33_X0Y105_IOB_X0Y106_I),
.O5(CLBLM_R_X11Y110_SLICE_X15Y110_CO5),
.O6(CLBLM_R_X11Y110_SLICE_X15Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hed84eded8484ed84)
  ) CLBLM_R_X11Y110_SLICE_X15Y110_BLUT (
.I0(CLBLM_R_X11Y108_SLICE_X15Y108_AO5),
.I1(CLBLM_R_X11Y110_SLICE_X14Y110_BO6),
.I2(CLBLM_R_X11Y108_SLICE_X15Y108_BO6),
.I3(CLBLM_L_X12Y108_SLICE_X16Y108_AO5),
.I4(CLBLM_R_X13Y108_SLICE_X19Y108_AO6),
.I5(CLBLM_L_X10Y107_SLICE_X13Y107_AO6),
.O5(CLBLM_R_X11Y110_SLICE_X15Y110_BO5),
.O6(CLBLM_R_X11Y110_SLICE_X15Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6969966996699696)
  ) CLBLM_R_X11Y110_SLICE_X15Y110_ALUT (
.I0(CLBLM_R_X11Y108_SLICE_X15Y108_AO5),
.I1(CLBLM_R_X11Y110_SLICE_X14Y110_BO6),
.I2(CLBLM_R_X11Y108_SLICE_X15Y108_BO6),
.I3(CLBLM_R_X13Y108_SLICE_X19Y108_AO6),
.I4(CLBLM_L_X12Y108_SLICE_X16Y108_AO5),
.I5(CLBLM_L_X10Y107_SLICE_X13Y107_AO6),
.O5(CLBLM_R_X11Y110_SLICE_X15Y110_AO5),
.O6(CLBLM_R_X11Y110_SLICE_X15Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6999666996669996)
  ) CLBLM_R_X11Y111_SLICE_X14Y111_DLUT (
.I0(CLBLM_R_X11Y111_SLICE_X14Y111_AO6),
.I1(CLBLM_L_X10Y110_SLICE_X12Y110_BO6),
.I2(CLBLM_R_X11Y111_SLICE_X15Y111_AO6),
.I3(CLBLM_R_X11Y111_SLICE_X14Y111_AO5),
.I4(CLBLM_R_X11Y111_SLICE_X14Y111_CO6),
.I5(CLBLM_L_X10Y110_SLICE_X13Y110_AO6),
.O5(CLBLM_R_X11Y111_SLICE_X14Y111_DO5),
.O6(CLBLM_R_X11Y111_SLICE_X14Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996a55a96965a5a)
  ) CLBLM_R_X11Y111_SLICE_X14Y111_CLUT (
.I0(CLBLM_R_X11Y109_SLICE_X14Y109_CO6),
.I1(LIOB33_X0Y107_IOB_X0Y107_I),
.I2(CLBLM_R_X13Y108_SLICE_X18Y108_CO6),
.I3(LIOB33_X0Y105_IOB_X0Y106_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(RIOB33_X105Y107_IOB_X1Y107_I),
.O5(CLBLM_R_X11Y111_SLICE_X14Y111_CO5),
.O6(CLBLM_R_X11Y111_SLICE_X14Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdf7c431dc734010)
  ) CLBLM_R_X11Y111_SLICE_X14Y111_BLUT (
.I0(CLBLM_R_X11Y111_SLICE_X14Y111_CO6),
.I1(CLBLM_L_X10Y110_SLICE_X12Y110_BO6),
.I2(CLBLM_R_X11Y111_SLICE_X15Y111_AO6),
.I3(CLBLM_L_X10Y110_SLICE_X13Y110_AO6),
.I4(CLBLM_R_X11Y111_SLICE_X14Y111_AO6),
.I5(CLBLM_R_X11Y111_SLICE_X14Y111_AO5),
.O5(CLBLM_R_X11Y111_SLICE_X14Y111_BO5),
.O6(CLBLM_R_X11Y111_SLICE_X14Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ffffff5555ffff)
  ) CLBLM_R_X11Y111_SLICE_X14Y111_ALUT (
.I0(LIOB33_X0Y107_IOB_X0Y108_I),
.I1(1'b1),
.I2(1'b1),
.I3(LIOB33_X0Y109_IOB_X0Y109_I),
.I4(RIOB33_X105Y103_IOB_X1Y104_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y111_SLICE_X14Y111_AO5),
.O6(CLBLM_R_X11Y111_SLICE_X14Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h2b8eaf0abbeeffaa)
  ) CLBLM_R_X11Y111_SLICE_X15Y111_DLUT (
.I0(CLBLM_R_X11Y111_SLICE_X15Y111_AO6),
.I1(LIOB33_X0Y107_IOB_X0Y107_I),
.I2(LIOB33_X0Y107_IOB_X0Y108_I),
.I3(CLBLM_L_X12Y110_SLICE_X16Y110_DO6),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(RIOB33_X105Y103_IOB_X1Y104_I),
.O5(CLBLM_R_X11Y111_SLICE_X15Y111_DO5),
.O6(CLBLM_R_X11Y111_SLICE_X15Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'he888b222eee8bbb2)
  ) CLBLM_R_X11Y111_SLICE_X15Y111_CLUT (
.I0(CLBLM_R_X11Y112_SLICE_X15Y112_AO5),
.I1(CLBLM_R_X11Y111_SLICE_X14Y111_AO5),
.I2(CLBLM_R_X11Y110_SLICE_X15Y110_DO6),
.I3(CLBLM_L_X12Y110_SLICE_X16Y110_AO5),
.I4(CLBLM_R_X11Y109_SLICE_X15Y109_DO6),
.I5(CLBLM_R_X11Y111_SLICE_X15Y111_BO6),
.O5(CLBLM_R_X11Y111_SLICE_X15Y111_CO5),
.O6(CLBLM_R_X11Y111_SLICE_X15Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7887887787787788)
  ) CLBLM_R_X11Y111_SLICE_X15Y111_BLUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(RIOB33_X105Y103_IOB_X1Y104_I),
.I3(CLBLM_L_X12Y108_SLICE_X17Y108_CO6),
.I4(LIOB33_X0Y107_IOB_X0Y107_I),
.I5(CLBLM_L_X12Y109_SLICE_X17Y109_BO6),
.O5(CLBLM_R_X11Y111_SLICE_X15Y111_BO5),
.O6(CLBLM_R_X11Y111_SLICE_X15Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6fcfffff060c66cc)
  ) CLBLM_R_X11Y111_SLICE_X15Y111_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X12Y108_SLICE_X17Y108_CO6),
.I2(RIOB33_X105Y103_IOB_X1Y104_I),
.I3(LIOB33_X0Y105_IOB_X0Y106_I),
.I4(LIOB33_X0Y107_IOB_X0Y107_I),
.I5(CLBLM_L_X12Y109_SLICE_X17Y109_BO6),
.O5(CLBLM_R_X11Y111_SLICE_X15Y111_AO5),
.O6(CLBLM_R_X11Y111_SLICE_X15Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6fcfffff060c66cc)
  ) CLBLM_R_X11Y112_SLICE_X14Y112_DLUT (
.I0(LIOB33_X0Y107_IOB_X0Y107_I),
.I1(CLBLM_L_X12Y111_SLICE_X16Y111_DO6),
.I2(LIOB33_X0Y107_IOB_X0Y108_I),
.I3(RIOB33_X105Y103_IOB_X1Y104_I),
.I4(RIOB33_X105Y103_IOB_X1Y103_I),
.I5(CLBLM_R_X11Y110_SLICE_X15Y110_DO6),
.O5(CLBLM_R_X11Y112_SLICE_X14Y112_DO5),
.O6(CLBLM_R_X11Y112_SLICE_X14Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'he888eee8d444ddd4)
  ) CLBLM_R_X11Y112_SLICE_X14Y112_CLUT (
.I0(CLBLM_R_X11Y110_SLICE_X14Y110_DO6),
.I1(CLBLM_R_X11Y112_SLICE_X15Y112_AO6),
.I2(CLBLM_L_X10Y109_SLICE_X13Y109_DO6),
.I3(CLBLM_L_X10Y111_SLICE_X13Y111_AO5),
.I4(CLBLM_L_X12Y111_SLICE_X16Y111_CO6),
.I5(CLBLM_L_X10Y113_SLICE_X13Y113_AO5),
.O5(CLBLM_R_X11Y112_SLICE_X14Y112_CO5),
.O6(CLBLM_R_X11Y112_SLICE_X14Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'he673198c2abfd540)
  ) CLBLM_R_X11Y112_SLICE_X14Y112_BLUT (
.I0(CLBLM_L_X10Y109_SLICE_X13Y109_DO6),
.I1(LIOB33_X0Y107_IOB_X0Y108_I),
.I2(RIOB33_X105Y101_IOB_X1Y101_I),
.I3(CLBLM_L_X12Y111_SLICE_X16Y111_CO6),
.I4(CLBLM_R_X11Y110_SLICE_X14Y110_DO6),
.I5(RIOB33_X105Y101_IOB_X1Y102_I),
.O5(CLBLM_R_X11Y112_SLICE_X14Y112_BO5),
.O6(CLBLM_R_X11Y112_SLICE_X14Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h693c96c3c3693c96)
  ) CLBLM_R_X11Y112_SLICE_X14Y112_ALUT (
.I0(CLBLM_L_X10Y109_SLICE_X13Y109_DO6),
.I1(CLBLM_L_X10Y113_SLICE_X13Y113_AO5),
.I2(CLBLM_R_X11Y112_SLICE_X15Y112_AO6),
.I3(CLBLM_L_X12Y111_SLICE_X16Y111_CO6),
.I4(CLBLM_R_X11Y110_SLICE_X14Y110_DO6),
.I5(CLBLM_L_X10Y111_SLICE_X13Y111_AO5),
.O5(CLBLM_R_X11Y112_SLICE_X14Y112_AO5),
.O6(CLBLM_R_X11Y112_SLICE_X14Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996969699666666)
  ) CLBLM_R_X11Y112_SLICE_X15Y112_DLUT (
.I0(CLBLM_R_X11Y111_SLICE_X15Y111_AO6),
.I1(CLBLM_L_X12Y110_SLICE_X16Y110_DO6),
.I2(LIOB33_X0Y107_IOB_X0Y108_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(LIOB33_X0Y107_IOB_X0Y107_I),
.I5(RIOB33_X105Y103_IOB_X1Y104_I),
.O5(CLBLM_R_X11Y112_SLICE_X15Y112_DO5),
.O6(CLBLM_R_X11Y112_SLICE_X15Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h9c63f00f39c6ff00)
  ) CLBLM_R_X11Y112_SLICE_X15Y112_CLUT (
.I0(RIOB33_X105Y103_IOB_X1Y103_I),
.I1(RIOB33_X105Y103_IOB_X1Y104_I),
.I2(CLBLM_R_X11Y110_SLICE_X15Y110_DO6),
.I3(CLBLM_R_X11Y109_SLICE_X15Y109_DO6),
.I4(LIOB33_X0Y107_IOB_X0Y108_I),
.I5(CLBLM_R_X11Y111_SLICE_X15Y111_BO6),
.O5(CLBLM_R_X11Y112_SLICE_X15Y112_CO5),
.O6(CLBLM_R_X11Y112_SLICE_X15Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h4bd2b42db42d4bd2)
  ) CLBLM_R_X11Y112_SLICE_X15Y112_BLUT (
.I0(CLBLM_L_X12Y110_SLICE_X16Y110_AO5),
.I1(CLBLM_R_X11Y111_SLICE_X15Y111_BO6),
.I2(CLBLM_R_X11Y109_SLICE_X15Y109_DO6),
.I3(CLBLM_R_X11Y110_SLICE_X15Y110_DO6),
.I4(CLBLM_R_X11Y111_SLICE_X14Y111_AO5),
.I5(CLBLM_R_X11Y112_SLICE_X15Y112_AO5),
.O5(CLBLM_R_X11Y112_SLICE_X15Y112_BO5),
.O6(CLBLM_R_X11Y112_SLICE_X15Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h7777777733ff33ff)
  ) CLBLM_R_X11Y112_SLICE_X15Y112_ALUT (
.I0(RIOB33_X105Y101_IOB_X1Y101_I),
.I1(LIOB33_X0Y109_IOB_X0Y109_I),
.I2(1'b1),
.I3(RIOB33_X105Y103_IOB_X1Y103_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y112_SLICE_X15Y112_AO5),
.O6(CLBLM_R_X11Y112_SLICE_X15Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h1f077f575f17ff77)
  ) CLBLM_R_X11Y113_SLICE_X14Y113_DLUT (
.I0(CLBLM_R_X11Y112_SLICE_X15Y112_BO6),
.I1(CLBLM_R_X11Y113_SLICE_X15Y113_AO6),
.I2(RIOB33_X105Y101_IOB_X1Y102_I),
.I3(CLBLM_R_X11Y114_SLICE_X14Y114_CO6),
.I4(LIOB33_X0Y109_IOB_X0Y110_I),
.I5(LIOB33_X0Y109_IOB_X0Y109_I),
.O5(CLBLM_R_X11Y113_SLICE_X14Y113_DO5),
.O6(CLBLM_R_X11Y113_SLICE_X14Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffd4d4ffd40000d4)
  ) CLBLM_R_X11Y113_SLICE_X14Y113_CLUT (
.I0(CLBLM_L_X12Y110_SLICE_X17Y110_AO6),
.I1(CLBLM_L_X12Y111_SLICE_X16Y111_AO6),
.I2(CLBLM_L_X10Y113_SLICE_X13Y113_AO5),
.I3(CLBLM_L_X12Y110_SLICE_X16Y110_AO5),
.I4(CLBLM_R_X11Y109_SLICE_X15Y109_CO6),
.I5(CLBLM_L_X10Y113_SLICE_X13Y113_AO6),
.O5(CLBLM_R_X11Y113_SLICE_X14Y113_CO5),
.O6(CLBLM_R_X11Y113_SLICE_X14Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha569695a9999aaaa)
  ) CLBLM_R_X11Y113_SLICE_X14Y113_BLUT (
.I0(CLBLM_R_X11Y109_SLICE_X15Y109_CO6),
.I1(CLBLM_L_X12Y111_SLICE_X16Y111_AO6),
.I2(RIOB33_X105Y103_IOB_X1Y103_I),
.I3(RIOB33_X105Y101_IOB_X1Y102_I),
.I4(CLBLM_L_X12Y110_SLICE_X17Y110_AO6),
.I5(LIOB33_X0Y107_IOB_X0Y108_I),
.O5(CLBLM_R_X11Y113_SLICE_X14Y113_BO5),
.O6(CLBLM_R_X11Y113_SLICE_X14Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6a9556a9956aa956)
  ) CLBLM_R_X11Y113_SLICE_X14Y113_ALUT (
.I0(CLBLM_R_X11Y109_SLICE_X15Y109_CO6),
.I1(CLBLM_L_X10Y113_SLICE_X13Y113_AO5),
.I2(CLBLM_L_X12Y111_SLICE_X16Y111_AO6),
.I3(CLBLM_L_X10Y113_SLICE_X13Y113_AO6),
.I4(CLBLM_L_X12Y110_SLICE_X17Y110_AO6),
.I5(CLBLM_L_X12Y110_SLICE_X16Y110_AO5),
.O5(CLBLM_R_X11Y113_SLICE_X14Y113_AO5),
.O6(CLBLM_R_X11Y113_SLICE_X14Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y113_SLICE_X15Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y113_SLICE_X15Y113_DO5),
.O6(CLBLM_R_X11Y113_SLICE_X15Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y113_SLICE_X15Y113_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y113_SLICE_X15Y113_CO5),
.O6(CLBLM_R_X11Y113_SLICE_X15Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y113_SLICE_X15Y113_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y113_SLICE_X15Y113_BO5),
.O6(CLBLM_R_X11Y113_SLICE_X15Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6999966696669666)
  ) CLBLM_R_X11Y113_SLICE_X15Y113_ALUT (
.I0(CLBLM_R_X11Y110_SLICE_X15Y110_DO6),
.I1(CLBLM_L_X12Y111_SLICE_X16Y111_DO6),
.I2(RIOB33_X105Y103_IOB_X1Y103_I),
.I3(LIOB33_X0Y107_IOB_X0Y108_I),
.I4(RIOB33_X105Y103_IOB_X1Y104_I),
.I5(LIOB33_X0Y107_IOB_X0Y107_I),
.O5(CLBLM_R_X11Y113_SLICE_X15Y113_AO5),
.O6(CLBLM_R_X11Y113_SLICE_X15Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h95a96a56aa66aa66)
  ) CLBLM_R_X11Y114_SLICE_X14Y114_DLUT (
.I0(CLBLM_R_X11Y112_SLICE_X15Y112_CO6),
.I1(CLBLM_R_X11Y113_SLICE_X15Y113_AO6),
.I2(RIOB33_X105Y101_IOB_X1Y102_I),
.I3(CLBLM_R_X11Y114_SLICE_X14Y114_CO6),
.I4(RIOB33_X105Y103_IOB_X1Y103_I),
.I5(LIOB33_X0Y109_IOB_X0Y109_I),
.O5(CLBLM_R_X11Y114_SLICE_X14Y114_DO5),
.O6(CLBLM_R_X11Y114_SLICE_X14Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h2abfbf2abf2abf2a)
  ) CLBLM_R_X11Y114_SLICE_X14Y114_CLUT (
.I0(CLBLM_L_X12Y111_SLICE_X16Y111_AO6),
.I1(LIOB33_X0Y107_IOB_X0Y108_I),
.I2(RIOB33_X105Y101_IOB_X1Y102_I),
.I3(CLBLM_R_X11Y110_SLICE_X15Y110_CO6),
.I4(RIOB33_X105Y103_IOB_X1Y103_I),
.I5(LIOB33_X0Y107_IOB_X0Y107_I),
.O5(CLBLM_R_X11Y114_SLICE_X14Y114_CO5),
.O6(CLBLM_R_X11Y114_SLICE_X14Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hb43c78f0d2961e5a)
  ) CLBLM_R_X11Y114_SLICE_X14Y114_BLUT (
.I0(CLBLM_R_X11Y113_SLICE_X15Y113_AO6),
.I1(RIOB33_X105Y101_IOB_X1Y102_I),
.I2(CLBLM_R_X11Y112_SLICE_X15Y112_BO6),
.I3(LIOB33_X0Y109_IOB_X0Y109_I),
.I4(LIOB33_X0Y109_IOB_X0Y110_I),
.I5(CLBLM_R_X11Y114_SLICE_X14Y114_CO6),
.O5(CLBLM_R_X11Y114_SLICE_X14Y114_BO5),
.O6(CLBLM_R_X11Y114_SLICE_X14Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6ac0953f953f6ac0)
  ) CLBLM_R_X11Y114_SLICE_X14Y114_ALUT (
.I0(LIOB33_X0Y107_IOB_X0Y108_I),
.I1(RIOB33_X105Y103_IOB_X1Y103_I),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(RIOB33_X105Y101_IOB_X1Y102_I),
.I4(CLBLM_L_X12Y111_SLICE_X16Y111_AO6),
.I5(CLBLM_R_X11Y110_SLICE_X15Y110_CO6),
.O5(CLBLM_R_X11Y114_SLICE_X14Y114_AO5),
.O6(CLBLM_R_X11Y114_SLICE_X14Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y114_SLICE_X15Y114_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y114_SLICE_X15Y114_DO5),
.O6(CLBLM_R_X11Y114_SLICE_X15Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y114_SLICE_X15Y114_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y114_SLICE_X15Y114_CO5),
.O6(CLBLM_R_X11Y114_SLICE_X15Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y114_SLICE_X15Y114_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y114_SLICE_X15Y114_BO5),
.O6(CLBLM_R_X11Y114_SLICE_X15Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y114_SLICE_X15Y114_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y114_SLICE_X15Y114_AO5),
.O6(CLBLM_R_X11Y114_SLICE_X15Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h2dd2b44bd22d4bb4)
  ) CLBLM_R_X13Y108_SLICE_X18Y108_DLUT (
.I0(CLBLM_R_X11Y106_SLICE_X15Y106_CO6),
.I1(CLBLM_R_X13Y108_SLICE_X18Y108_AO6),
.I2(CLBLM_L_X12Y109_SLICE_X16Y109_AO6),
.I3(CLBLM_R_X11Y106_SLICE_X14Y106_BO6),
.I4(CLBLM_L_X12Y108_SLICE_X17Y108_AO6),
.I5(CLBLM_R_X11Y109_SLICE_X15Y109_AO5),
.O5(CLBLM_R_X13Y108_SLICE_X18Y108_DO5),
.O6(CLBLM_R_X13Y108_SLICE_X18Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdd0f440d0fd40f4)
  ) CLBLM_R_X13Y108_SLICE_X18Y108_CLUT (
.I0(CLBLM_R_X11Y106_SLICE_X15Y106_CO6),
.I1(CLBLM_R_X13Y108_SLICE_X18Y108_AO6),
.I2(CLBLM_L_X12Y109_SLICE_X16Y109_AO6),
.I3(CLBLM_R_X11Y106_SLICE_X14Y106_BO6),
.I4(CLBLM_L_X12Y108_SLICE_X17Y108_AO6),
.I5(CLBLM_R_X11Y109_SLICE_X15Y109_AO5),
.O5(CLBLM_R_X13Y108_SLICE_X18Y108_CO5),
.O6(CLBLM_R_X13Y108_SLICE_X18Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996c33c996633cc)
  ) CLBLM_R_X13Y108_SLICE_X18Y108_BLUT (
.I0(LIOB33_X0Y101_IOB_X0Y102_I),
.I1(CLBLM_L_X12Y107_SLICE_X16Y107_BO6),
.I2(LIOB33_X0Y103_IOB_X0Y104_I),
.I3(CLBLM_R_X11Y107_SLICE_X15Y107_BO6),
.I4(RIOB33_X105Y107_IOB_X1Y107_I),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X13Y108_SLICE_X18Y108_BO5),
.O6(CLBLM_R_X13Y108_SLICE_X18Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h4d8ecf0cddeeffcc)
  ) CLBLM_R_X13Y108_SLICE_X18Y108_ALUT (
.I0(LIOB33_X0Y101_IOB_X0Y102_I),
.I1(CLBLM_R_X11Y107_SLICE_X15Y107_BO6),
.I2(LIOB33_X0Y103_IOB_X0Y104_I),
.I3(CLBLM_L_X12Y107_SLICE_X16Y107_BO6),
.I4(RIOB33_X105Y107_IOB_X1Y107_I),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X13Y108_SLICE_X18Y108_AO5),
.O6(CLBLM_R_X13Y108_SLICE_X18Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y108_SLICE_X19Y108_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y108_SLICE_X19Y108_DO5),
.O6(CLBLM_R_X13Y108_SLICE_X19Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y108_SLICE_X19Y108_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y108_SLICE_X19Y108_CO5),
.O6(CLBLM_R_X13Y108_SLICE_X19Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fff8fff07770888)
  ) CLBLM_R_X13Y108_SLICE_X19Y108_BLUT (
.I0(LIOB33_X0Y101_IOB_X0Y102_I),
.I1(RIOB33_X105Y103_IOB_X1Y104_I),
.I2(RIOB33_X105Y103_IOB_X1Y103_I),
.I3(LIOB33_X0Y103_IOB_X0Y104_I),
.I4(CLBLM_R_X11Y108_SLICE_X14Y108_CO6),
.I5(CLBLM_L_X10Y108_SLICE_X13Y108_DO6),
.O5(CLBLM_R_X13Y108_SLICE_X19Y108_BO5),
.O6(CLBLM_R_X13Y108_SLICE_X19Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h7887878787787878)
  ) CLBLM_R_X13Y108_SLICE_X19Y108_ALUT (
.I0(LIOB33_X0Y101_IOB_X0Y102_I),
.I1(RIOB33_X105Y103_IOB_X1Y104_I),
.I2(CLBLM_R_X11Y108_SLICE_X14Y108_CO6),
.I3(LIOB33_X0Y103_IOB_X0Y104_I),
.I4(RIOB33_X105Y103_IOB_X1Y103_I),
.I5(CLBLM_L_X10Y108_SLICE_X13Y108_DO6),
.O5(CLBLM_R_X13Y108_SLICE_X19Y108_AO5),
.O6(CLBLM_R_X13Y108_SLICE_X19Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y101_IOB_X0Y101_IBUF (
.I(LIOB33_X0Y101_IOB_X0Y101_IPAD),
.O(LIOB33_X0Y101_IOB_X0Y101_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y101_IOB_X0Y102_IBUF (
.I(LIOB33_X0Y101_IOB_X0Y102_IPAD),
.O(LIOB33_X0Y101_IOB_X0Y102_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y103_IOB_X0Y103_IBUF (
.I(LIOB33_X0Y103_IOB_X0Y103_IPAD),
.O(LIOB33_X0Y103_IOB_X0Y103_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y103_IOB_X0Y104_IBUF (
.I(LIOB33_X0Y103_IOB_X0Y104_IPAD),
.O(LIOB33_X0Y103_IOB_X0Y104_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y105_IOB_X0Y105_IBUF (
.I(LIOB33_X0Y105_IOB_X0Y105_IPAD),
.O(LIOB33_X0Y105_IOB_X0Y105_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y105_IOB_X0Y106_IBUF (
.I(LIOB33_X0Y105_IOB_X0Y106_IPAD),
.O(LIOB33_X0Y105_IOB_X0Y106_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y107_IOB_X0Y107_IBUF (
.I(LIOB33_X0Y107_IOB_X0Y107_IPAD),
.O(LIOB33_X0Y107_IOB_X0Y107_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y107_IOB_X0Y108_IBUF (
.I(LIOB33_X0Y107_IOB_X0Y108_IPAD),
.O(LIOB33_X0Y107_IOB_X0Y108_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y109_IOB_X0Y109_IBUF (
.I(LIOB33_X0Y109_IOB_X0Y109_IPAD),
.O(LIOB33_X0Y109_IOB_X0Y109_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y109_IOB_X0Y110_IBUF (
.I(LIOB33_X0Y109_IOB_X0Y110_IPAD),
.O(LIOB33_X0Y109_IOB_X0Y110_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y111_IOB_X0Y111_IBUF (
.I(LIOB33_X0Y111_IOB_X0Y111_IPAD),
.O(LIOB33_X0Y111_IOB_X0Y111_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y111_IOB_X0Y112_IBUF (
.I(LIOB33_X0Y111_IOB_X0Y112_IPAD),
.O(LIOB33_X0Y111_IOB_X0Y112_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y113_IOB_X0Y113_IBUF (
.I(LIOB33_X0Y113_IOB_X0Y113_IPAD),
.O(LIOB33_X0Y113_IOB_X0Y113_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y113_IOB_X0Y114_IBUF (
.I(LIOB33_X0Y113_IOB_X0Y114_IPAD),
.O(LIOB33_X0Y113_IOB_X0Y114_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y115_IOB_X0Y115_IBUF (
.I(LIOB33_X0Y115_IOB_X0Y115_IPAD),
.O(LIOB33_X0Y115_IOB_X0Y115_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y115_IOB_X0Y116_IBUF (
.I(LIOB33_X0Y115_IOB_X0Y116_IPAD),
.O(LIOB33_X0Y115_IOB_X0Y116_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y117_IOB_X0Y117_IBUF (
.I(LIOB33_X0Y117_IOB_X0Y117_IPAD),
.O(LIOB33_X0Y117_IOB_X0Y117_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y117_IOB_X0Y118_OBUF (
.I(CLBLL_L_X2Y112_SLICE_X0Y112_AO5),
.O(LIOB33_X0Y117_IOB_X0Y118_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y119_IOB_X0Y119_OBUF (
.I(CLBLL_L_X2Y112_SLICE_X0Y112_AO6),
.O(LIOB33_X0Y119_IOB_X0Y119_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y119_IOB_X0Y120_OBUF (
.I(CLBLL_L_X2Y109_SLICE_X0Y109_AO5),
.O(LIOB33_X0Y119_IOB_X0Y120_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y121_IOB_X0Y121_OBUF (
.I(CLBLL_L_X2Y108_SLICE_X0Y108_AO5),
.O(LIOB33_X0Y121_IOB_X0Y121_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y121_IOB_X0Y122_OBUF (
.I(CLBLL_L_X2Y108_SLICE_X1Y108_AO6),
.O(LIOB33_X0Y121_IOB_X0Y122_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y123_IOB_X0Y123_OBUF (
.I(CLBLL_L_X2Y108_SLICE_X0Y108_CO6),
.O(LIOB33_X0Y123_IOB_X0Y123_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y123_IOB_X0Y124_OBUF (
.I(CLBLL_L_X2Y107_SLICE_X1Y107_AO5),
.O(LIOB33_X0Y123_IOB_X0Y124_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y125_IOB_X0Y125_OBUF (
.I(CLBLM_R_X3Y107_SLICE_X2Y107_AO6),
.O(LIOB33_X0Y125_IOB_X0Y125_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y125_IOB_X0Y126_OBUF (
.I(CLBLM_R_X3Y108_SLICE_X3Y108_AO6),
.O(LIOB33_X0Y125_IOB_X0Y126_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y127_IOB_X0Y127_OBUF (
.I(CLBLL_L_X4Y109_SLICE_X4Y109_AO6),
.O(LIOB33_X0Y127_IOB_X0Y127_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y127_IOB_X0Y128_OBUF (
.I(CLBLM_R_X3Y110_SLICE_X3Y110_AO6),
.O(LIOB33_X0Y127_IOB_X0Y128_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y129_IOB_X0Y129_OBUF (
.I(CLBLM_R_X3Y110_SLICE_X3Y110_BO6),
.O(LIOB33_X0Y129_IOB_X0Y129_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y129_IOB_X0Y130_OBUF (
.I(CLBLL_L_X2Y109_SLICE_X0Y109_BO5),
.O(LIOB33_X0Y129_IOB_X0Y130_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y131_IOB_X0Y131_OBUF (
.I(CLBLL_L_X4Y111_SLICE_X4Y111_AO6),
.O(LIOB33_X0Y131_IOB_X0Y131_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y131_IOB_X0Y132_OBUF (
.I(CLBLM_R_X3Y114_SLICE_X3Y114_AO5),
.O(LIOB33_X0Y131_IOB_X0Y132_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y133_IOB_X0Y133_OBUF (
.I(CLBLL_L_X4Y112_SLICE_X4Y112_AO6),
.O(LIOB33_X0Y133_IOB_X0Y133_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y133_IOB_X0Y134_OBUF (
.I(1'b0),
.O(LIOB33_X0Y133_IOB_X0Y134_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y135_IOB_X0Y135_OBUF (
.I(CLBLM_R_X5Y114_SLICE_X6Y114_AO5),
.O(LIOB33_X0Y135_IOB_X0Y135_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y135_IOB_X0Y136_OBUF (
.I(CLBLM_R_X5Y114_SLICE_X6Y114_AO6),
.O(LIOB33_X0Y135_IOB_X0Y136_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y137_IOB_X0Y137_OBUF (
.I(CLBLL_L_X4Y116_SLICE_X5Y116_AO6),
.O(LIOB33_X0Y137_IOB_X0Y137_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y137_IOB_X0Y138_OBUF (
.I(CLBLL_L_X4Y116_SLICE_X5Y116_AO5),
.O(LIOB33_X0Y137_IOB_X0Y138_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y139_IOB_X0Y139_OBUF (
.I(CLBLL_L_X4Y116_SLICE_X5Y116_BO6),
.O(LIOB33_X0Y139_IOB_X0Y139_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y139_IOB_X0Y140_OBUF (
.I(CLBLL_L_X4Y116_SLICE_X5Y116_BO5),
.O(LIOB33_X0Y139_IOB_X0Y140_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y141_IOB_X0Y141_OBUF (
.I(CLBLM_R_X5Y116_SLICE_X7Y116_DO6),
.O(LIOB33_X0Y141_IOB_X0Y141_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y141_IOB_X0Y142_OBUF (
.I(CLBLL_L_X4Y116_SLICE_X4Y116_BO6),
.O(LIOB33_X0Y141_IOB_X0Y142_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y143_IOB_X0Y143_OBUF (
.I(CLBLL_L_X4Y115_SLICE_X4Y115_DO6),
.O(LIOB33_X0Y143_IOB_X0Y143_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y145_IOB_X0Y145_OBUF (
.I(CLBLL_L_X4Y114_SLICE_X4Y114_AO6),
.O(LIOB33_X0Y145_IOB_X0Y145_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y145_IOB_X0Y146_OBUF (
.I(CLBLL_L_X4Y113_SLICE_X4Y113_BO6),
.O(LIOB33_X0Y145_IOB_X0Y146_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y147_IOB_X0Y147_OBUF (
.I(CLBLM_R_X3Y113_SLICE_X3Y113_AO6),
.O(LIOB33_X0Y147_IOB_X0Y147_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y147_IOB_X0Y148_OBUF (
.I(CLBLM_R_X3Y113_SLICE_X3Y113_CO6),
.O(LIOB33_X0Y147_IOB_X0Y148_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_SING_X0Y100_IOB_X0Y100_IBUF (
.I(LIOB33_SING_X0Y100_IOB_X0Y100_IPAD),
.O(LIOB33_SING_X0Y100_IOB_X0Y100_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y149_IOB_X0Y149_OBUF (
.I(CLBLM_R_X3Y113_SLICE_X3Y113_AO5),
.O(LIOB33_SING_X0Y149_IOB_X0Y149_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y101_IOB_X1Y101_IBUF (
.I(RIOB33_X105Y101_IOB_X1Y101_IPAD),
.O(RIOB33_X105Y101_IOB_X1Y101_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y101_IOB_X1Y102_IBUF (
.I(RIOB33_X105Y101_IOB_X1Y102_IPAD),
.O(RIOB33_X105Y101_IOB_X1Y102_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y103_IOB_X1Y103_IBUF (
.I(RIOB33_X105Y103_IOB_X1Y103_IPAD),
.O(RIOB33_X105Y103_IOB_X1Y103_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y103_IOB_X1Y104_IBUF (
.I(RIOB33_X105Y103_IOB_X1Y104_IPAD),
.O(RIOB33_X105Y103_IOB_X1Y104_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y105_IOB_X1Y105_IBUF (
.I(RIOB33_X105Y105_IOB_X1Y105_IPAD),
.O(RIOB33_X105Y105_IOB_X1Y105_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y105_IOB_X1Y106_IBUF (
.I(RIOB33_X105Y105_IOB_X1Y106_IPAD),
.O(RIOB33_X105Y105_IOB_X1Y106_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y107_IOB_X1Y107_IBUF (
.I(RIOB33_X105Y107_IOB_X1Y107_IPAD),
.O(RIOB33_X105Y107_IOB_X1Y107_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y107_IOB_X1Y108_IBUF (
.I(RIOB33_X105Y107_IOB_X1Y108_IPAD),
.O(RIOB33_X105Y107_IOB_X1Y108_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y109_IOB_X1Y109_IBUF (
.I(RIOB33_X105Y109_IOB_X1Y109_IPAD),
.O(RIOB33_X105Y109_IOB_X1Y109_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y109_IOB_X1Y110_IBUF (
.I(RIOB33_X105Y109_IOB_X1Y110_IPAD),
.O(RIOB33_X105Y109_IOB_X1Y110_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y111_IOB_X1Y111_IBUF (
.I(RIOB33_X105Y111_IOB_X1Y111_IPAD),
.O(RIOB33_X105Y111_IOB_X1Y111_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y111_IOB_X1Y112_IBUF (
.I(RIOB33_X105Y111_IOB_X1Y112_IPAD),
.O(RIOB33_X105Y111_IOB_X1Y112_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y113_IOB_X1Y113_IBUF (
.I(RIOB33_X105Y113_IOB_X1Y113_IPAD),
.O(RIOB33_X105Y113_IOB_X1Y113_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_SING_X105Y100_IOB_X1Y100_IBUF (
.I(RIOB33_SING_X105Y100_IOB_X1Y100_IPAD),
.O(RIOB33_SING_X105Y100_IOB_X1Y100_I)
  );
  assign CLBLL_L_X2Y106_SLICE_X0Y106_A = CLBLL_L_X2Y106_SLICE_X0Y106_AO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_B = CLBLL_L_X2Y106_SLICE_X0Y106_BO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_C = CLBLL_L_X2Y106_SLICE_X0Y106_CO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_D = CLBLL_L_X2Y106_SLICE_X0Y106_DO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_AMUX = CLBLL_L_X2Y106_SLICE_X0Y106_AO5;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_BMUX = CLBLL_L_X2Y106_SLICE_X0Y106_BO5;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_A = CLBLL_L_X2Y106_SLICE_X1Y106_AO6;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_B = CLBLL_L_X2Y106_SLICE_X1Y106_BO6;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_C = CLBLL_L_X2Y106_SLICE_X1Y106_CO6;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_D = CLBLL_L_X2Y106_SLICE_X1Y106_DO6;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_AMUX = CLBLL_L_X2Y106_SLICE_X1Y106_AO6;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_A = CLBLL_L_X2Y107_SLICE_X0Y107_AO6;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_B = CLBLL_L_X2Y107_SLICE_X0Y107_BO6;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_C = CLBLL_L_X2Y107_SLICE_X0Y107_CO6;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_D = CLBLL_L_X2Y107_SLICE_X0Y107_DO6;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_AMUX = CLBLL_L_X2Y107_SLICE_X0Y107_AO5;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_A = CLBLL_L_X2Y107_SLICE_X1Y107_AO6;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_B = CLBLL_L_X2Y107_SLICE_X1Y107_BO6;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_C = CLBLL_L_X2Y107_SLICE_X1Y107_CO6;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_D = CLBLL_L_X2Y107_SLICE_X1Y107_DO6;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_AMUX = CLBLL_L_X2Y107_SLICE_X1Y107_AO5;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_CMUX = CLBLL_L_X2Y107_SLICE_X1Y107_CO6;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_A = CLBLL_L_X2Y108_SLICE_X0Y108_AO6;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_B = CLBLL_L_X2Y108_SLICE_X0Y108_BO6;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_C = CLBLL_L_X2Y108_SLICE_X0Y108_CO6;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_D = CLBLL_L_X2Y108_SLICE_X0Y108_DO6;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_AMUX = CLBLL_L_X2Y108_SLICE_X0Y108_AO5;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_A = CLBLL_L_X2Y108_SLICE_X1Y108_AO6;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_B = CLBLL_L_X2Y108_SLICE_X1Y108_BO6;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_C = CLBLL_L_X2Y108_SLICE_X1Y108_CO6;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_D = CLBLL_L_X2Y108_SLICE_X1Y108_DO6;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_AMUX = CLBLL_L_X2Y108_SLICE_X1Y108_AO5;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_BMUX = CLBLL_L_X2Y108_SLICE_X1Y108_BO5;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_CMUX = CLBLL_L_X2Y108_SLICE_X1Y108_CO6;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_A = CLBLL_L_X2Y109_SLICE_X0Y109_AO6;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_B = CLBLL_L_X2Y109_SLICE_X0Y109_BO6;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_C = CLBLL_L_X2Y109_SLICE_X0Y109_CO6;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_D = CLBLL_L_X2Y109_SLICE_X0Y109_DO6;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_AMUX = CLBLL_L_X2Y109_SLICE_X0Y109_AO5;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_BMUX = CLBLL_L_X2Y109_SLICE_X0Y109_BO5;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_CMUX = CLBLL_L_X2Y109_SLICE_X0Y109_CO6;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_A = CLBLL_L_X2Y109_SLICE_X1Y109_AO6;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_B = CLBLL_L_X2Y109_SLICE_X1Y109_BO6;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_C = CLBLL_L_X2Y109_SLICE_X1Y109_CO6;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_D = CLBLL_L_X2Y109_SLICE_X1Y109_DO6;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_A = CLBLL_L_X2Y110_SLICE_X0Y110_AO6;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_B = CLBLL_L_X2Y110_SLICE_X0Y110_BO6;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_C = CLBLL_L_X2Y110_SLICE_X0Y110_CO6;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_D = CLBLL_L_X2Y110_SLICE_X0Y110_DO6;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_A = CLBLL_L_X2Y110_SLICE_X1Y110_AO6;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_B = CLBLL_L_X2Y110_SLICE_X1Y110_BO6;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_C = CLBLL_L_X2Y110_SLICE_X1Y110_CO6;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_D = CLBLL_L_X2Y110_SLICE_X1Y110_DO6;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_A = CLBLL_L_X2Y111_SLICE_X0Y111_AO6;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_B = CLBLL_L_X2Y111_SLICE_X0Y111_BO6;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_C = CLBLL_L_X2Y111_SLICE_X0Y111_CO6;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_D = CLBLL_L_X2Y111_SLICE_X0Y111_DO6;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_A = CLBLL_L_X2Y111_SLICE_X1Y111_AO6;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_B = CLBLL_L_X2Y111_SLICE_X1Y111_BO6;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_C = CLBLL_L_X2Y111_SLICE_X1Y111_CO6;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_D = CLBLL_L_X2Y111_SLICE_X1Y111_DO6;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_A = CLBLL_L_X2Y112_SLICE_X0Y112_AO6;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_B = CLBLL_L_X2Y112_SLICE_X0Y112_BO6;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_C = CLBLL_L_X2Y112_SLICE_X0Y112_CO6;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_D = CLBLL_L_X2Y112_SLICE_X0Y112_DO6;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_AMUX = CLBLL_L_X2Y112_SLICE_X0Y112_AO5;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_A = CLBLL_L_X2Y112_SLICE_X1Y112_AO6;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_B = CLBLL_L_X2Y112_SLICE_X1Y112_BO6;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_C = CLBLL_L_X2Y112_SLICE_X1Y112_CO6;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_D = CLBLL_L_X2Y112_SLICE_X1Y112_DO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_A = CLBLL_L_X4Y105_SLICE_X4Y105_AO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_B = CLBLL_L_X4Y105_SLICE_X4Y105_BO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_C = CLBLL_L_X4Y105_SLICE_X4Y105_CO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_D = CLBLL_L_X4Y105_SLICE_X4Y105_DO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_AMUX = CLBLL_L_X4Y105_SLICE_X4Y105_AO5;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_A = CLBLL_L_X4Y105_SLICE_X5Y105_AO6;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_B = CLBLL_L_X4Y105_SLICE_X5Y105_BO6;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_C = CLBLL_L_X4Y105_SLICE_X5Y105_CO6;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_D = CLBLL_L_X4Y105_SLICE_X5Y105_DO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_A = CLBLL_L_X4Y106_SLICE_X4Y106_AO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_B = CLBLL_L_X4Y106_SLICE_X4Y106_BO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_C = CLBLL_L_X4Y106_SLICE_X4Y106_CO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_D = CLBLL_L_X4Y106_SLICE_X4Y106_DO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_AMUX = CLBLL_L_X4Y106_SLICE_X4Y106_AO5;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_A = CLBLL_L_X4Y106_SLICE_X5Y106_AO6;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_B = CLBLL_L_X4Y106_SLICE_X5Y106_BO6;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_C = CLBLL_L_X4Y106_SLICE_X5Y106_CO6;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_D = CLBLL_L_X4Y106_SLICE_X5Y106_DO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_A = CLBLL_L_X4Y107_SLICE_X4Y107_AO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_B = CLBLL_L_X4Y107_SLICE_X4Y107_BO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_C = CLBLL_L_X4Y107_SLICE_X4Y107_CO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_D = CLBLL_L_X4Y107_SLICE_X4Y107_DO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_A = CLBLL_L_X4Y107_SLICE_X5Y107_AO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_B = CLBLL_L_X4Y107_SLICE_X5Y107_BO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_C = CLBLL_L_X4Y107_SLICE_X5Y107_CO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_D = CLBLL_L_X4Y107_SLICE_X5Y107_DO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_A = CLBLL_L_X4Y108_SLICE_X4Y108_AO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_B = CLBLL_L_X4Y108_SLICE_X4Y108_BO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_C = CLBLL_L_X4Y108_SLICE_X4Y108_CO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_D = CLBLL_L_X4Y108_SLICE_X4Y108_DO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_A = CLBLL_L_X4Y108_SLICE_X5Y108_AO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_B = CLBLL_L_X4Y108_SLICE_X5Y108_BO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_C = CLBLL_L_X4Y108_SLICE_X5Y108_CO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_D = CLBLL_L_X4Y108_SLICE_X5Y108_DO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_AMUX = CLBLL_L_X4Y108_SLICE_X5Y108_AO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A = CLBLL_L_X4Y109_SLICE_X4Y109_AO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B = CLBLL_L_X4Y109_SLICE_X4Y109_BO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C = CLBLL_L_X4Y109_SLICE_X4Y109_CO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D = CLBLL_L_X4Y109_SLICE_X4Y109_DO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_AMUX = CLBLL_L_X4Y109_SLICE_X4Y109_AO5;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A = CLBLL_L_X4Y109_SLICE_X5Y109_AO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B = CLBLL_L_X4Y109_SLICE_X5Y109_BO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C = CLBLL_L_X4Y109_SLICE_X5Y109_CO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D = CLBLL_L_X4Y109_SLICE_X5Y109_DO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_A = CLBLL_L_X4Y110_SLICE_X4Y110_AO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_B = CLBLL_L_X4Y110_SLICE_X4Y110_BO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_C = CLBLL_L_X4Y110_SLICE_X4Y110_CO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_D = CLBLL_L_X4Y110_SLICE_X4Y110_DO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_AMUX = CLBLL_L_X4Y110_SLICE_X4Y110_AO5;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_BMUX = CLBLL_L_X4Y110_SLICE_X4Y110_BO5;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_A = CLBLL_L_X4Y110_SLICE_X5Y110_AO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_B = CLBLL_L_X4Y110_SLICE_X5Y110_BO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_C = CLBLL_L_X4Y110_SLICE_X5Y110_CO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_D = CLBLL_L_X4Y110_SLICE_X5Y110_DO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_A = CLBLL_L_X4Y111_SLICE_X4Y111_AO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_B = CLBLL_L_X4Y111_SLICE_X4Y111_BO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_C = CLBLL_L_X4Y111_SLICE_X4Y111_CO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_D = CLBLL_L_X4Y111_SLICE_X4Y111_DO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_AMUX = CLBLL_L_X4Y111_SLICE_X4Y111_AO5;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_A = CLBLL_L_X4Y111_SLICE_X5Y111_AO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_B = CLBLL_L_X4Y111_SLICE_X5Y111_BO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_C = CLBLL_L_X4Y111_SLICE_X5Y111_CO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_D = CLBLL_L_X4Y111_SLICE_X5Y111_DO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_BMUX = CLBLL_L_X4Y111_SLICE_X5Y111_BO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_A = CLBLL_L_X4Y112_SLICE_X4Y112_AO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_B = CLBLL_L_X4Y112_SLICE_X4Y112_BO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_C = CLBLL_L_X4Y112_SLICE_X4Y112_CO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_D = CLBLL_L_X4Y112_SLICE_X4Y112_DO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_A = CLBLL_L_X4Y112_SLICE_X5Y112_AO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_B = CLBLL_L_X4Y112_SLICE_X5Y112_BO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_C = CLBLL_L_X4Y112_SLICE_X5Y112_CO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_D = CLBLL_L_X4Y112_SLICE_X5Y112_DO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_AMUX = CLBLL_L_X4Y112_SLICE_X5Y112_AO5;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_BMUX = CLBLL_L_X4Y112_SLICE_X5Y112_BO5;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A = CLBLL_L_X4Y113_SLICE_X4Y113_AO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B = CLBLL_L_X4Y113_SLICE_X4Y113_BO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C = CLBLL_L_X4Y113_SLICE_X4Y113_CO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D = CLBLL_L_X4Y113_SLICE_X4Y113_DO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_AMUX = CLBLL_L_X4Y113_SLICE_X4Y113_AO5;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A = CLBLL_L_X4Y113_SLICE_X5Y113_AO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B = CLBLL_L_X4Y113_SLICE_X5Y113_BO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C = CLBLL_L_X4Y113_SLICE_X5Y113_CO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D = CLBLL_L_X4Y113_SLICE_X5Y113_DO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_AMUX = CLBLL_L_X4Y113_SLICE_X5Y113_AO5;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_BMUX = CLBLL_L_X4Y113_SLICE_X5Y113_BO5;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_CMUX = CLBLL_L_X4Y113_SLICE_X5Y113_CO6;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_A = CLBLL_L_X4Y114_SLICE_X4Y114_AO6;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_B = CLBLL_L_X4Y114_SLICE_X4Y114_BO6;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_C = CLBLL_L_X4Y114_SLICE_X4Y114_CO6;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_D = CLBLL_L_X4Y114_SLICE_X4Y114_DO6;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_A = CLBLL_L_X4Y114_SLICE_X5Y114_AO6;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_B = CLBLL_L_X4Y114_SLICE_X5Y114_BO6;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_C = CLBLL_L_X4Y114_SLICE_X5Y114_CO6;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_D = CLBLL_L_X4Y114_SLICE_X5Y114_DO6;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_AMUX = CLBLL_L_X4Y114_SLICE_X5Y114_AO5;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_A = CLBLL_L_X4Y115_SLICE_X4Y115_AO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_B = CLBLL_L_X4Y115_SLICE_X4Y115_BO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_C = CLBLL_L_X4Y115_SLICE_X4Y115_CO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_D = CLBLL_L_X4Y115_SLICE_X4Y115_DO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_AMUX = CLBLL_L_X4Y115_SLICE_X4Y115_AO5;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_A = CLBLL_L_X4Y115_SLICE_X5Y115_AO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_B = CLBLL_L_X4Y115_SLICE_X5Y115_BO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_C = CLBLL_L_X4Y115_SLICE_X5Y115_CO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_D = CLBLL_L_X4Y115_SLICE_X5Y115_DO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_AMUX = CLBLL_L_X4Y115_SLICE_X5Y115_AO5;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_A = CLBLL_L_X4Y116_SLICE_X4Y116_AO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_B = CLBLL_L_X4Y116_SLICE_X4Y116_BO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_C = CLBLL_L_X4Y116_SLICE_X4Y116_CO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_D = CLBLL_L_X4Y116_SLICE_X4Y116_DO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_AMUX = CLBLL_L_X4Y116_SLICE_X4Y116_AO5;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_A = CLBLL_L_X4Y116_SLICE_X5Y116_AO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_B = CLBLL_L_X4Y116_SLICE_X5Y116_BO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_C = CLBLL_L_X4Y116_SLICE_X5Y116_CO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_D = CLBLL_L_X4Y116_SLICE_X5Y116_DO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_AMUX = CLBLL_L_X4Y116_SLICE_X5Y116_AO5;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_BMUX = CLBLL_L_X4Y116_SLICE_X5Y116_BO5;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_CMUX = CLBLL_L_X4Y116_SLICE_X5Y116_CO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_DMUX = CLBLL_L_X4Y116_SLICE_X5Y116_DO6;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_A = CLBLM_L_X8Y104_SLICE_X10Y104_AO6;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_B = CLBLM_L_X8Y104_SLICE_X10Y104_BO6;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_C = CLBLM_L_X8Y104_SLICE_X10Y104_CO6;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_D = CLBLM_L_X8Y104_SLICE_X10Y104_DO6;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_A = CLBLM_L_X8Y104_SLICE_X11Y104_AO6;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_B = CLBLM_L_X8Y104_SLICE_X11Y104_BO6;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_C = CLBLM_L_X8Y104_SLICE_X11Y104_CO6;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_D = CLBLM_L_X8Y104_SLICE_X11Y104_DO6;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_A = CLBLM_L_X8Y105_SLICE_X10Y105_AO6;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_B = CLBLM_L_X8Y105_SLICE_X10Y105_BO6;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_C = CLBLM_L_X8Y105_SLICE_X10Y105_CO6;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_D = CLBLM_L_X8Y105_SLICE_X10Y105_DO6;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_AMUX = CLBLM_L_X8Y105_SLICE_X10Y105_AO5;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_BMUX = CLBLM_L_X8Y105_SLICE_X10Y105_BO6;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_A = CLBLM_L_X8Y105_SLICE_X11Y105_AO6;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_B = CLBLM_L_X8Y105_SLICE_X11Y105_BO6;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_C = CLBLM_L_X8Y105_SLICE_X11Y105_CO6;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_D = CLBLM_L_X8Y105_SLICE_X11Y105_DO6;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_A = CLBLM_L_X8Y106_SLICE_X10Y106_AO6;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_B = CLBLM_L_X8Y106_SLICE_X10Y106_BO6;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_C = CLBLM_L_X8Y106_SLICE_X10Y106_CO6;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_D = CLBLM_L_X8Y106_SLICE_X10Y106_DO6;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_A = CLBLM_L_X8Y106_SLICE_X11Y106_AO6;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_B = CLBLM_L_X8Y106_SLICE_X11Y106_BO6;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_C = CLBLM_L_X8Y106_SLICE_X11Y106_CO6;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_D = CLBLM_L_X8Y106_SLICE_X11Y106_DO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_A = CLBLM_L_X8Y107_SLICE_X10Y107_AO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_B = CLBLM_L_X8Y107_SLICE_X10Y107_BO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_C = CLBLM_L_X8Y107_SLICE_X10Y107_CO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_D = CLBLM_L_X8Y107_SLICE_X10Y107_DO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_AMUX = CLBLM_L_X8Y107_SLICE_X10Y107_AO5;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_A = CLBLM_L_X8Y107_SLICE_X11Y107_AO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_B = CLBLM_L_X8Y107_SLICE_X11Y107_BO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_C = CLBLM_L_X8Y107_SLICE_X11Y107_CO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_D = CLBLM_L_X8Y107_SLICE_X11Y107_DO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_AMUX = CLBLM_L_X8Y107_SLICE_X11Y107_AO5;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_A = CLBLM_L_X8Y108_SLICE_X10Y108_AO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_B = CLBLM_L_X8Y108_SLICE_X10Y108_BO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_C = CLBLM_L_X8Y108_SLICE_X10Y108_CO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_D = CLBLM_L_X8Y108_SLICE_X10Y108_DO6;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_A = CLBLM_L_X8Y108_SLICE_X11Y108_AO6;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_B = CLBLM_L_X8Y108_SLICE_X11Y108_BO6;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_C = CLBLM_L_X8Y108_SLICE_X11Y108_CO6;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_D = CLBLM_L_X8Y108_SLICE_X11Y108_DO6;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_AMUX = CLBLM_L_X8Y108_SLICE_X11Y108_AO5;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_A = CLBLM_L_X8Y109_SLICE_X10Y109_AO6;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_B = CLBLM_L_X8Y109_SLICE_X10Y109_BO6;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_C = CLBLM_L_X8Y109_SLICE_X10Y109_CO6;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_D = CLBLM_L_X8Y109_SLICE_X10Y109_DO6;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_A = CLBLM_L_X8Y109_SLICE_X11Y109_AO6;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_B = CLBLM_L_X8Y109_SLICE_X11Y109_BO6;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_C = CLBLM_L_X8Y109_SLICE_X11Y109_CO6;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_D = CLBLM_L_X8Y109_SLICE_X11Y109_DO6;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_AMUX = CLBLM_L_X8Y109_SLICE_X11Y109_AO5;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_A = CLBLM_L_X8Y110_SLICE_X10Y110_AO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_B = CLBLM_L_X8Y110_SLICE_X10Y110_BO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_C = CLBLM_L_X8Y110_SLICE_X10Y110_CO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_D = CLBLM_L_X8Y110_SLICE_X10Y110_DO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_AMUX = CLBLM_L_X8Y110_SLICE_X10Y110_AO5;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_A = CLBLM_L_X8Y110_SLICE_X11Y110_AO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_B = CLBLM_L_X8Y110_SLICE_X11Y110_BO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_C = CLBLM_L_X8Y110_SLICE_X11Y110_CO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_D = CLBLM_L_X8Y110_SLICE_X11Y110_DO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_BMUX = CLBLM_L_X8Y110_SLICE_X11Y110_BO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_A = CLBLM_L_X8Y111_SLICE_X10Y111_AO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_B = CLBLM_L_X8Y111_SLICE_X10Y111_BO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_C = CLBLM_L_X8Y111_SLICE_X10Y111_CO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_D = CLBLM_L_X8Y111_SLICE_X10Y111_DO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_AMUX = CLBLM_L_X8Y111_SLICE_X10Y111_AO5;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_A = CLBLM_L_X8Y111_SLICE_X11Y111_AO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_B = CLBLM_L_X8Y111_SLICE_X11Y111_BO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_C = CLBLM_L_X8Y111_SLICE_X11Y111_CO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_D = CLBLM_L_X8Y111_SLICE_X11Y111_DO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_A = CLBLM_L_X8Y112_SLICE_X10Y112_AO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_B = CLBLM_L_X8Y112_SLICE_X10Y112_BO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_C = CLBLM_L_X8Y112_SLICE_X10Y112_CO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_D = CLBLM_L_X8Y112_SLICE_X10Y112_DO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_AMUX = CLBLM_L_X8Y112_SLICE_X10Y112_AO5;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_A = CLBLM_L_X8Y112_SLICE_X11Y112_AO6;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_B = CLBLM_L_X8Y112_SLICE_X11Y112_BO6;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_C = CLBLM_L_X8Y112_SLICE_X11Y112_CO6;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_D = CLBLM_L_X8Y112_SLICE_X11Y112_DO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_A = CLBLM_L_X8Y113_SLICE_X10Y113_AO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_B = CLBLM_L_X8Y113_SLICE_X10Y113_BO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_C = CLBLM_L_X8Y113_SLICE_X10Y113_CO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_D = CLBLM_L_X8Y113_SLICE_X10Y113_DO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_AMUX = CLBLM_L_X8Y113_SLICE_X10Y113_AO5;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_A = CLBLM_L_X8Y113_SLICE_X11Y113_AO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_B = CLBLM_L_X8Y113_SLICE_X11Y113_BO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_C = CLBLM_L_X8Y113_SLICE_X11Y113_CO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_D = CLBLM_L_X8Y113_SLICE_X11Y113_DO6;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_A = CLBLM_L_X8Y114_SLICE_X10Y114_AO6;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_B = CLBLM_L_X8Y114_SLICE_X10Y114_BO6;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_C = CLBLM_L_X8Y114_SLICE_X10Y114_CO6;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_D = CLBLM_L_X8Y114_SLICE_X10Y114_DO6;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_A = CLBLM_L_X8Y114_SLICE_X11Y114_AO6;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_B = CLBLM_L_X8Y114_SLICE_X11Y114_BO6;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_C = CLBLM_L_X8Y114_SLICE_X11Y114_CO6;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_D = CLBLM_L_X8Y114_SLICE_X11Y114_DO6;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_A = CLBLM_L_X8Y115_SLICE_X10Y115_AO6;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_B = CLBLM_L_X8Y115_SLICE_X10Y115_BO6;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_C = CLBLM_L_X8Y115_SLICE_X10Y115_CO6;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_D = CLBLM_L_X8Y115_SLICE_X10Y115_DO6;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_AMUX = CLBLM_L_X8Y115_SLICE_X10Y115_AO5;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_CMUX = CLBLM_L_X8Y115_SLICE_X10Y115_CO6;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_A = CLBLM_L_X8Y115_SLICE_X11Y115_AO6;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_B = CLBLM_L_X8Y115_SLICE_X11Y115_BO6;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_C = CLBLM_L_X8Y115_SLICE_X11Y115_CO6;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_D = CLBLM_L_X8Y115_SLICE_X11Y115_DO6;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_A = CLBLM_L_X8Y116_SLICE_X10Y116_AO6;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_B = CLBLM_L_X8Y116_SLICE_X10Y116_BO6;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_C = CLBLM_L_X8Y116_SLICE_X10Y116_CO6;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_D = CLBLM_L_X8Y116_SLICE_X10Y116_DO6;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_AMUX = CLBLM_L_X8Y116_SLICE_X10Y116_AO5;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_A = CLBLM_L_X8Y116_SLICE_X11Y116_AO6;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_B = CLBLM_L_X8Y116_SLICE_X11Y116_BO6;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_C = CLBLM_L_X8Y116_SLICE_X11Y116_CO6;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_D = CLBLM_L_X8Y116_SLICE_X11Y116_DO6;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_A = CLBLM_L_X10Y105_SLICE_X12Y105_AO6;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_B = CLBLM_L_X10Y105_SLICE_X12Y105_BO6;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_C = CLBLM_L_X10Y105_SLICE_X12Y105_CO6;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_D = CLBLM_L_X10Y105_SLICE_X12Y105_DO6;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_CMUX = CLBLM_L_X10Y105_SLICE_X12Y105_CO6;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_A = CLBLM_L_X10Y105_SLICE_X13Y105_AO6;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_B = CLBLM_L_X10Y105_SLICE_X13Y105_BO6;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_C = CLBLM_L_X10Y105_SLICE_X13Y105_CO6;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_D = CLBLM_L_X10Y105_SLICE_X13Y105_DO6;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_AMUX = CLBLM_L_X10Y105_SLICE_X13Y105_AO5;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_A = CLBLM_L_X10Y106_SLICE_X12Y106_AO6;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_B = CLBLM_L_X10Y106_SLICE_X12Y106_BO6;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_C = CLBLM_L_X10Y106_SLICE_X12Y106_CO6;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_D = CLBLM_L_X10Y106_SLICE_X12Y106_DO6;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_AMUX = CLBLM_L_X10Y106_SLICE_X12Y106_AO5;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_A = CLBLM_L_X10Y106_SLICE_X13Y106_AO6;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_B = CLBLM_L_X10Y106_SLICE_X13Y106_BO6;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_C = CLBLM_L_X10Y106_SLICE_X13Y106_CO6;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_D = CLBLM_L_X10Y106_SLICE_X13Y106_DO6;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_AMUX = CLBLM_L_X10Y106_SLICE_X13Y106_AO5;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_A = CLBLM_L_X10Y107_SLICE_X12Y107_AO6;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_B = CLBLM_L_X10Y107_SLICE_X12Y107_BO6;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_C = CLBLM_L_X10Y107_SLICE_X12Y107_CO6;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_D = CLBLM_L_X10Y107_SLICE_X12Y107_DO6;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_A = CLBLM_L_X10Y107_SLICE_X13Y107_AO6;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_B = CLBLM_L_X10Y107_SLICE_X13Y107_BO6;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_C = CLBLM_L_X10Y107_SLICE_X13Y107_CO6;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_D = CLBLM_L_X10Y107_SLICE_X13Y107_DO6;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_BMUX = CLBLM_L_X10Y107_SLICE_X13Y107_BO6;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_CMUX = CLBLM_L_X10Y107_SLICE_X13Y107_CO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_A = CLBLM_L_X10Y108_SLICE_X12Y108_AO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_B = CLBLM_L_X10Y108_SLICE_X12Y108_BO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_C = CLBLM_L_X10Y108_SLICE_X12Y108_CO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_D = CLBLM_L_X10Y108_SLICE_X12Y108_DO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_AMUX = CLBLM_L_X10Y108_SLICE_X12Y108_AO5;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_A = CLBLM_L_X10Y108_SLICE_X13Y108_AO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_B = CLBLM_L_X10Y108_SLICE_X13Y108_BO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_C = CLBLM_L_X10Y108_SLICE_X13Y108_CO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_D = CLBLM_L_X10Y108_SLICE_X13Y108_DO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_AMUX = CLBLM_L_X10Y108_SLICE_X13Y108_AO5;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_CMUX = CLBLM_L_X10Y108_SLICE_X13Y108_CO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_A = CLBLM_L_X10Y109_SLICE_X12Y109_AO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_B = CLBLM_L_X10Y109_SLICE_X12Y109_BO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_C = CLBLM_L_X10Y109_SLICE_X12Y109_CO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_D = CLBLM_L_X10Y109_SLICE_X12Y109_DO6;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_A = CLBLM_L_X10Y109_SLICE_X13Y109_AO6;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_B = CLBLM_L_X10Y109_SLICE_X13Y109_BO6;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_C = CLBLM_L_X10Y109_SLICE_X13Y109_CO6;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_D = CLBLM_L_X10Y109_SLICE_X13Y109_DO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_A = CLBLM_L_X10Y110_SLICE_X12Y110_AO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_B = CLBLM_L_X10Y110_SLICE_X12Y110_BO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_C = CLBLM_L_X10Y110_SLICE_X12Y110_CO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_D = CLBLM_L_X10Y110_SLICE_X12Y110_DO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_AMUX = CLBLM_L_X10Y110_SLICE_X12Y110_AO5;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_BMUX = CLBLM_L_X10Y110_SLICE_X12Y110_BO5;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_A = CLBLM_L_X10Y110_SLICE_X13Y110_AO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_B = CLBLM_L_X10Y110_SLICE_X13Y110_BO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_C = CLBLM_L_X10Y110_SLICE_X13Y110_CO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_D = CLBLM_L_X10Y110_SLICE_X13Y110_DO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_AMUX = CLBLM_L_X10Y110_SLICE_X13Y110_AO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_A = CLBLM_L_X10Y111_SLICE_X12Y111_AO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_B = CLBLM_L_X10Y111_SLICE_X12Y111_BO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_C = CLBLM_L_X10Y111_SLICE_X12Y111_CO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_D = CLBLM_L_X10Y111_SLICE_X12Y111_DO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_AMUX = CLBLM_L_X10Y111_SLICE_X12Y111_AO5;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_A = CLBLM_L_X10Y111_SLICE_X13Y111_AO6;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_B = CLBLM_L_X10Y111_SLICE_X13Y111_BO6;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_C = CLBLM_L_X10Y111_SLICE_X13Y111_CO6;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_D = CLBLM_L_X10Y111_SLICE_X13Y111_DO6;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_AMUX = CLBLM_L_X10Y111_SLICE_X13Y111_AO5;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_A = CLBLM_L_X10Y112_SLICE_X12Y112_AO6;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_B = CLBLM_L_X10Y112_SLICE_X12Y112_BO6;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_C = CLBLM_L_X10Y112_SLICE_X12Y112_CO6;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_D = CLBLM_L_X10Y112_SLICE_X12Y112_DO6;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_AMUX = CLBLM_L_X10Y112_SLICE_X12Y112_AO5;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_A = CLBLM_L_X10Y112_SLICE_X13Y112_AO6;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_B = CLBLM_L_X10Y112_SLICE_X13Y112_BO6;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_C = CLBLM_L_X10Y112_SLICE_X13Y112_CO6;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_D = CLBLM_L_X10Y112_SLICE_X13Y112_DO6;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_AMUX = CLBLM_L_X10Y112_SLICE_X13Y112_AO5;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_DMUX = CLBLM_L_X10Y112_SLICE_X13Y112_DO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_A = CLBLM_L_X10Y113_SLICE_X12Y113_AO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_B = CLBLM_L_X10Y113_SLICE_X12Y113_BO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_C = CLBLM_L_X10Y113_SLICE_X12Y113_CO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_D = CLBLM_L_X10Y113_SLICE_X12Y113_DO6;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_A = CLBLM_L_X10Y113_SLICE_X13Y113_AO6;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_B = CLBLM_L_X10Y113_SLICE_X13Y113_BO6;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_C = CLBLM_L_X10Y113_SLICE_X13Y113_CO6;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_D = CLBLM_L_X10Y113_SLICE_X13Y113_DO6;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_AMUX = CLBLM_L_X10Y113_SLICE_X13Y113_AO5;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_A = CLBLM_L_X10Y114_SLICE_X12Y114_AO6;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_B = CLBLM_L_X10Y114_SLICE_X12Y114_BO6;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_C = CLBLM_L_X10Y114_SLICE_X12Y114_CO6;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_D = CLBLM_L_X10Y114_SLICE_X12Y114_DO6;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_A = CLBLM_L_X10Y114_SLICE_X13Y114_AO6;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_B = CLBLM_L_X10Y114_SLICE_X13Y114_BO6;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_C = CLBLM_L_X10Y114_SLICE_X13Y114_CO6;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_D = CLBLM_L_X10Y114_SLICE_X13Y114_DO6;
  assign CLBLM_L_X12Y105_SLICE_X16Y105_A = CLBLM_L_X12Y105_SLICE_X16Y105_AO6;
  assign CLBLM_L_X12Y105_SLICE_X16Y105_B = CLBLM_L_X12Y105_SLICE_X16Y105_BO6;
  assign CLBLM_L_X12Y105_SLICE_X16Y105_C = CLBLM_L_X12Y105_SLICE_X16Y105_CO6;
  assign CLBLM_L_X12Y105_SLICE_X16Y105_D = CLBLM_L_X12Y105_SLICE_X16Y105_DO6;
  assign CLBLM_L_X12Y105_SLICE_X16Y105_AMUX = CLBLM_L_X12Y105_SLICE_X16Y105_AO5;
  assign CLBLM_L_X12Y105_SLICE_X17Y105_A = CLBLM_L_X12Y105_SLICE_X17Y105_AO6;
  assign CLBLM_L_X12Y105_SLICE_X17Y105_B = CLBLM_L_X12Y105_SLICE_X17Y105_BO6;
  assign CLBLM_L_X12Y105_SLICE_X17Y105_C = CLBLM_L_X12Y105_SLICE_X17Y105_CO6;
  assign CLBLM_L_X12Y105_SLICE_X17Y105_D = CLBLM_L_X12Y105_SLICE_X17Y105_DO6;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_A = CLBLM_L_X12Y106_SLICE_X16Y106_AO6;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_B = CLBLM_L_X12Y106_SLICE_X16Y106_BO6;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_C = CLBLM_L_X12Y106_SLICE_X16Y106_CO6;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_D = CLBLM_L_X12Y106_SLICE_X16Y106_DO6;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_AMUX = CLBLM_L_X12Y106_SLICE_X16Y106_AO5;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_A = CLBLM_L_X12Y106_SLICE_X17Y106_AO6;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_B = CLBLM_L_X12Y106_SLICE_X17Y106_BO6;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_C = CLBLM_L_X12Y106_SLICE_X17Y106_CO6;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_D = CLBLM_L_X12Y106_SLICE_X17Y106_DO6;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_A = CLBLM_L_X12Y107_SLICE_X16Y107_AO6;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_B = CLBLM_L_X12Y107_SLICE_X16Y107_BO6;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_C = CLBLM_L_X12Y107_SLICE_X16Y107_CO6;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_D = CLBLM_L_X12Y107_SLICE_X16Y107_DO6;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_AMUX = CLBLM_L_X12Y107_SLICE_X16Y107_AO5;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_CMUX = CLBLM_L_X12Y107_SLICE_X16Y107_CO6;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_A = CLBLM_L_X12Y107_SLICE_X17Y107_AO6;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_B = CLBLM_L_X12Y107_SLICE_X17Y107_BO6;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_C = CLBLM_L_X12Y107_SLICE_X17Y107_CO6;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_D = CLBLM_L_X12Y107_SLICE_X17Y107_DO6;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_A = CLBLM_L_X12Y108_SLICE_X16Y108_AO6;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_B = CLBLM_L_X12Y108_SLICE_X16Y108_BO6;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_C = CLBLM_L_X12Y108_SLICE_X16Y108_CO6;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_D = CLBLM_L_X12Y108_SLICE_X16Y108_DO6;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_AMUX = CLBLM_L_X12Y108_SLICE_X16Y108_AO5;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_BMUX = CLBLM_L_X12Y108_SLICE_X16Y108_BO5;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_A = CLBLM_L_X12Y108_SLICE_X17Y108_AO6;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_B = CLBLM_L_X12Y108_SLICE_X17Y108_BO6;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_C = CLBLM_L_X12Y108_SLICE_X17Y108_CO6;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_D = CLBLM_L_X12Y108_SLICE_X17Y108_DO6;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_AMUX = CLBLM_L_X12Y108_SLICE_X17Y108_AO5;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_A = CLBLM_L_X12Y109_SLICE_X16Y109_AO6;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_B = CLBLM_L_X12Y109_SLICE_X16Y109_BO6;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_C = CLBLM_L_X12Y109_SLICE_X16Y109_CO6;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_D = CLBLM_L_X12Y109_SLICE_X16Y109_DO6;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_AMUX = CLBLM_L_X12Y109_SLICE_X16Y109_AO5;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_A = CLBLM_L_X12Y109_SLICE_X17Y109_AO6;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_B = CLBLM_L_X12Y109_SLICE_X17Y109_BO6;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_C = CLBLM_L_X12Y109_SLICE_X17Y109_CO6;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_D = CLBLM_L_X12Y109_SLICE_X17Y109_DO6;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_AMUX = CLBLM_L_X12Y109_SLICE_X17Y109_AO5;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_A = CLBLM_L_X12Y110_SLICE_X16Y110_AO6;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_B = CLBLM_L_X12Y110_SLICE_X16Y110_BO6;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_C = CLBLM_L_X12Y110_SLICE_X16Y110_CO6;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_D = CLBLM_L_X12Y110_SLICE_X16Y110_DO6;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_AMUX = CLBLM_L_X12Y110_SLICE_X16Y110_AO5;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_A = CLBLM_L_X12Y110_SLICE_X17Y110_AO6;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_B = CLBLM_L_X12Y110_SLICE_X17Y110_BO6;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_C = CLBLM_L_X12Y110_SLICE_X17Y110_CO6;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_D = CLBLM_L_X12Y110_SLICE_X17Y110_DO6;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_A = CLBLM_L_X12Y111_SLICE_X16Y111_AO6;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_B = CLBLM_L_X12Y111_SLICE_X16Y111_BO6;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_C = CLBLM_L_X12Y111_SLICE_X16Y111_CO6;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_D = CLBLM_L_X12Y111_SLICE_X16Y111_DO6;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_A = CLBLM_L_X12Y111_SLICE_X17Y111_AO6;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_B = CLBLM_L_X12Y111_SLICE_X17Y111_BO6;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_C = CLBLM_L_X12Y111_SLICE_X17Y111_CO6;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_D = CLBLM_L_X12Y111_SLICE_X17Y111_DO6;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_A = CLBLM_R_X3Y104_SLICE_X2Y104_AO6;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_B = CLBLM_R_X3Y104_SLICE_X2Y104_BO6;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_C = CLBLM_R_X3Y104_SLICE_X2Y104_CO6;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_D = CLBLM_R_X3Y104_SLICE_X2Y104_DO6;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_A = CLBLM_R_X3Y104_SLICE_X3Y104_AO6;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_B = CLBLM_R_X3Y104_SLICE_X3Y104_BO6;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_C = CLBLM_R_X3Y104_SLICE_X3Y104_CO6;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_D = CLBLM_R_X3Y104_SLICE_X3Y104_DO6;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_AMUX = CLBLM_R_X3Y104_SLICE_X3Y104_AO5;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_A = CLBLM_R_X3Y105_SLICE_X2Y105_AO6;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_B = CLBLM_R_X3Y105_SLICE_X2Y105_BO6;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_C = CLBLM_R_X3Y105_SLICE_X2Y105_CO6;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_D = CLBLM_R_X3Y105_SLICE_X2Y105_DO6;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_A = CLBLM_R_X3Y105_SLICE_X3Y105_AO6;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_B = CLBLM_R_X3Y105_SLICE_X3Y105_BO6;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_C = CLBLM_R_X3Y105_SLICE_X3Y105_CO6;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_D = CLBLM_R_X3Y105_SLICE_X3Y105_DO6;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_AMUX = CLBLM_R_X3Y105_SLICE_X3Y105_AO5;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_BMUX = CLBLM_R_X3Y105_SLICE_X3Y105_BO5;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_A = CLBLM_R_X3Y106_SLICE_X2Y106_AO6;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_B = CLBLM_R_X3Y106_SLICE_X2Y106_BO6;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_C = CLBLM_R_X3Y106_SLICE_X2Y106_CO6;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_D = CLBLM_R_X3Y106_SLICE_X2Y106_DO6;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_AMUX = CLBLM_R_X3Y106_SLICE_X2Y106_AO5;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_A = CLBLM_R_X3Y106_SLICE_X3Y106_AO6;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_B = CLBLM_R_X3Y106_SLICE_X3Y106_BO6;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_C = CLBLM_R_X3Y106_SLICE_X3Y106_CO6;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_D = CLBLM_R_X3Y106_SLICE_X3Y106_DO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_A = CLBLM_R_X3Y107_SLICE_X2Y107_AO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_B = CLBLM_R_X3Y107_SLICE_X2Y107_BO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_C = CLBLM_R_X3Y107_SLICE_X2Y107_CO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_D = CLBLM_R_X3Y107_SLICE_X2Y107_DO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_AMUX = CLBLM_R_X3Y107_SLICE_X2Y107_AO5;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_CMUX = CLBLM_R_X3Y107_SLICE_X2Y107_CO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_A = CLBLM_R_X3Y107_SLICE_X3Y107_AO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_B = CLBLM_R_X3Y107_SLICE_X3Y107_BO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_C = CLBLM_R_X3Y107_SLICE_X3Y107_CO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_D = CLBLM_R_X3Y107_SLICE_X3Y107_DO6;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_A = CLBLM_R_X3Y108_SLICE_X2Y108_AO6;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_B = CLBLM_R_X3Y108_SLICE_X2Y108_BO6;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_C = CLBLM_R_X3Y108_SLICE_X2Y108_CO6;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_D = CLBLM_R_X3Y108_SLICE_X2Y108_DO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_A = CLBLM_R_X3Y108_SLICE_X3Y108_AO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_B = CLBLM_R_X3Y108_SLICE_X3Y108_BO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_C = CLBLM_R_X3Y108_SLICE_X3Y108_CO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_D = CLBLM_R_X3Y108_SLICE_X3Y108_DO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_A = CLBLM_R_X3Y109_SLICE_X2Y109_AO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_B = CLBLM_R_X3Y109_SLICE_X2Y109_BO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_C = CLBLM_R_X3Y109_SLICE_X2Y109_CO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_D = CLBLM_R_X3Y109_SLICE_X2Y109_DO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_A = CLBLM_R_X3Y109_SLICE_X3Y109_AO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_B = CLBLM_R_X3Y109_SLICE_X3Y109_BO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_C = CLBLM_R_X3Y109_SLICE_X3Y109_CO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_D = CLBLM_R_X3Y109_SLICE_X3Y109_DO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_A = CLBLM_R_X3Y110_SLICE_X2Y110_AO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_B = CLBLM_R_X3Y110_SLICE_X2Y110_BO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_C = CLBLM_R_X3Y110_SLICE_X2Y110_CO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_D = CLBLM_R_X3Y110_SLICE_X2Y110_DO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_A = CLBLM_R_X3Y110_SLICE_X3Y110_AO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_B = CLBLM_R_X3Y110_SLICE_X3Y110_BO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_C = CLBLM_R_X3Y110_SLICE_X3Y110_CO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_D = CLBLM_R_X3Y110_SLICE_X3Y110_DO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_AMUX = CLBLM_R_X3Y110_SLICE_X3Y110_AO5;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_DMUX = CLBLM_R_X3Y110_SLICE_X3Y110_DO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_A = CLBLM_R_X3Y111_SLICE_X2Y111_AO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_B = CLBLM_R_X3Y111_SLICE_X2Y111_BO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_C = CLBLM_R_X3Y111_SLICE_X2Y111_CO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_D = CLBLM_R_X3Y111_SLICE_X2Y111_DO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_AMUX = CLBLM_R_X3Y111_SLICE_X2Y111_AO5;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_A = CLBLM_R_X3Y111_SLICE_X3Y111_AO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_B = CLBLM_R_X3Y111_SLICE_X3Y111_BO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_C = CLBLM_R_X3Y111_SLICE_X3Y111_CO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_D = CLBLM_R_X3Y111_SLICE_X3Y111_DO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_AMUX = CLBLM_R_X3Y111_SLICE_X3Y111_AO5;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_DMUX = CLBLM_R_X3Y111_SLICE_X3Y111_DO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_A = CLBLM_R_X3Y112_SLICE_X2Y112_AO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_B = CLBLM_R_X3Y112_SLICE_X2Y112_BO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_C = CLBLM_R_X3Y112_SLICE_X2Y112_CO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_D = CLBLM_R_X3Y112_SLICE_X2Y112_DO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_AMUX = CLBLM_R_X3Y112_SLICE_X2Y112_AO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_A = CLBLM_R_X3Y112_SLICE_X3Y112_AO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_B = CLBLM_R_X3Y112_SLICE_X3Y112_BO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_C = CLBLM_R_X3Y112_SLICE_X3Y112_CO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_D = CLBLM_R_X3Y112_SLICE_X3Y112_DO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_A = CLBLM_R_X3Y113_SLICE_X2Y113_AO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_B = CLBLM_R_X3Y113_SLICE_X2Y113_BO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_C = CLBLM_R_X3Y113_SLICE_X2Y113_CO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_D = CLBLM_R_X3Y113_SLICE_X2Y113_DO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_A = CLBLM_R_X3Y113_SLICE_X3Y113_AO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_B = CLBLM_R_X3Y113_SLICE_X3Y113_BO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_C = CLBLM_R_X3Y113_SLICE_X3Y113_CO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_D = CLBLM_R_X3Y113_SLICE_X3Y113_DO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_AMUX = CLBLM_R_X3Y113_SLICE_X3Y113_AO5;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_A = CLBLM_R_X3Y114_SLICE_X2Y114_AO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_B = CLBLM_R_X3Y114_SLICE_X2Y114_BO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_C = CLBLM_R_X3Y114_SLICE_X2Y114_CO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_D = CLBLM_R_X3Y114_SLICE_X2Y114_DO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_A = CLBLM_R_X3Y114_SLICE_X3Y114_AO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_B = CLBLM_R_X3Y114_SLICE_X3Y114_BO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_C = CLBLM_R_X3Y114_SLICE_X3Y114_CO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_D = CLBLM_R_X3Y114_SLICE_X3Y114_DO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_AMUX = CLBLM_R_X3Y114_SLICE_X3Y114_AO5;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_A = CLBLM_R_X5Y104_SLICE_X6Y104_AO6;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_B = CLBLM_R_X5Y104_SLICE_X6Y104_BO6;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_C = CLBLM_R_X5Y104_SLICE_X6Y104_CO6;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_D = CLBLM_R_X5Y104_SLICE_X6Y104_DO6;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_A = CLBLM_R_X5Y104_SLICE_X7Y104_AO6;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_B = CLBLM_R_X5Y104_SLICE_X7Y104_BO6;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_C = CLBLM_R_X5Y104_SLICE_X7Y104_CO6;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_D = CLBLM_R_X5Y104_SLICE_X7Y104_DO6;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_A = CLBLM_R_X5Y105_SLICE_X6Y105_AO6;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_B = CLBLM_R_X5Y105_SLICE_X6Y105_BO6;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_C = CLBLM_R_X5Y105_SLICE_X6Y105_CO6;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_D = CLBLM_R_X5Y105_SLICE_X6Y105_DO6;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_A = CLBLM_R_X5Y105_SLICE_X7Y105_AO6;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_B = CLBLM_R_X5Y105_SLICE_X7Y105_BO6;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_C = CLBLM_R_X5Y105_SLICE_X7Y105_CO6;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_D = CLBLM_R_X5Y105_SLICE_X7Y105_DO6;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_CMUX = CLBLM_R_X5Y105_SLICE_X7Y105_CO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_A = CLBLM_R_X5Y106_SLICE_X6Y106_AO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_B = CLBLM_R_X5Y106_SLICE_X6Y106_BO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_C = CLBLM_R_X5Y106_SLICE_X6Y106_CO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_D = CLBLM_R_X5Y106_SLICE_X6Y106_DO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_AMUX = CLBLM_R_X5Y106_SLICE_X6Y106_AO5;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_BMUX = CLBLM_R_X5Y106_SLICE_X6Y106_BO5;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_CMUX = CLBLM_R_X5Y106_SLICE_X6Y106_CO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_DMUX = CLBLM_R_X5Y106_SLICE_X6Y106_DO6;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_A = CLBLM_R_X5Y106_SLICE_X7Y106_AO6;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_B = CLBLM_R_X5Y106_SLICE_X7Y106_BO6;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_C = CLBLM_R_X5Y106_SLICE_X7Y106_CO6;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_D = CLBLM_R_X5Y106_SLICE_X7Y106_DO6;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_AMUX = CLBLM_R_X5Y106_SLICE_X7Y106_AO5;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_A = CLBLM_R_X5Y107_SLICE_X6Y107_AO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_B = CLBLM_R_X5Y107_SLICE_X6Y107_BO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_C = CLBLM_R_X5Y107_SLICE_X6Y107_CO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_D = CLBLM_R_X5Y107_SLICE_X6Y107_DO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_A = CLBLM_R_X5Y107_SLICE_X7Y107_AO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_B = CLBLM_R_X5Y107_SLICE_X7Y107_BO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_C = CLBLM_R_X5Y107_SLICE_X7Y107_CO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_D = CLBLM_R_X5Y107_SLICE_X7Y107_DO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_AMUX = CLBLM_R_X5Y107_SLICE_X7Y107_AO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_A = CLBLM_R_X5Y108_SLICE_X6Y108_AO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_B = CLBLM_R_X5Y108_SLICE_X6Y108_BO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_C = CLBLM_R_X5Y108_SLICE_X6Y108_CO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_D = CLBLM_R_X5Y108_SLICE_X6Y108_DO6;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_A = CLBLM_R_X5Y108_SLICE_X7Y108_AO6;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_B = CLBLM_R_X5Y108_SLICE_X7Y108_BO6;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_C = CLBLM_R_X5Y108_SLICE_X7Y108_CO6;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_D = CLBLM_R_X5Y108_SLICE_X7Y108_DO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_A = CLBLM_R_X5Y109_SLICE_X6Y109_AO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_B = CLBLM_R_X5Y109_SLICE_X6Y109_BO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_C = CLBLM_R_X5Y109_SLICE_X6Y109_CO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_D = CLBLM_R_X5Y109_SLICE_X6Y109_DO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_AMUX = CLBLM_R_X5Y109_SLICE_X6Y109_AO5;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_A = CLBLM_R_X5Y109_SLICE_X7Y109_AO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_B = CLBLM_R_X5Y109_SLICE_X7Y109_BO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_C = CLBLM_R_X5Y109_SLICE_X7Y109_CO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_D = CLBLM_R_X5Y109_SLICE_X7Y109_DO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_AMUX = CLBLM_R_X5Y109_SLICE_X7Y109_AO5;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_A = CLBLM_R_X5Y110_SLICE_X6Y110_AO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_B = CLBLM_R_X5Y110_SLICE_X6Y110_BO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_C = CLBLM_R_X5Y110_SLICE_X6Y110_CO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_D = CLBLM_R_X5Y110_SLICE_X6Y110_DO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_A = CLBLM_R_X5Y110_SLICE_X7Y110_AO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_B = CLBLM_R_X5Y110_SLICE_X7Y110_BO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_C = CLBLM_R_X5Y110_SLICE_X7Y110_CO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_D = CLBLM_R_X5Y110_SLICE_X7Y110_DO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_AMUX = CLBLM_R_X5Y110_SLICE_X7Y110_AO5;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_BMUX = CLBLM_R_X5Y110_SLICE_X7Y110_BO5;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_A = CLBLM_R_X5Y111_SLICE_X6Y111_AO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_B = CLBLM_R_X5Y111_SLICE_X6Y111_BO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_C = CLBLM_R_X5Y111_SLICE_X6Y111_CO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_D = CLBLM_R_X5Y111_SLICE_X6Y111_DO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_AMUX = CLBLM_R_X5Y111_SLICE_X6Y111_AO5;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_A = CLBLM_R_X5Y111_SLICE_X7Y111_AO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_B = CLBLM_R_X5Y111_SLICE_X7Y111_BO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_C = CLBLM_R_X5Y111_SLICE_X7Y111_CO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_D = CLBLM_R_X5Y111_SLICE_X7Y111_DO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_BMUX = CLBLM_R_X5Y111_SLICE_X7Y111_BO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_A = CLBLM_R_X5Y112_SLICE_X6Y112_AO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_B = CLBLM_R_X5Y112_SLICE_X6Y112_BO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_C = CLBLM_R_X5Y112_SLICE_X6Y112_CO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_D = CLBLM_R_X5Y112_SLICE_X6Y112_DO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_AMUX = CLBLM_R_X5Y112_SLICE_X6Y112_AO5;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_CMUX = CLBLM_R_X5Y112_SLICE_X6Y112_CO6;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_A = CLBLM_R_X5Y112_SLICE_X7Y112_AO6;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_B = CLBLM_R_X5Y112_SLICE_X7Y112_BO6;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_C = CLBLM_R_X5Y112_SLICE_X7Y112_CO6;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_D = CLBLM_R_X5Y112_SLICE_X7Y112_DO6;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_AMUX = CLBLM_R_X5Y112_SLICE_X7Y112_AO5;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_A = CLBLM_R_X5Y113_SLICE_X6Y113_AO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_B = CLBLM_R_X5Y113_SLICE_X6Y113_BO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_C = CLBLM_R_X5Y113_SLICE_X6Y113_CO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_D = CLBLM_R_X5Y113_SLICE_X6Y113_DO6;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_A = CLBLM_R_X5Y113_SLICE_X7Y113_AO6;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_B = CLBLM_R_X5Y113_SLICE_X7Y113_BO6;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_C = CLBLM_R_X5Y113_SLICE_X7Y113_CO6;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_D = CLBLM_R_X5Y113_SLICE_X7Y113_DO6;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_A = CLBLM_R_X5Y114_SLICE_X6Y114_AO6;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_B = CLBLM_R_X5Y114_SLICE_X6Y114_BO6;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_C = CLBLM_R_X5Y114_SLICE_X6Y114_CO6;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_D = CLBLM_R_X5Y114_SLICE_X6Y114_DO6;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_AMUX = CLBLM_R_X5Y114_SLICE_X6Y114_AO5;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_A = CLBLM_R_X5Y114_SLICE_X7Y114_AO6;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_B = CLBLM_R_X5Y114_SLICE_X7Y114_BO6;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_C = CLBLM_R_X5Y114_SLICE_X7Y114_CO6;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_D = CLBLM_R_X5Y114_SLICE_X7Y114_DO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_A = CLBLM_R_X5Y115_SLICE_X6Y115_AO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_B = CLBLM_R_X5Y115_SLICE_X6Y115_BO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_C = CLBLM_R_X5Y115_SLICE_X6Y115_CO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_D = CLBLM_R_X5Y115_SLICE_X6Y115_DO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_AMUX = CLBLM_R_X5Y115_SLICE_X6Y115_AO5;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_A = CLBLM_R_X5Y115_SLICE_X7Y115_AO6;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_B = CLBLM_R_X5Y115_SLICE_X7Y115_BO6;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_C = CLBLM_R_X5Y115_SLICE_X7Y115_CO6;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_D = CLBLM_R_X5Y115_SLICE_X7Y115_DO6;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_AMUX = CLBLM_R_X5Y115_SLICE_X7Y115_AO5;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_A = CLBLM_R_X5Y116_SLICE_X6Y116_AO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_B = CLBLM_R_X5Y116_SLICE_X6Y116_BO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_C = CLBLM_R_X5Y116_SLICE_X6Y116_CO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_D = CLBLM_R_X5Y116_SLICE_X6Y116_DO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_AMUX = CLBLM_R_X5Y116_SLICE_X6Y116_AO6;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_A = CLBLM_R_X5Y116_SLICE_X7Y116_AO6;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_B = CLBLM_R_X5Y116_SLICE_X7Y116_BO6;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_C = CLBLM_R_X5Y116_SLICE_X7Y116_CO6;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_D = CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_AMUX = CLBLM_R_X5Y116_SLICE_X7Y116_AO5;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_BMUX = CLBLM_R_X5Y116_SLICE_X7Y116_BO6;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_A = CLBLM_R_X7Y104_SLICE_X8Y104_AO6;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_B = CLBLM_R_X7Y104_SLICE_X8Y104_BO6;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_C = CLBLM_R_X7Y104_SLICE_X8Y104_CO6;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_D = CLBLM_R_X7Y104_SLICE_X8Y104_DO6;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_A = CLBLM_R_X7Y104_SLICE_X9Y104_AO6;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_B = CLBLM_R_X7Y104_SLICE_X9Y104_BO6;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_C = CLBLM_R_X7Y104_SLICE_X9Y104_CO6;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_D = CLBLM_R_X7Y104_SLICE_X9Y104_DO6;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_AMUX = CLBLM_R_X7Y104_SLICE_X9Y104_AO5;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_CMUX = CLBLM_R_X7Y104_SLICE_X9Y104_CO6;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_A = CLBLM_R_X7Y105_SLICE_X8Y105_AO6;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_B = CLBLM_R_X7Y105_SLICE_X8Y105_BO6;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_C = CLBLM_R_X7Y105_SLICE_X8Y105_CO6;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_D = CLBLM_R_X7Y105_SLICE_X8Y105_DO6;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_AMUX = CLBLM_R_X7Y105_SLICE_X8Y105_AO5;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_BMUX = CLBLM_R_X7Y105_SLICE_X8Y105_BO6;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_A = CLBLM_R_X7Y105_SLICE_X9Y105_AO6;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_B = CLBLM_R_X7Y105_SLICE_X9Y105_BO6;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_C = CLBLM_R_X7Y105_SLICE_X9Y105_CO6;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_D = CLBLM_R_X7Y105_SLICE_X9Y105_DO6;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_A = CLBLM_R_X7Y106_SLICE_X8Y106_AO6;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_B = CLBLM_R_X7Y106_SLICE_X8Y106_BO6;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_C = CLBLM_R_X7Y106_SLICE_X8Y106_CO6;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_D = CLBLM_R_X7Y106_SLICE_X8Y106_DO6;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_AMUX = CLBLM_R_X7Y106_SLICE_X8Y106_AO5;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_BMUX = CLBLM_R_X7Y106_SLICE_X8Y106_BO5;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_CMUX = CLBLM_R_X7Y106_SLICE_X8Y106_CO6;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_A = CLBLM_R_X7Y106_SLICE_X9Y106_AO6;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_B = CLBLM_R_X7Y106_SLICE_X9Y106_BO6;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_C = CLBLM_R_X7Y106_SLICE_X9Y106_CO6;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_D = CLBLM_R_X7Y106_SLICE_X9Y106_DO6;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_AMUX = CLBLM_R_X7Y106_SLICE_X9Y106_AO5;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_A = CLBLM_R_X7Y107_SLICE_X8Y107_AO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_B = CLBLM_R_X7Y107_SLICE_X8Y107_BO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_C = CLBLM_R_X7Y107_SLICE_X8Y107_CO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_D = CLBLM_R_X7Y107_SLICE_X8Y107_DO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_A = CLBLM_R_X7Y107_SLICE_X9Y107_AO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_B = CLBLM_R_X7Y107_SLICE_X9Y107_BO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_C = CLBLM_R_X7Y107_SLICE_X9Y107_CO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_D = CLBLM_R_X7Y107_SLICE_X9Y107_DO6;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_A = CLBLM_R_X7Y108_SLICE_X8Y108_AO6;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_B = CLBLM_R_X7Y108_SLICE_X8Y108_BO6;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_C = CLBLM_R_X7Y108_SLICE_X8Y108_CO6;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_D = CLBLM_R_X7Y108_SLICE_X8Y108_DO6;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_AMUX = CLBLM_R_X7Y108_SLICE_X8Y108_AO5;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_A = CLBLM_R_X7Y108_SLICE_X9Y108_AO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_B = CLBLM_R_X7Y108_SLICE_X9Y108_BO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_C = CLBLM_R_X7Y108_SLICE_X9Y108_CO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_D = CLBLM_R_X7Y108_SLICE_X9Y108_DO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_AMUX = CLBLM_R_X7Y108_SLICE_X9Y108_AO5;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_A = CLBLM_R_X7Y109_SLICE_X8Y109_AO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_B = CLBLM_R_X7Y109_SLICE_X8Y109_BO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_C = CLBLM_R_X7Y109_SLICE_X8Y109_CO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_D = CLBLM_R_X7Y109_SLICE_X8Y109_DO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_AMUX = CLBLM_R_X7Y109_SLICE_X8Y109_AO5;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_A = CLBLM_R_X7Y109_SLICE_X9Y109_AO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_B = CLBLM_R_X7Y109_SLICE_X9Y109_BO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_C = CLBLM_R_X7Y109_SLICE_X9Y109_CO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_D = CLBLM_R_X7Y109_SLICE_X9Y109_DO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_AMUX = CLBLM_R_X7Y109_SLICE_X9Y109_AO5;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_BMUX = CLBLM_R_X7Y109_SLICE_X9Y109_BO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_A = CLBLM_R_X7Y110_SLICE_X8Y110_AO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_B = CLBLM_R_X7Y110_SLICE_X8Y110_BO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_C = CLBLM_R_X7Y110_SLICE_X8Y110_CO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_D = CLBLM_R_X7Y110_SLICE_X8Y110_DO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_A = CLBLM_R_X7Y110_SLICE_X9Y110_AO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_B = CLBLM_R_X7Y110_SLICE_X9Y110_BO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_C = CLBLM_R_X7Y110_SLICE_X9Y110_CO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_D = CLBLM_R_X7Y110_SLICE_X9Y110_DO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_AMUX = CLBLM_R_X7Y110_SLICE_X9Y110_AO5;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_BMUX = CLBLM_R_X7Y110_SLICE_X9Y110_BO5;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_A = CLBLM_R_X7Y111_SLICE_X8Y111_AO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_B = CLBLM_R_X7Y111_SLICE_X8Y111_BO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_C = CLBLM_R_X7Y111_SLICE_X8Y111_CO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_D = CLBLM_R_X7Y111_SLICE_X8Y111_DO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_AMUX = CLBLM_R_X7Y111_SLICE_X8Y111_AO5;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_A = CLBLM_R_X7Y111_SLICE_X9Y111_AO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_B = CLBLM_R_X7Y111_SLICE_X9Y111_BO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_C = CLBLM_R_X7Y111_SLICE_X9Y111_CO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_D = CLBLM_R_X7Y111_SLICE_X9Y111_DO6;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_A = CLBLM_R_X7Y112_SLICE_X8Y112_AO6;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_B = CLBLM_R_X7Y112_SLICE_X8Y112_BO6;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_C = CLBLM_R_X7Y112_SLICE_X8Y112_CO6;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_D = CLBLM_R_X7Y112_SLICE_X8Y112_DO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_A = CLBLM_R_X7Y112_SLICE_X9Y112_AO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_B = CLBLM_R_X7Y112_SLICE_X9Y112_BO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_C = CLBLM_R_X7Y112_SLICE_X9Y112_CO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_D = CLBLM_R_X7Y112_SLICE_X9Y112_DO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_AMUX = CLBLM_R_X7Y112_SLICE_X9Y112_AO5;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_BMUX = CLBLM_R_X7Y112_SLICE_X9Y112_BO5;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_A = CLBLM_R_X7Y113_SLICE_X8Y113_AO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_B = CLBLM_R_X7Y113_SLICE_X8Y113_BO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_C = CLBLM_R_X7Y113_SLICE_X8Y113_CO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_D = CLBLM_R_X7Y113_SLICE_X8Y113_DO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_A = CLBLM_R_X7Y113_SLICE_X9Y113_AO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_B = CLBLM_R_X7Y113_SLICE_X9Y113_BO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_C = CLBLM_R_X7Y113_SLICE_X9Y113_CO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_D = CLBLM_R_X7Y113_SLICE_X9Y113_DO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_A = CLBLM_R_X7Y114_SLICE_X8Y114_AO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_B = CLBLM_R_X7Y114_SLICE_X8Y114_BO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_C = CLBLM_R_X7Y114_SLICE_X8Y114_CO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_D = CLBLM_R_X7Y114_SLICE_X8Y114_DO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_AMUX = CLBLM_R_X7Y114_SLICE_X8Y114_AO5;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_A = CLBLM_R_X7Y114_SLICE_X9Y114_AO6;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_B = CLBLM_R_X7Y114_SLICE_X9Y114_BO6;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_C = CLBLM_R_X7Y114_SLICE_X9Y114_CO6;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_D = CLBLM_R_X7Y114_SLICE_X9Y114_DO6;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_AMUX = CLBLM_R_X7Y114_SLICE_X9Y114_AO5;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_A = CLBLM_R_X7Y115_SLICE_X8Y115_AO6;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_B = CLBLM_R_X7Y115_SLICE_X8Y115_BO6;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_C = CLBLM_R_X7Y115_SLICE_X8Y115_CO6;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_D = CLBLM_R_X7Y115_SLICE_X8Y115_DO6;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_A = CLBLM_R_X7Y115_SLICE_X9Y115_AO6;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_B = CLBLM_R_X7Y115_SLICE_X9Y115_BO6;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_C = CLBLM_R_X7Y115_SLICE_X9Y115_CO6;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_D = CLBLM_R_X7Y115_SLICE_X9Y115_DO6;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_A = CLBLM_R_X7Y116_SLICE_X8Y116_AO6;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_B = CLBLM_R_X7Y116_SLICE_X8Y116_BO6;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_C = CLBLM_R_X7Y116_SLICE_X8Y116_CO6;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_D = CLBLM_R_X7Y116_SLICE_X8Y116_DO6;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_A = CLBLM_R_X7Y116_SLICE_X9Y116_AO6;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_B = CLBLM_R_X7Y116_SLICE_X9Y116_BO6;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_C = CLBLM_R_X7Y116_SLICE_X9Y116_CO6;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_D = CLBLM_R_X7Y116_SLICE_X9Y116_DO6;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_A = CLBLM_R_X11Y105_SLICE_X14Y105_AO6;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_B = CLBLM_R_X11Y105_SLICE_X14Y105_BO6;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_C = CLBLM_R_X11Y105_SLICE_X14Y105_CO6;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_D = CLBLM_R_X11Y105_SLICE_X14Y105_DO6;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_BMUX = CLBLM_R_X11Y105_SLICE_X14Y105_BO6;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_A = CLBLM_R_X11Y105_SLICE_X15Y105_AO6;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_B = CLBLM_R_X11Y105_SLICE_X15Y105_BO6;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_C = CLBLM_R_X11Y105_SLICE_X15Y105_CO6;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_D = CLBLM_R_X11Y105_SLICE_X15Y105_DO6;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_AMUX = CLBLM_R_X11Y105_SLICE_X15Y105_AO5;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_DMUX = CLBLM_R_X11Y105_SLICE_X15Y105_DO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_A = CLBLM_R_X11Y106_SLICE_X14Y106_AO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_B = CLBLM_R_X11Y106_SLICE_X14Y106_BO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_C = CLBLM_R_X11Y106_SLICE_X14Y106_CO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_D = CLBLM_R_X11Y106_SLICE_X14Y106_DO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_AMUX = CLBLM_R_X11Y106_SLICE_X14Y106_AO5;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_A = CLBLM_R_X11Y106_SLICE_X15Y106_AO6;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_B = CLBLM_R_X11Y106_SLICE_X15Y106_BO6;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_C = CLBLM_R_X11Y106_SLICE_X15Y106_CO6;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_D = CLBLM_R_X11Y106_SLICE_X15Y106_DO6;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_AMUX = CLBLM_R_X11Y106_SLICE_X15Y106_AO5;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_A = CLBLM_R_X11Y107_SLICE_X14Y107_AO6;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_B = CLBLM_R_X11Y107_SLICE_X14Y107_BO6;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_C = CLBLM_R_X11Y107_SLICE_X14Y107_CO6;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_D = CLBLM_R_X11Y107_SLICE_X14Y107_DO6;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_AMUX = CLBLM_R_X11Y107_SLICE_X14Y107_AO5;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_BMUX = CLBLM_R_X11Y107_SLICE_X14Y107_BO6;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_A = CLBLM_R_X11Y107_SLICE_X15Y107_AO6;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_B = CLBLM_R_X11Y107_SLICE_X15Y107_BO6;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_C = CLBLM_R_X11Y107_SLICE_X15Y107_CO6;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_D = CLBLM_R_X11Y107_SLICE_X15Y107_DO6;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_AMUX = CLBLM_R_X11Y107_SLICE_X15Y107_AO5;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_A = CLBLM_R_X11Y108_SLICE_X14Y108_AO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_B = CLBLM_R_X11Y108_SLICE_X14Y108_BO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_C = CLBLM_R_X11Y108_SLICE_X14Y108_CO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_D = CLBLM_R_X11Y108_SLICE_X14Y108_DO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_AMUX = CLBLM_R_X11Y108_SLICE_X14Y108_AO5;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_CMUX = CLBLM_R_X11Y108_SLICE_X14Y108_CO6;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_A = CLBLM_R_X11Y108_SLICE_X15Y108_AO6;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_B = CLBLM_R_X11Y108_SLICE_X15Y108_BO6;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_C = CLBLM_R_X11Y108_SLICE_X15Y108_CO6;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_D = CLBLM_R_X11Y108_SLICE_X15Y108_DO6;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_AMUX = CLBLM_R_X11Y108_SLICE_X15Y108_AO5;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_CMUX = CLBLM_R_X11Y108_SLICE_X15Y108_CO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_A = CLBLM_R_X11Y109_SLICE_X14Y109_AO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_B = CLBLM_R_X11Y109_SLICE_X14Y109_BO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_C = CLBLM_R_X11Y109_SLICE_X14Y109_CO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_D = CLBLM_R_X11Y109_SLICE_X14Y109_DO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_AMUX = CLBLM_R_X11Y109_SLICE_X14Y109_AO5;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_CMUX = CLBLM_R_X11Y109_SLICE_X14Y109_CO6;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_A = CLBLM_R_X11Y109_SLICE_X15Y109_AO6;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_B = CLBLM_R_X11Y109_SLICE_X15Y109_BO6;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_C = CLBLM_R_X11Y109_SLICE_X15Y109_CO6;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_D = CLBLM_R_X11Y109_SLICE_X15Y109_DO6;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_AMUX = CLBLM_R_X11Y109_SLICE_X15Y109_AO5;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_A = CLBLM_R_X11Y110_SLICE_X14Y110_AO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_B = CLBLM_R_X11Y110_SLICE_X14Y110_BO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_C = CLBLM_R_X11Y110_SLICE_X14Y110_CO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_D = CLBLM_R_X11Y110_SLICE_X14Y110_DO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_AMUX = CLBLM_R_X11Y110_SLICE_X14Y110_AO5;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_BMUX = CLBLM_R_X11Y110_SLICE_X14Y110_BO5;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_A = CLBLM_R_X11Y110_SLICE_X15Y110_AO6;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_B = CLBLM_R_X11Y110_SLICE_X15Y110_BO6;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_C = CLBLM_R_X11Y110_SLICE_X15Y110_CO6;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_D = CLBLM_R_X11Y110_SLICE_X15Y110_DO6;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_BMUX = CLBLM_R_X11Y110_SLICE_X15Y110_BO6;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_A = CLBLM_R_X11Y111_SLICE_X14Y111_AO6;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_B = CLBLM_R_X11Y111_SLICE_X14Y111_BO6;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_C = CLBLM_R_X11Y111_SLICE_X14Y111_CO6;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_D = CLBLM_R_X11Y111_SLICE_X14Y111_DO6;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_AMUX = CLBLM_R_X11Y111_SLICE_X14Y111_AO5;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_A = CLBLM_R_X11Y111_SLICE_X15Y111_AO6;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_B = CLBLM_R_X11Y111_SLICE_X15Y111_BO6;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_C = CLBLM_R_X11Y111_SLICE_X15Y111_CO6;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_D = CLBLM_R_X11Y111_SLICE_X15Y111_DO6;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_A = CLBLM_R_X11Y112_SLICE_X14Y112_AO6;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_B = CLBLM_R_X11Y112_SLICE_X14Y112_BO6;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_C = CLBLM_R_X11Y112_SLICE_X14Y112_CO6;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_D = CLBLM_R_X11Y112_SLICE_X14Y112_DO6;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_A = CLBLM_R_X11Y112_SLICE_X15Y112_AO6;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_B = CLBLM_R_X11Y112_SLICE_X15Y112_BO6;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_C = CLBLM_R_X11Y112_SLICE_X15Y112_CO6;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_D = CLBLM_R_X11Y112_SLICE_X15Y112_DO6;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_AMUX = CLBLM_R_X11Y112_SLICE_X15Y112_AO5;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_A = CLBLM_R_X11Y113_SLICE_X14Y113_AO6;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_B = CLBLM_R_X11Y113_SLICE_X14Y113_BO6;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_C = CLBLM_R_X11Y113_SLICE_X14Y113_CO6;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_D = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_BMUX = CLBLM_R_X11Y113_SLICE_X14Y113_BO6;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_A = CLBLM_R_X11Y113_SLICE_X15Y113_AO6;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_B = CLBLM_R_X11Y113_SLICE_X15Y113_BO6;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_C = CLBLM_R_X11Y113_SLICE_X15Y113_CO6;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_D = CLBLM_R_X11Y113_SLICE_X15Y113_DO6;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_AMUX = CLBLM_R_X11Y113_SLICE_X15Y113_AO6;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_A = CLBLM_R_X11Y114_SLICE_X14Y114_AO6;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_B = CLBLM_R_X11Y114_SLICE_X14Y114_BO6;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_C = CLBLM_R_X11Y114_SLICE_X14Y114_CO6;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_D = CLBLM_R_X11Y114_SLICE_X14Y114_DO6;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_A = CLBLM_R_X11Y114_SLICE_X15Y114_AO6;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_B = CLBLM_R_X11Y114_SLICE_X15Y114_BO6;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_C = CLBLM_R_X11Y114_SLICE_X15Y114_CO6;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_D = CLBLM_R_X11Y114_SLICE_X15Y114_DO6;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_A = CLBLM_R_X13Y108_SLICE_X18Y108_AO6;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_B = CLBLM_R_X13Y108_SLICE_X18Y108_BO6;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_C = CLBLM_R_X13Y108_SLICE_X18Y108_CO6;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_D = CLBLM_R_X13Y108_SLICE_X18Y108_DO6;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_A = CLBLM_R_X13Y108_SLICE_X19Y108_AO6;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_B = CLBLM_R_X13Y108_SLICE_X19Y108_BO6;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_C = CLBLM_R_X13Y108_SLICE_X19Y108_CO6;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_D = CLBLM_R_X13Y108_SLICE_X19Y108_DO6;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_AMUX = CLBLM_R_X13Y108_SLICE_X19Y108_AO6;
  assign LIOI3_X0Y101_ILOGIC_X0Y102_O = LIOB33_X0Y101_IOB_X0Y102_I;
  assign LIOI3_X0Y101_ILOGIC_X0Y101_O = LIOB33_X0Y101_IOB_X0Y101_I;
  assign LIOI3_X0Y103_ILOGIC_X0Y104_O = LIOB33_X0Y103_IOB_X0Y104_I;
  assign LIOI3_X0Y103_ILOGIC_X0Y103_O = LIOB33_X0Y103_IOB_X0Y103_I;
  assign LIOI3_X0Y105_ILOGIC_X0Y106_O = LIOB33_X0Y105_IOB_X0Y106_I;
  assign LIOI3_X0Y105_ILOGIC_X0Y105_O = LIOB33_X0Y105_IOB_X0Y105_I;
  assign LIOI3_X0Y109_ILOGIC_X0Y110_O = LIOB33_X0Y109_IOB_X0Y110_I;
  assign LIOI3_X0Y109_ILOGIC_X0Y109_O = LIOB33_X0Y109_IOB_X0Y109_I;
  assign LIOI3_X0Y111_ILOGIC_X0Y112_O = LIOB33_X0Y111_IOB_X0Y112_I;
  assign LIOI3_X0Y111_ILOGIC_X0Y111_O = LIOB33_X0Y111_IOB_X0Y111_I;
  assign LIOI3_X0Y115_ILOGIC_X0Y116_O = LIOB33_X0Y115_IOB_X0Y116_I;
  assign LIOI3_X0Y115_ILOGIC_X0Y115_O = LIOB33_X0Y115_IOB_X0Y115_I;
  assign LIOI3_X0Y117_ILOGIC_X0Y117_O = LIOB33_X0Y117_IOB_X0Y117_I;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_OQ = CLBLL_L_X2Y112_SLICE_X0Y112_AO5;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_TQ = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_OQ = CLBLL_L_X2Y108_SLICE_X1Y108_AO6;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_TQ = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_OQ = CLBLL_L_X2Y108_SLICE_X0Y108_AO5;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_TQ = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_OQ = CLBLL_L_X2Y107_SLICE_X1Y107_AO5;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_TQ = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_OQ = CLBLL_L_X2Y108_SLICE_X0Y108_CO6;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_TQ = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_OQ = CLBLM_R_X3Y108_SLICE_X3Y108_AO6;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_TQ = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_OQ = CLBLM_R_X3Y107_SLICE_X2Y107_AO6;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_TQ = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_OQ = CLBLM_R_X3Y110_SLICE_X3Y110_AO6;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_TQ = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_OQ = CLBLL_L_X4Y109_SLICE_X4Y109_AO6;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_TQ = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_OQ = CLBLL_L_X2Y109_SLICE_X0Y109_BO5;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_TQ = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_OQ = CLBLM_R_X3Y110_SLICE_X3Y110_BO6;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_TQ = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_OQ = 1'b0;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_TQ = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_OQ = CLBLL_L_X4Y112_SLICE_X4Y112_AO6;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_TQ = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_OQ = CLBLM_R_X5Y114_SLICE_X6Y114_AO6;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_TQ = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_OQ = CLBLM_R_X5Y114_SLICE_X6Y114_AO5;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_TQ = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_OQ = CLBLL_L_X4Y116_SLICE_X5Y116_BO5;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_TQ = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_OQ = CLBLL_L_X4Y116_SLICE_X5Y116_BO6;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_TQ = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_OQ = CLBLL_L_X4Y116_SLICE_X4Y116_BO6;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_TQ = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_OQ = CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_TQ = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_OQ = CLBLL_L_X4Y113_SLICE_X4Y113_BO6;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_TQ = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_OQ = CLBLL_L_X4Y114_SLICE_X4Y114_AO6;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_TQ = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_OQ = CLBLM_R_X3Y113_SLICE_X3Y113_CO6;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_TQ = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_OQ = CLBLM_R_X3Y113_SLICE_X3Y113_AO6;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_TQ = 1'b1;
  assign LIOI3_SING_X0Y100_ILOGIC_X0Y100_O = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_OQ = CLBLM_R_X3Y113_SLICE_X3Y113_AO5;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y108_O = LIOB33_X0Y107_IOB_X0Y108_I;
  assign LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y107_O = LIOB33_X0Y107_IOB_X0Y107_I;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_OQ = CLBLL_L_X2Y109_SLICE_X0Y109_AO5;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_OQ = CLBLL_L_X2Y112_SLICE_X0Y112_AO6;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_OQ = CLBLM_R_X3Y114_SLICE_X3Y114_AO5;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_OQ = CLBLL_L_X4Y111_SLICE_X4Y111_AO6;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_OQ = CLBLL_L_X4Y116_SLICE_X4Y116_CO6;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_OQ = CLBLL_L_X4Y115_SLICE_X4Y115_DO6;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y114_O = LIOB33_X0Y113_IOB_X0Y114_I;
  assign LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y113_O = LIOB33_X0Y113_IOB_X0Y113_I;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_OQ = CLBLL_L_X4Y116_SLICE_X5Y116_AO5;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_OQ = CLBLL_L_X4Y116_SLICE_X5Y116_AO6;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_TQ = 1'b1;
  assign RIOI3_X105Y101_ILOGIC_X1Y102_O = RIOB33_X105Y101_IOB_X1Y102_I;
  assign RIOI3_X105Y101_ILOGIC_X1Y101_O = RIOB33_X105Y101_IOB_X1Y101_I;
  assign RIOI3_X105Y103_ILOGIC_X1Y104_O = RIOB33_X105Y103_IOB_X1Y104_I;
  assign RIOI3_X105Y103_ILOGIC_X1Y103_O = RIOB33_X105Y103_IOB_X1Y103_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y106_O = RIOB33_X105Y105_IOB_X1Y106_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y105_O = RIOB33_X105Y105_IOB_X1Y105_I;
  assign RIOI3_X105Y109_ILOGIC_X1Y110_O = RIOB33_X105Y109_IOB_X1Y110_I;
  assign RIOI3_X105Y109_ILOGIC_X1Y109_O = RIOB33_X105Y109_IOB_X1Y109_I;
  assign RIOI3_X105Y111_ILOGIC_X1Y112_O = RIOB33_X105Y111_IOB_X1Y112_I;
  assign RIOI3_X105Y111_ILOGIC_X1Y111_O = RIOB33_X105Y111_IOB_X1Y111_I;
  assign RIOI3_SING_X105Y100_ILOGIC_X1Y100_O = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_O = RIOB33_X105Y107_IOB_X1Y108_I;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_O = RIOB33_X105Y107_IOB_X1Y107_I;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_O = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_A4 = CLBLM_L_X8Y109_SLICE_X10Y109_AO6;
  assign LIOB33_X0Y147_IOB_X0Y147_O = CLBLM_R_X3Y113_SLICE_X3Y113_AO6;
  assign LIOB33_X0Y147_IOB_X0Y148_O = CLBLM_R_X3Y113_SLICE_X3Y113_CO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_A5 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_A6 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_B6 = CLBLL_L_X2Y106_SLICE_X1Y106_CO6;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_A1 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_A2 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_A3 = CLBLM_R_X11Y108_SLICE_X14Y108_CO6;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_A4 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_A5 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_A6 = CLBLM_L_X10Y108_SLICE_X13Y108_DO6;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_B1 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_B2 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_B3 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_B4 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_B5 = CLBLM_R_X11Y108_SLICE_X14Y108_CO6;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_B6 = CLBLM_L_X10Y108_SLICE_X13Y108_DO6;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_C1 = 1'b1;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_C2 = 1'b1;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_C3 = 1'b1;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_C4 = 1'b1;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_C5 = 1'b1;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_C6 = 1'b1;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_D1 = 1'b1;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_D2 = 1'b1;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_D3 = 1'b1;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_D4 = 1'b1;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_D5 = 1'b1;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_D6 = 1'b1;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_A1 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_A2 = CLBLM_R_X11Y107_SLICE_X15Y107_BO6;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_A3 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_A4 = CLBLM_L_X12Y107_SLICE_X16Y107_BO6;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_A5 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_A6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_B1 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_B2 = CLBLM_L_X12Y107_SLICE_X16Y107_BO6;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_B3 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_B4 = CLBLM_R_X11Y107_SLICE_X15Y107_BO6;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_B5 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_C1 = CLBLM_R_X11Y106_SLICE_X15Y106_CO6;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_C2 = CLBLM_R_X13Y108_SLICE_X18Y108_AO6;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_C3 = CLBLM_L_X12Y109_SLICE_X16Y109_AO6;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_C4 = CLBLM_R_X11Y106_SLICE_X14Y106_BO6;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_C5 = CLBLM_L_X12Y108_SLICE_X17Y108_AO6;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_C6 = CLBLM_R_X11Y109_SLICE_X15Y109_AO5;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_D1 = CLBLM_R_X11Y106_SLICE_X15Y106_CO6;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_D2 = CLBLM_R_X13Y108_SLICE_X18Y108_AO6;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_D3 = CLBLM_L_X12Y109_SLICE_X16Y109_AO6;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_D4 = CLBLM_R_X11Y106_SLICE_X14Y106_BO6;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_D5 = CLBLM_L_X12Y108_SLICE_X17Y108_AO6;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_D6 = CLBLM_R_X11Y109_SLICE_X15Y109_AO5;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_A1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_A2 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_A3 = 1'b1;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_A4 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_A5 = 1'b1;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_A6 = 1'b1;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_B1 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_B2 = CLBLM_R_X11Y105_SLICE_X14Y105_AO6;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_B3 = CLBLM_L_X10Y105_SLICE_X12Y105_CO6;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_B4 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_B5 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_B6 = CLBLM_L_X10Y106_SLICE_X12Y106_AO5;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_C1 = CLBLM_L_X10Y105_SLICE_X13Y105_AO6;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_C2 = CLBLM_L_X10Y106_SLICE_X12Y106_AO5;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_C3 = CLBLM_R_X11Y105_SLICE_X14Y105_BO6;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_C4 = CLBLM_L_X10Y105_SLICE_X13Y105_AO5;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_C5 = CLBLM_R_X11Y105_SLICE_X14Y105_CO6;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_C6 = CLBLM_R_X11Y105_SLICE_X14Y105_AO6;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_D1 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_D2 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_D3 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_D4 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_D5 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_D6 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_A1 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_A2 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_A3 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_A4 = CLBLM_R_X11Y105_SLICE_X14Y105_AO6;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_A5 = CLBLM_L_X10Y105_SLICE_X12Y105_CO6;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_A6 = CLBLM_L_X10Y106_SLICE_X12Y106_AO5;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_B1 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_B2 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_B3 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_B4 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_B5 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_B6 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_C1 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_C2 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_C3 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_C4 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_C5 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_C6 = CLBLM_L_X10Y105_SLICE_X12Y105_BO6;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_D1 = 1'b1;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_D2 = 1'b1;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_D3 = 1'b1;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_D4 = 1'b1;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_D5 = 1'b1;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_D6 = 1'b1;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_A1 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_A2 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_A3 = 1'b1;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_A4 = CLBLM_L_X10Y106_SLICE_X13Y106_BO6;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_A5 = CLBLM_R_X11Y105_SLICE_X15Y105_BO6;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_A6 = 1'b1;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_B1 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_B2 = CLBLM_L_X10Y106_SLICE_X12Y106_BO6;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_B3 = CLBLM_R_X11Y105_SLICE_X14Y105_AO6;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_B4 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_B5 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_B6 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_C1 = CLBLM_R_X11Y105_SLICE_X15Y105_BO6;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_C2 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_C3 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_C4 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_C5 = CLBLM_L_X10Y105_SLICE_X13Y105_BO6;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_C6 = CLBLM_L_X10Y106_SLICE_X13Y106_BO6;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_D1 = CLBLM_R_X11Y105_SLICE_X15Y105_BO6;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_D2 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_D3 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_D4 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_D5 = CLBLM_L_X10Y105_SLICE_X13Y105_BO6;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_D6 = CLBLM_L_X10Y106_SLICE_X13Y106_BO6;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_A1 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_A2 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_A3 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_A4 = CLBLM_L_X10Y106_SLICE_X12Y106_BO6;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_A5 = CLBLM_L_X8Y105_SLICE_X11Y105_AO6;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_A6 = 1'b1;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_B1 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_B2 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_B3 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_B4 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_B5 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_B6 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_C1 = 1'b1;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_C2 = 1'b1;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_C3 = 1'b1;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_C4 = 1'b1;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_C5 = 1'b1;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_C6 = 1'b1;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_D1 = 1'b1;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_D2 = 1'b1;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_D3 = 1'b1;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_D4 = 1'b1;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_D5 = 1'b1;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_D6 = 1'b1;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_A1 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_A2 = CLBLM_L_X10Y107_SLICE_X12Y107_BO6;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_A3 = CLBLM_L_X8Y105_SLICE_X10Y105_CO6;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_A4 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_A5 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_A6 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_B2 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_B3 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_B4 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_B5 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_B6 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_C1 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_C2 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_C3 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_C5 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_C6 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_D1 = 1'b1;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_D2 = 1'b1;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_D3 = 1'b1;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_D4 = 1'b1;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_D5 = 1'b1;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_D6 = 1'b1;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_A1 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_A2 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_A3 = CLBLM_L_X8Y105_SLICE_X10Y105_CO6;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_A4 = CLBLM_L_X10Y107_SLICE_X12Y107_BO6;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_A5 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_A6 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_B1 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_B2 = CLBLM_L_X10Y107_SLICE_X13Y107_BO6;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_B3 = CLBLM_L_X10Y107_SLICE_X13Y107_CO6;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_B4 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_B5 = CLBLM_L_X10Y108_SLICE_X12Y108_DO6;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_B6 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_C1 = CLBLM_L_X10Y108_SLICE_X12Y108_AO6;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_C2 = CLBLM_L_X8Y107_SLICE_X11Y107_AO5;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_C3 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_C4 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_C5 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_C6 = CLBLM_L_X10Y107_SLICE_X12Y107_BO6;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_D1 = CLBLM_L_X10Y108_SLICE_X12Y108_DO6;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_D2 = CLBLM_L_X10Y107_SLICE_X13Y107_CO6;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_D3 = CLBLM_L_X10Y107_SLICE_X13Y107_BO6;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_D4 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_D5 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_D6 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_T1 = 1'b1;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_A4 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_A5 = 1'b1;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_A6 = 1'b1;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_A1 = 1'b1;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_A2 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_A3 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_A4 = 1'b1;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_A5 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_A6 = 1'b1;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_C1 = CLBLM_L_X12Y108_SLICE_X16Y108_BO5;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_B1 = CLBLM_L_X10Y108_SLICE_X12Y108_DO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_B2 = CLBLM_L_X10Y107_SLICE_X13Y107_BO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_B3 = CLBLM_R_X11Y107_SLICE_X14Y107_AO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_B4 = CLBLM_L_X10Y107_SLICE_X13Y107_CO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_B5 = CLBLM_L_X10Y108_SLICE_X13Y108_AO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_B6 = CLBLM_L_X10Y108_SLICE_X13Y108_AO5;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_C2 = CLBLM_R_X11Y107_SLICE_X14Y107_CO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_C1 = CLBLM_L_X12Y108_SLICE_X16Y108_AO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_C2 = CLBLM_R_X11Y108_SLICE_X15Y108_AO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_C3 = CLBLM_L_X8Y105_SLICE_X10Y105_CO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_C4 = CLBLM_R_X11Y107_SLICE_X14Y107_BO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_C5 = CLBLM_L_X10Y108_SLICE_X13Y108_DO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_C6 = CLBLM_L_X10Y108_SLICE_X13Y108_BO6;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_C5 = CLBLM_R_X11Y107_SLICE_X15Y107_DO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_D1 = CLBLM_L_X10Y108_SLICE_X13Y108_AO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_D2 = CLBLM_L_X10Y107_SLICE_X13Y107_BO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_D3 = CLBLM_L_X10Y108_SLICE_X12Y108_DO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_D4 = CLBLM_L_X10Y108_SLICE_X13Y108_AO5;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_D5 = CLBLM_R_X11Y107_SLICE_X14Y107_AO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_D6 = CLBLM_L_X10Y107_SLICE_X13Y107_CO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_A1 = 1'b1;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_A2 = CLBLM_L_X10Y107_SLICE_X13Y107_CO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_A3 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_A4 = CLBLM_L_X10Y107_SLICE_X13Y107_BO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_A5 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_A6 = 1'b1;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_B1 = CLBLM_L_X12Y108_SLICE_X16Y108_AO5;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_B2 = CLBLM_L_X8Y107_SLICE_X10Y107_AO5;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_B3 = CLBLM_L_X10Y108_SLICE_X13Y108_CO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_B4 = CLBLM_L_X8Y108_SLICE_X11Y108_CO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_B5 = CLBLM_L_X10Y107_SLICE_X12Y107_AO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_B6 = CLBLM_L_X8Y108_SLICE_X11Y108_AO5;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_C1 = CLBLM_L_X10Y107_SLICE_X12Y107_AO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_C2 = CLBLM_L_X10Y108_SLICE_X13Y108_CO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_C3 = CLBLM_L_X12Y108_SLICE_X16Y108_AO5;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_C4 = CLBLM_L_X8Y108_SLICE_X11Y108_AO5;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_C5 = CLBLM_L_X8Y107_SLICE_X10Y107_AO5;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_C6 = CLBLM_L_X8Y108_SLICE_X11Y108_CO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_A1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_D1 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_D2 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_D3 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_D4 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_D5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_D6 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_B2 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_B3 = CLBLM_R_X7Y109_SLICE_X9Y109_AO5;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_B6 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_C3 = CLBLM_L_X8Y110_SLICE_X10Y110_CO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_C4 = CLBLM_L_X8Y110_SLICE_X10Y110_BO6;
  assign LIOI3_X0Y101_ILOGIC_X0Y102_D = LIOB33_X0Y101_IOB_X0Y102_I;
  assign LIOI3_X0Y101_ILOGIC_X0Y101_D = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_A1 = CLBLM_L_X10Y109_SLICE_X12Y109_CO6;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_A2 = CLBLM_R_X11Y110_SLICE_X15Y110_AO6;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_A3 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_A4 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_A5 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_A6 = CLBLM_L_X10Y109_SLICE_X13Y109_CO6;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_B1 = CLBLM_L_X10Y109_SLICE_X12Y109_CO6;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_B2 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_B3 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_B4 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_B5 = CLBLM_R_X11Y109_SLICE_X15Y109_BO6;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_B6 = CLBLM_L_X10Y109_SLICE_X13Y109_CO6;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_C1 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_C2 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_C3 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_C4 = CLBLM_R_X11Y108_SLICE_X14Y108_DO6;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_C5 = CLBLM_L_X10Y107_SLICE_X13Y107_AO6;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_C6 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_D1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_D2 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_D3 = CLBLM_R_X11Y110_SLICE_X15Y110_AO6;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_D4 = CLBLM_L_X10Y109_SLICE_X13Y109_CO6;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_D5 = CLBLM_L_X10Y109_SLICE_X12Y109_CO6;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_D6 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_A1 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_A2 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_A3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_A4 = CLBLM_R_X11Y109_SLICE_X14Y109_AO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_A5 = CLBLM_L_X10Y106_SLICE_X13Y106_AO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_A6 = CLBLM_L_X10Y106_SLICE_X13Y106_DO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_B1 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_B2 = CLBLM_R_X11Y109_SLICE_X14Y109_AO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_B3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_B4 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_B5 = CLBLM_L_X10Y106_SLICE_X13Y106_AO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_B6 = CLBLM_L_X10Y106_SLICE_X13Y106_DO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_C1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_C2 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_C3 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_C4 = CLBLM_L_X10Y107_SLICE_X12Y107_CO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_C5 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_C6 = CLBLM_L_X8Y108_SLICE_X11Y108_CO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_D1 = CLBLM_L_X10Y107_SLICE_X12Y107_AO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_D2 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_D3 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_D4 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_D5 = CLBLM_L_X10Y108_SLICE_X13Y108_CO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_D6 = CLBLM_L_X8Y108_SLICE_X11Y108_CO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_A1 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_A2 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_A3 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_A4 = 1'b1;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_A5 = 1'b1;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_A6 = 1'b1;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_B1 = CLBLM_R_X5Y106_SLICE_X6Y106_CO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_B2 = CLBLL_L_X4Y105_SLICE_X4Y105_AO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_B3 = CLBLM_R_X7Y106_SLICE_X8Y106_CO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_B4 = CLBLM_R_X7Y106_SLICE_X8Y106_AO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_B5 = CLBLM_R_X5Y104_SLICE_X6Y104_AO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_B6 = CLBLL_L_X4Y105_SLICE_X4Y105_AO5;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_C1 = CLBLM_R_X5Y104_SLICE_X6Y104_AO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_C2 = CLBLM_R_X7Y106_SLICE_X8Y106_CO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_C3 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_C4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_C5 = CLBLM_R_X5Y106_SLICE_X6Y106_CO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_C6 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_D1 = CLBLL_L_X4Y105_SLICE_X4Y105_AO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_D2 = CLBLM_R_X5Y104_SLICE_X6Y104_AO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_D3 = CLBLM_R_X7Y106_SLICE_X8Y106_CO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_D4 = CLBLL_L_X4Y105_SLICE_X4Y105_AO5;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_D5 = CLBLM_R_X5Y106_SLICE_X6Y106_CO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_D6 = CLBLM_R_X7Y106_SLICE_X8Y106_AO6;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_D1 = CLBLL_L_X4Y116_SLICE_X5Y116_AO5;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_A1 = CLBLM_R_X7Y105_SLICE_X8Y105_BO6;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_A2 = CLBLL_L_X4Y105_SLICE_X4Y105_BO6;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_A3 = CLBLM_R_X3Y104_SLICE_X3Y104_CO6;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_A4 = CLBLL_L_X4Y105_SLICE_X4Y105_DO6;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_A5 = CLBLM_R_X7Y105_SLICE_X8Y105_AO6;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_A6 = CLBLM_R_X3Y105_SLICE_X3Y105_BO5;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_B1 = 1'b1;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_B2 = 1'b1;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_B3 = 1'b1;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_B4 = 1'b1;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_B5 = 1'b1;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_B6 = 1'b1;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_C1 = 1'b1;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_C2 = 1'b1;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_C3 = 1'b1;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_C4 = 1'b1;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_C5 = 1'b1;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_C6 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_D6 = 1'b1;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_D1 = 1'b1;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_D2 = 1'b1;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_D3 = 1'b1;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_D4 = 1'b1;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_D5 = 1'b1;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_D6 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_T1 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_A5 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_A6 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_D1 = CLBLL_L_X4Y116_SLICE_X5Y116_AO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_A1 = CLBLM_L_X10Y110_SLICE_X12Y110_AO5;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_A2 = CLBLM_L_X12Y109_SLICE_X16Y109_AO5;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_A3 = CLBLM_R_X11Y109_SLICE_X14Y109_DO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_A4 = CLBLM_R_X11Y109_SLICE_X14Y109_BO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_A5 = CLBLM_L_X10Y106_SLICE_X13Y106_DO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_A6 = CLBLM_R_X13Y108_SLICE_X18Y108_CO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_B1 = CLBLM_L_X8Y110_SLICE_X11Y110_CO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_B2 = CLBLM_L_X10Y111_SLICE_X13Y111_AO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_B3 = CLBLM_L_X10Y109_SLICE_X13Y109_AO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_B4 = CLBLM_R_X11Y110_SLICE_X14Y110_CO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_B5 = CLBLM_L_X8Y109_SLICE_X11Y109_AO5;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_B6 = CLBLM_L_X10Y111_SLICE_X13Y111_AO5;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_C1 = 1'b1;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_C1 = CLBLM_L_X10Y109_SLICE_X13Y109_AO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_C2 = CLBLM_R_X11Y110_SLICE_X14Y110_CO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_C3 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_C4 = CLBLM_L_X8Y110_SLICE_X11Y110_CO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_C5 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_C6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_C2 = 1'b1;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_D1 = CLBLM_L_X8Y109_SLICE_X11Y109_AO5;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_D2 = CLBLM_L_X10Y111_SLICE_X13Y111_AO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_D3 = CLBLM_L_X8Y110_SLICE_X11Y110_CO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_D4 = CLBLM_L_X10Y111_SLICE_X13Y111_AO5;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_D5 = CLBLM_L_X10Y109_SLICE_X13Y109_AO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_D6 = CLBLM_R_X11Y110_SLICE_X14Y110_CO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_A1 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_A2 = 1'b1;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_A3 = 1'b1;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_A4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_A5 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_A6 = 1'b1;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_B2 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_B3 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_B4 = 1'b1;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_B5 = 1'b1;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_B6 = 1'b1;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_C1 = CLBLM_L_X8Y106_SLICE_X11Y106_AO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_C2 = CLBLM_L_X10Y106_SLICE_X13Y106_DO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_C3 = CLBLM_L_X10Y110_SLICE_X12Y110_AO5;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_C4 = CLBLM_L_X8Y110_SLICE_X10Y110_AO5;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_C5 = CLBLM_L_X10Y106_SLICE_X13Y106_CO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_C6 = CLBLM_R_X11Y109_SLICE_X14Y109_BO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_A1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_A2 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_A3 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_A4 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_A5 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_A6 = 1'b1;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_D1 = CLBLM_L_X10Y110_SLICE_X12Y110_AO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_D2 = CLBLM_R_X11Y110_SLICE_X14Y110_AO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_D3 = CLBLM_L_X10Y108_SLICE_X12Y108_BO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_B1 = CLBLM_R_X3Y105_SLICE_X3Y105_DO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_B2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_B3 = CLBLM_R_X3Y106_SLICE_X2Y106_BO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_B4 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_B5 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_B6 = CLBLM_R_X3Y106_SLICE_X3Y106_AO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_C1 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_C2 = CLBLL_L_X4Y105_SLICE_X4Y105_CO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_C3 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_C4 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_C5 = CLBLM_R_X5Y106_SLICE_X6Y106_AO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_C6 = CLBLM_R_X3Y105_SLICE_X3Y105_AO5;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_D1 = CLBLM_R_X3Y106_SLICE_X2Y106_BO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_D2 = CLBLM_R_X3Y105_SLICE_X3Y105_DO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_D3 = CLBLM_R_X3Y106_SLICE_X2Y106_AO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_D4 = CLBLM_R_X5Y106_SLICE_X6Y106_BO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_D5 = CLBLL_L_X4Y106_SLICE_X4Y106_AO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_D6 = CLBLM_R_X3Y106_SLICE_X3Y106_AO6;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_A1 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_A2 = CLBLM_R_X3Y104_SLICE_X3Y104_CO6;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_A3 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_A4 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_A5 = CLBLL_L_X4Y105_SLICE_X4Y105_CO6;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_A6 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_B1 = CLBLM_R_X3Y106_SLICE_X3Y106_BO6;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_B2 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_B3 = CLBLL_L_X4Y105_SLICE_X5Y105_AO6;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_B4 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_B5 = CLBLL_L_X4Y106_SLICE_X5Y106_AO6;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_B6 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_C1 = CLBLM_R_X3Y104_SLICE_X3Y104_CO6;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_C2 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_C3 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_C4 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_C5 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_C6 = CLBLL_L_X4Y105_SLICE_X4Y105_CO6;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_D1 = CLBLL_L_X4Y106_SLICE_X5Y106_AO6;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_D2 = CLBLL_L_X4Y106_SLICE_X4Y106_AO5;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_D3 = CLBLM_R_X5Y106_SLICE_X6Y106_BO5;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_D4 = CLBLM_R_X3Y106_SLICE_X3Y106_BO6;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_D5 = CLBLM_R_X5Y106_SLICE_X6Y106_BO6;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_D6 = CLBLL_L_X4Y105_SLICE_X5Y105_AO6;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_A1 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_A2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_A3 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_A4 = 1'b1;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_A5 = 1'b1;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_A6 = 1'b1;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_B1 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_B2 = CLBLM_L_X10Y111_SLICE_X12Y111_BO6;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_B4 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_B5 = CLBLM_R_X11Y111_SLICE_X14Y111_BO6;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_B6 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_C1 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_C2 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_C3 = CLBLM_R_X11Y109_SLICE_X14Y109_CO6;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_C5 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_C6 = CLBLM_R_X13Y108_SLICE_X18Y108_CO6;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_D1 = CLBLM_R_X11Y111_SLICE_X15Y111_AO6;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_D2 = CLBLM_L_X10Y110_SLICE_X13Y110_AO6;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_D3 = CLBLM_R_X11Y111_SLICE_X14Y111_CO6;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_D4 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_D5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_D6 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_A1 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_A2 = 1'b1;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_A3 = CLBLM_L_X10Y109_SLICE_X12Y109_AO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_A4 = CLBLM_L_X10Y111_SLICE_X13Y111_CO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_A6 = 1'b1;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_B1 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_B2 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_B3 = CLBLM_L_X10Y109_SLICE_X12Y109_AO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_B4 = CLBLM_L_X10Y111_SLICE_X13Y111_CO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_B6 = CLBLM_L_X10Y110_SLICE_X12Y110_CO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_C1 = CLBLM_L_X10Y109_SLICE_X12Y109_AO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_C2 = CLBLM_L_X10Y111_SLICE_X13Y111_CO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_C3 = CLBLM_L_X10Y110_SLICE_X12Y110_CO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_C4 = CLBLM_L_X8Y111_SLICE_X10Y111_AO5;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_C5 = CLBLM_L_X10Y110_SLICE_X12Y110_BO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_C6 = CLBLM_L_X10Y110_SLICE_X12Y110_BO5;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_A1 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_A2 = CLBLL_L_X4Y106_SLICE_X4Y106_CO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_A3 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_A4 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_A5 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_A6 = CLBLM_R_X3Y106_SLICE_X3Y106_BO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_D1 = CLBLM_L_X10Y111_SLICE_X12Y111_AO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_D2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_B1 = CLBLL_L_X4Y106_SLICE_X4Y106_DO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_B2 = CLBLL_L_X4Y106_SLICE_X5Y106_BO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_B3 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_B4 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_B5 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_B6 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_D6 = CLBLM_L_X10Y111_SLICE_X12Y111_BO6;
  assign LIOI3_X0Y103_ILOGIC_X0Y103_D = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_C1 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_C2 = CLBLM_R_X3Y106_SLICE_X3Y106_BO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_C3 = CLBLL_L_X4Y106_SLICE_X4Y106_CO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_C4 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_C5 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_C6 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_D1 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_D2 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_D3 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_D4 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_D5 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_D6 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_A5 = 1'b1;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_A1 = 1'b1;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_A2 = CLBLM_L_X12Y105_SLICE_X16Y105_CO6;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_A3 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_A4 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_A5 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_A1 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_A2 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_A3 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_A4 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_A5 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_A6 = 1'b1;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_A6 = 1'b1;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_B4 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_B1 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_B2 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_B3 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_B4 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_B5 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_B6 = 1'b1;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_B6 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_C3 = CLBLM_R_X11Y105_SLICE_X14Y105_BO6;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_C4 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_C1 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_C2 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_C3 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_C4 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_C5 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_C6 = 1'b1;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_C5 = CLBLM_L_X12Y105_SLICE_X16Y105_AO5;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_C6 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_D1 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_D2 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_D3 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_D4 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_D1 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_D2 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_D3 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_D4 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_D5 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_D6 = 1'b1;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_A1 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_A2 = CLBLM_R_X11Y105_SLICE_X15Y105_DO6;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_A3 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_A4 = CLBLM_L_X12Y105_SLICE_X16Y105_CO6;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_A5 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_A6 = CLBLM_L_X10Y105_SLICE_X13Y105_DO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_C2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_B1 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_B2 = CLBLM_R_X11Y105_SLICE_X15Y105_DO6;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_B3 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_B4 = CLBLM_L_X12Y105_SLICE_X16Y105_CO6;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_B5 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_C3 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_C4 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_B6 = CLBLM_L_X10Y105_SLICE_X13Y105_DO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_C5 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_C2 = CLBLM_R_X11Y105_SLICE_X15Y105_AO5;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_C1 = CLBLM_R_X7Y109_SLICE_X9Y109_AO6;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_C4 = CLBLM_R_X11Y106_SLICE_X14Y106_AO6;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_C5 = CLBLM_R_X11Y107_SLICE_X14Y107_DO6;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_C6 = CLBLM_L_X12Y105_SLICE_X16Y105_CO6;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_C3 = CLBLM_L_X12Y105_SLICE_X16Y105_DO6;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_D1 = CLBLM_R_X7Y109_SLICE_X9Y109_AO6;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_D2 = CLBLM_R_X11Y105_SLICE_X15Y105_AO5;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_D3 = CLBLM_R_X11Y107_SLICE_X14Y107_DO6;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_D4 = CLBLM_R_X11Y106_SLICE_X14Y106_AO6;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_D5 = CLBLM_L_X12Y105_SLICE_X16Y105_DO6;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_D6 = CLBLM_L_X12Y105_SLICE_X16Y105_CO6;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_A1 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_A2 = 1'b1;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_A3 = 1'b1;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_A4 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_A5 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_A6 = 1'b1;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_B1 = CLBLM_R_X11Y113_SLICE_X14Y113_CO6;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_B2 = CLBLM_R_X11Y111_SLICE_X15Y111_CO6;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_B3 = CLBLM_R_X11Y111_SLICE_X14Y111_DO6;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_B4 = CLBLM_L_X10Y112_SLICE_X13Y112_DO6;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_B5 = CLBLM_R_X11Y112_SLICE_X15Y112_BO6;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_B6 = CLBLM_L_X10Y112_SLICE_X13Y112_AO5;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_C1 = CLBLM_L_X10Y112_SLICE_X13Y112_AO6;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_C2 = CLBLM_R_X11Y112_SLICE_X15Y112_BO6;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_C3 = CLBLM_R_X11Y113_SLICE_X14Y113_CO6;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_C4 = CLBLM_L_X10Y112_SLICE_X13Y112_AO5;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_C5 = CLBLM_R_X11Y113_SLICE_X14Y113_AO6;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_C6 = CLBLM_R_X11Y112_SLICE_X14Y112_CO6;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_D1 = 1'b1;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_D2 = 1'b1;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_D3 = 1'b1;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_D4 = 1'b1;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_D5 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_D6 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_A1 = CLBLM_L_X10Y111_SLICE_X12Y111_DO6;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_A2 = CLBLM_L_X10Y112_SLICE_X12Y112_DO6;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_A3 = 1'b1;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_A4 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_A5 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_A6 = 1'b1;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_B1 = CLBLM_L_X10Y110_SLICE_X13Y110_DO6;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_B2 = CLBLM_R_X11Y112_SLICE_X14Y112_AO6;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_B3 = CLBLM_L_X10Y112_SLICE_X13Y112_AO6;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_B4 = CLBLM_R_X11Y113_SLICE_X14Y113_AO6;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_B5 = CLBLM_L_X8Y112_SLICE_X10Y112_AO6;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_B6 = CLBLM_R_X11Y112_SLICE_X14Y112_CO6;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_C1 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_C2 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_C3 = CLBLM_R_X11Y112_SLICE_X14Y112_DO6;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_C4 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_C5 = CLBLM_R_X11Y112_SLICE_X15Y112_DO6;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_C6 = CLBLM_L_X10Y111_SLICE_X13Y111_DO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_A1 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_A2 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_A3 = CLBLL_L_X4Y108_SLICE_X5Y108_AO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_A4 = CLBLL_L_X4Y107_SLICE_X4Y107_BO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_A5 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_A6 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_D1 = CLBLM_R_X11Y111_SLICE_X14Y111_DO6;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_D2 = CLBLM_R_X11Y112_SLICE_X14Y112_DO6;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_D3 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_D4 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_D5 = CLBLM_R_X11Y112_SLICE_X15Y112_DO6;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_D6 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_B1 = CLBLM_R_X5Y107_SLICE_X7Y107_AO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_B2 = CLBLL_L_X4Y108_SLICE_X5Y108_BO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_B3 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_B4 = CLBLL_L_X4Y107_SLICE_X4Y107_BO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_B5 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_B6 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_C1 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_C2 = CLBLL_L_X4Y108_SLICE_X5Y108_AO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_C3 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_C4 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_C5 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_C6 = CLBLL_L_X4Y107_SLICE_X4Y107_BO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_D1 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_D2 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_D3 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_D4 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_D5 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_D6 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_A1 = CLBLM_R_X5Y107_SLICE_X6Y107_AO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_A2 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_A3 = CLBLM_R_X5Y106_SLICE_X7Y106_BO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_A4 = CLBLL_L_X4Y107_SLICE_X4Y107_CO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_A5 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_A6 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_A1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_A2 = 1'b1;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_A3 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_B1 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_B2 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_B3 = CLBLM_R_X5Y106_SLICE_X7Y106_BO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_B4 = CLBLL_L_X4Y106_SLICE_X5Y106_DO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_B5 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_B6 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_B1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_B2 = CLBLM_L_X12Y105_SLICE_X16Y105_BO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_C1 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_C2 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_C3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_C4 = CLBLM_R_X5Y108_SLICE_X6Y108_DO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_C5 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_C6 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_C1 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_C2 = CLBLM_R_X11Y106_SLICE_X14Y106_CO6;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_C3 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_C4 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_C5 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_C6 = CLBLM_L_X12Y105_SLICE_X16Y105_BO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_D1 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_D2 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_D3 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_D4 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_D5 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_D6 = 1'b1;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_D4 = CLBLM_R_X11Y105_SLICE_X14Y105_DO6;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_D5 = CLBLM_L_X12Y108_SLICE_X17Y108_AO5;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_D6 = CLBLM_R_X11Y107_SLICE_X15Y107_BO6;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_D3 = CLBLM_R_X11Y106_SLICE_X14Y106_DO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_A1 = 1'b1;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_A2 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_A3 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_A4 = 1'b1;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_A5 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_A6 = 1'b1;
  assign RIOI3_X105Y103_ILOGIC_X1Y104_D = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_B1 = CLBLM_R_X11Y105_SLICE_X14Y105_DO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_B2 = CLBLM_R_X11Y105_SLICE_X14Y105_CO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_B3 = CLBLM_R_X11Y106_SLICE_X15Y106_AO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_B4 = CLBLM_L_X10Y105_SLICE_X13Y105_AO5;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_B5 = CLBLM_R_X11Y105_SLICE_X14Y105_BO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_B6 = CLBLM_R_X11Y106_SLICE_X14Y106_CO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_C1 = CLBLM_R_X7Y109_SLICE_X9Y109_AO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_C2 = CLBLM_R_X11Y106_SLICE_X15Y106_AO5;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_C3 = CLBLM_R_X11Y107_SLICE_X14Y107_DO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_C4 = CLBLM_R_X11Y106_SLICE_X14Y106_AO5;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_C5 = CLBLM_L_X12Y107_SLICE_X17Y107_AO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_C6 = CLBLM_L_X12Y106_SLICE_X16Y106_BO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_D1 = CLBLM_R_X7Y109_SLICE_X9Y109_AO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_D2 = CLBLM_R_X11Y106_SLICE_X15Y106_AO5;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_D3 = CLBLM_R_X11Y107_SLICE_X14Y107_DO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_D4 = CLBLM_R_X11Y106_SLICE_X14Y106_AO5;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_D5 = CLBLM_L_X12Y107_SLICE_X17Y107_AO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_D6 = CLBLM_L_X12Y106_SLICE_X16Y106_BO6;
  assign RIOI3_X105Y103_ILOGIC_X1Y103_D = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_B5 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_B6 = CLBLM_L_X10Y107_SLICE_X13Y107_AO6;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_A1 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_A2 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_A3 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_A4 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_A5 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_A6 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_B1 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_B2 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_B3 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_B4 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_B5 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_B6 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_C1 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_C2 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_C3 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_C4 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_C5 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_C6 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_D1 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_D2 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_D3 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_D4 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_D5 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_D6 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_A1 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_A2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_A3 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_A4 = CLBLM_L_X10Y109_SLICE_X13Y109_BO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_A5 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_A6 = CLBLM_L_X8Y110_SLICE_X11Y110_CO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_B1 = CLBLM_L_X10Y113_SLICE_X12Y113_DO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_B2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_B3 = CLBLM_R_X11Y112_SLICE_X14Y112_BO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_B4 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_B5 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_B6 = CLBLM_L_X10Y113_SLICE_X12Y113_CO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_C1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_C2 = CLBLM_L_X10Y109_SLICE_X13Y109_DO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_C3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_C4 = CLBLM_L_X12Y111_SLICE_X16Y111_BO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_C5 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_C6 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A1 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A3 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A4 = CLBLM_R_X3Y108_SLICE_X3Y108_BO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A5 = CLBLL_L_X4Y108_SLICE_X4Y108_AO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A6 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B3 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B4 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B5 = CLBLL_L_X4Y108_SLICE_X4Y108_AO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B6 = CLBLL_L_X4Y109_SLICE_X4Y109_CO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B1 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B2 = CLBLM_R_X3Y108_SLICE_X3Y108_BO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_D1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_D2 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_D3 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_D4 = CLBLM_L_X8Y110_SLICE_X11Y110_CO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_D5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_D6 = CLBLM_L_X10Y109_SLICE_X13Y109_BO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C2 = CLBLL_L_X4Y107_SLICE_X4Y107_BO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C3 = CLBLM_R_X5Y107_SLICE_X7Y107_AO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C1 = CLBLL_L_X4Y108_SLICE_X5Y108_BO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C5 = CLBLL_L_X4Y110_SLICE_X4Y110_AO5;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C4 = CLBLL_L_X4Y109_SLICE_X4Y109_AO5;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C6 = CLBLL_L_X4Y110_SLICE_X4Y110_AO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D1 = CLBLL_L_X4Y108_SLICE_X5Y108_BO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D2 = CLBLL_L_X4Y110_SLICE_X4Y110_AO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D3 = CLBLM_R_X5Y107_SLICE_X7Y107_AO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D4 = CLBLL_L_X4Y109_SLICE_X4Y109_AO5;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D5 = CLBLL_L_X4Y110_SLICE_X4Y110_AO5;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D6 = CLBLL_L_X4Y107_SLICE_X4Y107_BO6;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_C3 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A1 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A2 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A3 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A4 = CLBLL_L_X4Y108_SLICE_X4Y108_CO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A5 = CLBLM_R_X5Y108_SLICE_X6Y108_BO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A6 = CLBLM_R_X5Y109_SLICE_X6Y109_BO6;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_A1 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_A2 = 1'b1;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_A3 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B1 = CLBLM_R_X5Y109_SLICE_X6Y109_CO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B2 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B3 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B4 = CLBLL_L_X4Y108_SLICE_X4Y108_CO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B5 = CLBLM_R_X5Y108_SLICE_X6Y108_BO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B6 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_A5 = 1'b1;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_A6 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C1 = CLBLM_R_X5Y108_SLICE_X6Y108_BO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C3 = CLBLM_R_X5Y109_SLICE_X6Y109_CO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C4 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C5 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C6 = CLBLL_L_X4Y108_SLICE_X4Y108_CO6;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_B3 = CLBLM_R_X11Y106_SLICE_X15Y106_AO5;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_B4 = CLBLM_L_X12Y107_SLICE_X16Y107_CO6;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_B5 = CLBLM_L_X12Y107_SLICE_X17Y107_BO6;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_B6 = CLBLM_R_X11Y107_SLICE_X15Y107_AO5;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_C1 = CLBLM_L_X12Y107_SLICE_X17Y107_BO6;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_C2 = CLBLM_L_X12Y107_SLICE_X16Y107_CO6;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D1 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D2 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D3 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D4 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D5 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D6 = 1'b1;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_D1 = CLBLM_L_X12Y107_SLICE_X17Y107_AO6;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_D2 = CLBLM_R_X11Y106_SLICE_X15Y106_AO5;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_D3 = CLBLM_L_X12Y107_SLICE_X17Y107_BO6;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_D4 = CLBLM_R_X11Y107_SLICE_X15Y107_AO5;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_D5 = CLBLM_R_X11Y107_SLICE_X15Y107_AO6;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_D6 = CLBLM_L_X12Y107_SLICE_X16Y107_CO6;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_A1 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_A2 = 1'b1;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_A3 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_A4 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_A5 = 1'b1;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_A6 = 1'b1;
  assign LIOI3_X0Y105_ILOGIC_X0Y106_D = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_B1 = CLBLM_R_X11Y108_SLICE_X14Y108_BO6;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_B2 = CLBLM_L_X12Y107_SLICE_X17Y107_BO6;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_B3 = CLBLM_R_X11Y107_SLICE_X15Y107_AO6;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_B4 = CLBLM_L_X10Y108_SLICE_X12Y108_DO6;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_B5 = CLBLM_R_X11Y107_SLICE_X14Y107_AO6;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_B6 = CLBLM_R_X11Y107_SLICE_X14Y107_AO5;
  assign LIOI3_X0Y105_ILOGIC_X0Y105_D = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_D3 = CLBLM_L_X10Y112_SLICE_X13Y112_CO6;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_C1 = CLBLM_R_X11Y107_SLICE_X14Y107_AO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_C6 = 1'b1;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_C2 = CLBLM_R_X11Y107_SLICE_X15Y107_AO6;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_C3 = CLBLM_R_X11Y108_SLICE_X14Y108_BO6;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_C4 = CLBLM_R_X11Y107_SLICE_X14Y107_AO5;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_C5 = CLBLM_L_X12Y107_SLICE_X17Y107_BO6;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_C6 = CLBLM_L_X10Y108_SLICE_X12Y108_DO6;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_D1 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_D2 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_D3 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_D4 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_D5 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_D6 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y114_D = LIOB33_X0Y113_IOB_X0Y114_I;
  assign LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y113_D = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_A1 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_A2 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_A3 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_A4 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_A5 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_A6 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_B1 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_B2 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_B3 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_B4 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_B5 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_B6 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_A1 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_A2 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_A3 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_C4 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_C5 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_C6 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_A4 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_A5 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_A6 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_C1 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_C2 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_B1 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_B2 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_B3 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_B4 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_B5 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_B6 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_D5 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_D6 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_D1 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_D2 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_C1 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_C2 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_C3 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_C4 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_C5 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_C6 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_A1 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_A2 = CLBLM_R_X11Y114_SLICE_X14Y114_AO6;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_A3 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_A4 = CLBLM_L_X10Y114_SLICE_X12Y114_BO6;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_A5 = CLBLM_R_X11Y113_SLICE_X14Y113_AO6;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_A6 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_D1 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_D2 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_D3 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_D4 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_B4 = CLBLM_L_X10Y109_SLICE_X13Y109_DO6;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_B5 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_B6 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_D5 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_A1 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_A2 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_A1 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_A2 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_A3 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_A4 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_A3 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_A4 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_A6 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_B1 = CLBLM_R_X7Y110_SLICE_X9Y110_BO5;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_B2 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_C1 = CLBLM_R_X11Y113_SLICE_X14Y113_AO6;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_B1 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_B2 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_B3 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_B4 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_B5 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_B6 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_B4 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_C1 = CLBLL_L_X4Y109_SLICE_X5Y109_AO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_B3 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_B5 = CLBLM_R_X5Y109_SLICE_X7Y109_DO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_B6 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_C6 = CLBLL_L_X4Y109_SLICE_X4Y109_BO6;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_C3 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_C4 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_C5 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_C6 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_D2 = CLBLM_R_X11Y114_SLICE_X14Y114_AO6;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_D3 = CLBLM_R_X11Y113_SLICE_X14Y113_BO6;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_D4 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_D6 = CLBLM_L_X10Y114_SLICE_X12Y114_BO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_D1 = CLBLM_R_X5Y110_SLICE_X6Y110_BO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_D2 = CLBLM_R_X3Y111_SLICE_X2Y111_AO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_D3 = CLBLL_L_X4Y109_SLICE_X4Y109_BO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_D4 = CLBLL_L_X4Y109_SLICE_X5Y109_CO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_D5 = CLBLL_L_X4Y111_SLICE_X4Y111_AO5;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_D6 = CLBLL_L_X4Y110_SLICE_X4Y110_BO6;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_D1 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_D2 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_D3 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_D4 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_D5 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_D6 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_A1 = CLBLM_R_X3Y110_SLICE_X3Y110_DO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_A2 = CLBLM_R_X5Y109_SLICE_X7Y109_AO5;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_A3 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_A4 = CLBLM_R_X5Y108_SLICE_X7Y108_AO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_A5 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_A6 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_B1 = CLBLM_R_X3Y110_SLICE_X3Y110_DO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_B2 = CLBLM_R_X5Y109_SLICE_X7Y109_AO5;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_B3 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_B4 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_B5 = CLBLM_R_X5Y108_SLICE_X7Y108_AO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_B6 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_A1 = 1'b1;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_A2 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_A3 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_C1 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_C2 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_C3 = CLBLM_R_X5Y108_SLICE_X6Y108_DO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_C4 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_C5 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_C6 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_B1 = CLBLM_R_X11Y107_SLICE_X15Y107_DO6;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_B2 = CLBLM_R_X11Y107_SLICE_X14Y107_BO6;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_B3 = CLBLM_L_X10Y108_SLICE_X13Y108_DO6;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_B4 = CLBLM_L_X12Y108_SLICE_X16Y108_BO5;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_B5 = CLBLM_R_X11Y108_SLICE_X15Y108_AO6;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_B6 = CLBLM_R_X11Y107_SLICE_X14Y107_CO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_D1 = CLBLM_R_X5Y109_SLICE_X7Y109_CO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_D2 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_D3 = CLBLM_R_X5Y110_SLICE_X6Y110_AO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_D4 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_D5 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_D6 = CLBLL_L_X4Y110_SLICE_X5Y110_BO6;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_C3 = CLBLM_R_X11Y106_SLICE_X14Y106_DO6;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_C4 = CLBLM_L_X12Y108_SLICE_X17Y108_AO5;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_C6 = CLBLM_R_X11Y107_SLICE_X15Y107_BO6;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_D1 = CLBLM_R_X11Y107_SLICE_X15Y107_CO6;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_D2 = CLBLM_R_X11Y108_SLICE_X14Y108_AO5;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_D3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_D4 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_D5 = CLBLM_L_X12Y107_SLICE_X16Y107_AO6;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_D6 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_A1 = CLBLM_L_X10Y108_SLICE_X12Y108_DO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_A2 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_A3 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_A4 = CLBLM_R_X11Y108_SLICE_X14Y108_BO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_A5 = 1'b1;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_A6 = 1'b1;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_B1 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_B2 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_B3 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_B4 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_B6 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_C1 = CLBLM_L_X12Y107_SLICE_X17Y107_BO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_C2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_C3 = CLBLM_L_X10Y108_SLICE_X12Y108_DO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_C4 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_C5 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_C6 = CLBLM_R_X11Y108_SLICE_X14Y108_BO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_D1 = CLBLM_R_X11Y108_SLICE_X14Y108_AO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_D2 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_D3 = CLBLM_L_X10Y108_SLICE_X12Y108_AO5;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_D4 = CLBLM_R_X11Y108_SLICE_X14Y108_CO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_D5 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_D6 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_A1 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_A2 = CLBLM_L_X10Y105_SLICE_X12Y105_BO6;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_A3 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_A4 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_A5 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_A6 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_B1 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_B2 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_B3 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_B4 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_B5 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_B6 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_C1 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_C2 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_C3 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_C4 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_C5 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_C6 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_D1 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_D2 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_D3 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_D4 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_D5 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_D6 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_A1 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_A2 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_A3 = CLBLL_L_X4Y111_SLICE_X5Y111_AO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_A4 = CLBLL_L_X4Y110_SLICE_X4Y110_CO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_A5 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_A6 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_A1 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_A3 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_A4 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_A5 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_B3 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_B4 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_B5 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_B6 = CLBLM_R_X5Y109_SLICE_X7Y109_DO6;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_A6 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_A2 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_B1 = CLBLM_R_X3Y111_SLICE_X3Y111_AO5;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_C2 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_C3 = CLBLM_R_X7Y110_SLICE_X9Y110_BO5;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_B1 = CLBLM_L_X10Y107_SLICE_X13Y107_BO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_C5 = CLBLM_R_X3Y111_SLICE_X3Y111_AO5;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_B2 = CLBLM_L_X8Y105_SLICE_X10Y105_AO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_C1 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_B3 = CLBLM_L_X8Y104_SLICE_X10Y104_AO6;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_B4 = CLBLM_L_X8Y107_SLICE_X10Y107_BO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_C4 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_B5 = CLBLM_L_X10Y108_SLICE_X13Y108_AO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_C6 = CLBLM_R_X5Y109_SLICE_X7Y109_DO6;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_B6 = CLBLM_L_X8Y105_SLICE_X10Y105_AO5;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_D1 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_D2 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_D3 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_C1 = CLBLM_L_X10Y108_SLICE_X13Y108_AO6;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_C2 = CLBLM_L_X8Y104_SLICE_X10Y104_AO6;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_C3 = CLBLM_L_X8Y105_SLICE_X10Y105_AO5;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_C4 = CLBLM_L_X8Y105_SLICE_X10Y105_AO6;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_C5 = CLBLM_L_X10Y107_SLICE_X13Y107_BO6;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_C6 = CLBLM_L_X8Y107_SLICE_X10Y107_BO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_D4 = CLBLL_L_X4Y110_SLICE_X5Y110_CO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_D5 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_D6 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_D1 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_D2 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_D3 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_D4 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_D5 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_D6 = CLBLM_L_X10Y105_SLICE_X12Y105_BO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_A1 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_A2 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_A3 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_A4 = CLBLL_L_X4Y109_SLICE_X5Y109_BO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_A5 = CLBLM_R_X5Y109_SLICE_X7Y109_BO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_A6 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_B1 = CLBLM_R_X7Y110_SLICE_X9Y110_DO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_B2 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_B3 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_B4 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_B5 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_B6 = CLBLM_R_X5Y110_SLICE_X7Y110_DO6;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_A1 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_A2 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_A3 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_C1 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_C2 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_C3 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_C4 = CLBLM_R_X7Y110_SLICE_X9Y110_DO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_C5 = CLBLM_R_X5Y110_SLICE_X7Y110_DO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_C6 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_A4 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_A5 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_A6 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_B1 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_B2 = CLBLM_R_X13Y108_SLICE_X19Y108_AO6;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_B3 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_B4 = CLBLM_R_X11Y108_SLICE_X15Y108_BO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_D1 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_D2 = CLBLM_R_X5Y109_SLICE_X7Y109_CO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_D3 = CLBLM_R_X5Y110_SLICE_X6Y110_AO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_D4 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_D5 = CLBLL_L_X4Y110_SLICE_X5Y110_BO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_D6 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_C1 = CLBLM_R_X13Y108_SLICE_X18Y108_DO6;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_C2 = CLBLM_L_X12Y109_SLICE_X17Y109_BO6;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_C3 = CLBLM_L_X12Y109_SLICE_X17Y109_AO5;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_C4 = CLBLM_R_X11Y110_SLICE_X14Y110_AO5;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_C5 = CLBLM_L_X12Y109_SLICE_X16Y109_CO6;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_C6 = CLBLM_L_X12Y109_SLICE_X17Y109_CO6;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_D1 = CLBLM_R_X13Y108_SLICE_X18Y108_DO6;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_D2 = CLBLM_L_X12Y109_SLICE_X17Y109_BO6;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_D3 = CLBLM_R_X11Y109_SLICE_X14Y109_DO6;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_D4 = CLBLM_R_X13Y108_SLICE_X18Y108_CO6;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_D5 = CLBLM_L_X12Y109_SLICE_X17Y109_AO5;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_D6 = CLBLM_L_X12Y109_SLICE_X16Y109_AO5;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_T1 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_A1 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_A2 = CLBLM_R_X11Y105_SLICE_X15Y105_CO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_A3 = CLBLM_R_X11Y106_SLICE_X15Y106_BO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_A4 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_A5 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_A6 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_B1 = CLBLM_R_X11Y109_SLICE_X15Y109_AO5;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_B2 = CLBLM_R_X11Y105_SLICE_X15Y105_CO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_B3 = CLBLM_R_X11Y109_SLICE_X15Y109_AO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_B4 = CLBLM_L_X10Y106_SLICE_X13Y106_AO5;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_B5 = CLBLM_R_X11Y106_SLICE_X15Y106_BO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_B6 = CLBLM_L_X10Y105_SLICE_X13Y105_CO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_C1 = CLBLM_R_X11Y106_SLICE_X15Y106_BO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_C2 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_C3 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_C4 = CLBLM_R_X11Y105_SLICE_X15Y105_CO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_C5 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_C6 = CLBLM_L_X10Y105_SLICE_X13Y105_CO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_D1 = CLBLM_R_X11Y106_SLICE_X15Y106_BO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_D2 = CLBLM_R_X11Y109_SLICE_X15Y109_AO5;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_D3 = CLBLM_R_X11Y109_SLICE_X15Y109_AO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_D4 = CLBLM_L_X10Y106_SLICE_X13Y106_AO5;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_D5 = CLBLM_L_X10Y105_SLICE_X13Y105_CO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_D6 = CLBLM_R_X11Y105_SLICE_X15Y105_CO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_D1 = 1'b1;
  assign LIOI3_X0Y109_ILOGIC_X0Y110_D = LIOB33_X0Y109_IOB_X0Y110_I;
  assign LIOI3_X0Y109_ILOGIC_X0Y109_D = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_A1 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_A2 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_A3 = CLBLM_L_X8Y105_SLICE_X11Y105_AO6;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_A4 = CLBLM_L_X10Y105_SLICE_X12Y105_AO6;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_A5 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_A6 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_B1 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_B2 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_B3 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_B4 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_B5 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_B6 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_C1 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_C2 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_C3 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_C4 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_C5 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_C6 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_D1 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_A1 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_A2 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_A3 = CLBLM_R_X5Y111_SLICE_X6Y111_BO6;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_D5 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_D6 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_A4 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_A5 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_A6 = CLBLM_R_X3Y111_SLICE_X3Y111_CO6;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_D2 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_D3 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_B3 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_B4 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_B5 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_B6 = CLBLL_L_X4Y112_SLICE_X4Y112_CO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_B1 = CLBLM_R_X3Y111_SLICE_X2Y111_DO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_B2 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_A1 = CLBLM_R_X7Y106_SLICE_X9Y106_CO6;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_A2 = CLBLM_R_X7Y105_SLICE_X8Y105_DO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_C1 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_C2 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_C3 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_C4 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_C5 = CLBLL_L_X4Y111_SLICE_X4Y111_DO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_C6 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_B1 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_B2 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_B3 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_B4 = CLBLM_L_X8Y105_SLICE_X10Y105_DO6;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_B5 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_B6 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_D1 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_D2 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_D3 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_D4 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_D5 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_D6 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_C1 = CLBLM_L_X10Y105_SLICE_X12Y105_AO6;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_C2 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_C3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_C4 = CLBLM_L_X10Y106_SLICE_X12Y106_AO6;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_C5 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_C6 = CLBLM_L_X8Y106_SLICE_X10Y106_BO6;
  assign RIOI3_X105Y111_ILOGIC_X1Y111_D = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_D1 = CLBLM_L_X10Y105_SLICE_X12Y105_AO6;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_D2 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_D3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_D4 = CLBLM_L_X10Y106_SLICE_X12Y106_AO6;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_D5 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_D6 = CLBLM_L_X8Y106_SLICE_X10Y106_BO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_A1 = CLBLL_L_X4Y111_SLICE_X5Y111_DO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_A2 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_A3 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_A4 = CLBLM_R_X3Y111_SLICE_X2Y111_BO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_A5 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_A6 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_B1 = CLBLM_R_X5Y111_SLICE_X7Y111_DO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_B2 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_B4 = CLBLL_L_X4Y111_SLICE_X4Y111_BO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_B5 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_B6 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_B2 = CLBLM_R_X7Y110_SLICE_X9Y110_BO5;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_C1 = CLBLL_L_X4Y112_SLICE_X5Y112_AO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_C2 = CLBLM_R_X5Y111_SLICE_X7Y111_CO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_C3 = CLBLL_L_X4Y111_SLICE_X4Y111_BO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_C4 = CLBLM_R_X7Y111_SLICE_X8Y111_DO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_C5 = CLBLM_R_X5Y111_SLICE_X7Y111_DO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_C6 = CLBLL_L_X4Y112_SLICE_X5Y112_DO6;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_A1 = CLBLM_R_X11Y108_SLICE_X15Y108_AO5;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_A2 = CLBLM_R_X11Y110_SLICE_X14Y110_BO6;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_A3 = CLBLM_R_X11Y108_SLICE_X15Y108_BO6;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_A4 = CLBLM_R_X13Y108_SLICE_X19Y108_AO6;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_A5 = CLBLM_L_X12Y108_SLICE_X16Y108_AO5;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_A6 = CLBLM_L_X10Y107_SLICE_X13Y107_AO6;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_B1 = CLBLM_R_X11Y108_SLICE_X15Y108_AO5;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_D1 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_D2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_D3 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_D4 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_D5 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_D6 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_B3 = CLBLM_R_X11Y108_SLICE_X15Y108_BO6;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_B4 = CLBLM_L_X12Y108_SLICE_X16Y108_AO5;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_B6 = CLBLM_L_X10Y107_SLICE_X13Y107_AO6;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_C1 = CLBLM_L_X12Y110_SLICE_X17Y110_BO6;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_C2 = CLBLM_L_X12Y110_SLICE_X17Y110_CO6;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_C3 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_C4 = CLBLM_L_X12Y108_SLICE_X16Y108_CO6;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_C5 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_C6 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_D1 = CLBLM_L_X12Y110_SLICE_X17Y110_BO6;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_D2 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_D3 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_D4 = CLBLM_L_X12Y108_SLICE_X16Y108_CO6;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_D5 = CLBLM_L_X12Y109_SLICE_X17Y109_CO6;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_D6 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_A1 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_A2 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_A3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_A4 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_A5 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_A6 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_B1 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_B2 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_B3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_B4 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_B5 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_B6 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_C1 = CLBLM_L_X12Y109_SLICE_X16Y109_BO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_C2 = CLBLM_R_X11Y110_SLICE_X15Y110_AO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_C3 = CLBLM_R_X11Y110_SLICE_X15Y110_BO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_C4 = CLBLM_R_X11Y110_SLICE_X14Y110_AO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_C5 = CLBLM_R_X11Y110_SLICE_X14Y110_BO5;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_C6 = CLBLM_L_X10Y108_SLICE_X12Y108_CO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_D1 = CLBLM_L_X12Y109_SLICE_X16Y109_BO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_D2 = CLBLM_L_X12Y109_SLICE_X17Y109_CO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_D3 = CLBLM_R_X11Y110_SLICE_X15Y110_BO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_D4 = CLBLM_R_X11Y110_SLICE_X14Y110_AO5;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_D5 = CLBLM_R_X11Y110_SLICE_X14Y110_BO5;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_D6 = CLBLM_L_X12Y109_SLICE_X16Y109_CO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_A1 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_A2 = CLBLM_L_X8Y107_SLICE_X10Y107_BO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_A3 = 1'b1;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_A4 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_A5 = CLBLM_L_X8Y104_SLICE_X10Y104_AO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_A6 = 1'b1;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_B1 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_B2 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_B3 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_B4 = CLBLM_L_X8Y107_SLICE_X10Y107_DO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_B5 = CLBLM_L_X8Y107_SLICE_X11Y107_AO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_B6 = CLBLM_R_X7Y106_SLICE_X9Y106_AO5;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_C3 = 1'b1;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_C1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_C2 = CLBLM_L_X10Y107_SLICE_X13Y107_BO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_C3 = CLBLM_L_X10Y107_SLICE_X12Y107_DO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_C4 = CLBLL_L_X2Y107_SLICE_X0Y107_CO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_C5 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_C6 = CLBLM_L_X12Y107_SLICE_X16Y107_AO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A1 = CLBLL_L_X4Y110_SLICE_X5Y110_DO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A2 = CLBLL_L_X4Y111_SLICE_X4Y111_CO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A3 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A4 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A5 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A6 = 1'b1;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_D4 = 1'b1;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_D5 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B1 = CLBLL_L_X4Y115_SLICE_X4Y115_CO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B2 = CLBLL_L_X4Y113_SLICE_X5Y113_BO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B3 = CLBLM_R_X3Y112_SLICE_X2Y112_BO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B4 = CLBLM_R_X3Y112_SLICE_X2Y112_AO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B5 = CLBLL_L_X4Y112_SLICE_X4Y112_BO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B6 = CLBLL_L_X4Y113_SLICE_X5Y113_DO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_D6 = 1'b1;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_A1 = 1'b1;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_A2 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C2 = CLBLM_R_X3Y112_SLICE_X2Y112_BO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C3 = CLBLL_L_X4Y113_SLICE_X5Y113_DO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C4 = CLBLL_L_X4Y113_SLICE_X5Y113_BO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C5 = CLBLL_L_X4Y115_SLICE_X4Y115_CO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_A3 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_A4 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_A5 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_A6 = 1'b1;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_B1 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_B2 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_B3 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_B4 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D1 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D2 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D3 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D4 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D5 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D6 = 1'b1;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_B5 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_B6 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_C1 = CLBLM_L_X8Y107_SLICE_X10Y107_AO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_C2 = CLBLM_L_X8Y105_SLICE_X10Y105_BO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_C3 = CLBLM_L_X10Y108_SLICE_X13Y108_BO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_C4 = CLBLM_L_X12Y108_SLICE_X16Y108_AO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_C5 = CLBLM_R_X7Y104_SLICE_X9Y104_DO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_C6 = CLBLM_L_X8Y105_SLICE_X10Y105_CO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_D1 = CLBLM_L_X8Y104_SLICE_X10Y104_AO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_D2 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_D3 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_D4 = CLBLM_L_X10Y107_SLICE_X13Y107_BO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_D5 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_D6 = CLBLM_L_X8Y107_SLICE_X10Y107_BO6;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_D3 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_D4 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A1 = CLBLL_L_X4Y113_SLICE_X4Y113_AO5;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A2 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A3 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A4 = CLBLL_L_X4Y112_SLICE_X5Y112_BO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A6 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B1 = CLBLL_L_X4Y113_SLICE_X4Y113_AO5;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B2 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B4 = CLBLL_L_X4Y112_SLICE_X5Y112_BO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B5 = CLBLL_L_X4Y113_SLICE_X5Y113_CO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B6 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C1 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C2 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C3 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C4 = CLBLL_L_X4Y112_SLICE_X5Y112_AO5;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C5 = CLBLL_L_X4Y110_SLICE_X5Y110_DO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C6 = CLBLL_L_X4Y111_SLICE_X4Y111_CO6;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_A1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_A2 = CLBLM_L_X12Y108_SLICE_X17Y108_CO6;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_A3 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_A4 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_A5 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_A6 = CLBLM_L_X12Y109_SLICE_X17Y109_BO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D1 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D2 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D3 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D4 = CLBLL_L_X4Y112_SLICE_X5Y112_AO5;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D5 = CLBLL_L_X4Y110_SLICE_X5Y110_DO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D6 = CLBLL_L_X4Y111_SLICE_X4Y111_CO6;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_B1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_B2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_B3 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_B4 = CLBLM_L_X12Y108_SLICE_X17Y108_CO6;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_B5 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_B6 = CLBLM_L_X12Y109_SLICE_X17Y109_BO6;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_C1 = CLBLM_R_X11Y112_SLICE_X15Y112_AO5;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_C2 = CLBLM_R_X11Y111_SLICE_X14Y111_AO5;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_C3 = CLBLM_R_X11Y110_SLICE_X15Y110_DO6;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_C4 = CLBLM_L_X12Y110_SLICE_X16Y110_AO5;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_C5 = CLBLM_R_X11Y109_SLICE_X15Y109_DO6;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_C6 = CLBLM_R_X11Y111_SLICE_X15Y111_BO6;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_D1 = CLBLM_R_X11Y111_SLICE_X15Y111_AO6;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_D2 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_D3 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_D4 = CLBLM_L_X12Y110_SLICE_X16Y110_DO6;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_D5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_D6 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_A1 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_A2 = 1'b1;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_A3 = 1'b1;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_A4 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_A5 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_A6 = 1'b1;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_B1 = CLBLM_R_X11Y111_SLICE_X14Y111_CO6;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_B2 = CLBLM_L_X10Y110_SLICE_X12Y110_BO6;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_B3 = CLBLM_R_X11Y111_SLICE_X15Y111_AO6;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_B4 = CLBLM_L_X10Y110_SLICE_X13Y110_AO6;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_B5 = CLBLM_R_X11Y111_SLICE_X14Y111_AO6;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_B6 = CLBLM_R_X11Y111_SLICE_X14Y111_AO5;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_C1 = CLBLM_R_X11Y109_SLICE_X14Y109_CO6;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_C2 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_B1 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_C3 = CLBLM_R_X13Y108_SLICE_X18Y108_CO6;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_C4 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_C5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_C6 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_B2 = CLBLM_L_X12Y111_SLICE_X16Y111_BO6;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_B3 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_D1 = CLBLM_R_X11Y111_SLICE_X14Y111_AO6;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_D2 = CLBLM_L_X10Y110_SLICE_X12Y110_BO6;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_D3 = CLBLM_R_X11Y111_SLICE_X15Y111_AO6;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_D4 = CLBLM_R_X11Y111_SLICE_X14Y111_AO5;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_D5 = CLBLM_R_X11Y111_SLICE_X14Y111_CO6;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_D6 = CLBLM_L_X10Y110_SLICE_X13Y110_AO6;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_C2 = CLBLM_R_X11Y114_SLICE_X14Y114_AO6;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_C3 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_C4 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_C5 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_B2 = CLBLM_R_X11Y110_SLICE_X14Y110_BO6;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_C6 = CLBLM_L_X10Y114_SLICE_X12Y114_BO6;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_B5 = CLBLM_R_X13Y108_SLICE_X19Y108_AO6;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_A1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_A2 = 1'b1;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_A3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_A4 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_A5 = 1'b1;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_A6 = 1'b1;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_B1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_B2 = CLBLM_L_X8Y107_SLICE_X11Y107_BO6;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_B3 = CLBLM_L_X8Y106_SLICE_X10Y106_AO6;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_B4 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_B5 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_B6 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_D1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_C1 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_C2 = CLBLM_L_X8Y107_SLICE_X10Y107_DO6;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_C3 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_C4 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_C5 = CLBLM_R_X7Y104_SLICE_X9Y104_DO6;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_C6 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_A1 = CLBLL_L_X4Y115_SLICE_X4Y115_CO6;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_A2 = CLBLL_L_X4Y113_SLICE_X5Y113_BO6;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_A3 = CLBLM_R_X3Y112_SLICE_X2Y112_AO6;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_A4 = CLBLL_L_X4Y113_SLICE_X5Y113_DO6;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_A5 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_A6 = 1'b1;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_D1 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_B1 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_B2 = 1'b1;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_D4 = CLBLM_L_X8Y106_SLICE_X10Y106_AO6;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_D5 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_B3 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_D5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_D6 = CLBLM_L_X8Y107_SLICE_X11Y107_BO6;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_B4 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_B5 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_B6 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_C1 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_C2 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_C3 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_C4 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_C5 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_C6 = 1'b1;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_A1 = CLBLM_R_X7Y108_SLICE_X9Y108_AO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_A2 = CLBLM_L_X8Y107_SLICE_X10Y107_AO5;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_A3 = CLBLM_L_X8Y108_SLICE_X11Y108_AO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_A4 = CLBLM_L_X8Y108_SLICE_X10Y108_BO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_A5 = CLBLM_L_X8Y106_SLICE_X10Y106_AO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_A6 = CLBLM_L_X8Y107_SLICE_X10Y107_CO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_B2 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_B3 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_B4 = CLBLM_L_X8Y107_SLICE_X10Y107_DO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_B5 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_B6 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_B1 = CLBLM_R_X7Y104_SLICE_X9Y104_DO6;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_D1 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_D2 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_D3 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_D4 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_D5 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_D6 = 1'b1;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_C1 = CLBLM_L_X8Y106_SLICE_X10Y106_AO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_C2 = CLBLM_L_X8Y107_SLICE_X10Y107_AO5;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_C3 = CLBLM_L_X8Y108_SLICE_X11Y108_AO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_C4 = CLBLM_L_X8Y107_SLICE_X10Y107_CO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_C5 = CLBLM_R_X7Y108_SLICE_X9Y108_AO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_C6 = CLBLM_L_X8Y108_SLICE_X10Y108_BO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_D1 = CLBLM_L_X8Y106_SLICE_X10Y106_AO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_D2 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_D3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_D4 = CLBLM_L_X8Y107_SLICE_X10Y107_CO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_D5 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_D6 = CLBLM_L_X8Y108_SLICE_X10Y108_BO6;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_A1 = CLBLM_R_X7Y111_SLICE_X8Y111_DO6;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_A2 = CLBLM_R_X5Y111_SLICE_X7Y111_CO6;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_A3 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_A4 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_A5 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_A6 = 1'b1;
  assign LIOI3_X0Y111_ILOGIC_X0Y112_D = LIOB33_X0Y111_IOB_X0Y112_I;
  assign LIOI3_X0Y111_ILOGIC_X0Y111_D = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_B1 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_B2 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_B3 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_B4 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_B5 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_B6 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_A6 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_C1 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_C2 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_C3 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_C4 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_C5 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_C6 = 1'b1;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_A1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_A2 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_A3 = 1'b1;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_A4 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_D1 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_D2 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_D3 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_D4 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_D5 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_D6 = 1'b1;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_A5 = 1'b1;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_A6 = 1'b1;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_B1 = CLBLM_L_X12Y110_SLICE_X16Y110_AO5;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_B3 = 1'b1;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_B2 = CLBLM_R_X11Y111_SLICE_X15Y111_BO6;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_B3 = CLBLM_R_X11Y109_SLICE_X15Y109_DO6;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_B4 = CLBLM_R_X11Y110_SLICE_X15Y110_DO6;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_B5 = CLBLM_R_X11Y111_SLICE_X14Y111_AO5;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_B6 = CLBLM_R_X11Y112_SLICE_X15Y112_AO5;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_C1 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_C2 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_C3 = CLBLM_R_X11Y110_SLICE_X15Y110_DO6;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_C4 = CLBLM_R_X11Y109_SLICE_X15Y109_DO6;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_C5 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_C6 = CLBLM_R_X11Y111_SLICE_X15Y111_BO6;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_D1 = CLBLM_R_X11Y111_SLICE_X15Y111_AO6;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_D2 = CLBLM_L_X12Y110_SLICE_X16Y110_DO6;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_D3 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_D4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_D5 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_D6 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_A1 = CLBLM_L_X10Y109_SLICE_X13Y109_DO6;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_A2 = CLBLM_L_X10Y113_SLICE_X13Y113_AO5;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_A3 = CLBLM_R_X11Y112_SLICE_X15Y112_AO6;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_A4 = CLBLM_L_X12Y111_SLICE_X16Y111_CO6;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_A5 = CLBLM_R_X11Y110_SLICE_X14Y110_DO6;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_A6 = CLBLM_L_X10Y111_SLICE_X13Y111_AO5;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_B1 = CLBLM_L_X10Y109_SLICE_X13Y109_DO6;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_B2 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_B3 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_B4 = CLBLM_L_X12Y111_SLICE_X16Y111_CO6;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_B5 = CLBLM_R_X11Y110_SLICE_X14Y110_DO6;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_B6 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_C1 = CLBLM_R_X11Y110_SLICE_X14Y110_DO6;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_C2 = CLBLM_R_X11Y112_SLICE_X15Y112_AO6;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_C3 = CLBLM_L_X10Y109_SLICE_X13Y109_DO6;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_C4 = CLBLM_L_X10Y111_SLICE_X13Y111_AO5;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_C5 = CLBLM_L_X12Y111_SLICE_X16Y111_CO6;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_C6 = CLBLM_L_X10Y113_SLICE_X13Y113_AO5;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_D1 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_D2 = CLBLM_L_X12Y111_SLICE_X16Y111_DO6;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_D3 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_D4 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_D5 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_D6 = CLBLM_R_X11Y110_SLICE_X15Y110_DO6;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_A1 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_A2 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_A3 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_A4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_A5 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_A6 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_B1 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_B2 = CLBLM_L_X10Y107_SLICE_X12Y107_CO6;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_B3 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_B4 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_B5 = CLBLM_L_X8Y108_SLICE_X11Y108_CO6;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_B6 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_C1 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_A1 = CLBLL_L_X4Y114_SLICE_X5Y114_AO5;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_A2 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_A3 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_C5 = CLBLM_L_X8Y109_SLICE_X11Y109_DO6;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_C6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_A4 = CLBLL_L_X4Y112_SLICE_X5Y112_CO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_A5 = CLBLL_L_X4Y112_SLICE_X5Y112_BO5;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_A6 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_C2 = CLBLM_R_X7Y109_SLICE_X9Y109_DO6;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_C3 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_C4 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_B1 = CLBLM_R_X5Y115_SLICE_X7Y115_AO5;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_B2 = CLBLL_L_X4Y116_SLICE_X5Y116_DO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_B3 = CLBLL_L_X4Y113_SLICE_X5Y113_AO5;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_B4 = CLBLL_L_X4Y114_SLICE_X4Y114_BO6;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_D3 = CLBLM_L_X10Y109_SLICE_X12Y109_DO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_B5 = CLBLL_L_X4Y112_SLICE_X5Y112_BO5;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_D5 = CLBLM_L_X8Y108_SLICE_X11Y108_DO6;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_D6 = CLBLM_L_X8Y109_SLICE_X11Y109_BO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_B6 = CLBLL_L_X4Y114_SLICE_X5Y114_AO5;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_D1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_C1 = CLBLL_L_X4Y115_SLICE_X4Y115_AO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_C2 = CLBLM_R_X5Y115_SLICE_X7Y115_AO5;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_C3 = CLBLL_L_X4Y113_SLICE_X5Y113_BO5;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_C4 = CLBLL_L_X4Y115_SLICE_X4Y115_AO5;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_C5 = CLBLL_L_X4Y113_SLICE_X5Y113_AO5;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_C6 = CLBLL_L_X4Y116_SLICE_X5Y116_DO6;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_A1 = CLBLM_L_X10Y106_SLICE_X13Y106_CO6;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_A2 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_A3 = CLBLM_L_X8Y106_SLICE_X11Y106_AO6;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_A4 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_A5 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_A6 = CLBLM_L_X8Y106_SLICE_X10Y106_DO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_D1 = CLBLL_L_X4Y115_SLICE_X4Y115_AO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_D2 = CLBLL_L_X4Y113_SLICE_X5Y113_AO5;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_D3 = CLBLM_R_X5Y115_SLICE_X7Y115_AO5;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_C5 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_D4 = CLBLL_L_X4Y115_SLICE_X4Y115_AO5;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_D5 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_D6 = CLBLL_L_X4Y116_SLICE_X5Y116_DO6;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_B1 = CLBLM_L_X10Y106_SLICE_X13Y106_CO6;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_B2 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_B3 = CLBLM_L_X8Y106_SLICE_X11Y106_AO6;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_B4 = CLBLM_L_X8Y106_SLICE_X10Y106_DO6;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_B5 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_B6 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_C1 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_C2 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_C3 = CLBLM_L_X8Y109_SLICE_X11Y109_DO6;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_C4 = CLBLM_R_X7Y109_SLICE_X9Y109_DO6;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_C5 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_C6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_D1 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_D2 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_D3 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_D4 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_D5 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_A1 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_A2 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_A3 = CLBLM_R_X7Y114_SLICE_X9Y114_DO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_A4 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_A5 = CLBLM_R_X7Y114_SLICE_X8Y114_BO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_A6 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_D6 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_B1 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_B2 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_B3 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_B4 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_B5 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_B6 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_C1 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_C2 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_C3 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_C4 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_C5 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_C6 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_D1 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_D2 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_D3 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_D4 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_D5 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_D6 = 1'b1;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_A1 = CLBLM_R_X11Y110_SLICE_X15Y110_DO6;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_A2 = CLBLM_L_X12Y111_SLICE_X16Y111_DO6;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_A3 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_B1 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_D5 = 1'b1;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_B2 = 1'b1;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_B3 = 1'b1;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_B4 = 1'b1;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_B5 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_D6 = 1'b1;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_B6 = 1'b1;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_C1 = 1'b1;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_C2 = 1'b1;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_C3 = 1'b1;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_C4 = 1'b1;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_C5 = 1'b1;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_C6 = 1'b1;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_D1 = 1'b1;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_D2 = 1'b1;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_D3 = 1'b1;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_D4 = 1'b1;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_D5 = 1'b1;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_D6 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_D4 = 1'b1;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_A1 = CLBLM_R_X11Y109_SLICE_X15Y109_CO6;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_A2 = CLBLM_L_X10Y113_SLICE_X13Y113_AO5;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_A3 = CLBLM_L_X12Y111_SLICE_X16Y111_AO6;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_A4 = CLBLM_L_X10Y113_SLICE_X13Y113_AO6;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_A5 = CLBLM_L_X12Y110_SLICE_X17Y110_AO6;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_A6 = CLBLM_L_X12Y110_SLICE_X16Y110_AO5;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_B1 = CLBLM_R_X11Y109_SLICE_X15Y109_CO6;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_B2 = CLBLM_L_X12Y111_SLICE_X16Y111_AO6;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_B3 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_B4 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_B5 = CLBLM_L_X12Y110_SLICE_X17Y110_AO6;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_B6 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_C1 = CLBLM_L_X12Y110_SLICE_X17Y110_AO6;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_C2 = CLBLM_L_X12Y111_SLICE_X16Y111_AO6;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_C3 = CLBLM_L_X10Y113_SLICE_X13Y113_AO5;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_C4 = CLBLM_L_X12Y110_SLICE_X16Y110_AO5;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_C5 = CLBLM_R_X11Y109_SLICE_X15Y109_CO6;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_C6 = CLBLM_L_X10Y113_SLICE_X13Y113_AO6;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_D1 = CLBLM_R_X11Y112_SLICE_X15Y112_BO6;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_D2 = CLBLM_R_X11Y113_SLICE_X15Y113_AO6;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_D3 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_D4 = CLBLM_R_X11Y114_SLICE_X14Y114_CO6;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_D5 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_D6 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_A3 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_A4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_A5 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_A6 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_B6 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_C4 = CLBLM_R_X5Y112_SLICE_X6Y112_AO5;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_C5 = CLBLM_R_X3Y114_SLICE_X3Y114_AO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_A1 = CLBLM_L_X8Y110_SLICE_X11Y110_BO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_A2 = CLBLM_L_X10Y111_SLICE_X13Y111_AO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_A3 = CLBLM_R_X7Y109_SLICE_X9Y109_DO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_A4 = CLBLM_L_X8Y109_SLICE_X11Y109_AO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_A5 = CLBLM_L_X10Y110_SLICE_X12Y110_DO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_A6 = CLBLM_R_X7Y109_SLICE_X8Y109_AO5;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_C6 = CLBLM_R_X5Y113_SLICE_X6Y113_BO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_B1 = CLBLM_L_X8Y108_SLICE_X11Y108_DO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_B2 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_B3 = CLBLM_L_X8Y109_SLICE_X11Y109_BO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_B4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_B5 = CLBLM_L_X10Y108_SLICE_X12Y108_BO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_B6 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_A1 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_A2 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_A3 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_A4 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_C1 = CLBLM_L_X10Y108_SLICE_X12Y108_BO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_C2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_A5 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_A6 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_C3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_C5 = CLBLM_L_X8Y108_SLICE_X11Y108_DO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_B1 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_B2 = CLBLL_L_X4Y116_SLICE_X5Y116_DO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_B3 = CLBLM_R_X5Y115_SLICE_X7Y115_DO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_B4 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_B5 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_B6 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_D1 = CLBLM_L_X8Y109_SLICE_X11Y109_AO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_C1 = CLBLL_L_X4Y115_SLICE_X4Y115_BO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_C2 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_C3 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_C4 = CLBLL_L_X4Y113_SLICE_X5Y113_BO5;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_C5 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_C6 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_D2 = CLBLM_R_X7Y109_SLICE_X8Y109_AO5;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_D3 = CLBLM_L_X10Y110_SLICE_X12Y110_DO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_D4 = CLBLM_R_X7Y109_SLICE_X9Y109_DO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_D5 = CLBLM_L_X10Y111_SLICE_X13Y111_AO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_D6 = CLBLM_L_X8Y110_SLICE_X11Y110_BO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_A1 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_A2 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_D1 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_D2 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_D3 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_D4 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_D5 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_D6 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_A3 = CLBLM_L_X8Y106_SLICE_X11Y106_AO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_A4 = CLBLM_L_X10Y106_SLICE_X13Y106_CO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_A5 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_A6 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_B1 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_B2 = CLBLM_L_X10Y109_SLICE_X12Y109_BO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_B3 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_B4 = CLBLM_L_X8Y109_SLICE_X10Y109_BO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_B5 = CLBLM_L_X8Y110_SLICE_X10Y110_AO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_B6 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_C1 = CLBLM_L_X8Y110_SLICE_X10Y110_AO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_C2 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_C3 = CLBLM_L_X10Y109_SLICE_X12Y109_BO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_C4 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_C5 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_C6 = CLBLM_L_X8Y109_SLICE_X10Y109_BO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_A1 = CLBLM_R_X5Y115_SLICE_X6Y115_DO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_A2 = CLBLM_R_X5Y114_SLICE_X6Y114_CO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_D3 = CLBLM_L_X8Y110_SLICE_X11Y110_BO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_A3 = CLBLM_R_X5Y115_SLICE_X6Y115_CO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_D4 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_D5 = CLBLM_L_X10Y110_SLICE_X12Y110_DO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_D6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_A4 = CLBLM_R_X7Y116_SLICE_X8Y116_BO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_A5 = CLBLL_L_X4Y116_SLICE_X5Y116_CO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_A6 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_D2 = CLBLM_R_X7Y109_SLICE_X9Y109_DO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_B1 = CLBLM_R_X5Y116_SLICE_X7Y116_BO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_B2 = CLBLM_R_X5Y116_SLICE_X6Y116_AO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_B3 = CLBLM_R_X5Y116_SLICE_X7Y116_AO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_B4 = CLBLM_R_X7Y116_SLICE_X8Y116_CO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_B5 = CLBLM_R_X5Y115_SLICE_X7Y115_BO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_B6 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_C1 = CLBLM_R_X7Y116_SLICE_X9Y116_AO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_C2 = CLBLM_R_X7Y116_SLICE_X8Y116_AO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_C3 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_C4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_C5 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_C6 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_D1 = CLBLM_R_X7Y114_SLICE_X8Y114_CO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_D2 = CLBLL_L_X4Y116_SLICE_X4Y116_AO5;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_D3 = CLBLM_R_X5Y116_SLICE_X6Y116_DO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_D4 = CLBLL_L_X4Y115_SLICE_X5Y115_AO5;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_D5 = CLBLM_R_X5Y116_SLICE_X7Y116_AO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_D6 = CLBLM_R_X5Y115_SLICE_X7Y115_AO6;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_A1 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_A2 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_A3 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_A4 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_A5 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_A6 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_B1 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_B2 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_B3 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_B4 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_B5 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_B6 = 1'b1;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_A1 = 1'b1;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_A2 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_A3 = 1'b1;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_A4 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_A5 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_A6 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_C1 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_C2 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_C3 = 1'b1;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_B1 = CLBLM_L_X8Y105_SLICE_X10Y105_AO6;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_B2 = CLBLM_R_X7Y104_SLICE_X9Y104_AO6;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_B3 = CLBLM_R_X7Y104_SLICE_X8Y104_AO6;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_B4 = CLBLM_L_X8Y104_SLICE_X10Y104_AO6;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_B5 = CLBLM_R_X7Y104_SLICE_X9Y104_CO6;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_B6 = CLBLM_R_X7Y104_SLICE_X9Y104_AO5;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_D1 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_D2 = 1'b1;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_C1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_C2 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_C3 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_C4 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_C5 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_C6 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_D3 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_D4 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_A1 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_A2 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_A3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_A4 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_A5 = CLBLM_L_X12Y111_SLICE_X16Y111_AO6;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_A6 = CLBLM_R_X11Y110_SLICE_X15Y110_CO6;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_D1 = CLBLM_R_X7Y104_SLICE_X9Y104_CO6;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_D2 = CLBLM_R_X7Y104_SLICE_X9Y104_AO6;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_D3 = CLBLM_L_X8Y105_SLICE_X10Y105_AO6;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_D4 = CLBLM_R_X7Y104_SLICE_X9Y104_AO5;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_D5 = CLBLM_R_X7Y104_SLICE_X8Y104_AO6;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_D6 = CLBLM_L_X8Y104_SLICE_X10Y104_AO6;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_B1 = CLBLM_R_X11Y113_SLICE_X15Y113_AO6;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_B2 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_B3 = CLBLM_R_X11Y112_SLICE_X15Y112_BO6;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_B4 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_B5 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_A1 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_A2 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_A3 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_A4 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_A5 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_A6 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_C1 = CLBLM_L_X12Y111_SLICE_X16Y111_AO6;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_C2 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_C3 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_B1 = 1'b1;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_B2 = 1'b1;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_B3 = 1'b1;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_B4 = 1'b1;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_B5 = 1'b1;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_B6 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_D1 = CLBLM_R_X11Y112_SLICE_X15Y112_CO6;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_D2 = CLBLM_R_X11Y113_SLICE_X15Y113_AO6;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_D3 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_C1 = 1'b1;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_C2 = 1'b1;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_C3 = 1'b1;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_C4 = 1'b1;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_C5 = 1'b1;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_C6 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_D4 = CLBLM_R_X11Y114_SLICE_X14Y114_CO6;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_D5 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_D6 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_D1 = 1'b1;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_D2 = 1'b1;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_D3 = 1'b1;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_D4 = 1'b1;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_D5 = 1'b1;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_D6 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_A1 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_A2 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_A3 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_A4 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_A5 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_A6 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_B1 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_B2 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_B3 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_B4 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_B5 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_B6 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_C1 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_C2 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_C3 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_C4 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_C5 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_C6 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_D1 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_D2 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_D3 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_D4 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_D5 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_D6 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_A1 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_A2 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_A3 = CLBLM_L_X8Y110_SLICE_X10Y110_AO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_A4 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_A5 = CLBLM_L_X10Y109_SLICE_X12Y109_BO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_A6 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_B1 = CLBLM_L_X10Y111_SLICE_X12Y111_AO5;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_B2 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_B3 = CLBLM_L_X8Y110_SLICE_X10Y110_BO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_B4 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_B5 = CLBLM_L_X8Y111_SLICE_X10Y111_AO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_C1 = CLBLM_R_X7Y109_SLICE_X8Y109_CO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_C2 = CLBLM_L_X8Y112_SLICE_X10Y112_AO5;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_C3 = CLBLM_L_X8Y110_SLICE_X11Y110_DO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_C4 = CLBLM_R_X7Y110_SLICE_X9Y110_AO5;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_C5 = CLBLM_L_X8Y110_SLICE_X11Y110_AO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_C6 = CLBLM_L_X10Y110_SLICE_X13Y110_BO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_D1 = CLBLM_L_X8Y111_SLICE_X10Y111_AO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_D2 = CLBLM_L_X8Y110_SLICE_X10Y110_BO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_D3 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_D4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_D5 = CLBLM_L_X10Y111_SLICE_X12Y111_AO5;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_D6 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_D5 = CLBLL_L_X4Y114_SLICE_X5Y114_AO6;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_A1 = CLBLM_R_X7Y104_SLICE_X9Y104_DO6;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_A2 = CLBLM_R_X7Y104_SLICE_X9Y104_BO6;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_A3 = CLBLM_R_X7Y105_SLICE_X8Y105_AO5;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_A4 = CLBLM_R_X7Y105_SLICE_X8Y105_DO6;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_A5 = CLBLM_L_X8Y107_SLICE_X10Y107_AO6;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_A6 = CLBLM_L_X8Y105_SLICE_X10Y105_BO6;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_B1 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_B2 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_B3 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_B4 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_B5 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_B6 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_C1 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_C2 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_C3 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_C4 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_C5 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_C6 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_D1 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_D2 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_D3 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_D4 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_D5 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_D6 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_A1 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_A2 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_A3 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_A4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_A5 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_A6 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_B1 = CLBLM_R_X7Y106_SLICE_X8Y106_CO6;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_B2 = CLBLM_R_X7Y104_SLICE_X9Y104_AO6;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_B3 = CLBLM_R_X7Y106_SLICE_X8Y106_AO6;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_B4 = CLBLM_R_X7Y104_SLICE_X8Y104_AO6;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_B5 = CLBLM_R_X5Y105_SLICE_X7Y105_AO6;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_B6 = CLBLM_R_X7Y106_SLICE_X8Y106_AO5;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_C1 = CLBLM_R_X7Y105_SLICE_X8Y105_AO6;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_C2 = CLBLL_L_X4Y105_SLICE_X4Y105_DO6;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_C3 = CLBLM_R_X7Y105_SLICE_X8Y105_DO6;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_C4 = CLBLM_R_X7Y105_SLICE_X8Y105_AO5;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_C5 = CLBLM_R_X7Y105_SLICE_X8Y105_BO6;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_C6 = CLBLM_R_X7Y104_SLICE_X9Y104_BO6;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_D1 = CLBLM_R_X5Y105_SLICE_X7Y105_AO6;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_D2 = CLBLM_R_X7Y104_SLICE_X9Y104_AO6;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_D3 = CLBLM_R_X7Y106_SLICE_X8Y106_AO6;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_D4 = CLBLM_R_X7Y106_SLICE_X8Y106_AO5;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_D5 = CLBLM_R_X7Y106_SLICE_X8Y106_CO6;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_D6 = CLBLM_R_X7Y104_SLICE_X8Y104_AO6;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_A1 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_A2 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_A3 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_A4 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_A5 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_A6 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_B1 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_B2 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_B3 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_B4 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_B5 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_B6 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_C1 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_C2 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_C3 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_C4 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_C5 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_C6 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_D1 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_D2 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_D3 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_D4 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_D5 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_D6 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_A1 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_A2 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_A3 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_A4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_A5 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_A6 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_B1 = CLBLM_L_X10Y110_SLICE_X13Y110_CO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_B2 = CLBLM_L_X8Y109_SLICE_X11Y109_CO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_B3 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_B4 = CLBLM_L_X10Y113_SLICE_X12Y113_AO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_B5 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_B6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_C1 = CLBLM_L_X8Y112_SLICE_X10Y112_AO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_C2 = CLBLM_L_X10Y110_SLICE_X13Y110_BO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_C3 = CLBLM_R_X11Y112_SLICE_X14Y112_AO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_C4 = CLBLM_L_X8Y112_SLICE_X10Y112_AO5;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_C5 = CLBLM_L_X10Y110_SLICE_X13Y110_DO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_C6 = CLBLM_L_X8Y110_SLICE_X11Y110_DO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_D1 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_D2 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_D3 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_D4 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_D5 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_D6 = 1'b1;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_D1 = CLBLL_L_X2Y112_SLICE_X0Y112_AO5;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_T1 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_A1 = CLBLM_R_X7Y104_SLICE_X8Y104_AO6;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_A2 = CLBLM_R_X7Y104_SLICE_X9Y104_CO6;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_A3 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_A4 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_A5 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_A6 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_B1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_B2 = CLBLM_R_X7Y105_SLICE_X8Y105_DO6;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_B3 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_B4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_B5 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_B6 = CLBLM_R_X7Y106_SLICE_X9Y106_CO6;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_C1 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_C2 = CLBLM_R_X7Y104_SLICE_X9Y104_CO6;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_C3 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_C4 = CLBLM_R_X7Y104_SLICE_X8Y104_AO6;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_C5 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_C6 = CLBLM_L_X8Y104_SLICE_X10Y104_AO6;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_D1 = CLBLM_R_X7Y106_SLICE_X9Y106_AO6;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_D2 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_D3 = CLBLM_R_X7Y106_SLICE_X8Y106_BO5;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_D4 = CLBLM_R_X7Y106_SLICE_X9Y106_CO6;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_D5 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_D6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_A1 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_A2 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_A3 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_A4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_A5 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_A6 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_B1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_B2 = CLBLM_R_X5Y105_SLICE_X7Y105_AO6;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_B3 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_B4 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_B5 = CLBLM_R_X7Y106_SLICE_X8Y106_CO6;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_B6 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_C1 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_C2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_C3 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_C4 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_C5 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_C6 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_D1 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_D2 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_D3 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_D4 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_D5 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_D6 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_A1 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_A2 = CLBLM_L_X10Y112_SLICE_X12Y112_CO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_A3 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_A4 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_A5 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_A6 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_B1 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_B2 = CLBLM_L_X10Y112_SLICE_X12Y112_CO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_B3 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_B4 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_B5 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_B6 = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign LIOI3_X0Y117_ILOGIC_X0Y117_D = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_C1 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_C2 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_C3 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_C4 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_C5 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_C6 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_D1 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_D2 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_D3 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_D4 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_D5 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_D6 = 1'b1;
  assign RIOI3_X105Y101_ILOGIC_X1Y102_D = RIOB33_X105Y101_IOB_X1Y102_I;
  assign RIOI3_X105Y101_ILOGIC_X1Y101_D = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_A1 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_A2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_A3 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_A4 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_A5 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_A6 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_B1 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_B2 = CLBLM_L_X10Y113_SLICE_X12Y113_AO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_B3 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_B4 = CLBLM_L_X8Y109_SLICE_X11Y109_CO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_B5 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_B6 = CLBLM_L_X10Y110_SLICE_X13Y110_BO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_C1 = CLBLM_L_X8Y114_SLICE_X11Y114_AO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_C2 = CLBLM_L_X8Y113_SLICE_X10Y113_AO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_C3 = CLBLM_L_X8Y114_SLICE_X11Y114_BO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_C4 = CLBLM_L_X8Y113_SLICE_X10Y113_AO5;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_C5 = CLBLM_L_X8Y113_SLICE_X10Y113_DO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_C6 = CLBLM_L_X10Y114_SLICE_X12Y114_AO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_D1 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_D2 = CLBLM_L_X10Y113_SLICE_X12Y113_AO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_D3 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_D4 = CLBLM_L_X10Y110_SLICE_X13Y110_BO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_D5 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_D6 = CLBLM_L_X8Y109_SLICE_X11Y109_CO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_A1 = CLBLM_R_X7Y106_SLICE_X9Y106_BO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_A2 = CLBLM_R_X7Y108_SLICE_X9Y108_AO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_A3 = CLBLM_R_X7Y105_SLICE_X9Y105_AO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_A4 = CLBLM_R_X5Y106_SLICE_X7Y106_AO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_A5 = CLBLM_R_X5Y105_SLICE_X6Y105_AO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_A6 = CLBLM_R_X7Y108_SLICE_X9Y108_AO5;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_B1 = CLBLM_R_X7Y105_SLICE_X9Y105_AO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_B2 = CLBLM_R_X7Y108_SLICE_X9Y108_AO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_B3 = CLBLM_R_X5Y105_SLICE_X6Y105_AO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_B4 = CLBLM_R_X7Y106_SLICE_X9Y106_BO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_B5 = CLBLM_R_X5Y106_SLICE_X7Y106_AO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_B6 = CLBLM_R_X7Y108_SLICE_X9Y108_AO5;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_C1 = CLBLM_R_X5Y105_SLICE_X6Y105_AO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_C2 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_C3 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_C4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_C5 = CLBLM_R_X7Y105_SLICE_X9Y105_AO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_C6 = CLBLM_R_X7Y106_SLICE_X9Y106_BO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_D1 = CLBLM_R_X5Y105_SLICE_X6Y105_AO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_D2 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_D3 = CLBLM_R_X7Y106_SLICE_X9Y106_DO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_D4 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_D5 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_D6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_A1 = 1'b1;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_A2 = 1'b1;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_A3 = 1'b1;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_A4 = 1'b1;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_A5 = 1'b1;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_A6 = 1'b1;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_B1 = 1'b1;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_B2 = 1'b1;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_B3 = 1'b1;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_B4 = 1'b1;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_B5 = 1'b1;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_B6 = 1'b1;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_C1 = 1'b1;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_C2 = 1'b1;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_C3 = 1'b1;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_C4 = 1'b1;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_C5 = 1'b1;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_C6 = 1'b1;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_D1 = 1'b1;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_D2 = 1'b1;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_D3 = 1'b1;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_D4 = 1'b1;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_D5 = 1'b1;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_D6 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_A1 = CLBLM_R_X11Y112_SLICE_X14Y112_AO6;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_A2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_A3 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_A4 = CLBLM_L_X10Y113_SLICE_X12Y113_DO6;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_A5 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_A6 = CLBLM_L_X10Y113_SLICE_X12Y113_CO6;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_B1 = CLBLM_R_X11Y112_SLICE_X14Y112_AO6;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_B2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_B3 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_B4 = CLBLM_L_X10Y113_SLICE_X12Y113_DO6;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_B5 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_B6 = CLBLM_L_X10Y113_SLICE_X12Y113_CO6;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_C1 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_C2 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_C3 = CLBLM_R_X11Y114_SLICE_X14Y114_DO6;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_C4 = CLBLM_L_X10Y114_SLICE_X12Y114_CO6;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_C5 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_C6 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_D1 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_D2 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_D3 = CLBLM_R_X11Y114_SLICE_X14Y114_DO6;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_D4 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_D5 = CLBLM_L_X10Y114_SLICE_X12Y114_CO6;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_D6 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_A1 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_A2 = CLBLM_L_X8Y113_SLICE_X11Y113_BO6;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_A3 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_A4 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_A5 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_A6 = CLBLM_L_X10Y112_SLICE_X12Y112_AO6;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_B1 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_B2 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_B3 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_B4 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_B5 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_B6 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_C4 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_C1 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_C2 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_C3 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_C4 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_C5 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_C6 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_A1 = CLBLL_L_X2Y106_SLICE_X1Y106_CO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_A2 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_A3 = CLBLL_L_X2Y106_SLICE_X1Y106_AO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_A4 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_A5 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_A6 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_C6 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_D1 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_D2 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_D3 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_D4 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_D5 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_D6 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_B1 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_B2 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_B3 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_B4 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_B5 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_C1 = CLBLL_L_X2Y106_SLICE_X1Y106_CO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_C2 = CLBLL_L_X2Y106_SLICE_X1Y106_AO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_C3 = CLBLM_R_X3Y105_SLICE_X2Y105_AO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_C4 = CLBLM_R_X3Y104_SLICE_X3Y104_AO5;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_C5 = CLBLL_L_X2Y106_SLICE_X0Y106_BO5;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_C6 = CLBLL_L_X2Y107_SLICE_X0Y107_AO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_D1 = CLBLL_L_X2Y106_SLICE_X1Y106_CO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_D2 = CLBLL_L_X2Y106_SLICE_X1Y106_AO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_D3 = CLBLM_R_X3Y105_SLICE_X2Y105_AO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_D4 = CLBLL_L_X2Y107_SLICE_X0Y107_AO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_D5 = CLBLL_L_X2Y106_SLICE_X0Y106_BO5;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_D6 = CLBLM_R_X3Y104_SLICE_X3Y104_AO5;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_D3 = CLBLL_L_X4Y112_SLICE_X5Y112_CO6;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_A1 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_A2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_A3 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_A4 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_A5 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_A6 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_A2 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_A3 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_A4 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_A5 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_A6 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_D6 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_B3 = CLBLM_R_X7Y107_SLICE_X9Y107_BO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_B4 = CLBLM_L_X8Y108_SLICE_X10Y108_CO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_B5 = CLBLM_L_X10Y110_SLICE_X12Y110_AO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_B6 = CLBLM_L_X10Y108_SLICE_X12Y108_BO6;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_B1 = CLBLM_R_X3Y105_SLICE_X2Y105_AO6;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_B2 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_B3 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_B4 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_B5 = CLBLL_L_X2Y106_SLICE_X1Y106_AO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_C4 = CLBLM_L_X8Y108_SLICE_X10Y108_DO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_C5 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_C1 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_C2 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_C3 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_C4 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_C5 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_C6 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_D2 = 1'b1;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_D3 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_D1 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_D3 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_D1 = CLBLM_R_X3Y104_SLICE_X3Y104_DO6;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_D2 = CLBLL_L_X2Y106_SLICE_X0Y106_CO6;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_D3 = CLBLL_L_X2Y106_SLICE_X0Y106_DO6;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_D4 = CLBLL_L_X2Y108_SLICE_X1Y108_AO5;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_D5 = CLBLL_L_X2Y107_SLICE_X0Y107_DO6;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_D6 = CLBLM_R_X3Y105_SLICE_X3Y105_BO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_D2 = CLBLM_R_X7Y108_SLICE_X8Y108_CO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_D6 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_A1 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_A2 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_A3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_A4 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_A5 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_A6 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_B1 = CLBLM_R_X5Y106_SLICE_X7Y106_DO6;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_B2 = CLBLM_L_X8Y108_SLICE_X10Y108_AO6;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_B3 = CLBLM_R_X7Y107_SLICE_X9Y107_AO6;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_B4 = CLBLM_R_X7Y107_SLICE_X9Y107_BO6;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_B5 = CLBLM_R_X7Y108_SLICE_X8Y108_AO6;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_B6 = CLBLM_R_X7Y108_SLICE_X8Y108_AO5;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_C1 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_C2 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_C3 = CLBLM_R_X5Y106_SLICE_X7Y106_DO6;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_C4 = CLBLM_R_X7Y107_SLICE_X9Y107_CO6;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_C5 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_C6 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_D1 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_D2 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_D3 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_D4 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_D5 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_D6 = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_D1 = CLBLL_L_X2Y108_SLICE_X1Y108_AO6;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_T1 = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_D1 = CLBLL_L_X2Y108_SLICE_X0Y108_AO5;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_T1 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_B6 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_A1 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_A2 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_A3 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_A4 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_A5 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_A6 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_C5 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_B1 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_B2 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_B3 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_B4 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_B5 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_B6 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_C1 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_C2 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_C3 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_C4 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_C5 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_C6 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_D1 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_D2 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_D3 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_D4 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_D5 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_D6 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_A1 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_A2 = CLBLM_L_X8Y114_SLICE_X11Y114_CO6;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_A3 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_A4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_A5 = CLBLM_L_X8Y115_SLICE_X10Y115_CO6;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_A6 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_B1 = CLBLM_R_X11Y114_SLICE_X14Y114_BO6;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_B2 = CLBLM_L_X10Y114_SLICE_X12Y114_AO6;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_B3 = CLBLM_L_X8Y114_SLICE_X11Y114_AO6;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_B4 = CLBLM_L_X8Y116_SLICE_X10Y116_AO6;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_B5 = CLBLM_L_X8Y113_SLICE_X10Y113_AO6;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_B6 = CLBLM_L_X10Y114_SLICE_X12Y114_CO6;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_C1 = CLBLM_L_X8Y114_SLICE_X11Y114_AO6;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_A1 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_A2 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_C4 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_C5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_A3 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_A4 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_C6 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_A5 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_A6 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_C2 = CLBLM_L_X10Y114_SLICE_X12Y114_DO6;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_B1 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_B2 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_B3 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_B4 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_B5 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_B6 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_D1 = CLBLM_L_X8Y115_SLICE_X10Y115_AO6;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_D2 = CLBLM_L_X8Y114_SLICE_X11Y114_AO6;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_C1 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_C2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_C3 = CLBLL_L_X2Y108_SLICE_X1Y108_BO5;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_C4 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_C5 = CLBLL_L_X2Y106_SLICE_X0Y106_AO6;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_C6 = CLBLL_L_X2Y106_SLICE_X1Y106_BO6;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_D4 = CLBLM_L_X10Y114_SLICE_X12Y114_AO6;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_D5 = CLBLM_L_X8Y113_SLICE_X10Y113_AO6;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_D6 = CLBLM_L_X8Y116_SLICE_X10Y116_AO6;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_D1 = CLBLL_L_X2Y107_SLICE_X0Y107_AO6;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_D2 = CLBLL_L_X2Y106_SLICE_X1Y106_AO6;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_D3 = CLBLL_L_X2Y106_SLICE_X0Y106_BO6;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_D4 = CLBLL_L_X2Y110_SLICE_X0Y110_AO6;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_D5 = CLBLL_L_X2Y107_SLICE_X0Y107_AO5;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_D6 = CLBLL_L_X2Y107_SLICE_X0Y107_BO6;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_A1 = CLBLM_R_X3Y107_SLICE_X2Y107_BO6;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_A2 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_A3 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_A4 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_A5 = CLBLL_L_X2Y107_SLICE_X1Y107_CO6;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_A6 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_A1 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_A2 = CLBLM_R_X5Y108_SLICE_X7Y108_BO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_A3 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_B1 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_B2 = CLBLL_L_X2Y107_SLICE_X0Y107_BO6;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_B3 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_B4 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_B1 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_B2 = CLBLM_L_X8Y108_SLICE_X10Y108_DO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_B3 = CLBLM_R_X7Y107_SLICE_X9Y107_BO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_B4 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_B5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_B6 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_B5 = CLBLL_L_X2Y110_SLICE_X0Y110_AO6;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_B6 = CLBLL_L_X2Y106_SLICE_X1Y106_AO6;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_C1 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_C2 = CLBLL_L_X2Y107_SLICE_X0Y107_CO6;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_C3 = CLBLL_L_X2Y108_SLICE_X1Y108_DO6;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_C4 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_C5 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_C6 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_C1 = CLBLM_R_X7Y108_SLICE_X9Y108_CO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_C2 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_C3 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_C4 = CLBLM_R_X7Y108_SLICE_X8Y108_CO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_C5 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_C6 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_D1 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_D2 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_D3 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_D4 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_D5 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_D6 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_D1 = CLBLM_R_X7Y107_SLICE_X9Y107_BO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_D2 = CLBLM_L_X8Y108_SLICE_X10Y108_DO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_D3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_D4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_D5 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_D6 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_A1 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_A2 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_A3 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_A4 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_A5 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_A6 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_B1 = CLBLM_R_X7Y108_SLICE_X9Y108_BO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_B2 = CLBLM_R_X7Y109_SLICE_X9Y109_BO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_B3 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_B4 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_B5 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_B6 = CLBLM_R_X7Y108_SLICE_X8Y108_CO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_C1 = CLBLM_R_X7Y109_SLICE_X8Y109_AO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_C2 = CLBLM_R_X5Y109_SLICE_X6Y109_AO5;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_C3 = CLBLM_R_X7Y109_SLICE_X9Y109_BO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_C4 = CLBLM_R_X7Y109_SLICE_X8Y109_AO5;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_C5 = CLBLM_R_X7Y108_SLICE_X8Y108_CO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_C6 = CLBLM_R_X7Y108_SLICE_X9Y108_BO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_D1 = CLBLM_R_X7Y109_SLICE_X8Y109_AO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_D2 = CLBLM_R_X5Y109_SLICE_X6Y109_AO5;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_D3 = CLBLM_R_X7Y109_SLICE_X9Y109_BO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_D4 = CLBLM_R_X7Y109_SLICE_X8Y109_AO5;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_D5 = CLBLM_R_X7Y108_SLICE_X8Y108_CO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_D6 = CLBLM_R_X7Y108_SLICE_X9Y108_BO6;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_A1 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_A2 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_A3 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_A4 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_A5 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_A6 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_B1 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_B2 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_B3 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_B4 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_B5 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_B6 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_C1 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_C2 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_C3 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_C4 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_C5 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_C6 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_D1 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_D2 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_D3 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_D4 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_D5 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_D6 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_A1 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_A2 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_A3 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_A4 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_A5 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_A6 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_B1 = CLBLM_L_X10Y112_SLICE_X13Y112_BO6;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_B2 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_B3 = CLBLM_L_X10Y114_SLICE_X12Y114_CO6;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_B4 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_B5 = CLBLM_R_X11Y114_SLICE_X14Y114_BO6;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_B6 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_A1 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_A2 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_A3 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_C1 = CLBLM_R_X11Y114_SLICE_X14Y114_BO6;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_C2 = CLBLM_L_X8Y116_SLICE_X10Y116_AO6;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_C3 = CLBLM_L_X10Y114_SLICE_X12Y114_CO6;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_C4 = CLBLM_L_X8Y116_SLICE_X10Y116_AO5;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_C5 = CLBLM_L_X10Y112_SLICE_X13Y112_BO6;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_C6 = CLBLM_R_X7Y114_SLICE_X9Y114_AO6;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_A4 = CLBLL_L_X2Y108_SLICE_X0Y108_BO6;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_A5 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_A6 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_B1 = CLBLL_L_X2Y109_SLICE_X0Y109_DO6;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_B6 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_B2 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_B3 = CLBLL_L_X2Y110_SLICE_X0Y110_AO6;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_B4 = CLBLL_L_X2Y109_SLICE_X0Y109_CO6;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_B5 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_D1 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_D2 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_D3 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_D4 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_D5 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_D6 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_C1 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_C2 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_C3 = CLBLL_L_X2Y108_SLICE_X1Y108_DO6;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_C4 = CLBLL_L_X2Y107_SLICE_X0Y107_CO6;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_C5 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_C6 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_D1 = CLBLL_L_X2Y110_SLICE_X0Y110_AO6;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_D2 = CLBLL_L_X2Y109_SLICE_X0Y109_BO6;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_D3 = CLBLL_L_X2Y108_SLICE_X0Y108_AO6;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_D4 = CLBLL_L_X2Y107_SLICE_X0Y107_AO5;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_D5 = CLBLL_L_X2Y109_SLICE_X0Y109_DO6;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_D6 = CLBLL_L_X2Y109_SLICE_X0Y109_CO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C1 = CLBLL_L_X4Y112_SLICE_X4Y112_BO6;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_A1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_A2 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_A3 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_A4 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_A5 = CLBLL_L_X2Y108_SLICE_X1Y108_CO6;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_A6 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_B1 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_B2 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_A3 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_A4 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_A5 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_A6 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_B3 = CLBLL_L_X2Y107_SLICE_X0Y107_BO6;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_B4 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_B5 = CLBLL_L_X2Y110_SLICE_X0Y110_AO6;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_B6 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_A2 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C6 = CLBLM_R_X3Y112_SLICE_X2Y112_AO6;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_C1 = CLBLL_L_X2Y109_SLICE_X0Y109_AO6;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_C2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_C3 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_C4 = CLBLL_L_X2Y107_SLICE_X1Y107_BO6;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_C5 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_C6 = CLBLL_L_X2Y108_SLICE_X1Y108_BO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_B1 = CLBLM_L_X8Y110_SLICE_X10Y110_CO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_C1 = CLBLM_R_X7Y110_SLICE_X9Y110_AO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_C2 = CLBLM_R_X7Y109_SLICE_X9Y109_AO5;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_B4 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_B5 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_C5 = CLBLM_L_X10Y111_SLICE_X12Y111_CO6;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_D1 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_D2 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_D3 = CLBLL_L_X2Y108_SLICE_X0Y108_DO6;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_D4 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_D5 = CLBLL_L_X2Y107_SLICE_X1Y107_BO6;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_D6 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_C6 = CLBLM_R_X5Y110_SLICE_X7Y110_BO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_D1 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_D2 = CLBLM_L_X8Y109_SLICE_X10Y109_CO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_D3 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_D4 = CLBLM_L_X8Y110_SLICE_X10Y110_DO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_D5 = CLBLM_R_X7Y108_SLICE_X9Y108_DO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_D6 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_A1 = CLBLM_R_X5Y109_SLICE_X6Y109_DO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_A2 = CLBLM_L_X8Y110_SLICE_X11Y110_AO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_A3 = CLBLM_R_X7Y109_SLICE_X8Y109_CO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_A4 = CLBLM_R_X7Y110_SLICE_X9Y110_AO5;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_A5 = CLBLM_R_X5Y110_SLICE_X7Y110_BO5;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_A6 = CLBLM_R_X7Y109_SLICE_X8Y109_DO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_B1 = CLBLM_R_X7Y108_SLICE_X9Y108_DO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_B2 = CLBLM_L_X8Y110_SLICE_X11Y110_AO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_B3 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_B4 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_B5 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_B6 = CLBLM_L_X8Y109_SLICE_X10Y109_CO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_C1 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_C2 = CLBLM_R_X7Y108_SLICE_X9Y108_DO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_C3 = CLBLM_L_X8Y110_SLICE_X11Y110_AO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_C4 = CLBLM_L_X8Y109_SLICE_X10Y109_CO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_C5 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_C6 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_D1 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_D2 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_D3 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_D4 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_D5 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_D6 = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_D1 = CLBLL_L_X2Y107_SLICE_X1Y107_AO5;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_T1 = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_D1 = CLBLL_L_X2Y108_SLICE_X0Y108_CO6;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_A1 = CLBLL_L_X2Y109_SLICE_X0Y109_DO6;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_A2 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_A3 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_A4 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_A5 = CLBLL_L_X2Y109_SLICE_X0Y109_CO6;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_A6 = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_T1 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_B1 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_B2 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_B3 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_B4 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_B5 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_B6 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_C1 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_C2 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_C3 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_C4 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_C5 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_C6 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_D1 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_D2 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_D3 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_D4 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_D5 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_D6 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_A1 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_A2 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_A3 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_A4 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_A5 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_A6 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_B1 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_B2 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_B3 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_B4 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_B5 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_B6 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_A1 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_A2 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_A3 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_C1 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_C2 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_C3 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_C4 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_C5 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_C6 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_A4 = CLBLM_L_X10Y111_SLICE_X13Y111_BO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_A5 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_A6 = CLBLM_L_X8Y111_SLICE_X10Y111_BO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_B5 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_B6 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_B1 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_B2 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_B3 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_B4 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_D1 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_D2 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_D3 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_D4 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_D5 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_D6 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_C1 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_C2 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_C3 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_C4 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_C5 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_D1 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_D2 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_D3 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_D4 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_D5 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_D6 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_A1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_A2 = CLBLM_L_X8Y111_SLICE_X10Y111_DO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_A3 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_A4 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_A5 = CLBLM_R_X7Y110_SLICE_X9Y110_BO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_A6 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_B1 = CLBLM_R_X7Y112_SLICE_X9Y112_BO5;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_B2 = CLBLM_R_X5Y110_SLICE_X7Y110_AO5;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_B3 = CLBLM_L_X10Y111_SLICE_X13Y111_BO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_B4 = CLBLM_L_X8Y111_SLICE_X10Y111_BO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_B5 = CLBLM_R_X7Y111_SLICE_X8Y111_AO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_B6 = CLBLM_R_X7Y110_SLICE_X9Y110_CO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_C1 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_C2 = CLBLM_R_X7Y110_SLICE_X9Y110_CO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_C3 = CLBLM_L_X10Y111_SLICE_X13Y111_BO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_C4 = CLBLM_L_X8Y111_SLICE_X10Y111_BO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_C5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_C6 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_D1 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_D2 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_D3 = CLBLM_L_X10Y111_SLICE_X13Y111_BO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_D4 = CLBLM_R_X7Y111_SLICE_X8Y111_AO5;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_D5 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_D6 = CLBLM_L_X8Y111_SLICE_X10Y111_BO6;
  assign RIOI3_X105Y105_ILOGIC_X1Y106_D = RIOB33_X105Y105_IOB_X1Y106_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y105_D = RIOB33_X105Y105_IOB_X1Y105_I;
  assign LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y108_D = LIOB33_X0Y107_IOB_X0Y108_I;
  assign LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y107_D = LIOB33_X0Y107_IOB_X0Y107_I;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_D = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_A1 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_A2 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_A3 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_A4 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_A5 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_A6 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_B1 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_B2 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_B3 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_B4 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_B5 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_B6 = 1'b1;
  assign RIOI3_SING_X105Y100_ILOGIC_X1Y100_D = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_C1 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_C2 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_C3 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_C4 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_C5 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_C6 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_D1 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_D2 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_D3 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_D4 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_D5 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_D6 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_A1 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_A2 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_A3 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_A4 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_A5 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_A6 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_B1 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_B2 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_B3 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_B4 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_B5 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_B6 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_C1 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_C2 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_C3 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_C4 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_C5 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_C6 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_A1 = CLBLM_L_X10Y112_SLICE_X12Y112_AO5;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_A2 = CLBLM_L_X10Y112_SLICE_X12Y112_DO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_A3 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_B1 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_B2 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_A4 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_A5 = CLBLM_L_X10Y112_SLICE_X12Y112_AO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_B5 = CLBLM_R_X7Y111_SLICE_X9Y111_AO6;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_D1 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_D2 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_D3 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_D4 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_D5 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_D6 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_B4 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_B6 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_C1 = CLBLM_L_X8Y112_SLICE_X10Y112_BO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_C2 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_C3 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_C4 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_C5 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_C6 = CLBLM_R_X7Y110_SLICE_X8Y110_BO6;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_B6 = CLBLM_L_X8Y114_SLICE_X11Y114_DO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_D1 = CLBLM_R_X7Y111_SLICE_X9Y111_AO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_D2 = CLBLM_L_X10Y112_SLICE_X12Y112_AO5;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_D3 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_D4 = CLBLM_L_X10Y112_SLICE_X12Y112_DO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_D5 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_D6 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_A1 = CLBLM_L_X8Y113_SLICE_X10Y113_AO5;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_A2 = CLBLM_R_X7Y110_SLICE_X8Y110_BO6;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_A3 = CLBLM_R_X5Y111_SLICE_X6Y111_AO5;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_A4 = CLBLM_L_X8Y113_SLICE_X10Y113_BO6;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_A5 = CLBLM_R_X5Y112_SLICE_X7Y112_AO6;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_A6 = CLBLM_L_X8Y112_SLICE_X10Y112_CO6;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_B1 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_B2 = CLBLM_R_X7Y110_SLICE_X8Y110_BO6;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_B3 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_B4 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_B5 = CLBLM_L_X8Y112_SLICE_X10Y112_BO6;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_B6 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_C3 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_C1 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_C2 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_C3 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_C4 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_C5 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_C6 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_C4 = CLBLM_R_X7Y112_SLICE_X9Y112_AO5;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_C5 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_C6 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_D1 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_D2 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_D3 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_D4 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_D5 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_D6 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_D5 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_D6 = CLBLM_R_X7Y112_SLICE_X9Y112_AO5;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_A1 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_A2 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_A3 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_A4 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_A5 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_A6 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_B1 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_B2 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_B3 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_B4 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_B5 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_B6 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_C1 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_C2 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_C3 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_C4 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_C5 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_C6 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_C3 = CLBLM_R_X7Y116_SLICE_X8Y116_CO6;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_D1 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_D2 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_D3 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_D4 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_D5 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_D6 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_A1 = CLBLL_L_X4Y111_SLICE_X4Y111_DO6;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_A2 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_A3 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_A4 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_A5 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_A6 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_B1 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_B2 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_B3 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_B4 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_B5 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_B6 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_C1 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_C2 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_C3 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_C4 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_C5 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_C6 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_A1 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_A2 = CLBLM_L_X10Y113_SLICE_X12Y113_BO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_A3 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_A4 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_A5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_A6 = CLBLM_L_X8Y113_SLICE_X10Y113_DO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_C4 = CLBLM_L_X8Y113_SLICE_X11Y113_BO6;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_D1 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_D2 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_D3 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_D4 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_D5 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_D6 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_B1 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_B2 = CLBLM_R_X7Y113_SLICE_X9Y113_AO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_B3 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_B4 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_B5 = CLBLM_R_X7Y112_SLICE_X9Y112_CO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_B6 = CLBLM_L_X8Y113_SLICE_X10Y113_CO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_C1 = CLBLM_R_X7Y113_SLICE_X9Y113_AO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_C2 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_C3 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_C4 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_C5 = CLBLM_R_X7Y113_SLICE_X9Y113_DO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_C6 = CLBLM_R_X7Y112_SLICE_X9Y112_CO6;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_D1 = CLBLM_R_X3Y107_SLICE_X2Y107_AO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_D1 = CLBLM_L_X8Y113_SLICE_X10Y113_AO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_D2 = CLBLM_L_X10Y112_SLICE_X12Y112_BO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_D3 = CLBLM_R_X5Y115_SLICE_X6Y115_AO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_D4 = CLBLM_L_X8Y113_SLICE_X10Y113_DO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_D5 = CLBLM_L_X8Y113_SLICE_X10Y113_AO5;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_D6 = CLBLM_L_X8Y114_SLICE_X11Y114_BO6;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_D2 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_D3 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_T1 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_A1 = CLBLM_L_X8Y113_SLICE_X10Y113_AO5;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_A2 = CLBLM_L_X8Y113_SLICE_X10Y113_DO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_A3 = CLBLM_R_X5Y111_SLICE_X6Y111_AO5;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_A4 = CLBLM_L_X8Y114_SLICE_X11Y114_BO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_A5 = CLBLM_R_X7Y110_SLICE_X8Y110_BO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_A6 = CLBLM_L_X8Y113_SLICE_X10Y113_BO6;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_D1 = CLBLL_L_X2Y109_SLICE_X0Y109_AO5;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_B1 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_B2 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_B3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_B4 = CLBLM_L_X10Y113_SLICE_X12Y113_BO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_B5 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_B6 = CLBLM_L_X8Y113_SLICE_X10Y113_DO6;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_T1 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_C1 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_C2 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_C3 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_C4 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_C5 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_C6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_D1 = CLBLL_L_X2Y112_SLICE_X0Y112_AO6;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_T1 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_D1 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_D2 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_D3 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_D4 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_D5 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_D6 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_C1 = CLBLM_R_X7Y116_SLICE_X9Y116_CO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_C2 = CLBLM_R_X7Y113_SLICE_X9Y113_CO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_C3 = CLBLM_R_X7Y116_SLICE_X8Y116_AO6;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_A1 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_A2 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_A3 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_A4 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_A5 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_A6 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_B1 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_B2 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_B3 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_B4 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_B5 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_B6 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_C1 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_C2 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_C3 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_C4 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_C5 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_C6 = 1'b1;
  assign RIOI3_X105Y109_ILOGIC_X1Y110_D = RIOB33_X105Y109_IOB_X1Y110_I;
  assign RIOI3_X105Y109_ILOGIC_X1Y109_D = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_D1 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_D2 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_D3 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_D4 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_D5 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_D6 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_D4 = CLBLM_R_X5Y115_SLICE_X6Y115_DO6;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_A1 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_A2 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_A3 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_A4 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_A5 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_A6 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_B1 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_B2 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_B3 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_B4 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_B5 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_B6 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_C1 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_C2 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_C3 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_C4 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_C5 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_C6 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_A1 = CLBLM_L_X8Y114_SLICE_X11Y114_DO6;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_A2 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_A3 = CLBLM_L_X8Y113_SLICE_X11Y113_AO6;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_A4 = CLBLM_L_X8Y114_SLICE_X10Y114_AO6;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_D1 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_D2 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_D3 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_D4 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_D5 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_D6 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_A5 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_A6 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_B1 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_B2 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_B3 = CLBLM_L_X8Y113_SLICE_X11Y113_AO6;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_B4 = CLBLM_L_X8Y114_SLICE_X10Y114_AO6;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_B5 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_A1 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_A2 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_A3 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_A4 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_A5 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_A6 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_C1 = CLBLM_R_X7Y112_SLICE_X9Y112_BO6;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_C2 = CLBLM_R_X7Y114_SLICE_X8Y114_AO5;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_B1 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_B2 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_B3 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_B4 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_B5 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_B6 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_D1 = CLBLM_R_X7Y112_SLICE_X9Y112_BO6;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_D2 = CLBLM_R_X7Y114_SLICE_X8Y114_AO5;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_C1 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_C2 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_C3 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_C4 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_C5 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_C6 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_D3 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_D4 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_A1 = CLBLM_R_X7Y112_SLICE_X9Y112_DO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_A2 = CLBLM_R_X7Y111_SLICE_X8Y111_CO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_A3 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_A4 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_A5 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_A6 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_D1 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_D2 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_D3 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_D4 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_D5 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_D6 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_B1 = CLBLM_R_X7Y112_SLICE_X9Y112_DO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_B6 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_B2 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_B3 = CLBLM_L_X8Y113_SLICE_X11Y113_BO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_B4 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_B5 = CLBLM_R_X7Y112_SLICE_X9Y112_AO6;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_A1 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_A2 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_A3 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_C3 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_A4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_A5 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_A6 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_C1 = CLBLM_R_X7Y114_SLICE_X8Y114_AO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_C2 = CLBLM_R_X7Y112_SLICE_X9Y112_AO6;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_B1 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_B2 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_B3 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_B4 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_B5 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_B6 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_D1 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_D2 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_D3 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_C1 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_C2 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_C3 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_C4 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_C5 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_C6 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_D4 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_D5 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_D6 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_D1 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_D2 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_D3 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_D4 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_D5 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_D6 = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_D1 = CLBLM_R_X3Y108_SLICE_X3Y108_AO6;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_A1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_A2 = CLBLM_L_X10Y114_SLICE_X12Y114_DO6;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_A3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_A4 = CLBLM_L_X8Y114_SLICE_X11Y114_AO6;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_A5 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_A6 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_B1 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_B2 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_B3 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_B4 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_B5 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_B6 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_A1 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_A2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_A3 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_A4 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_A5 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_A6 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_C1 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_C2 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_C3 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_B1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_B2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_B3 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_B4 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_B5 = CLBLM_R_X5Y105_SLICE_X7Y105_CO6;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_B6 = CLBLL_L_X4Y105_SLICE_X4Y105_DO6;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_D1 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_D2 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_C1 = CLBLM_R_X5Y105_SLICE_X7Y105_AO6;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_C2 = CLBLM_R_X7Y106_SLICE_X8Y106_CO6;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_C3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_C4 = CLBLM_R_X7Y104_SLICE_X8Y104_AO6;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_C5 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_C6 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_D3 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_D4 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_A1 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_A2 = CLBLM_L_X8Y115_SLICE_X10Y115_BO6;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_A3 = CLBLM_R_X7Y115_SLICE_X9Y115_AO6;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_A4 = CLBLM_R_X7Y113_SLICE_X8Y113_BO6;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_A5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_A6 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_D1 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_D2 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_D3 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_D4 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_D5 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_D6 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_B1 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_B2 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_B3 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_B4 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_B5 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_A1 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_A2 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_A3 = CLBLM_R_X5Y105_SLICE_X7Y105_CO6;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_A4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_A5 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_A6 = CLBLL_L_X4Y105_SLICE_X4Y105_DO6;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_C1 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_C2 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_C3 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_B1 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_B2 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_B3 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_B4 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_B5 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_B6 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_D1 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_D2 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_D3 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_C1 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_C2 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_C3 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_C4 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_C5 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_C6 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_D4 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_D5 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_D6 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_D1 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_D2 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_D3 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_D4 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_D5 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_D6 = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_D1 = CLBLM_R_X3Y110_SLICE_X3Y110_AO6;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_T1 = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_D1 = CLBLL_L_X4Y109_SLICE_X4Y109_AO6;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_D1 = CLBLM_R_X3Y114_SLICE_X3Y114_AO5;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_D1 = CLBLL_L_X4Y111_SLICE_X4Y111_AO6;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_T1 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_A1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_A2 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_A3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_A4 = CLBLM_L_X8Y116_SLICE_X10Y116_BO6;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_A5 = CLBLM_L_X8Y114_SLICE_X11Y114_CO6;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_A6 = CLBLM_L_X8Y115_SLICE_X10Y115_CO6;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_B1 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_B2 = CLBLM_L_X8Y115_SLICE_X10Y115_AO5;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_B3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_B4 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_B5 = CLBLM_L_X8Y116_SLICE_X10Y116_BO6;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_B6 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_A1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_A2 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_A3 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_A4 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_A5 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_A6 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_C1 = CLBLM_L_X8Y114_SLICE_X11Y114_CO6;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_C2 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_C3 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_B1 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_B2 = CLBLM_R_X7Y105_SLICE_X8Y105_CO6;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_B3 = CLBLM_R_X5Y105_SLICE_X7Y105_BO6;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_B4 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_B5 = CLBLL_L_X4Y106_SLICE_X5Y106_CO6;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_B6 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_D1 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_D3 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_C1 = CLBLM_R_X5Y105_SLICE_X7Y105_BO6;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_C2 = CLBLM_R_X7Y105_SLICE_X8Y105_CO6;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_C3 = CLBLM_R_X5Y106_SLICE_X6Y106_BO5;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_C4 = CLBLM_R_X5Y106_SLICE_X7Y106_AO5;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_C5 = CLBLL_L_X4Y106_SLICE_X5Y106_CO6;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_C6 = CLBLM_R_X7Y108_SLICE_X9Y108_AO5;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_D4 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_D5 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_A1 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_A2 = CLBLM_R_X7Y113_SLICE_X8Y113_BO6;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_A3 = CLBLM_L_X8Y115_SLICE_X10Y115_DO6;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_A4 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_A5 = CLBLM_R_X7Y115_SLICE_X9Y115_AO6;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_A6 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_D1 = CLBLM_R_X5Y105_SLICE_X7Y105_BO6;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_D2 = CLBLM_R_X7Y105_SLICE_X8Y105_CO6;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_D3 = CLBLM_R_X5Y106_SLICE_X6Y106_BO5;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_D4 = CLBLM_R_X5Y106_SLICE_X7Y106_AO5;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_D5 = CLBLL_L_X4Y106_SLICE_X5Y106_CO6;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_D6 = CLBLM_R_X7Y108_SLICE_X9Y108_AO5;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_B1 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_B2 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_B3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_B4 = CLBLM_R_X7Y114_SLICE_X9Y114_AO5;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_B5 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_A1 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_A2 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_A3 = CLBLM_R_X5Y104_SLICE_X6Y104_AO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_A4 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_A5 = CLBLM_R_X5Y106_SLICE_X6Y106_CO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_A6 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_C1 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_C2 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_C3 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_B1 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_B2 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_B3 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_B4 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_B5 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_B6 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_D1 = CLBLM_L_X8Y115_SLICE_X10Y115_DO6;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_D2 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_D3 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_C1 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_C2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_C3 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_C4 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_C5 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_C6 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_D4 = CLBLM_R_X7Y115_SLICE_X9Y115_AO6;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_D5 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_D6 = CLBLM_R_X7Y113_SLICE_X8Y113_BO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_D1 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_D2 = CLBLM_R_X5Y105_SLICE_X7Y105_CO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_D3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_D4 = CLBLM_R_X5Y106_SLICE_X6Y106_AO5;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_D5 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_D6 = CLBLM_R_X7Y106_SLICE_X8Y106_BO6;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_A4 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign LIOB33_X0Y117_IOB_X0Y118_O = CLBLL_L_X2Y112_SLICE_X0Y112_AO5;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_A5 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_A6 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_A1 = CLBLM_R_X5Y106_SLICE_X7Y106_DO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_A2 = CLBLM_R_X7Y108_SLICE_X8Y108_AO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_A3 = CLBLM_R_X3Y107_SLICE_X2Y107_AO5;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_A4 = CLBLM_R_X7Y107_SLICE_X9Y107_AO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_A5 = CLBLL_L_X4Y106_SLICE_X5Y106_DO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_A6 = CLBLM_R_X5Y106_SLICE_X7Y106_CO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_B1 = CLBLM_R_X7Y107_SLICE_X9Y107_CO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_B2 = CLBLM_R_X5Y106_SLICE_X7Y106_DO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_B3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_B4 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_B5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_B6 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_C1 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_C2 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_C3 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_C4 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_C5 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_C6 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_D1 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_D2 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_D3 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_D4 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_D5 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_D6 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_A1 = CLBLL_L_X4Y106_SLICE_X5Y106_CO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_A2 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_A3 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_A4 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_A5 = CLBLM_R_X5Y106_SLICE_X6Y106_DO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_A6 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_B1 = CLBLM_R_X5Y107_SLICE_X6Y107_DO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_B2 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_B3 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_B4 = CLBLM_R_X7Y107_SLICE_X9Y107_CO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_B5 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_B6 = CLBLM_R_X5Y107_SLICE_X6Y107_CO6;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_C4 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_C5 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_C1 = CLBLM_R_X5Y105_SLICE_X6Y105_AO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_C2 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_C3 = CLBLM_R_X7Y106_SLICE_X9Y106_DO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_C4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_C5 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_C6 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_C6 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_D1 = CLBLM_R_X5Y106_SLICE_X6Y106_DO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_D2 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_D3 = CLBLL_L_X4Y106_SLICE_X5Y106_CO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_D4 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_D5 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_D6 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_D5 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_D6 = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_D1 = CLBLL_L_X2Y109_SLICE_X0Y109_BO5;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_T1 = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_D1 = CLBLM_R_X3Y110_SLICE_X3Y110_BO6;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_D1 = CLBLL_L_X4Y116_SLICE_X4Y116_CO6;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_B6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_D1 = CLBLL_L_X4Y115_SLICE_X4Y115_DO6;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_T1 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_C4 = 1'b1;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_A1 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_A2 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_A3 = CLBLM_R_X5Y109_SLICE_X7Y109_AO6;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_A4 = CLBLL_L_X4Y108_SLICE_X5Y108_CO6;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_A5 = CLBLM_L_X8Y106_SLICE_X10Y106_CO6;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_A6 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_C5 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_C6 = 1'b1;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_B1 = CLBLM_R_X5Y108_SLICE_X7Y108_DO6;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_B2 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_B3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_B4 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_B5 = CLBLM_L_X8Y106_SLICE_X10Y106_CO6;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_B6 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_C1 = CLBLM_R_X5Y109_SLICE_X7Y109_AO6;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_C2 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_C3 = CLBLL_L_X4Y108_SLICE_X5Y108_CO6;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_C4 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_C5 = CLBLM_L_X8Y106_SLICE_X10Y106_CO6;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_C6 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_D2 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_D1 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_D2 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_D3 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_D4 = CLBLM_L_X8Y105_SLICE_X10Y105_DO6;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_D5 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_D6 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_D4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_A1 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_A2 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_A3 = CLBLL_L_X4Y106_SLICE_X5Y106_DO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_A4 = CLBLM_R_X5Y106_SLICE_X7Y106_BO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_A5 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_A6 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_B1 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_B2 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_B3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_B4 = CLBLM_R_X5Y108_SLICE_X6Y108_AO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_B5 = CLBLM_R_X5Y107_SLICE_X6Y107_BO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_B6 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_C1 = CLBLM_R_X5Y107_SLICE_X6Y107_BO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_C2 = CLBLM_R_X5Y108_SLICE_X6Y108_AO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_C3 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_C4 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_C5 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_C6 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign RIOI3_X105Y111_ILOGIC_X1Y112_D = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_D1 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_D2 = CLBLM_L_X8Y105_SLICE_X10Y105_DO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_D3 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_D4 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_D5 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_D6 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_A1 = CLBLM_R_X5Y108_SLICE_X7Y108_DO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_A2 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_A3 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_A4 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_A5 = CLBLM_R_X5Y110_SLICE_X6Y110_CO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_A6 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_B1 = CLBLM_R_X7Y109_SLICE_X9Y109_CO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_B2 = CLBLM_R_X7Y109_SLICE_X8Y109_BO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_B3 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_B4 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_B5 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_B6 = CLBLM_R_X5Y108_SLICE_X6Y108_CO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_C1 = CLBLM_R_X5Y108_SLICE_X7Y108_CO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_C2 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_C3 = CLBLM_L_X8Y109_SLICE_X10Y109_AO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_C4 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_C5 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_C6 = CLBLM_R_X5Y108_SLICE_X7Y108_BO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_D1 = CLBLM_R_X5Y108_SLICE_X7Y108_CO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_D2 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_D3 = CLBLM_L_X8Y109_SLICE_X10Y109_AO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_D4 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_D5 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_D6 = CLBLM_R_X5Y108_SLICE_X7Y108_BO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_A1 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_A2 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_A3 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_A4 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_A5 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_A6 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_B1 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_B2 = CLBLM_R_X5Y107_SLICE_X7Y107_BO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_B3 = CLBLM_R_X7Y108_SLICE_X8Y108_BO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_B4 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_B5 = CLBLM_R_X5Y108_SLICE_X6Y108_AO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_B6 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_C1 = CLBLM_R_X5Y109_SLICE_X6Y109_AO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_C2 = CLBLM_R_X7Y109_SLICE_X8Y109_AO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_C3 = CLBLM_R_X7Y108_SLICE_X8Y108_BO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_C4 = CLBLL_L_X4Y110_SLICE_X4Y110_AO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_C5 = CLBLM_R_X5Y108_SLICE_X6Y108_AO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_C6 = CLBLM_R_X5Y107_SLICE_X7Y107_BO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_D1 = CLBLM_R_X5Y109_SLICE_X6Y109_AO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_D2 = CLBLL_L_X4Y110_SLICE_X4Y110_AO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_D3 = CLBLM_R_X7Y108_SLICE_X8Y108_BO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_D4 = CLBLM_R_X7Y109_SLICE_X8Y109_AO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_D5 = CLBLM_R_X5Y108_SLICE_X6Y108_AO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_D6 = CLBLM_R_X5Y107_SLICE_X7Y107_BO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_A1 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_A2 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_A3 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_A4 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_A5 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_A6 = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_D1 = 1'b0;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_B1 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_B2 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_B3 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_B4 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_B5 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_B6 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_C1 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_C2 = CLBLM_R_X7Y109_SLICE_X9Y109_CO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_C3 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_C4 = CLBLM_R_X5Y108_SLICE_X6Y108_CO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_C5 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_C6 = CLBLM_R_X7Y109_SLICE_X8Y109_DO6;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_T1 = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_D1 = CLBLL_L_X4Y112_SLICE_X4Y112_AO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_D1 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_D2 = CLBLM_R_X7Y109_SLICE_X9Y109_CO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_D3 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_D4 = CLBLM_R_X5Y108_SLICE_X6Y108_CO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_D5 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_D6 = CLBLM_R_X7Y109_SLICE_X8Y109_DO6;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_T1 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_A1 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_A2 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_A3 = CLBLM_R_X5Y108_SLICE_X7Y108_AO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_A4 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_A5 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_A6 = CLBLM_R_X5Y110_SLICE_X6Y110_CO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_B1 = CLBLM_R_X5Y109_SLICE_X6Y109_DO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_B2 = CLBLM_R_X5Y110_SLICE_X7Y110_BO5;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_B3 = CLBLM_R_X5Y109_SLICE_X6Y109_CO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_B4 = CLBLM_R_X7Y109_SLICE_X8Y109_DO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_B5 = CLBLL_L_X4Y109_SLICE_X4Y109_DO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_B6 = CLBLM_R_X3Y110_SLICE_X3Y110_AO5;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_C1 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_C2 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_C3 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_C4 = CLBLM_R_X5Y108_SLICE_X6Y108_DO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_C5 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_C6 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_D1 = CLBLM_R_X3Y111_SLICE_X2Y111_AO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_D2 = CLBLM_R_X5Y110_SLICE_X7Y110_CO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_D3 = CLBLM_R_X5Y110_SLICE_X7Y110_AO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_D4 = CLBLM_R_X5Y111_SLICE_X6Y111_AO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_D5 = CLBLL_L_X4Y109_SLICE_X5Y109_BO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_D6 = CLBLM_R_X7Y110_SLICE_X8Y110_AO6;
  assign LIOB33_X0Y119_IOB_X0Y120_O = CLBLL_L_X2Y109_SLICE_X0Y109_AO5;
  assign LIOB33_X0Y119_IOB_X0Y119_O = CLBLL_L_X2Y112_SLICE_X0Y112_AO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_A1 = CLBLM_R_X5Y111_SLICE_X6Y111_AO5;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_A2 = CLBLM_R_X5Y110_SLICE_X7Y110_DO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_A3 = CLBLM_R_X5Y111_SLICE_X6Y111_AO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_A4 = CLBLM_R_X7Y110_SLICE_X8Y110_BO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_A5 = CLBLM_R_X7Y110_SLICE_X8Y110_CO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_A6 = CLBLM_L_X8Y113_SLICE_X10Y113_BO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_B1 = CLBLM_R_X5Y111_SLICE_X6Y111_AO5;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_B2 = CLBLM_R_X5Y110_SLICE_X7Y110_DO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_B3 = CLBLM_R_X5Y111_SLICE_X6Y111_AO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_B4 = CLBLM_R_X5Y112_SLICE_X7Y112_AO5;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_B5 = CLBLM_R_X7Y110_SLICE_X8Y110_CO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_B6 = CLBLM_L_X8Y111_SLICE_X10Y111_CO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_C1 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_C2 = CLBLM_R_X7Y110_SLICE_X9Y110_BO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_C3 = CLBLM_L_X8Y111_SLICE_X10Y111_DO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_C4 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_C5 = CLBLL_L_X4Y110_SLICE_X4Y110_BO5;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_C6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_D1 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_D2 = CLBLM_R_X7Y110_SLICE_X9Y110_BO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_D3 = CLBLM_L_X8Y111_SLICE_X10Y111_DO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_D4 = CLBLL_L_X4Y110_SLICE_X4Y110_BO5;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_D5 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_D6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_A1 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_A2 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_A3 = 1'b1;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_A4 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_A5 = 1'b1;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_A6 = 1'b1;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_B1 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_B2 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_B3 = CLBLM_R_X5Y111_SLICE_X7Y111_AO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_B4 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_B5 = CLBLL_L_X4Y111_SLICE_X5Y111_BO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_B6 = CLBLM_R_X5Y111_SLICE_X6Y111_CO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_C1 = CLBLL_L_X4Y109_SLICE_X5Y109_BO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_C2 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_C3 = CLBLM_R_X5Y109_SLICE_X7Y109_BO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_C4 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_C5 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_C6 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_D1 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_D2 = CLBLL_L_X4Y111_SLICE_X5Y111_BO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_D3 = CLBLM_R_X5Y111_SLICE_X7Y111_BO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_D4 = CLBLM_R_X5Y111_SLICE_X6Y111_CO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_D5 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_D6 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_C4 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_C5 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_C6 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_D5 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_D6 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_A1 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_A2 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_A3 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_A4 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_A5 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_A6 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_B1 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_B2 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_B3 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_B4 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_B5 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_B6 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_C1 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_C2 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_C3 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_C4 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_C5 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_C6 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_D1 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_D2 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_D3 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_D4 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_D5 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_D6 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_A1 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_A2 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_A3 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_A4 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_A5 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_A6 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_B1 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_B2 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_B3 = CLBLM_R_X7Y112_SLICE_X8Y112_AO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_B4 = CLBLM_R_X7Y112_SLICE_X8Y112_BO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_B5 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_B6 = CLBLL_L_X4Y111_SLICE_X5Y111_CO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_C1 = CLBLM_R_X5Y112_SLICE_X6Y112_AO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_C2 = CLBLL_L_X4Y113_SLICE_X5Y113_AO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_C3 = CLBLM_R_X3Y111_SLICE_X3Y111_CO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_C4 = CLBLM_R_X5Y111_SLICE_X6Y111_DO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_C5 = CLBLM_R_X5Y112_SLICE_X6Y112_DO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_C6 = CLBLM_R_X5Y112_SLICE_X6Y112_BO6;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_C4 = CLBLM_L_X8Y115_SLICE_X10Y115_CO6;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_C5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_C6 = CLBLM_L_X8Y116_SLICE_X10Y116_CO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_D1 = CLBLL_L_X4Y111_SLICE_X5Y111_BO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_D2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_D3 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_D4 = CLBLM_R_X5Y111_SLICE_X6Y111_CO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_D5 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_D6 = CLBLM_R_X5Y111_SLICE_X7Y111_BO6;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_B6 = CLBLM_R_X11Y114_SLICE_X14Y114_CO6;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_D1 = CLBLM_R_X5Y114_SLICE_X6Y114_AO6;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_T1 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_D2 = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_D1 = CLBLM_R_X5Y114_SLICE_X6Y114_AO5;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_C4 = CLBLM_R_X11Y110_SLICE_X15Y110_CO6;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_C5 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_D6 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_C6 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_T1 = 1'b1;
  assign LIOI3_X0Y115_ILOGIC_X0Y116_D = LIOB33_X0Y115_IOB_X0Y116_I;
  assign LIOI3_X0Y115_ILOGIC_X0Y115_D = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_B6 = CLBLM_R_X7Y116_SLICE_X9Y116_BO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_C4 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_C6 = CLBLM_L_X8Y109_SLICE_X11Y109_BO6;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_A1 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_A2 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_A3 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_A4 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_A5 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_A6 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_C4 = CLBLM_R_X7Y116_SLICE_X9Y116_BO6;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_B1 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_B2 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_B3 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_B4 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_B5 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_B6 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_C5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_C6 = CLBLM_R_X7Y114_SLICE_X9Y114_AO5;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_C1 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_C2 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_C3 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_C4 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_C5 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_C6 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_D1 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_D2 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_D3 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_D4 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_D5 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_D6 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_A1 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_A2 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_A3 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_A4 = CLBLM_R_X5Y111_SLICE_X6Y111_DO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_A5 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_A6 = CLBLM_R_X5Y113_SLICE_X6Y113_CO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_B1 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_B2 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_B3 = CLBLM_R_X7Y112_SLICE_X8Y112_BO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_B4 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_B5 = CLBLM_R_X7Y112_SLICE_X8Y112_AO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_B6 = CLBLL_L_X4Y111_SLICE_X5Y111_CO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_C1 = CLBLM_R_X7Y112_SLICE_X8Y112_BO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_C2 = CLBLL_L_X4Y111_SLICE_X5Y111_CO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_C3 = CLBLM_R_X7Y113_SLICE_X8Y113_AO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_C4 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_C5 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_C6 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_D1 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_D2 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_D3 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_D4 = CLBLM_R_X7Y113_SLICE_X9Y113_BO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_D5 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_D6 = CLBLM_R_X5Y113_SLICE_X6Y113_BO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_D1 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_A1 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_A2 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_A3 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_A4 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_A5 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_A6 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_B1 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_B2 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_B3 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_B4 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_B5 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_B6 = 1'b1;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_A1 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_A2 = 1'b1;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_A3 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_A4 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_A5 = 1'b1;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_A6 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_C1 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_C2 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_C3 = 1'b1;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_B1 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_B2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_B3 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_B4 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_B5 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_B6 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_D1 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_D2 = 1'b1;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_C1 = CLBLM_R_X3Y104_SLICE_X3Y104_AO6;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_C2 = CLBLM_R_X3Y105_SLICE_X2Y105_AO6;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_C3 = CLBLM_R_X5Y104_SLICE_X6Y104_AO6;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_C4 = CLBLM_R_X3Y104_SLICE_X3Y104_AO5;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_C5 = CLBLL_L_X4Y105_SLICE_X4Y105_AO6;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_C6 = CLBLM_R_X3Y104_SLICE_X3Y104_BO6;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_D3 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_D4 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_A1 = CLBLM_R_X5Y113_SLICE_X6Y113_DO6;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_A2 = CLBLM_R_X5Y115_SLICE_X6Y115_BO6;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_A3 = CLBLM_R_X5Y112_SLICE_X6Y112_CO6;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_A4 = CLBLM_R_X5Y114_SLICE_X6Y114_BO6;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_A5 = CLBLM_R_X5Y113_SLICE_X6Y113_AO6;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_A6 = 1'b1;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_D1 = CLBLM_R_X3Y104_SLICE_X3Y104_AO6;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_D2 = CLBLM_R_X3Y105_SLICE_X2Y105_AO6;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_D3 = CLBLM_R_X5Y104_SLICE_X6Y104_AO6;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_D4 = CLBLM_R_X3Y104_SLICE_X3Y104_AO5;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_D5 = CLBLL_L_X4Y105_SLICE_X4Y105_AO6;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_D6 = CLBLM_R_X3Y104_SLICE_X3Y104_BO6;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_B1 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_B2 = CLBLM_R_X5Y113_SLICE_X6Y113_BO6;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_B3 = CLBLM_R_X7Y113_SLICE_X9Y113_BO6;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_B4 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_B5 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_A1 = 1'b1;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_A2 = 1'b1;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_A3 = 1'b1;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_A4 = 1'b1;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_A5 = 1'b1;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_A6 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_C1 = CLBLM_R_X5Y113_SLICE_X6Y113_AO6;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_C2 = CLBLM_R_X5Y112_SLICE_X6Y112_CO6;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_C3 = CLBLM_R_X5Y115_SLICE_X6Y115_BO6;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_B1 = 1'b1;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_B2 = 1'b1;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_B3 = 1'b1;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_B4 = 1'b1;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_B5 = 1'b1;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_B6 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_D1 = CLBLM_R_X5Y113_SLICE_X6Y113_AO6;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_D2 = CLBLM_R_X5Y112_SLICE_X6Y112_CO6;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_D3 = CLBLM_R_X5Y115_SLICE_X6Y115_BO6;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_C1 = 1'b1;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_C2 = 1'b1;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_C3 = 1'b1;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_C4 = 1'b1;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_C5 = 1'b1;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_C6 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_D4 = CLBLM_R_X5Y116_SLICE_X6Y116_CO6;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_D5 = CLBLM_R_X5Y113_SLICE_X6Y113_DO6;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_D6 = CLBLM_R_X5Y114_SLICE_X6Y114_BO6;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_D1 = 1'b1;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_D2 = 1'b1;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_D3 = 1'b1;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_D4 = 1'b1;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_D5 = 1'b1;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_D6 = 1'b1;
  assign LIOB33_SING_X0Y149_IOB_X0Y149_O = CLBLM_R_X3Y113_SLICE_X3Y113_AO5;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_D1 = CLBLL_L_X4Y116_SLICE_X5Y116_BO5;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_T1 = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_D1 = CLBLL_L_X4Y116_SLICE_X5Y116_BO6;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_T1 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_A1 = CLBLL_L_X4Y114_SLICE_X5Y114_AO6;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_A2 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_A3 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_A4 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_A5 = CLBLM_R_X7Y114_SLICE_X9Y114_CO6;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_A6 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_B1 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_B2 = CLBLM_R_X7Y114_SLICE_X8Y114_CO6;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_B3 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_B4 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_B5 = CLBLM_R_X7Y114_SLICE_X9Y114_DO6;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_B6 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_A1 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_A2 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_A3 = CLBLM_R_X3Y105_SLICE_X2Y105_AO6;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_A4 = CLBLM_R_X3Y104_SLICE_X3Y104_BO6;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_C5 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_A5 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_A6 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_C1 = CLBLM_R_X7Y114_SLICE_X9Y114_DO6;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_C2 = CLBLM_R_X7Y114_SLICE_X8Y114_CO6;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_C3 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_B1 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_B2 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_B3 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_B4 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_B5 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_B6 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_D1 = CLBLM_R_X7Y114_SLICE_X9Y114_CO6;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_D2 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_C1 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_C2 = CLBLM_R_X5Y104_SLICE_X6Y104_AO6;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_C3 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_C4 = CLBLM_R_X3Y105_SLICE_X2Y105_AO6;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_C5 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_C6 = CLBLM_R_X3Y104_SLICE_X3Y104_BO6;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_D4 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_A1 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_A2 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_A3 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_A4 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_A5 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_A6 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_D1 = CLBLM_R_X3Y104_SLICE_X3Y104_CO6;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_D2 = CLBLL_L_X4Y105_SLICE_X4Y105_BO6;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_D3 = CLBLM_R_X3Y104_SLICE_X3Y104_DO6;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_D4 = CLBLL_L_X2Y106_SLICE_X0Y106_CO6;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_D5 = CLBLM_R_X3Y105_SLICE_X3Y105_BO5;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_D6 = CLBLM_R_X3Y105_SLICE_X3Y105_BO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_B1 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_B2 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_B3 = CLBLM_R_X7Y115_SLICE_X8Y115_AO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_B4 = CLBLM_R_X7Y113_SLICE_X9Y113_CO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_B5 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_A1 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_A2 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_A3 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_A4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_A5 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_C4 = CLBLM_R_X7Y113_SLICE_X9Y113_CO6;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_A6 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_C6 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_C1 = CLBLM_R_X7Y115_SLICE_X8Y115_AO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_C2 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_C3 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_B1 = CLBLL_L_X2Y106_SLICE_X0Y106_AO5;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_B2 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_B3 = CLBLM_R_X3Y105_SLICE_X3Y105_AO6;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_B4 = CLBLM_R_X3Y105_SLICE_X3Y105_CO6;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_B5 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_B6 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_D1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_D2 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_D3 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_C1 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_C2 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_C3 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_C4 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_C5 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_C6 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_D4 = CLBLM_R_X7Y116_SLICE_X8Y116_AO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_D5 = CLBLM_R_X7Y116_SLICE_X9Y116_AO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_D6 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_D1 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_D2 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_D3 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_D4 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_D5 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_D6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_D = RIOB33_X105Y107_IOB_X1Y108_I;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_D = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_A1 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_A2 = CLBLM_R_X7Y114_SLICE_X9Y114_BO6;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_A3 = CLBLL_L_X4Y115_SLICE_X5Y115_AO6;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_A4 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_A5 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_A6 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_B1 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_B2 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_B3 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_B4 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_B5 = CLBLM_R_X7Y114_SLICE_X8Y114_BO6;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_B6 = CLBLM_R_X7Y114_SLICE_X9Y114_BO6;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_A1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_A2 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_A3 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_C4 = CLBLM_R_X5Y116_SLICE_X7Y116_AO5;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_C5 = CLBLL_L_X4Y115_SLICE_X5Y115_AO6;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_C6 = CLBLM_R_X5Y115_SLICE_X7Y115_BO6;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_A4 = CLBLL_L_X2Y106_SLICE_X0Y106_CO6;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_A5 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_A6 = CLBLM_R_X3Y105_SLICE_X3Y105_CO6;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_C1 = CLBLM_R_X7Y114_SLICE_X9Y114_BO6;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_C2 = CLBLM_R_X5Y116_SLICE_X6Y116_AO6;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_B1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_B2 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_B3 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_B4 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_B5 = CLBLL_L_X2Y106_SLICE_X0Y106_CO6;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_B6 = CLBLM_R_X3Y105_SLICE_X3Y105_CO6;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_D5 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_D6 = CLBLM_R_X5Y115_SLICE_X7Y115_CO6;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_D1 = CLBLM_R_X5Y115_SLICE_X7Y115_AO6;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_D2 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_C1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_C2 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_C3 = CLBLL_L_X2Y106_SLICE_X0Y106_CO6;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_C4 = CLBLM_R_X3Y105_SLICE_X3Y105_CO6;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_C5 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_C6 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_A1 = CLBLM_R_X5Y115_SLICE_X6Y115_CO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_A2 = CLBLM_R_X7Y116_SLICE_X8Y116_AO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_A3 = CLBLM_R_X7Y116_SLICE_X9Y116_CO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_A4 = CLBLM_R_X7Y116_SLICE_X8Y116_BO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_A5 = CLBLM_R_X5Y114_SLICE_X6Y114_CO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_A6 = CLBLM_R_X5Y115_SLICE_X6Y115_AO5;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_D1 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_D2 = CLBLM_R_X3Y105_SLICE_X3Y105_CO6;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_D3 = CLBLL_L_X2Y106_SLICE_X0Y106_CO6;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_D4 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_D5 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_D6 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_B6 = CLBLM_R_X5Y115_SLICE_X6Y115_AO5;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_B1 = CLBLM_R_X7Y116_SLICE_X8Y116_DO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_B2 = CLBLM_R_X7Y116_SLICE_X8Y116_AO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_B3 = CLBLM_R_X7Y113_SLICE_X9Y113_CO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_B4 = CLBLL_L_X4Y116_SLICE_X4Y116_AO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_B5 = CLBLM_R_X7Y116_SLICE_X9Y116_CO6;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_A1 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_C4 = CLBLM_R_X5Y115_SLICE_X6Y115_AO5;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_C5 = CLBLM_R_X7Y116_SLICE_X8Y116_DO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_C6 = CLBLL_L_X4Y116_SLICE_X4Y116_AO6;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_A2 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_A3 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_A4 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_A5 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_A6 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_B1 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_B2 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_B3 = CLBLL_L_X2Y106_SLICE_X1Y106_BO6;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_B4 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_B5 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_B6 = CLBLL_L_X2Y107_SLICE_X0Y107_DO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_D1 = CLBLM_R_X7Y116_SLICE_X8Y116_BO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_D2 = CLBLM_R_X5Y114_SLICE_X6Y114_DO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_D3 = CLBLM_R_X5Y116_SLICE_X7Y116_BO6;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_C1 = CLBLL_L_X2Y106_SLICE_X1Y106_BO6;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_C2 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_C3 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_C4 = CLBLL_L_X2Y107_SLICE_X0Y107_DO6;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_C5 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_C6 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_D5 = CLBLM_R_X7Y116_SLICE_X8Y116_CO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_D6 = CLBLM_R_X5Y116_SLICE_X6Y116_BO6;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_D1 = CLBLM_R_X3Y106_SLICE_X2Y106_AO6;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_D2 = CLBLL_L_X2Y107_SLICE_X1Y107_AO6;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_D3 = CLBLM_R_X3Y106_SLICE_X2Y106_CO6;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_D4 = CLBLM_R_X3Y106_SLICE_X2Y106_AO5;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_D5 = CLBLL_L_X2Y108_SLICE_X1Y108_DO6;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_D6 = CLBLL_L_X2Y106_SLICE_X1Y106_DO6;
  assign LIOB33_X0Y121_IOB_X0Y122_O = CLBLL_L_X2Y108_SLICE_X1Y108_AO6;
  assign LIOB33_X0Y121_IOB_X0Y121_O = CLBLL_L_X2Y108_SLICE_X0Y108_AO5;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_A1 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_A2 = CLBLL_L_X4Y107_SLICE_X4Y107_AO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_A3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_A4 = CLBLM_R_X3Y107_SLICE_X3Y107_BO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_A5 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_A6 = CLBLL_L_X4Y106_SLICE_X5Y106_BO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_B1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_B2 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_B3 = CLBLM_R_X3Y106_SLICE_X2Y106_BO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_B4 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_B5 = CLBLM_R_X3Y105_SLICE_X2Y105_BO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_B6 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_D1 = CLBLL_L_X4Y116_SLICE_X4Y116_BO6;
  assign LIOI3_X0Y103_ILOGIC_X0Y104_D = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_C1 = CLBLM_L_X8Y107_SLICE_X11Y107_CO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_C2 = CLBLL_L_X4Y106_SLICE_X4Y106_BO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_C3 = CLBLM_R_X3Y108_SLICE_X3Y108_CO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_C4 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_C5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_C6 = CLBLM_R_X3Y106_SLICE_X3Y106_CO6;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_T1 = 1'b1;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_D1 = CLBLM_L_X8Y107_SLICE_X11Y107_CO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_D2 = CLBLM_R_X3Y106_SLICE_X3Y106_DO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_D3 = CLBLL_L_X4Y106_SLICE_X4Y106_AO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_D4 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_D5 = CLBLL_L_X4Y106_SLICE_X4Y106_BO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_D6 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_D1 = CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_A1 = 1'b1;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_A2 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_A3 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_A4 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_A5 = CLBLM_R_X3Y107_SLICE_X2Y107_CO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_A6 = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_T1 = 1'b1;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_B1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_B2 = CLBLM_R_X3Y105_SLICE_X2Y105_BO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_B3 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_B4 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_B5 = CLBLM_R_X3Y106_SLICE_X2Y106_BO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_B6 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_C1 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_C2 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_C3 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_C4 = CLBLL_L_X4Y106_SLICE_X4Y106_BO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_C5 = CLBLL_L_X2Y107_SLICE_X1Y107_CO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_C6 = CLBLM_R_X3Y107_SLICE_X2Y107_BO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_D1 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_D2 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_D3 = CLBLL_L_X4Y106_SLICE_X4Y106_BO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_D4 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_D5 = CLBLM_R_X3Y106_SLICE_X2Y106_DO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_D6 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign LIOB33_X0Y123_IOB_X0Y124_O = CLBLL_L_X2Y107_SLICE_X1Y107_AO5;
  assign LIOB33_X0Y123_IOB_X0Y123_O = CLBLL_L_X2Y108_SLICE_X0Y108_CO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_A1 = CLBLM_R_X3Y107_SLICE_X2Y107_DO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_A2 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_A3 = CLBLM_R_X3Y107_SLICE_X3Y107_AO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_A4 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_A5 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_A6 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_B1 = CLBLM_R_X3Y107_SLICE_X2Y107_DO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_B2 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_B3 = CLBLM_R_X3Y107_SLICE_X3Y107_AO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_B4 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_B5 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_B6 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_C1 = CLBLM_R_X3Y107_SLICE_X3Y107_AO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_C2 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_C3 = CLBLM_R_X3Y107_SLICE_X2Y107_DO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_C4 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_C5 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_C6 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_D1 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_D2 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_D3 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_D4 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_D5 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_D6 = 1'b1;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_B1 = CLBLM_L_X12Y105_SLICE_X16Y105_AO5;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_B2 = CLBLM_R_X11Y105_SLICE_X14Y105_BO6;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_A1 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_A2 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_A3 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_A4 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_A5 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_A6 = 1'b1;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_B3 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_B1 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_B2 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_B3 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_B4 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_B5 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_B6 = 1'b1;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_B5 = CLBLM_R_X11Y105_SLICE_X15Y105_AO6;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_C1 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_C2 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_C3 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_C4 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_C5 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_C6 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_D1 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_D2 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_D3 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_D4 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_D5 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_D6 = 1'b1;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_C1 = CLBLM_R_X11Y105_SLICE_X15Y105_AO6;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_C2 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_D5 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_D6 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign LIOB33_X0Y125_IOB_X0Y126_O = CLBLM_R_X3Y108_SLICE_X3Y108_AO6;
  assign LIOB33_X0Y125_IOB_X0Y125_O = CLBLM_R_X3Y107_SLICE_X2Y107_AO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_A1 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_A2 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_A3 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_A4 = CLBLL_L_X4Y108_SLICE_X4Y108_AO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_A5 = CLBLL_L_X4Y108_SLICE_X4Y108_BO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_A6 = CLBLM_R_X3Y108_SLICE_X3Y108_BO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_B1 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_B2 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_B3 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_B4 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_B5 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_B6 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_C1 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_C2 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_C3 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_C4 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_C5 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_C6 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_D1 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_D2 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_D3 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_D4 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_D5 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_D6 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_A1 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_A2 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_A3 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_A4 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_A5 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_A6 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_B1 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_B2 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_B3 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_B4 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_B5 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_B6 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_C1 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_C2 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_C3 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_C4 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_C5 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_C6 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_D1 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_D2 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_D3 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_D4 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_D5 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_D6 = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_D1 = CLBLL_L_X4Y113_SLICE_X4Y113_BO6;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_T1 = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_D1 = CLBLL_L_X4Y114_SLICE_X4Y114_AO6;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_T1 = 1'b1;
  assign LIOB33_X0Y127_IOB_X0Y128_O = CLBLM_R_X3Y110_SLICE_X3Y110_AO6;
  assign LIOB33_X0Y127_IOB_X0Y127_O = CLBLL_L_X4Y109_SLICE_X4Y109_AO6;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_D3 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_D4 = CLBLM_R_X5Y116_SLICE_X7Y116_CO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_A1 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_A2 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_A3 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_A4 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_A5 = CLBLM_R_X3Y109_SLICE_X3Y109_AO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_A6 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_B1 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_B2 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_B3 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_B4 = CLBLL_L_X4Y109_SLICE_X5Y109_AO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_B5 = CLBLL_L_X4Y109_SLICE_X4Y109_BO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_B6 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_C1 = CLBLM_R_X3Y108_SLICE_X3Y108_CO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_C2 = CLBLM_R_X5Y109_SLICE_X7Y109_CO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_C3 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_C4 = CLBLM_R_X3Y107_SLICE_X3Y107_DO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_C5 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_C6 = CLBLM_R_X5Y110_SLICE_X6Y110_AO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_D1 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_D2 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_D3 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_D4 = CLBLL_L_X4Y110_SLICE_X5Y110_CO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_D5 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_D6 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_A1 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_A2 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_A3 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_A4 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_A5 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_A6 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_B1 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_B2 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_B3 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_B4 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_B5 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_B6 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_C1 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_C2 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_C3 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_C4 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_C5 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_C6 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_C5 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_D1 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_D2 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_D3 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_D4 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_D5 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_D6 = 1'b1;
  assign CLBLM_L_X12Y105_SLICE_X17Y105_A1 = 1'b1;
  assign CLBLM_L_X12Y105_SLICE_X17Y105_A2 = 1'b1;
  assign CLBLM_L_X12Y105_SLICE_X17Y105_A3 = 1'b1;
  assign CLBLM_L_X12Y105_SLICE_X17Y105_A4 = 1'b1;
  assign CLBLM_L_X12Y105_SLICE_X17Y105_A5 = 1'b1;
  assign CLBLM_L_X12Y105_SLICE_X17Y105_A6 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_C6 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_L_X12Y105_SLICE_X17Y105_B1 = 1'b1;
  assign CLBLM_L_X12Y105_SLICE_X17Y105_B2 = 1'b1;
  assign CLBLM_L_X12Y105_SLICE_X17Y105_B3 = 1'b1;
  assign CLBLM_L_X12Y105_SLICE_X17Y105_B4 = 1'b1;
  assign CLBLM_L_X12Y105_SLICE_X17Y105_B5 = 1'b1;
  assign CLBLM_L_X12Y105_SLICE_X17Y105_B6 = 1'b1;
  assign CLBLM_L_X12Y105_SLICE_X17Y105_C1 = 1'b1;
  assign CLBLM_L_X12Y105_SLICE_X17Y105_C2 = 1'b1;
  assign CLBLM_L_X12Y105_SLICE_X17Y105_C3 = 1'b1;
  assign CLBLM_L_X12Y105_SLICE_X17Y105_C4 = 1'b1;
  assign CLBLM_L_X12Y105_SLICE_X17Y105_C5 = 1'b1;
  assign CLBLM_L_X12Y105_SLICE_X17Y105_C6 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_C4 = 1'b1;
  assign CLBLM_L_X12Y105_SLICE_X17Y105_D1 = 1'b1;
  assign CLBLM_L_X12Y105_SLICE_X17Y105_D2 = 1'b1;
  assign CLBLM_L_X12Y105_SLICE_X17Y105_D3 = 1'b1;
  assign CLBLM_L_X12Y105_SLICE_X17Y105_D4 = 1'b1;
  assign CLBLM_L_X12Y105_SLICE_X17Y105_D5 = 1'b1;
  assign CLBLM_L_X12Y105_SLICE_X17Y105_D6 = 1'b1;
  assign CLBLM_L_X12Y105_SLICE_X16Y105_A1 = CLBLM_L_X12Y105_SLICE_X16Y105_DO6;
  assign CLBLM_L_X12Y105_SLICE_X16Y105_A2 = CLBLM_R_X11Y107_SLICE_X14Y107_DO6;
  assign CLBLM_L_X12Y105_SLICE_X16Y105_A3 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_L_X12Y105_SLICE_X16Y105_A4 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X12Y105_SLICE_X16Y105_A5 = 1'b1;
  assign CLBLM_L_X12Y105_SLICE_X16Y105_A6 = 1'b1;
  assign CLBLM_L_X12Y105_SLICE_X16Y105_B1 = CLBLM_L_X12Y105_SLICE_X16Y105_DO6;
  assign CLBLM_L_X12Y105_SLICE_X16Y105_B2 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_L_X12Y105_SLICE_X16Y105_B3 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_L_X12Y105_SLICE_X16Y105_B4 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X12Y105_SLICE_X16Y105_B5 = CLBLM_R_X11Y107_SLICE_X14Y107_DO6;
  assign CLBLM_L_X12Y105_SLICE_X16Y105_B6 = CLBLM_L_X12Y105_SLICE_X16Y105_CO6;
  assign CLBLM_L_X12Y105_SLICE_X16Y105_C1 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X12Y105_SLICE_X16Y105_C2 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_L_X12Y105_SLICE_X16Y105_C3 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_L_X12Y105_SLICE_X16Y105_C4 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_L_X12Y105_SLICE_X16Y105_C5 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_L_X12Y105_SLICE_X16Y105_C6 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign LIOB33_X0Y129_IOB_X0Y129_O = CLBLM_R_X3Y110_SLICE_X3Y110_BO6;
  assign LIOB33_X0Y129_IOB_X0Y130_O = CLBLL_L_X2Y109_SLICE_X0Y109_BO5;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_C6 = 1'b1;
  assign CLBLM_L_X12Y105_SLICE_X16Y105_D1 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X12Y105_SLICE_X16Y105_D2 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_L_X12Y105_SLICE_X16Y105_D3 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_L_X12Y105_SLICE_X16Y105_D4 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_L_X12Y105_SLICE_X16Y105_D5 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_L_X12Y105_SLICE_X16Y105_D6 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_A1 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_A2 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_A3 = CLBLM_R_X5Y110_SLICE_X6Y110_AO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_A4 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_A5 = CLBLM_R_X5Y109_SLICE_X7Y109_CO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_A6 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_B1 = CLBLM_R_X7Y111_SLICE_X8Y111_BO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_B2 = CLBLM_R_X3Y112_SLICE_X3Y112_AO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_B3 = CLBLL_L_X4Y110_SLICE_X4Y110_DO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_B4 = CLBLM_R_X5Y110_SLICE_X6Y110_DO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_B5 = CLBLM_R_X3Y111_SLICE_X3Y111_AO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_B6 = CLBLM_R_X3Y107_SLICE_X3Y107_CO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_C1 = CLBLL_L_X4Y113_SLICE_X4Y113_AO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_C2 = CLBLM_R_X3Y112_SLICE_X3Y112_AO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_C3 = CLBLM_R_X7Y111_SLICE_X8Y111_BO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_C4 = CLBLM_R_X3Y110_SLICE_X3Y110_CO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_C5 = CLBLL_L_X4Y110_SLICE_X4Y110_DO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_C6 = CLBLM_R_X5Y110_SLICE_X6Y110_DO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_D1 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_D2 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_D3 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_D4 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_D5 = CLBLL_L_X4Y110_SLICE_X5Y110_CO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_D6 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_A1 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_A2 = CLBLM_R_X3Y111_SLICE_X3Y111_DO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_A3 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_A4 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_A5 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_A6 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_B1 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_B2 = CLBLM_R_X3Y111_SLICE_X3Y111_DO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_B3 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_B4 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_B5 = CLBLL_L_X4Y110_SLICE_X5Y110_AO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_B6 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_C1 = CLBLL_L_X4Y110_SLICE_X5Y110_AO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_C2 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_C3 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_C4 = CLBLM_R_X3Y111_SLICE_X2Y111_AO5;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_C5 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_C6 = CLBLL_L_X2Y111_SLICE_X1Y111_AO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_D1 = CLBLL_L_X4Y110_SLICE_X5Y110_AO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_D2 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_D3 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_D4 = CLBLM_R_X3Y111_SLICE_X2Y111_AO5;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_D5 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_D6 = CLBLL_L_X2Y111_SLICE_X1Y111_AO6;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_A1 = 1'b1;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_A2 = 1'b1;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_A3 = 1'b1;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_A4 = 1'b1;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_A5 = 1'b1;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_A6 = 1'b1;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_B1 = 1'b1;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_B2 = 1'b1;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_B3 = 1'b1;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_B4 = 1'b1;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_B5 = 1'b1;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_B6 = 1'b1;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_C1 = 1'b1;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_C2 = 1'b1;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_C3 = 1'b1;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_C4 = 1'b1;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_C5 = 1'b1;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_C6 = 1'b1;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_D1 = 1'b1;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_D2 = 1'b1;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_D3 = 1'b1;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_D4 = 1'b1;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_D5 = 1'b1;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_D6 = 1'b1;
  assign LIOB33_X0Y131_IOB_X0Y131_O = CLBLL_L_X4Y111_SLICE_X4Y111_AO6;
  assign LIOB33_X0Y131_IOB_X0Y132_O = CLBLM_R_X3Y114_SLICE_X3Y114_AO5;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_A1 = 1'b1;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_A2 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_A3 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_A4 = CLBLM_L_X12Y106_SLICE_X16Y106_BO6;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_A5 = CLBLM_L_X12Y107_SLICE_X17Y107_AO6;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_A6 = 1'b1;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_B1 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_B2 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_B3 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_B4 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_B5 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_B6 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_C1 = CLBLM_L_X12Y105_SLICE_X16Y105_BO6;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_C2 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_C3 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_C4 = CLBLM_L_X12Y106_SLICE_X16Y106_AO5;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_C5 = CLBLM_L_X12Y105_SLICE_X16Y105_AO6;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_C6 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_D1 = 1'b1;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_D2 = 1'b1;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_D3 = 1'b1;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_D4 = 1'b1;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_D5 = 1'b1;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_D6 = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_D1 = CLBLM_R_X3Y113_SLICE_X3Y113_CO6;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_T1 = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_D1 = CLBLM_R_X3Y113_SLICE_X3Y113_AO6;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_T1 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_A1 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_A2 = CLBLM_R_X3Y111_SLICE_X2Y111_DO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_A3 = CLBLL_L_X4Y112_SLICE_X4Y112_CO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_A4 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_A5 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_A6 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_B1 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_B2 = CLBLM_R_X3Y111_SLICE_X2Y111_DO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_B3 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_B4 = CLBLL_L_X4Y112_SLICE_X4Y112_CO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_B5 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_B6 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_C1 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_C2 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_C3 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_C4 = CLBLL_L_X4Y111_SLICE_X4Y111_DO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_C5 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_C6 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_D1 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_D2 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_D3 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_D4 = CLBLM_R_X3Y112_SLICE_X3Y112_CO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_D5 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_D6 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_A1 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_A2 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_A3 = CLBLL_L_X4Y111_SLICE_X5Y111_DO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_A4 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_A5 = CLBLM_R_X3Y111_SLICE_X2Y111_BO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_A6 = CLBLM_R_X3Y111_SLICE_X2Y111_CO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_B1 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_B2 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_B3 = CLBLL_L_X4Y111_SLICE_X5Y111_DO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_B4 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_B5 = CLBLM_R_X3Y111_SLICE_X2Y111_BO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_B6 = CLBLM_R_X3Y111_SLICE_X2Y111_CO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_C1 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_C2 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_C3 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_C4 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_C5 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_C6 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_D1 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_D2 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_D3 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_D4 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_D5 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_D6 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_A1 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_A2 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_A3 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_A4 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_A5 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_A6 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign LIOB33_X0Y133_IOB_X0Y134_O = 1'b0;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_B1 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_B2 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_B4 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_B5 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_B6 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign LIOB33_X0Y133_IOB_X0Y133_O = CLBLL_L_X4Y112_SLICE_X4Y112_AO6;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_C1 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_C2 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_C3 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_C4 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_C5 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_C6 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_D1 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_D2 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_D3 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_D4 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_D5 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_D6 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_A1 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_A2 = CLBLM_L_X12Y107_SLICE_X17Y107_BO6;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_A3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_A4 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_A5 = CLBLM_L_X12Y107_SLICE_X16Y107_CO6;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_A6 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_B1 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_B2 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_B3 = CLBLM_L_X12Y107_SLICE_X17Y107_AO6;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_B4 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_B5 = CLBLM_L_X12Y106_SLICE_X16Y106_BO6;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_B6 = CLBLM_R_X11Y107_SLICE_X14Y107_DO6;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_C1 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_C2 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_C3 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_C4 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_C5 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_C6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_D1 = CLBLM_L_X12Y106_SLICE_X16Y106_AO6;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_D2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_D3 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_D4 = CLBLM_L_X12Y107_SLICE_X16Y107_AO5;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_D5 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_D6 = CLBLM_L_X12Y107_SLICE_X16Y107_BO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_A1 = CLBLM_R_X3Y112_SLICE_X3Y112_DO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_A2 = CLBLL_L_X4Y113_SLICE_X4Y113_CO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_A3 = CLBLM_R_X3Y112_SLICE_X3Y112_BO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_A4 = CLBLM_R_X3Y113_SLICE_X3Y113_BO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_A5 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_A6 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_B1 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_B2 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_B3 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_B4 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_B5 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_B6 = CLBLM_R_X3Y112_SLICE_X3Y112_CO6;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_A4 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_C1 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_C2 = CLBLL_L_X4Y113_SLICE_X4Y113_CO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_C3 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_C4 = CLBLM_R_X3Y112_SLICE_X3Y112_BO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_C5 = CLBLM_R_X3Y113_SLICE_X3Y113_DO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_C6 = CLBLM_R_X3Y113_SLICE_X3Y113_BO6;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_A5 = 1'b1;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_A6 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_D1 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_D2 = CLBLM_R_X3Y112_SLICE_X3Y112_CO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_D3 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_D4 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_D5 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_D6 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_A1 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_A2 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_A3 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_A4 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_A5 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_A6 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_B1 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_B2 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_B3 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_B4 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_B5 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_B6 = 1'b1;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_B3 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_B4 = CLBLM_R_X11Y106_SLICE_X14Y106_CO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_C1 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_C2 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_C3 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_C4 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_C5 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_C6 = 1'b1;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_B5 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_B6 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign LIOB33_X0Y135_IOB_X0Y135_O = CLBLM_R_X5Y114_SLICE_X6Y114_AO5;
  assign LIOB33_X0Y135_IOB_X0Y136_O = CLBLM_R_X5Y114_SLICE_X6Y114_AO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_D1 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_D2 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_D3 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_D4 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_D5 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_D6 = 1'b1;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_A1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_A2 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_A3 = 1'b1;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_A5 = 1'b1;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_A6 = 1'b1;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_B1 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_B2 = CLBLM_R_X11Y107_SLICE_X14Y107_CO6;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_B3 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_B4 = CLBLM_R_X11Y107_SLICE_X15Y107_CO6;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_B6 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_C1 = CLBLM_R_X11Y106_SLICE_X15Y106_CO6;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_C2 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_C4 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_C5 = CLBLM_R_X13Y108_SLICE_X18Y108_AO6;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_C6 = CLBLM_R_X11Y106_SLICE_X14Y106_BO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_D4 = CLBLM_L_X10Y108_SLICE_X12Y108_CO6;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_D1 = CLBLM_R_X11Y107_SLICE_X14Y107_CO6;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_D3 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_D2 = CLBLM_R_X11Y107_SLICE_X15Y107_CO6;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_D5 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_D6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_D5 = CLBLM_R_X11Y110_SLICE_X15Y110_AO6;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_D4 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_D6 = CLBLM_L_X8Y108_SLICE_X10Y108_CO6;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_A1 = 1'b1;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_A2 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_A3 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_A4 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_A5 = 1'b1;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_A6 = 1'b1;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_B1 = 1'b1;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_B2 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_B3 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_B4 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_B5 = 1'b1;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_B6 = 1'b1;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_C1 = CLBLM_R_X13Y108_SLICE_X19Y108_BO6;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_C2 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_C3 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_C4 = CLBLM_R_X11Y108_SLICE_X15Y108_DO6;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_C5 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_C6 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_A1 = 1'b1;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_D1 = CLBLM_R_X11Y106_SLICE_X15Y106_AO6;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_D1 = CLBLM_R_X13Y108_SLICE_X19Y108_BO6;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_D2 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_D3 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_D4 = CLBLM_R_X11Y108_SLICE_X15Y108_DO6;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_D5 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_D6 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_D2 = CLBLM_R_X11Y106_SLICE_X14Y106_CO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_B1 = CLBLM_R_X7Y108_SLICE_X8Y108_AO5;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_B2 = CLBLM_L_X8Y108_SLICE_X10Y108_AO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_C1 = CLBLM_L_X8Y108_SLICE_X11Y108_BO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_C2 = CLBLM_R_X7Y107_SLICE_X9Y107_DO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_C3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_C6 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_A1 = CLBLM_R_X7Y113_SLICE_X9Y113_BO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_A2 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_A3 = CLBLM_R_X3Y111_SLICE_X3Y111_BO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_A4 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_A5 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_A6 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_B1 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_B2 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_B3 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_B4 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_B5 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_B6 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_C1 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_C2 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_C3 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_C4 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_C5 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_C6 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_D1 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_D2 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_D3 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_D4 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_D5 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_D6 = 1'b1;
  assign LIOB33_X0Y137_IOB_X0Y137_O = CLBLL_L_X4Y116_SLICE_X5Y116_AO6;
  assign LIOB33_X0Y137_IOB_X0Y138_O = CLBLL_L_X4Y116_SLICE_X5Y116_AO5;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_A1 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_A2 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_A3 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_A4 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_A5 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_A6 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_D4 = CLBLM_R_X7Y108_SLICE_X9Y108_CO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_D5 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_B1 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_B2 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_B3 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_B4 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_B5 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_B6 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_C1 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_C2 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_C3 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_C4 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_C5 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_C6 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_D1 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_D2 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_D3 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_D4 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_D5 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_D6 = 1'b1;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_A1 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_A2 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_A3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_A4 = 1'b1;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_A5 = 1'b1;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_A6 = 1'b1;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_B1 = CLBLM_R_X11Y106_SLICE_X15Y106_DO6;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_B2 = CLBLM_L_X12Y108_SLICE_X17Y108_BO6;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_B3 = CLBLM_L_X12Y108_SLICE_X16Y108_BO6;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_B4 = CLBLM_L_X12Y108_SLICE_X17Y108_AO6;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_B5 = CLBLM_L_X12Y109_SLICE_X17Y109_AO6;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_B6 = CLBLM_R_X13Y108_SLICE_X18Y108_BO6;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_C1 = CLBLM_L_X12Y109_SLICE_X17Y109_AO6;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_C2 = CLBLM_L_X12Y108_SLICE_X16Y108_BO6;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_C3 = CLBLM_R_X11Y106_SLICE_X15Y106_DO6;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_C4 = CLBLM_R_X13Y108_SLICE_X18Y108_BO6;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_C5 = CLBLM_L_X12Y108_SLICE_X17Y108_AO6;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_C6 = CLBLM_L_X12Y108_SLICE_X17Y108_BO6;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_D1 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_D2 = CLBLM_L_X12Y106_SLICE_X16Y106_CO6;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_D3 = CLBLM_R_X13Y108_SLICE_X18Y108_AO6;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_D4 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_D5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_D6 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_A1 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_A2 = 1'b1;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_A3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_A4 = 1'b1;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_A6 = 1'b1;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_B1 = CLBLM_L_X12Y108_SLICE_X17Y108_DO6;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_B2 = CLBLM_R_X13Y108_SLICE_X19Y108_BO6;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_B3 = CLBLM_R_X11Y108_SLICE_X15Y108_CO6;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_B4 = CLBLM_L_X12Y110_SLICE_X16Y110_AO6;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_B5 = CLBLM_L_X12Y108_SLICE_X16Y108_BO6;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_B6 = CLBLM_R_X11Y108_SLICE_X15Y108_AO5;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_C1 = CLBLM_R_X11Y108_SLICE_X15Y108_CO6;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_C2 = CLBLM_R_X13Y108_SLICE_X19Y108_BO6;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_C3 = CLBLM_L_X12Y108_SLICE_X17Y108_DO6;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_C4 = CLBLM_L_X12Y108_SLICE_X16Y108_BO6;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_C5 = CLBLM_R_X11Y108_SLICE_X15Y108_AO5;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_C6 = CLBLM_L_X12Y110_SLICE_X16Y110_AO6;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_D1 = CLBLM_R_X11Y108_SLICE_X15Y108_CO6;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_D2 = CLBLM_R_X13Y108_SLICE_X19Y108_BO6;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_D3 = CLBLM_L_X12Y108_SLICE_X17Y108_DO6;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_D4 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_D5 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_D6 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign LIOB33_X0Y139_IOB_X0Y140_O = CLBLL_L_X4Y116_SLICE_X5Y116_BO5;
  assign LIOB33_X0Y139_IOB_X0Y139_O = CLBLL_L_X4Y116_SLICE_X5Y116_BO6;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_A1 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_A2 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_A3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_A4 = CLBLM_L_X12Y110_SLICE_X17Y110_BO6;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_A5 = CLBLM_L_X12Y109_SLICE_X17Y109_CO6;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_A6 = CLBLM_L_X12Y108_SLICE_X16Y108_CO6;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_B1 = CLBLM_L_X12Y107_SLICE_X16Y107_DO6;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_B2 = CLBLM_L_X12Y108_SLICE_X17Y108_BO6;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_B3 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_B4 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_B6 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_C1 = CLBLM_R_X13Y108_SLICE_X18Y108_BO6;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_C2 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_C3 = CLBLM_R_X11Y106_SLICE_X15Y106_DO6;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_C5 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_C6 = CLBLM_L_X12Y108_SLICE_X17Y108_BO6;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_D1 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_D2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_D3 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_D4 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_D5 = CLBLM_R_X13Y108_SLICE_X18Y108_AO6;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_D6 = CLBLM_L_X12Y106_SLICE_X16Y106_CO6;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_A1 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_A2 = 1'b1;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_A3 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_A4 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_A5 = 1'b1;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_A6 = 1'b1;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_B1 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_B2 = CLBLM_L_X10Y107_SLICE_X13Y107_AO6;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_B3 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_B4 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_B5 = CLBLM_R_X11Y108_SLICE_X14Y108_DO6;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_B6 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_C1 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_C2 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_C3 = CLBLM_L_X12Y107_SLICE_X16Y107_DO6;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_C5 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_C6 = CLBLM_L_X12Y108_SLICE_X17Y108_BO6;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_D1 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_D2 = CLBLM_R_X11Y109_SLICE_X14Y109_AO5;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_D3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_D4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_D5 = CLBLM_R_X11Y109_SLICE_X14Y109_CO6;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_D6 = CLBLM_L_X12Y109_SLICE_X17Y109_DO6;
  assign LIOB33_X0Y141_IOB_X0Y142_O = CLBLL_L_X4Y116_SLICE_X4Y116_BO6;
  assign LIOB33_X0Y141_IOB_X0Y141_O = CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_A1 = 1'b1;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_A2 = 1'b1;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_A3 = 1'b1;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_A4 = 1'b1;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_A5 = 1'b1;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_A6 = 1'b1;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_B1 = 1'b1;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_B2 = 1'b1;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_B3 = 1'b1;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_B4 = 1'b1;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_B5 = 1'b1;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_B6 = 1'b1;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_C1 = 1'b1;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_C2 = 1'b1;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_C3 = 1'b1;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_C4 = 1'b1;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_C5 = 1'b1;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_C6 = 1'b1;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_D1 = 1'b1;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_D2 = 1'b1;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_D3 = 1'b1;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_D4 = 1'b1;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_D5 = 1'b1;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_D6 = 1'b1;
  assign LIOI3_SING_X0Y100_ILOGIC_X0Y100_D = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_A1 = CLBLM_L_X12Y110_SLICE_X16Y110_BO6;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_A2 = CLBLM_L_X12Y109_SLICE_X16Y109_BO6;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_A3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_A4 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_A5 = CLBLM_L_X12Y108_SLICE_X16Y108_DO6;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_A6 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_B1 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_B2 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_B3 = CLBLM_L_X12Y109_SLICE_X16Y109_DO6;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_B4 = CLBLM_L_X12Y110_SLICE_X16Y110_BO6;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_B5 = CLBLM_L_X12Y108_SLICE_X16Y108_DO6;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_B6 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_C1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_C2 = CLBLM_L_X12Y108_SLICE_X16Y108_DO6;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_C3 = CLBLM_L_X12Y109_SLICE_X16Y109_BO6;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_C4 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_C5 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_C6 = CLBLM_L_X12Y110_SLICE_X16Y110_BO6;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_D1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_D2 = CLBLM_L_X12Y110_SLICE_X16Y110_CO6;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_D3 = CLBLM_L_X12Y108_SLICE_X17Y108_CO6;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_D4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_D5 = CLBLM_L_X12Y110_SLICE_X17Y110_DO6;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_D6 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign LIOB33_X0Y143_IOB_X0Y143_O = CLBLL_L_X4Y115_SLICE_X4Y115_DO6;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_D1 = CLBLM_R_X3Y113_SLICE_X3Y113_AO5;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_T1 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_B6 = 1'b1;
  assign LIOB33_X0Y145_IOB_X0Y146_O = CLBLL_L_X4Y113_SLICE_X4Y113_BO6;
  assign LIOB33_X0Y145_IOB_X0Y145_O = CLBLL_L_X4Y114_SLICE_X4Y114_AO6;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_B1 = CLBLM_R_X11Y107_SLICE_X15Y107_AO6;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_B2 = CLBLM_L_X12Y107_SLICE_X17Y107_AO6;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_C4 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_C5 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_D3 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_C6 = CLBLM_L_X12Y107_SLICE_X17Y107_AO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_D4 = CLBLM_R_X11Y111_SLICE_X15Y111_DO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_D5 = LIOB33_X0Y109_IOB_X0Y109_I;
endmodule
