module top(
  input LIOB33_SING_X0Y50_IOB_X0Y50_IPAD,
  input LIOB33_X0Y51_IOB_X0Y51_IPAD,
  input LIOB33_X0Y51_IOB_X0Y52_IPAD,
  input LIOB33_X0Y53_IOB_X0Y53_IPAD,
  input LIOB33_X0Y53_IOB_X0Y54_IPAD,
  input LIOB33_X0Y55_IOB_X0Y55_IPAD,
  input LIOB33_X0Y55_IOB_X0Y56_IPAD,
  input LIOB33_X0Y57_IOB_X0Y57_IPAD,
  input LIOB33_X0Y57_IOB_X0Y58_IPAD,
  input LIOB33_X0Y59_IOB_X0Y59_IPAD,
  input LIOB33_X0Y59_IOB_X0Y60_IPAD,
  input LIOB33_X0Y61_IOB_X0Y61_IPAD,
  input LIOB33_X0Y61_IOB_X0Y62_IPAD,
  input LIOB33_X0Y63_IOB_X0Y63_IPAD,
  input LIOB33_X0Y77_IOB_X0Y78_IPAD,
  input RIOB33_SING_X105Y100_IOB_X1Y100_IPAD,
  input RIOB33_SING_X105Y149_IOB_X1Y149_IPAD,
  input RIOB33_X105Y101_IOB_X1Y101_IPAD,
  input RIOB33_X105Y101_IOB_X1Y102_IPAD,
  input RIOB33_X105Y103_IOB_X1Y103_IPAD,
  input RIOB33_X105Y103_IOB_X1Y104_IPAD,
  input RIOB33_X105Y105_IOB_X1Y105_IPAD,
  input RIOB33_X105Y105_IOB_X1Y106_IPAD,
  input RIOB33_X105Y107_IOB_X1Y107_IPAD,
  input RIOB33_X105Y107_IOB_X1Y108_IPAD,
  input RIOB33_X105Y109_IOB_X1Y109_IPAD,
  input RIOB33_X105Y109_IOB_X1Y110_IPAD,
  input RIOB33_X105Y111_IOB_X1Y111_IPAD,
  input RIOB33_X105Y111_IOB_X1Y112_IPAD,
  input RIOB33_X105Y113_IOB_X1Y113_IPAD,
  input RIOB33_X105Y113_IOB_X1Y114_IPAD,
  input RIOB33_X105Y115_IOB_X1Y115_IPAD,
  input RIOB33_X105Y115_IOB_X1Y116_IPAD,
  input RIOB33_X105Y117_IOB_X1Y117_IPAD,
  input RIOB33_X105Y117_IOB_X1Y118_IPAD,
  input RIOB33_X105Y119_IOB_X1Y119_IPAD,
  input RIOB33_X105Y119_IOB_X1Y120_IPAD,
  input RIOB33_X105Y121_IOB_X1Y121_IPAD,
  input RIOB33_X105Y121_IOB_X1Y122_IPAD,
  input RIOB33_X105Y123_IOB_X1Y123_IPAD,
  input RIOB33_X105Y123_IOB_X1Y124_IPAD,
  input RIOB33_X105Y125_IOB_X1Y125_IPAD,
  input RIOB33_X105Y125_IOB_X1Y126_IPAD,
  input RIOB33_X105Y127_IOB_X1Y127_IPAD,
  input RIOB33_X105Y127_IOB_X1Y128_IPAD,
  input RIOB33_X105Y129_IOB_X1Y129_IPAD,
  input RIOB33_X105Y129_IOB_X1Y130_IPAD,
  input RIOB33_X105Y131_IOB_X1Y131_IPAD,
  input RIOB33_X105Y131_IOB_X1Y132_IPAD,
  input RIOB33_X105Y133_IOB_X1Y133_IPAD,
  input RIOB33_X105Y133_IOB_X1Y134_IPAD,
  input RIOB33_X105Y135_IOB_X1Y135_IPAD,
  input RIOB33_X105Y135_IOB_X1Y136_IPAD,
  input RIOB33_X105Y137_IOB_X1Y137_IPAD,
  input RIOB33_X105Y137_IOB_X1Y138_IPAD,
  input RIOB33_X105Y139_IOB_X1Y139_IPAD,
  input RIOB33_X105Y139_IOB_X1Y140_IPAD,
  input RIOB33_X105Y141_IOB_X1Y141_IPAD,
  input RIOB33_X105Y141_IOB_X1Y142_IPAD,
  input RIOB33_X105Y143_IOB_X1Y143_IPAD,
  input RIOB33_X105Y143_IOB_X1Y144_IPAD,
  input RIOB33_X105Y145_IOB_X1Y145_IPAD,
  input RIOB33_X105Y145_IOB_X1Y146_IPAD,
  input RIOB33_X105Y147_IOB_X1Y147_IPAD,
  input RIOB33_X105Y147_IOB_X1Y148_IPAD,
  output LIOB33_SING_X0Y100_IOB_X0Y100_OPAD,
  output LIOB33_SING_X0Y149_IOB_X0Y149_OPAD,
  output LIOB33_SING_X0Y150_IOB_X0Y150_OPAD,
  output LIOB33_SING_X0Y199_IOB_X0Y199_OPAD,
  output LIOB33_X0Y101_IOB_X0Y101_OPAD,
  output LIOB33_X0Y101_IOB_X0Y102_OPAD,
  output LIOB33_X0Y103_IOB_X0Y103_OPAD,
  output LIOB33_X0Y103_IOB_X0Y104_OPAD,
  output LIOB33_X0Y105_IOB_X0Y105_OPAD,
  output LIOB33_X0Y105_IOB_X0Y106_OPAD,
  output LIOB33_X0Y107_IOB_X0Y107_OPAD,
  output LIOB33_X0Y107_IOB_X0Y108_OPAD,
  output LIOB33_X0Y109_IOB_X0Y109_OPAD,
  output LIOB33_X0Y109_IOB_X0Y110_OPAD,
  output LIOB33_X0Y111_IOB_X0Y111_OPAD,
  output LIOB33_X0Y111_IOB_X0Y112_OPAD,
  output LIOB33_X0Y113_IOB_X0Y113_OPAD,
  output LIOB33_X0Y113_IOB_X0Y114_OPAD,
  output LIOB33_X0Y115_IOB_X0Y115_OPAD,
  output LIOB33_X0Y115_IOB_X0Y116_OPAD,
  output LIOB33_X0Y117_IOB_X0Y117_OPAD,
  output LIOB33_X0Y117_IOB_X0Y118_OPAD,
  output LIOB33_X0Y119_IOB_X0Y119_OPAD,
  output LIOB33_X0Y119_IOB_X0Y120_OPAD,
  output LIOB33_X0Y121_IOB_X0Y121_OPAD,
  output LIOB33_X0Y121_IOB_X0Y122_OPAD,
  output LIOB33_X0Y123_IOB_X0Y123_OPAD,
  output LIOB33_X0Y123_IOB_X0Y124_OPAD,
  output LIOB33_X0Y125_IOB_X0Y125_OPAD,
  output LIOB33_X0Y125_IOB_X0Y126_OPAD,
  output LIOB33_X0Y127_IOB_X0Y127_OPAD,
  output LIOB33_X0Y127_IOB_X0Y128_OPAD,
  output LIOB33_X0Y129_IOB_X0Y129_OPAD,
  output LIOB33_X0Y129_IOB_X0Y130_OPAD,
  output LIOB33_X0Y131_IOB_X0Y131_OPAD,
  output LIOB33_X0Y131_IOB_X0Y132_OPAD,
  output LIOB33_X0Y133_IOB_X0Y133_OPAD,
  output LIOB33_X0Y133_IOB_X0Y134_OPAD,
  output LIOB33_X0Y135_IOB_X0Y135_OPAD,
  output LIOB33_X0Y135_IOB_X0Y136_OPAD,
  output LIOB33_X0Y137_IOB_X0Y137_OPAD,
  output LIOB33_X0Y137_IOB_X0Y138_OPAD,
  output LIOB33_X0Y139_IOB_X0Y139_OPAD,
  output LIOB33_X0Y139_IOB_X0Y140_OPAD,
  output LIOB33_X0Y141_IOB_X0Y141_OPAD,
  output LIOB33_X0Y141_IOB_X0Y142_OPAD,
  output LIOB33_X0Y143_IOB_X0Y143_OPAD,
  output LIOB33_X0Y145_IOB_X0Y145_OPAD,
  output LIOB33_X0Y145_IOB_X0Y146_OPAD,
  output LIOB33_X0Y147_IOB_X0Y147_OPAD,
  output LIOB33_X0Y147_IOB_X0Y148_OPAD,
  output LIOB33_X0Y151_IOB_X0Y151_OPAD,
  output LIOB33_X0Y151_IOB_X0Y152_OPAD,
  output LIOB33_X0Y153_IOB_X0Y153_OPAD,
  output LIOB33_X0Y153_IOB_X0Y154_OPAD,
  output LIOB33_X0Y155_IOB_X0Y155_OPAD,
  output LIOB33_X0Y155_IOB_X0Y156_OPAD,
  output LIOB33_X0Y157_IOB_X0Y157_OPAD,
  output LIOB33_X0Y157_IOB_X0Y158_OPAD,
  output LIOB33_X0Y159_IOB_X0Y159_OPAD,
  output LIOB33_X0Y159_IOB_X0Y160_OPAD,
  output LIOB33_X0Y161_IOB_X0Y161_OPAD,
  output LIOB33_X0Y161_IOB_X0Y162_OPAD,
  output LIOB33_X0Y163_IOB_X0Y163_OPAD,
  output LIOB33_X0Y163_IOB_X0Y164_OPAD,
  output LIOB33_X0Y165_IOB_X0Y165_OPAD,
  output LIOB33_X0Y165_IOB_X0Y166_OPAD,
  output LIOB33_X0Y167_IOB_X0Y167_OPAD,
  output LIOB33_X0Y167_IOB_X0Y168_OPAD,
  output LIOB33_X0Y169_IOB_X0Y169_OPAD,
  output LIOB33_X0Y169_IOB_X0Y170_OPAD,
  output LIOB33_X0Y171_IOB_X0Y171_OPAD,
  output LIOB33_X0Y171_IOB_X0Y172_OPAD,
  output LIOB33_X0Y173_IOB_X0Y173_OPAD,
  output LIOB33_X0Y173_IOB_X0Y174_OPAD,
  output LIOB33_X0Y175_IOB_X0Y175_OPAD,
  output LIOB33_X0Y175_IOB_X0Y176_OPAD,
  output LIOB33_X0Y177_IOB_X0Y177_OPAD,
  output LIOB33_X0Y177_IOB_X0Y178_OPAD,
  output LIOB33_X0Y179_IOB_X0Y179_OPAD,
  output LIOB33_X0Y179_IOB_X0Y180_OPAD,
  output LIOB33_X0Y181_IOB_X0Y181_OPAD,
  output LIOB33_X0Y181_IOB_X0Y182_OPAD,
  output LIOB33_X0Y183_IOB_X0Y183_OPAD,
  output LIOB33_X0Y183_IOB_X0Y184_OPAD,
  output LIOB33_X0Y185_IOB_X0Y185_OPAD,
  output LIOB33_X0Y185_IOB_X0Y186_OPAD,
  output LIOB33_X0Y187_IOB_X0Y187_OPAD,
  output LIOB33_X0Y187_IOB_X0Y188_OPAD,
  output LIOB33_X0Y189_IOB_X0Y189_OPAD,
  output LIOB33_X0Y189_IOB_X0Y190_OPAD,
  output LIOB33_X0Y191_IOB_X0Y191_OPAD,
  output LIOB33_X0Y191_IOB_X0Y192_OPAD,
  output LIOB33_X0Y193_IOB_X0Y193_OPAD,
  output LIOB33_X0Y193_IOB_X0Y194_OPAD,
  output LIOB33_X0Y195_IOB_X0Y195_OPAD,
  output LIOB33_X0Y195_IOB_X0Y196_OPAD,
  output LIOB33_X0Y197_IOB_X0Y197_OPAD,
  output LIOB33_X0Y197_IOB_X0Y198_OPAD,
  output LIOB33_X0Y63_IOB_X0Y64_OPAD,
  output LIOB33_X0Y65_IOB_X0Y65_OPAD,
  output LIOB33_X0Y65_IOB_X0Y66_OPAD,
  output RIOB33_SING_X105Y150_IOB_X1Y150_OPAD,
  output RIOB33_SING_X105Y199_IOB_X1Y199_OPAD,
  output RIOB33_X105Y151_IOB_X1Y151_OPAD,
  output RIOB33_X105Y151_IOB_X1Y152_OPAD,
  output RIOB33_X105Y153_IOB_X1Y153_OPAD,
  output RIOB33_X105Y153_IOB_X1Y154_OPAD,
  output RIOB33_X105Y155_IOB_X1Y155_OPAD,
  output RIOB33_X105Y155_IOB_X1Y156_OPAD,
  output RIOB33_X105Y157_IOB_X1Y157_OPAD,
  output RIOB33_X105Y157_IOB_X1Y158_OPAD,
  output RIOB33_X105Y159_IOB_X1Y159_OPAD,
  output RIOB33_X105Y159_IOB_X1Y160_OPAD,
  output RIOB33_X105Y161_IOB_X1Y161_OPAD,
  output RIOB33_X105Y161_IOB_X1Y162_OPAD,
  output RIOB33_X105Y163_IOB_X1Y163_OPAD,
  output RIOB33_X105Y163_IOB_X1Y164_OPAD,
  output RIOB33_X105Y165_IOB_X1Y165_OPAD,
  output RIOB33_X105Y165_IOB_X1Y166_OPAD,
  output RIOB33_X105Y167_IOB_X1Y167_OPAD,
  output RIOB33_X105Y167_IOB_X1Y168_OPAD,
  output RIOB33_X105Y169_IOB_X1Y169_OPAD,
  output RIOB33_X105Y169_IOB_X1Y170_OPAD,
  output RIOB33_X105Y171_IOB_X1Y171_OPAD,
  output RIOB33_X105Y171_IOB_X1Y172_OPAD,
  output RIOB33_X105Y173_IOB_X1Y173_OPAD,
  output RIOB33_X105Y173_IOB_X1Y174_OPAD,
  output RIOB33_X105Y175_IOB_X1Y175_OPAD,
  output RIOB33_X105Y175_IOB_X1Y176_OPAD,
  output RIOB33_X105Y177_IOB_X1Y177_OPAD,
  output RIOB33_X105Y177_IOB_X1Y178_OPAD,
  output RIOB33_X105Y179_IOB_X1Y179_OPAD,
  output RIOB33_X105Y179_IOB_X1Y180_OPAD,
  output RIOB33_X105Y181_IOB_X1Y181_OPAD,
  output RIOB33_X105Y181_IOB_X1Y182_OPAD,
  output RIOB33_X105Y183_IOB_X1Y183_OPAD,
  output RIOB33_X105Y183_IOB_X1Y184_OPAD,
  output RIOB33_X105Y185_IOB_X1Y185_OPAD,
  output RIOB33_X105Y185_IOB_X1Y186_OPAD,
  output RIOB33_X105Y187_IOB_X1Y187_OPAD,
  output RIOB33_X105Y187_IOB_X1Y188_OPAD,
  output RIOB33_X105Y189_IOB_X1Y189_OPAD,
  output RIOB33_X105Y189_IOB_X1Y190_OPAD,
  output RIOB33_X105Y191_IOB_X1Y191_OPAD,
  output RIOB33_X105Y191_IOB_X1Y192_OPAD,
  output RIOB33_X105Y193_IOB_X1Y193_OPAD,
  output RIOB33_X105Y193_IOB_X1Y194_OPAD,
  output RIOB33_X105Y195_IOB_X1Y195_OPAD,
  output RIOB33_X105Y195_IOB_X1Y196_OPAD,
  output RIOB33_X105Y197_IOB_X1Y197_OPAD,
  output RIOB33_X105Y197_IOB_X1Y198_OPAD
  );
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_A;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_A1;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_A2;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_A3;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_A4;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_A5;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_A6;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_AO5;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_AO6;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_A_CY;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_A_XOR;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_B;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_B1;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_B2;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_B3;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_B4;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_B5;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_B6;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_BO5;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_BO6;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_B_CY;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_B_XOR;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_C;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_C1;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_C2;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_C3;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_C4;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_C5;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_C6;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_CO5;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_CO6;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_C_CY;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_C_XOR;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_D;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_D1;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_D2;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_D3;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_D4;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_D5;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_D6;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_DO5;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_DO6;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_D_CY;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X0Y143_D_XOR;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_A;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_A1;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_A2;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_A3;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_A4;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_A5;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_A6;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_AO5;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_AO6;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_AQ;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_A_CY;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_A_XOR;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_B;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_B1;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_B2;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_B3;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_B4;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_B5;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_B6;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_BO5;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_BO6;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_BQ;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_B_CY;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_B_XOR;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_C;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_C1;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_C2;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_C3;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_C4;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_C5;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_C6;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_CLK;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_CO5;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_CO6;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_CQ;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_C_CY;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_C_XOR;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_D;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_D1;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_D2;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_D3;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_D4;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_D5;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_D6;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_DO5;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_DO6;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_DQ;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_D_CY;
  wire [0:0] CLBLL_L_X2Y143_SLICE_X1Y143_D_XOR;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_A;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_A1;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_A2;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_A3;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_A4;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_A5;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_A6;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_AO5;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_AO6;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_AQ;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_AX;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_A_CY;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_A_XOR;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_B;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_B1;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_B2;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_B3;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_B4;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_B5;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_B6;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_BO5;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_BO6;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_B_CY;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_B_XOR;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_C;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_C1;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_C2;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_C3;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_C4;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_C5;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_C6;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_CLK;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_CO5;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_CO6;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_C_CY;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_C_XOR;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_D;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_D1;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_D2;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_D3;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_D4;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_D5;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_D6;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_DO5;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_DO6;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_D_CY;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_D_XOR;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X0Y144_SR;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_A;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_A1;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_A2;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_A3;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_A4;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_A5;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_A5Q;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_A6;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_AMUX;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_AO5;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_AO6;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_AQ;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_A_CY;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_A_XOR;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_B;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_B1;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_B2;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_B3;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_B4;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_B5;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_B5Q;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_B6;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_BMUX;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_BO5;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_BO6;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_BQ;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_B_CY;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_B_XOR;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_C;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_C1;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_C2;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_C3;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_C4;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_C5;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_C6;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_CLK;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_CO5;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_CO6;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_C_CY;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_C_XOR;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_D;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_D1;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_D2;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_D3;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_D4;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_D5;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_D6;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_DO5;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_DO6;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_D_CY;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_D_XOR;
  wire [0:0] CLBLL_L_X2Y144_SLICE_X1Y144_SR;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_A;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_A1;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_A2;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_A3;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_A4;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_A5;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_A6;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_AO5;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_AO6;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_A_CY;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_A_XOR;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_B;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_B1;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_B2;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_B3;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_B4;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_B5;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_B6;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_BO5;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_BO6;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_B_CY;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_B_XOR;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_C;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_C1;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_C2;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_C3;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_C4;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_C5;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_C6;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_CO5;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_CO6;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_C_CY;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_C_XOR;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_D;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_D1;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_D2;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_D3;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_D4;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_D5;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_D6;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_DO5;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_DO6;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_D_CY;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X0Y145_D_XOR;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_A;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_A1;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_A2;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_A3;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_A4;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_A5;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_A5Q;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_A6;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_AMUX;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_AO5;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_AO6;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_AQ;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_A_CY;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_A_XOR;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_B;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_B1;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_B2;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_B3;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_B4;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_B5;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_B6;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_BO5;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_BO6;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_B_CY;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_B_XOR;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_C;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_C1;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_C2;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_C3;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_C4;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_C5;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_C6;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_CLK;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_CO5;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_CO6;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_C_CY;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_C_XOR;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_D;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_D1;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_D2;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_D3;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_D4;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_D5;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_D6;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_DO5;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_DO6;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_D_CY;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_D_XOR;
  wire [0:0] CLBLL_L_X2Y145_SLICE_X1Y145_SR;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_A;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_A1;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_A2;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_A3;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_A4;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_A5;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_A6;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_AO5;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_AO6;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_A_CY;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_A_XOR;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_B;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_B1;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_B2;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_B3;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_B4;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_B5;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_B6;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_BO5;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_BO6;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_B_CY;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_B_XOR;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_C;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_C1;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_C2;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_C3;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_C4;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_C5;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_C6;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_CO5;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_CO6;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_C_CY;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_C_XOR;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_D;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_D1;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_D2;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_D3;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_D4;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_D5;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_D6;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_DO5;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_DO6;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_D_CY;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X0Y146_D_XOR;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_A;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_A1;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_A2;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_A3;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_A4;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_A5;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_A5Q;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_A6;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_AMUX;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_AO5;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_AO6;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_AQ;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_A_CY;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_A_XOR;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_B;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_B1;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_B2;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_B3;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_B4;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_B5;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_B6;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_BO5;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_BO6;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_B_CY;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_B_XOR;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_C;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_C1;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_C2;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_C3;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_C4;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_C5;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_C6;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_CLK;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_CO5;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_CO6;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_C_CY;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_C_XOR;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_D;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_D1;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_D2;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_D3;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_D4;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_D5;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_D6;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_DO5;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_DO6;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_D_CY;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_D_XOR;
  wire [0:0] CLBLL_L_X2Y146_SLICE_X1Y146_SR;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_A;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_A1;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_A2;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_A3;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_A4;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_A5;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_A6;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_AO5;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_AO6;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_AQ;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_A_CY;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_A_XOR;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_B;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_B1;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_B2;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_B3;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_B4;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_B5;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_B5Q;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_B6;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_BMUX;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_BO5;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_BO6;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_BQ;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_B_CY;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_B_XOR;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_C;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_C1;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_C2;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_C3;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_C4;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_C5;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_C6;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_CLK;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_CO5;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_CO6;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_C_CY;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_C_XOR;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_D;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_D1;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_D2;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_D3;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_D4;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_D5;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_D6;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_DO5;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_DO6;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_D_CY;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X0Y147_D_XOR;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_A;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_A1;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_A2;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_A3;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_A4;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_A5;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_A5Q;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_A6;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_AMUX;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_AO5;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_AO6;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_AQ;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_A_CY;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_A_XOR;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_B;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_B1;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_B2;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_B3;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_B4;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_B5;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_B6;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_BO5;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_BO6;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_B_CY;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_B_XOR;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_C;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_C1;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_C2;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_C3;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_C4;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_C5;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_C6;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_CLK;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_CO5;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_CO6;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_C_CY;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_C_XOR;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_D;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_D1;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_D2;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_D3;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_D4;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_D5;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_D6;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_DO5;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_DO6;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_D_CY;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_D_XOR;
  wire [0:0] CLBLL_L_X2Y147_SLICE_X1Y147_SR;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_A;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_A1;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_A2;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_A3;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_A4;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_A5;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_A5Q;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_A6;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_AMUX;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_AO5;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_AO6;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_AQ;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_A_CY;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_A_XOR;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_B;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_B1;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_B2;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_B3;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_B4;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_B5;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_B5Q;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_B6;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_BMUX;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_BO5;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_BO6;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_BQ;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_B_CY;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_B_XOR;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_C;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_C1;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_C2;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_C3;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_C4;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_C5;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_C6;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_CLK;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_CO5;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_CO6;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_C_CY;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_C_XOR;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_D;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_D1;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_D2;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_D3;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_D4;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_D5;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_D6;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_DO5;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_DO6;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_D_CY;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X0Y148_D_XOR;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_A;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_A1;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_A2;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_A3;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_A4;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_A5;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_A5Q;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_A6;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_AMUX;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_AO5;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_AO6;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_AQ;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_A_CY;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_A_XOR;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_B;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_B1;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_B2;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_B3;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_B4;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_B5;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_B6;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_BMUX;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_BO5;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_BO6;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_B_CY;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_B_XOR;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_C;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_C1;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_C2;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_C3;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_C4;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_C5;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_C6;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_CLK;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_CO5;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_CO6;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_C_CY;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_C_XOR;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_D;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_D1;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_D2;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_D3;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_D4;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_D5;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_D6;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_DO5;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_DO6;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_D_CY;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_D_XOR;
  wire [0:0] CLBLL_L_X2Y148_SLICE_X1Y148_SR;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_A;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_A1;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_A2;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_A3;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_A4;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_A5;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_A6;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_AO5;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_AO6;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_AQ;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_A_CY;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_A_XOR;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_B;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_B1;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_B2;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_B3;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_B4;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_B5;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_B6;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_BO5;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_BO6;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_B_CY;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_B_XOR;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_C;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_C1;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_C2;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_C3;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_C4;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_C5;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_C6;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_CLK;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_CO5;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_CO6;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_C_CY;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_C_XOR;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_D;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_D1;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_D2;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_D3;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_D4;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_D5;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_D6;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_DO5;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_DO6;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_D_CY;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X0Y149_D_XOR;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_A;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_A1;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_A2;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_A3;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_A4;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_A5;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_A5Q;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_A6;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_AMUX;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_AO5;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_AO6;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_AQ;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_A_CY;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_A_XOR;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_B;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_B1;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_B2;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_B3;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_B4;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_B5;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_B6;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_BO5;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_BO6;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_BQ;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_B_CY;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_B_XOR;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_C;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_C1;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_C2;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_C3;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_C4;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_C5;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_C6;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_CLK;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_CO5;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_CO6;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_CQ;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_C_CY;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_C_XOR;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_D;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_D1;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_D2;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_D3;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_D4;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_D5;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_D6;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_DO5;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_DO6;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_DQ;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_D_CY;
  wire [0:0] CLBLL_L_X2Y149_SLICE_X1Y149_D_XOR;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_A;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_A1;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_A2;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_A3;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_A4;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_A5;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_A6;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_AO5;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_AO6;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_A_CY;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_A_XOR;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_B;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_B1;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_B2;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_B3;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_B4;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_B5;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_B6;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_BO5;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_BO6;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_B_CY;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_B_XOR;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_C;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_C1;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_C2;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_C3;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_C4;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_C5;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_C6;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_CO5;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_CO6;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_C_CY;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_C_XOR;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_D;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_D1;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_D2;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_D3;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_D4;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_D5;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_D6;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_DO5;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_DO6;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_D_CY;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X0Y150_D_XOR;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_A;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_A1;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_A2;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_A3;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_A4;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_A5;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_A5Q;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_A6;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_AMUX;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_AO5;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_AO6;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_AQ;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_AX;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_A_CY;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_A_XOR;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_B;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_B1;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_B2;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_B3;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_B4;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_B5;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_B6;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_BMUX;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_BO5;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_BO6;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_B_CY;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_B_XOR;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_C;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_C1;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_C2;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_C3;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_C4;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_C5;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_C5Q;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_C6;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_CLK;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_CMUX;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_CO5;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_CO6;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_CQ;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_C_CY;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_C_XOR;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_D;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_D1;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_D2;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_D3;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_D4;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_D5;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_D6;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_DMUX;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_DO5;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_DO6;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_D_CY;
  wire [0:0] CLBLL_L_X2Y150_SLICE_X1Y150_D_XOR;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_A;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_A1;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_A2;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_A3;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_A4;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_A5;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_A6;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_AO5;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_AO6;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_A_CY;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_A_XOR;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_B;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_B1;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_B2;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_B3;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_B4;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_B5;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_B6;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_BO5;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_BO6;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_B_CY;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_B_XOR;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_C;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_C1;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_C2;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_C3;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_C4;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_C5;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_C6;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_CO5;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_CO6;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_C_CY;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_C_XOR;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_D;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_D1;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_D2;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_D3;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_D4;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_D5;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_D6;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_DO5;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_DO6;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_D_CY;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X0Y151_D_XOR;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_A;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_A1;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_A2;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_A3;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_A4;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_A5;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_A6;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_AO5;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_AO6;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_AQ;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_A_CY;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_A_XOR;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_B;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_B1;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_B2;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_B3;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_B4;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_B5;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_B6;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_BO5;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_BO6;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_BQ;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_B_CY;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_B_XOR;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_C;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_C1;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_C2;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_C3;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_C4;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_C5;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_C6;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_CLK;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_CO5;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_CO6;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_C_CY;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_C_XOR;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_D;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_D1;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_D2;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_D3;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_D4;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_D5;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_D6;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_DO5;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_DO6;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_D_CY;
  wire [0:0] CLBLL_L_X2Y151_SLICE_X1Y151_D_XOR;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_A;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_A1;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_A2;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_A3;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_A4;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_A5;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_A6;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_AO5;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_AO6;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_A_CY;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_A_XOR;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_B;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_B1;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_B2;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_B3;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_B4;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_B5;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_B6;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_BO5;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_BO6;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_B_CY;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_B_XOR;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_C;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_C1;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_C2;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_C3;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_C4;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_C5;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_C6;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_CO5;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_CO6;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_C_CY;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_C_XOR;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_D;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_D1;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_D2;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_D3;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_D4;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_D5;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_D6;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_DO5;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_DO6;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_D_CY;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X0Y152_D_XOR;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_A;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_A1;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_A2;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_A3;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_A4;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_A5;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_A6;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_AO5;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_AO6;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_A_CY;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_A_XOR;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_B;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_B1;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_B2;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_B3;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_B4;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_B5;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_B6;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_BO5;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_BO6;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_B_CY;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_B_XOR;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_C;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_C1;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_C2;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_C3;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_C4;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_C5;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_C6;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_CO5;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_CO6;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_C_CY;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_C_XOR;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_D;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_D1;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_D2;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_D3;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_D4;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_D5;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_D6;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_DO5;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_DO6;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_D_CY;
  wire [0:0] CLBLL_L_X2Y152_SLICE_X1Y152_D_XOR;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_A;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_A1;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_A2;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_A3;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_A4;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_A5;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_A6;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_AO5;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_AO6;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_A_CY;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_A_XOR;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_B;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_B1;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_B2;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_B3;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_B4;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_B5;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_B6;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_BO5;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_BO6;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_B_CY;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_B_XOR;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_C;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_C1;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_C2;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_C3;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_C4;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_C5;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_C6;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_CO5;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_CO6;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_C_CY;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_C_XOR;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_D;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_D1;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_D2;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_D3;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_D4;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_D5;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_D6;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_DO5;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_DO6;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_D_CY;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_D_XOR;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_A;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_A1;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_A2;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_A3;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_A4;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_A5;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_A6;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_AO5;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_AO6;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_AQ;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_AX;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_A_CY;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_A_XOR;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_B;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_B1;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_B2;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_B3;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_B4;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_B5;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_B6;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_BO5;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_BO6;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_B_CY;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_B_XOR;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_C;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_C1;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_C2;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_C3;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_C4;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_C5;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_C6;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_CLK;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_CO5;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_CO6;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_C_CY;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_C_XOR;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_D;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_D1;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_D2;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_D3;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_D4;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_D5;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_D6;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_DO5;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_DO6;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_D_CY;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_D_XOR;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X0Y166_A;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X0Y166_A1;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X0Y166_A2;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X0Y166_A3;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X0Y166_A4;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X0Y166_A5;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X0Y166_A6;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X0Y166_AO5;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X0Y166_AO6;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X0Y166_A_CY;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X0Y166_A_XOR;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X0Y166_B;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X0Y166_B1;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X0Y166_B2;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X0Y166_B3;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X0Y166_B4;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X0Y166_B5;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X0Y166_B6;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X0Y166_BO5;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X0Y166_BO6;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X0Y166_B_CY;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X0Y166_B_XOR;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X0Y166_C;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X0Y166_C1;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X0Y166_C2;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X0Y166_C3;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X0Y166_C4;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X0Y166_C5;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X0Y166_C6;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X0Y166_CO5;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X0Y166_CO6;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X0Y166_C_CY;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X0Y166_C_XOR;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X0Y166_D;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X0Y166_D1;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X0Y166_D2;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X0Y166_D3;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X0Y166_D4;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X0Y166_D5;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X0Y166_D6;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X0Y166_DO5;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X0Y166_DO6;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X0Y166_D_CY;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X0Y166_D_XOR;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X1Y166_A;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X1Y166_A1;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X1Y166_A2;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X1Y166_A3;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X1Y166_A4;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X1Y166_A5;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X1Y166_A6;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X1Y166_AO5;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X1Y166_AO6;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X1Y166_A_CY;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X1Y166_A_XOR;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X1Y166_B;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X1Y166_B1;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X1Y166_B2;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X1Y166_B3;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X1Y166_B4;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X1Y166_B5;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X1Y166_B6;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X1Y166_BO5;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X1Y166_BO6;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X1Y166_B_CY;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X1Y166_B_XOR;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X1Y166_C;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X1Y166_C1;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X1Y166_C2;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X1Y166_C3;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X1Y166_C4;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X1Y166_C5;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X1Y166_C6;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X1Y166_CO5;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X1Y166_CO6;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X1Y166_C_CY;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X1Y166_C_XOR;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X1Y166_D;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X1Y166_D1;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X1Y166_D2;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X1Y166_D3;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X1Y166_D4;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X1Y166_D5;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X1Y166_D6;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X1Y166_DO5;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X1Y166_DO6;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X1Y166_D_CY;
  wire [0:0] CLBLL_L_X2Y166_SLICE_X1Y166_D_XOR;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_A;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_A1;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_A2;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_A3;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_A4;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_A5;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_A6;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_AO5;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_AO6;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_A_CY;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_A_XOR;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_B;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_B1;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_B2;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_B3;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_B4;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_B5;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_B6;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_BO5;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_BO6;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_B_CY;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_B_XOR;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_C;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_C1;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_C2;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_C3;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_C4;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_C5;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_C6;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_CO5;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_CO6;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_C_CY;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_C_XOR;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_D;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_D1;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_D2;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_D3;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_D4;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_D5;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_D6;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_DO5;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_DO6;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_D_CY;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_D_XOR;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_A;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_A1;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_A2;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_A3;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_A4;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_A5;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_A6;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_AO5;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_AO6;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_A_CY;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_A_XOR;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_B;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_B1;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_B2;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_B3;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_B4;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_B5;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_B6;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_BO5;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_BO6;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_B_CY;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_B_XOR;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_C;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_C1;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_C2;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_C3;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_C4;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_C5;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_C6;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_CO5;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_CO6;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_C_CY;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_C_XOR;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_D;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_D1;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_D2;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_D3;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_D4;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_D5;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_D6;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_DO5;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_DO6;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_D_CY;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_D_XOR;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_A;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_A1;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_A2;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_A3;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_A4;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_A5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_A6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_AO5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_AO6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_A_CY;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_A_XOR;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_B;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_B1;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_B2;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_B3;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_B4;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_B5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_B6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_BO5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_BO6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_B_CY;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_B_XOR;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_C;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_C1;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_C2;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_C3;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_C4;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_C5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_C6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_CO5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_CO6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_C_CY;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_C_XOR;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_D;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_D1;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_D2;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_D3;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_D4;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_D5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_D6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_DO5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_DO6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_D_CY;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_D_XOR;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_A;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_A1;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_A2;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_A3;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_A4;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_A5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_A6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_AO5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_AO6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_AQ;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_A_CY;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_A_XOR;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_B;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_B1;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_B2;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_B3;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_B4;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_B5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_B6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_BO5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_BO6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_B_CY;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_B_XOR;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_C;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_C1;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_C2;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_C3;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_C4;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_C5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_C6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_CLK;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_CO5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_CO6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_C_CY;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_C_XOR;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_D;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_D1;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_D2;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_D3;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_D4;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_D5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_D6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_DO5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_DO6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_D_CY;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_D_XOR;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_SR;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_A;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_A1;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_A2;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_A3;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_A4;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_A5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_A6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_AO5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_AO6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_AQ;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_AX;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_A_CY;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_A_XOR;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_B;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_B1;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_B2;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_B3;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_B4;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_B5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_B6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_BO5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_BO6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_B_CY;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_B_XOR;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_C;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_C1;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_C2;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_C3;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_C4;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_C5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_C6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_CLK;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_CO5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_CO6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_C_CY;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_C_XOR;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_D;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_D1;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_D2;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_D3;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_D4;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_D5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_D6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_DO5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_DO6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_D_CY;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_D_XOR;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_SR;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_A;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_A1;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_A2;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_A3;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_A4;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_A5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_A5Q;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_A6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_AMUX;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_AO5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_AO6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_AQ;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_A_CY;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_A_XOR;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_B;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_B1;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_B2;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_B3;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_B4;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_B5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_B6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_BMUX;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_BO5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_BO6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_B_CY;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_B_XOR;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_C;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_C1;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_C2;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_C3;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_C4;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_C5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_C6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_CLK;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_CO5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_CO6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_C_CY;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_C_XOR;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_D;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_D1;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_D2;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_D3;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_D4;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_D5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_D6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_DO5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_DO6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_D_CY;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_D_XOR;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_SR;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_A;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_A1;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_A2;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_A3;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_A4;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_A5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_A5Q;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_A6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_AMUX;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_AO5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_AO6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_AQ;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_AX;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_A_CY;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_A_XOR;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_B;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_B1;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_B2;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_B3;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_B4;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_B5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_B6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_BMUX;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_BO5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_BO6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_B_CY;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_B_XOR;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_C;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_C1;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_C2;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_C3;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_C4;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_C5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_C6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_CLK;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_CMUX;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_CO5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_CO6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_C_CY;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_C_XOR;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_D;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_D1;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_D2;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_D3;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_D4;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_D5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_D6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_DMUX;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_DO5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_DO6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_D_CY;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_D_XOR;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_SR;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_A;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_A1;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_A2;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_A3;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_A4;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_A5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_A5Q;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_A6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_AMUX;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_AO5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_AO6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_AQ;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_AX;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_A_CY;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_A_XOR;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_B;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_B1;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_B2;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_B3;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_B4;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_B5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_B6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_BO5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_BO6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_BQ;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_B_CY;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_B_XOR;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_C;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_C1;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_C2;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_C3;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_C4;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_C5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_C6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_CLK;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_CO5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_CO6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_CQ;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_C_CY;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_C_XOR;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_D;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_D1;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_D2;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_D3;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_D4;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_D5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_D6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_DO5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_DO6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_D_CY;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_D_XOR;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_A;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_A1;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_A2;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_A3;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_A4;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_A5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_A6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_AO5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_AO6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_AQ;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_A_CY;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_A_XOR;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_B;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_B1;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_B2;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_B3;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_B4;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_B5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_B6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_BO5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_BO6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_BQ;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_B_CY;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_B_XOR;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_C;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_C1;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_C2;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_C3;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_C4;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_C5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_C6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_CLK;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_CO5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_CO6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_CQ;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_C_CY;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_C_XOR;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_D;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_D1;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_D2;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_D3;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_D4;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_D5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_D6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_DO5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_DO6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_DQ;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_D_CY;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_D_XOR;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_A;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_A1;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_A2;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_A3;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_A4;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_A5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_A6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_AO5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_AO6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_AQ;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_A_CY;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_A_XOR;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_B;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_B1;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_B2;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_B3;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_B4;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_B5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_B6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_BO5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_BO6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_BQ;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_B_CY;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_B_XOR;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_C;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_C1;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_C2;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_C3;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_C4;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_C5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_C5Q;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_C6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_CLK;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_CMUX;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_CO5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_CO6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_CQ;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_C_CY;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_C_XOR;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_D;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_D1;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_D2;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_D3;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_D4;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_D5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_D6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_DO5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_DO6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_DQ;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_D_CY;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_D_XOR;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_A;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_A1;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_A2;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_A3;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_A4;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_A5;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_A6;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_AO5;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_AO6;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_AQ;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_AX;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_A_CY;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_A_XOR;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_B;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_B1;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_B2;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_B3;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_B4;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_B5;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_B6;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_BMUX;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_BO5;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_BO6;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_B_CY;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_B_XOR;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_C;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_C1;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_C2;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_C3;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_C4;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_C5;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_C6;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_CLK;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_CO5;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_CO6;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_C_CY;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_C_XOR;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_D;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_D1;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_D2;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_D3;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_D4;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_D5;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_D6;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_DO5;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_DO6;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_D_CY;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_D_XOR;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X4Y144_SR;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_A;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_A1;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_A2;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_A3;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_A4;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_A5;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_A6;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_AO5;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_AO6;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_AQ;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_A_CY;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_A_XOR;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_B;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_B1;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_B2;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_B3;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_B4;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_B5;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_B5Q;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_B6;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_BMUX;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_BO5;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_BO6;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_BQ;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_B_CY;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_B_XOR;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_C;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_C1;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_C2;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_C3;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_C4;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_C5;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_C5Q;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_C6;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_CLK;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_CMUX;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_CO5;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_CO6;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_CQ;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_C_CY;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_C_XOR;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_D;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_D1;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_D2;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_D3;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_D4;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_D5;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_D5Q;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_D6;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_DMUX;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_DO5;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_DO6;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_DQ;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_D_CY;
  wire [0:0] CLBLL_L_X4Y144_SLICE_X5Y144_D_XOR;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_A;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_A1;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_A2;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_A3;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_A4;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_A5;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_A5Q;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_A6;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_AMUX;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_AO5;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_AO6;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_AQ;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_A_CY;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_A_XOR;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_B;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_B1;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_B2;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_B3;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_B4;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_B5;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_B6;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_BO5;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_BO6;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_B_CY;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_B_XOR;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_C;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_C1;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_C2;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_C3;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_C4;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_C5;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_C6;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_CLK;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_CO5;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_CO6;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_C_CY;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_C_XOR;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_D;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_D1;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_D2;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_D3;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_D4;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_D5;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_D6;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_DO5;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_DO6;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_D_CY;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_D_XOR;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X4Y145_SR;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_A;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_A1;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_A2;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_A3;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_A4;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_A5;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_A6;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_AO5;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_AO6;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_AQ;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_AX;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_A_CY;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_A_XOR;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_B;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_B1;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_B2;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_B3;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_B4;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_B5;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_B6;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_BO5;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_BO6;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_BQ;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_BX;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_B_CY;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_B_XOR;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_C;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_C1;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_C2;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_C3;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_C4;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_C5;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_C6;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_CE;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_CLK;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_CO5;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_CO6;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_C_CY;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_C_XOR;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_D;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_D1;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_D2;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_D3;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_D4;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_D5;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_D6;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_DO5;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_DO6;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_D_CY;
  wire [0:0] CLBLL_L_X4Y145_SLICE_X5Y145_D_XOR;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_A;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_A1;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_A2;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_A3;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_A4;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_A5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_A6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_AO5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_AO6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_AQ;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_A_CY;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_A_XOR;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_B;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_B1;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_B2;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_B3;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_B4;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_B5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_B6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_BO5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_BO6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_BQ;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_B_CY;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_B_XOR;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_C;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_C1;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_C2;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_C3;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_C4;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_C5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_C6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_CLK;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_CO5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_CO6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_CQ;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_C_CY;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_C_XOR;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_D;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_D1;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_D2;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_D3;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_D4;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_D5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_D6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_DO5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_DO6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_DQ;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_D_CY;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_D_XOR;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_A;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_A1;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_A2;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_A3;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_A4;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_A5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_A5Q;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_A6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_AMUX;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_AO5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_AO6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_AQ;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_A_CY;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_A_XOR;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_B;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_B1;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_B2;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_B3;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_B4;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_B5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_B5Q;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_B6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_BMUX;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_BO5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_BO6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_BQ;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_B_CY;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_B_XOR;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_C;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_C1;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_C2;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_C3;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_C4;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_C5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_C6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_CLK;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_CMUX;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_CO5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_CO6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_C_CY;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_C_XOR;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_D;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_D1;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_D2;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_D3;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_D4;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_D5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_D6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_DO5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_DO6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_D_CY;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_D_XOR;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_SR;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_A;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_A1;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_A2;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_A3;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_A4;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_A5;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_A6;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_AO5;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_AO6;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_AQ;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_A_CY;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_A_XOR;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_B;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_B1;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_B2;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_B3;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_B4;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_B5;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_B6;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_BO5;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_BO6;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_BQ;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_B_CY;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_B_XOR;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_C;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_C1;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_C2;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_C3;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_C4;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_C5;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_C5Q;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_C6;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_CLK;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_CMUX;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_CO5;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_CO6;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_CQ;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_C_CY;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_C_XOR;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_D;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_D1;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_D2;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_D3;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_D4;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_D5;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_D5Q;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_D6;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_DMUX;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_DO5;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_DO6;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_DQ;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_D_CY;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_D_XOR;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_A;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_A1;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_A2;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_A3;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_A4;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_A5;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_A6;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_AO5;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_AO6;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_AQ;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_A_CY;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_A_XOR;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_B;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_B1;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_B2;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_B3;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_B4;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_B5;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_B5Q;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_B6;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_BMUX;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_BO5;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_BO6;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_BQ;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_B_CY;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_B_XOR;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_C;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_C1;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_C2;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_C3;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_C4;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_C5;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_C5Q;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_C6;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_CLK;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_CMUX;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_CO5;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_CO6;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_CQ;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_C_CY;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_C_XOR;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_D;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_D1;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_D2;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_D3;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_D4;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_D5;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_D6;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_DO5;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_DO6;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_DQ;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_D_CY;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_D_XOR;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_A;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_A1;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_A2;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_A3;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_A4;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_A5;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_A5Q;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_A6;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_AMUX;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_AO5;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_AO6;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_AQ;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_A_CY;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_A_XOR;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_B;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_B1;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_B2;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_B3;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_B4;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_B5;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_B6;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_BMUX;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_BO5;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_BO6;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_BQ;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_BX;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_B_CY;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_B_XOR;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_C;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_C1;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_C2;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_C3;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_C4;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_C5;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_C6;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_CLK;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_CMUX;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_CO5;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_CO6;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_C_CY;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_C_XOR;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_D;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_D1;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_D2;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_D3;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_D4;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_D5;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_D6;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_DO5;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_DO6;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_D_CY;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_D_XOR;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_SR;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_A;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_A1;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_A2;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_A3;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_A4;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_A5;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_A6;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_AO5;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_AO6;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_AQ;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_A_CY;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_A_XOR;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_B;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_B1;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_B2;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_B3;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_B4;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_B5;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_B5Q;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_B6;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_BMUX;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_BO5;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_BO6;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_BQ;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_B_CY;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_B_XOR;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_C;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_C1;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_C2;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_C3;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_C4;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_C5;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_C6;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_CLK;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_CO5;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_CO6;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_CQ;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_C_CY;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_C_XOR;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_D;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_D1;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_D2;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_D3;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_D4;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_D5;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_D6;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_DO5;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_DO6;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_DQ;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_D_CY;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_D_XOR;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_A;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_A1;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_A2;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_A3;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_A4;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_A5;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_A6;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_AO5;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_AO6;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_AQ;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_A_CY;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_A_XOR;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_B;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_B1;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_B2;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_B3;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_B4;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_B5;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_B5Q;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_B6;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_BMUX;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_BO5;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_BO6;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_BQ;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_B_CY;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_B_XOR;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_C;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_C1;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_C2;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_C3;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_C4;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_C5;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_C5Q;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_C6;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_CLK;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_CMUX;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_CO5;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_CO6;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_CQ;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_C_CY;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_C_XOR;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_D;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_D1;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_D2;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_D3;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_D4;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_D5;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_D5Q;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_D6;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_DMUX;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_DO5;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_DO6;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_DQ;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_D_CY;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_D_XOR;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_A;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_A1;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_A2;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_A3;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_A4;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_A5;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_A6;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_AO5;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_AO6;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_AQ;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_A_CY;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_A_XOR;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_B;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_B1;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_B2;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_B3;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_B4;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_B5;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_B6;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_BO5;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_BO6;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_BQ;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_B_CY;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_B_XOR;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_C;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_C1;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_C2;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_C3;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_C4;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_C5;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_C6;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_CLK;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_CO5;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_CO6;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_CQ;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_C_CY;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_C_XOR;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_D;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_D1;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_D2;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_D3;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_D4;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_D5;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_D6;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_DO5;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_DO6;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_DQ;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_D_CY;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_D_XOR;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_A;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_A1;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_A2;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_A3;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_A4;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_A5;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_A6;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_AMUX;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_AO5;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_AO6;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_AQ;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_AX;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_A_CY;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_A_XOR;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_B;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_B1;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_B2;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_B3;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_B4;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_B5;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_B6;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_BMUX;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_BO5;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_BO6;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_B_CY;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_B_XOR;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_C;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_C1;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_C2;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_C3;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_C4;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_C5;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_C6;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_CE;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_CLK;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_CO5;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_CO6;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_C_CY;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_C_XOR;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_D;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_D1;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_D2;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_D3;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_D4;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_D5;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_D6;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_DO5;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_DO6;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_D_CY;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_D_XOR;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_A;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_A1;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_A2;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_A3;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_A4;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_A5;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_A6;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_AO5;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_AO6;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_AQ;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_A_CY;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_A_XOR;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_B;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_B1;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_B2;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_B3;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_B4;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_B5;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_B6;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_BO5;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_BO6;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_BQ;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_B_CY;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_B_XOR;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_C;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_C1;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_C2;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_C3;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_C4;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_C5;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_C5Q;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_C6;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_CLK;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_CMUX;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_CO5;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_CO6;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_CQ;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_C_CY;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_C_XOR;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_D;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_D1;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_D2;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_D3;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_D4;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_D5;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_D5Q;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_D6;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_DMUX;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_DO5;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_DO6;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_DQ;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_D_CY;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_D_XOR;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_A;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_A1;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_A2;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_A3;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_A4;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_A5;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_A6;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_AMUX;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_AO5;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_AO6;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_AQ;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_AX;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_A_CY;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_A_XOR;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_B;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_B1;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_B2;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_B3;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_B4;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_B5;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_B6;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_BMUX;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_BO5;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_BO6;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_B_CY;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_B_XOR;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_C;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_C1;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_C2;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_C3;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_C4;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_C5;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_C6;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_CLK;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_CO5;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_CO6;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_C_CY;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_C_XOR;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_D;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_D1;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_D2;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_D3;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_D4;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_D5;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_D6;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_DO5;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_DO6;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_D_CY;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_D_XOR;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_SR;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_A;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_A1;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_A2;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_A3;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_A4;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_A5;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_A5Q;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_A6;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_AMUX;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_AO5;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_AO6;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_AQ;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_AX;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_A_CY;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_A_XOR;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_B;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_B1;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_B2;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_B3;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_B4;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_B5;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_B6;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_BO5;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_BO6;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_BQ;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_B_CY;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_B_XOR;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_C;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_C1;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_C2;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_C3;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_C4;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_C5;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_C6;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_CLK;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_CO5;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_CO6;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_CQ;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_C_CY;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_C_XOR;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_D;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_D1;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_D2;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_D3;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_D4;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_D5;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_D6;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_DO5;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_DO6;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_DQ;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_D_CY;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_D_XOR;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_A;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_A1;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_A2;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_A3;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_A4;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_A5;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_A6;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_AO5;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_AO6;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_AQ;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_A_CY;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_A_XOR;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_B;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_B1;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_B2;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_B3;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_B4;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_B5;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_B6;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_BO5;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_BO6;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_BQ;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_B_CY;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_B_XOR;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_C;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_C1;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_C2;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_C3;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_C4;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_C5;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_C5Q;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_C6;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_CLK;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_CMUX;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_CO5;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_CO6;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_CQ;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_C_CY;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_C_XOR;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_D;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_D1;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_D2;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_D3;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_D4;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_D5;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_D6;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_DO5;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_DO6;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_DQ;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_D_CY;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_D_XOR;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_A;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_A1;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_A2;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_A3;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_A4;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_A5;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_A6;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_AO5;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_AO6;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_AQ;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_A_CY;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_A_XOR;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_B;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_B1;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_B2;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_B3;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_B4;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_B5;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_B5Q;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_B6;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_BMUX;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_BO5;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_BO6;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_BQ;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_B_CY;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_B_XOR;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_C;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_C1;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_C2;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_C3;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_C4;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_C5;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_C5Q;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_C6;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_CLK;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_CMUX;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_CO5;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_CO6;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_CQ;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_C_CY;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_C_XOR;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_D;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_D1;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_D2;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_D3;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_D4;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_D5;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_D6;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_DO5;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_DO6;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_DQ;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_D_CY;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_D_XOR;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_A;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_A1;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_A2;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_A3;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_A4;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_A5;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_A5Q;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_A6;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_AMUX;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_AO5;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_AO6;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_AQ;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_AX;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_A_CY;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_A_XOR;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_B;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_B1;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_B2;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_B3;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_B4;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_B5;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_B6;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_BO5;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_BO6;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_BQ;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_B_CY;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_B_XOR;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_C;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_C1;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_C2;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_C3;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_C4;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_C5;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_C6;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_CLK;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_CO5;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_CO6;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_CQ;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_C_CY;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_C_XOR;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_D;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_D1;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_D2;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_D3;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_D4;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_D5;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_D6;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_DMUX;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_DO5;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_DO6;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_D_CY;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_D_XOR;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_A;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_A1;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_A2;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_A3;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_A4;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_A5;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_A6;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_AO5;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_AO6;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_AQ;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_A_CY;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_A_XOR;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_B;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_B1;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_B2;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_B3;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_B4;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_B5;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_B6;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_BO5;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_BO6;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_BQ;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_B_CY;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_B_XOR;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_C;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_C1;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_C2;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_C3;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_C4;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_C5;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_C6;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_CLK;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_CO5;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_CO6;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_C_CY;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_C_XOR;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_D;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_D1;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_D2;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_D3;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_D4;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_D5;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_D6;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_DMUX;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_DO5;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_DO6;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_D_CY;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_D_XOR;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_A;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_A1;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_A2;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_A3;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_A4;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_A5;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_A6;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_AMUX;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_AO5;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_AO6;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_AQ;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_A_CY;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_A_XOR;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_B;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_B1;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_B2;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_B3;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_B4;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_B5;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_B6;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_BMUX;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_BO5;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_BO6;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_B_CY;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_B_XOR;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_C;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_C1;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_C2;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_C3;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_C4;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_C5;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_C6;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_CLK;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_CO5;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_CO6;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_C_CY;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_C_XOR;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_D;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_D1;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_D2;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_D3;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_D4;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_D5;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_D6;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_DO5;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_DO6;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_D_CY;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_D_XOR;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_A;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_A1;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_A2;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_A3;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_A4;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_A5;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_A6;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_AO5;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_AO6;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_A_CY;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_A_XOR;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_B;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_B1;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_B2;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_B3;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_B4;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_B5;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_B6;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_BO5;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_BO6;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_B_CY;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_B_XOR;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_C;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_C1;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_C2;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_C3;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_C4;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_C5;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_C6;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_CO5;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_CO6;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_C_CY;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_C_XOR;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_D;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_D1;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_D2;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_D3;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_D4;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_D5;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_D6;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_DO5;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_DO6;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_D_CY;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_D_XOR;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_A;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_A1;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_A2;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_A3;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_A4;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_A5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_A6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_AO5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_AO6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_A_CY;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_A_XOR;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_B;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_B1;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_B2;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_B3;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_B4;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_B5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_B6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_BO5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_BO6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_B_CY;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_B_XOR;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_C;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_C1;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_C2;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_C3;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_C4;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_C5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_C6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_CO5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_CO6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_C_CY;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_C_XOR;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_D;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_D1;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_D2;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_D3;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_D4;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_D5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_D6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_DO5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_DO6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_D_CY;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_D_XOR;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_A;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_A1;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_A2;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_A3;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_A4;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_A5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_A6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_AO5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_AO6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_A_CY;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_A_XOR;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_B;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_B1;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_B2;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_B3;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_B4;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_B5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_B6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_BO5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_BO6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_B_CY;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_B_XOR;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_C;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_C1;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_C2;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_C3;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_C4;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_C5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_C6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_CO5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_CO6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_C_CY;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_C_XOR;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_D;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_D1;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_D2;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_D3;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_D4;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_D5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_D6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_DO5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_DO6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_D_CY;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_D_XOR;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_A;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_A1;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_A2;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_A3;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_A4;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_A5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_A6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_AMUX;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_AO5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_AO6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_AQ;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_A_CY;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_A_XOR;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_B;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_B1;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_B2;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_B3;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_B4;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_B5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_B6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_BMUX;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_BO5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_BO6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_B_CY;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_B_XOR;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_C;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_C1;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_C2;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_C3;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_C4;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_C5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_C6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_CLK;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_CO5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_CO6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_C_CY;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_C_XOR;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_D;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_D1;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_D2;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_D3;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_D4;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_D5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_D6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_DO5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_DO6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_D_CY;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_D_XOR;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_A;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_A1;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_A2;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_A3;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_A4;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_A5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_A6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_AO5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_AO6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_AQ;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_A_CY;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_A_XOR;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_B;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_B1;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_B2;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_B3;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_B4;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_B5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_B6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_BO5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_BO6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_B_CY;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_B_XOR;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_C;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_C1;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_C2;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_C3;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_C4;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_C5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_C6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_CLK;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_CO5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_CO6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_C_CY;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_C_XOR;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_D;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_D1;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_D2;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_D3;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_D4;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_D5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_D6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_DO5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_DO6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_D_CY;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_D_XOR;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_A;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_A1;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_A2;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_A3;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_A4;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_A5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_A6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_AMUX;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_AO5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_AO6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_AQ;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_AX;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_A_CY;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_A_XOR;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_B;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_B1;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_B2;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_B3;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_B4;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_B5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_B6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_BMUX;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_BO5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_BO6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_B_CY;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_B_XOR;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_C;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_C1;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_C2;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_C3;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_C4;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_C5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_C6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_CE;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_CLK;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_CMUX;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_CO5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_CO6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_C_CY;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_C_XOR;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_D;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_D1;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_D2;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_D3;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_D4;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_D5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_D6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_DMUX;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_DO5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_DO6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_D_CY;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X12Y143_D_XOR;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_A;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_A1;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_A2;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_A3;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_A4;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_A5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_A6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_AO5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_AO6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_A_CY;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_A_XOR;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_B;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_B1;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_B2;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_B3;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_B4;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_B5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_B6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_BO5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_BO6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_B_CY;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_B_XOR;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_C;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_C1;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_C2;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_C3;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_C4;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_C5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_C6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_CO5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_CO6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_C_CY;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_C_XOR;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_D;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_D1;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_D2;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_D3;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_D4;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_D5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_D6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_DO5;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_DO6;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_D_CY;
  wire [0:0] CLBLM_L_X10Y143_SLICE_X13Y143_D_XOR;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_A;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_A1;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_A2;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_A3;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_A4;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_A5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_A6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_AMUX;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_AO5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_AO6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_A_CY;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_A_XOR;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_B;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_B1;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_B2;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_B3;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_B4;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_B5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_B6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_BO5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_BO6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_B_CY;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_B_XOR;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_C;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_C1;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_C2;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_C3;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_C4;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_C5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_C6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_CO5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_CO6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_C_CY;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_C_XOR;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_D;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_D1;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_D2;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_D3;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_D4;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_D5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_D6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_DO5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_DO6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_D_CY;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_D_XOR;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_A;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_A1;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_A2;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_A3;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_A4;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_A5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_A6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_AO5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_AO6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_A_CY;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_A_XOR;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_B;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_B1;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_B2;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_B3;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_B4;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_B5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_B6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_BMUX;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_BO5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_BO6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_B_CY;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_B_XOR;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_C;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_C1;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_C2;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_C3;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_C4;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_C5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_C6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_CO5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_CO6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_C_CY;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_C_XOR;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_D;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_D1;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_D2;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_D3;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_D4;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_D5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_D6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_DMUX;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_DO5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_DO6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_D_CY;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_D_XOR;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_A;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_A1;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_A2;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_A3;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_A4;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_A5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_A6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_AMUX;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_AO5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_AO6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_AQ;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_AX;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_A_CY;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_A_XOR;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_B;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_B1;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_B2;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_B3;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_B4;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_B5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_B6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_BO5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_BO6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_B_CY;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_B_XOR;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_C;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_C1;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_C2;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_C3;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_C4;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_C5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_C6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_CE;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_CLK;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_CMUX;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_CO5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_CO6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_C_CY;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_C_XOR;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_D;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_D1;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_D2;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_D3;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_D4;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_D5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_D6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_DO5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_DO6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_D_CY;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_D_XOR;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_A;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_A1;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_A2;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_A3;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_A4;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_A5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_A6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_AMUX;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_AO5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_AO6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_A_CY;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_A_XOR;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_B;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_B1;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_B2;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_B3;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_B4;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_B5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_B6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_BMUX;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_BO5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_BO6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_B_CY;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_B_XOR;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_C;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_C1;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_C2;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_C3;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_C4;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_C5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_C6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_CO5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_CO6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_C_CY;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_C_XOR;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_D;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_D1;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_D2;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_D3;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_D4;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_D5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_D6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_DO5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_DO6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_D_CY;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_D_XOR;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_A;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_A1;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_A2;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_A3;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_A4;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_A5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_A6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_AMUX;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_AO5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_AO6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_AQ;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_AX;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_A_CY;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_A_XOR;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_B;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_B1;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_B2;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_B3;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_B4;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_B5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_B6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_BMUX;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_BO5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_BO6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_B_CY;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_B_XOR;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_C;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_C1;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_C2;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_C3;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_C4;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_C5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_C6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_CLK;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_CMUX;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_CO5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_CO6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_C_CY;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_C_XOR;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_D;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_D1;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_D2;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_D3;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_D4;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_D5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_D6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_DO5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_DO6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_D_CY;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_D_XOR;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_SR;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_A;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_A1;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_A2;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_A3;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_A4;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_A5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_A6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_AO5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_AO6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_AQ;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_A_CY;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_A_XOR;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_B;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_B1;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_B2;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_B3;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_B4;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_B5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_B6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_BMUX;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_BO5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_BO6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_B_CY;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_B_XOR;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_C;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_C1;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_C2;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_C3;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_C4;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_C5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_C6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_CLK;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_CO5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_CO6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_C_CY;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_C_XOR;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_D;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_D1;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_D2;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_D3;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_D4;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_D5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_D6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_DMUX;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_DO5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_DO6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_D_CY;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_D_XOR;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_SR;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_A;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_A1;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_A2;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_A3;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_A4;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_A5;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_A6;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_AO5;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_AO6;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_AQ;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_A_CY;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_A_XOR;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_B;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_B1;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_B2;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_B3;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_B4;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_B5;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_B5Q;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_B6;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_BMUX;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_BO5;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_BO6;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_BQ;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_B_CY;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_B_XOR;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_C;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_C1;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_C2;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_C3;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_C4;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_C5;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_C5Q;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_C6;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_CLK;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_CMUX;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_CO5;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_CO6;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_CQ;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_C_CY;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_C_XOR;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_D;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_D1;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_D2;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_D3;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_D4;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_D5;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_D6;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_DMUX;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_DO5;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_DO6;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_D_CY;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_D_XOR;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_A;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_A1;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_A2;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_A3;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_A4;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_A5;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_A5Q;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_A6;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_AMUX;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_AO5;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_AO6;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_AQ;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_A_CY;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_A_XOR;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_B;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_B1;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_B2;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_B3;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_B4;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_B5;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_B5Q;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_B6;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_BMUX;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_BO5;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_BO6;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_BQ;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_B_CY;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_B_XOR;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_C;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_C1;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_C2;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_C3;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_C4;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_C5;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_C6;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_CLK;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_CO5;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_CO6;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_CQ;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_C_CY;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_C_XOR;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_D;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_D1;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_D2;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_D3;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_D4;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_D5;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_D6;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_DO5;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_DO6;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_DQ;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_D_CY;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_D_XOR;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_A;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_A1;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_A2;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_A3;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_A4;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_A5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_A5Q;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_A6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_AMUX;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_AO5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_AO6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_AQ;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_A_CY;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_A_XOR;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_B;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_B1;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_B2;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_B3;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_B4;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_B5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_B6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_BMUX;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_BO5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_BO6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_B_CY;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_B_XOR;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_C;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_C1;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_C2;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_C3;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_C4;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_C5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_C6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_CLK;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_CO5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_CO6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_C_CY;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_C_XOR;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_D;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_D1;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_D2;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_D3;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_D4;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_D5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_D6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_DO5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_DO6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_D_CY;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_D_XOR;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_SR;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_A;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_A1;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_A2;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_A3;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_A4;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_A5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_A6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_AMUX;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_AO5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_AO6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_AQ;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_AX;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_A_CY;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_A_XOR;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_B;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_B1;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_B2;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_B3;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_B4;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_B5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_B6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_BMUX;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_BO5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_BO6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_B_CY;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_B_XOR;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_C;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_C1;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_C2;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_C3;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_C4;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_C5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_C6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_CLK;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_CO5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_CO6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_C_CY;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_C_XOR;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_D;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_D1;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_D2;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_D3;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_D4;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_D5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_D6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_DO5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_DO6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_D_CY;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_D_XOR;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_SR;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_A;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_A1;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_A2;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_A3;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_A4;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_A5;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_A5Q;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_A6;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_AMUX;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_AO5;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_AO6;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_AQ;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_A_CY;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_A_XOR;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_B;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_B1;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_B2;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_B3;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_B4;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_B5;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_B5Q;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_B6;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_BMUX;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_BO5;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_BO6;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_BQ;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_B_CY;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_B_XOR;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_C;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_C1;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_C2;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_C3;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_C4;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_C5;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_C6;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_CLK;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_CO5;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_CO6;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_CQ;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_C_CY;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_C_XOR;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_D;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_D1;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_D2;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_D3;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_D4;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_D5;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_D6;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_DO5;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_DO6;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_DQ;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_D_CY;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_D_XOR;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_A;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_A1;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_A2;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_A3;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_A4;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_A5;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_A5Q;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_A6;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_AMUX;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_AO5;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_AO6;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_AQ;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_AX;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_A_CY;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_A_XOR;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_B;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_B1;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_B2;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_B3;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_B4;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_B5;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_B6;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_BMUX;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_BO5;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_BO6;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_B_CY;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_B_XOR;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_C;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_C1;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_C2;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_C3;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_C4;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_C5;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_C6;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_CLK;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_CO5;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_CO6;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_C_CY;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_C_XOR;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_D;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_D1;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_D2;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_D3;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_D4;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_D5;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_D6;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_DO5;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_DO6;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_D_CY;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_D_XOR;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_SR;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_A;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_A1;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_A2;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_A3;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_A4;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_A5;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_A5Q;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_A6;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_AMUX;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_AO5;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_AO6;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_AQ;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_A_CY;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_A_XOR;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_B;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_B1;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_B2;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_B3;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_B4;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_B5;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_B6;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_BO5;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_BO6;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_BQ;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_B_CY;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_B_XOR;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_C;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_C1;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_C2;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_C3;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_C4;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_C5;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_C6;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_CLK;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_CO5;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_CO6;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_CQ;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_C_CY;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_C_XOR;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_D;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_D1;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_D2;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_D3;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_D4;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_D5;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_D6;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_DMUX;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_DO5;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_DO6;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_D_CY;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_D_XOR;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_A;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_A1;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_A2;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_A3;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_A4;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_A5;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_A5Q;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_A6;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_AMUX;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_AO5;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_AO6;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_AQ;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_A_CY;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_A_XOR;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_B;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_B1;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_B2;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_B3;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_B4;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_B5;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_B5Q;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_B6;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_BMUX;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_BO5;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_BO6;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_BQ;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_BX;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_B_CY;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_B_XOR;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_C;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_C1;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_C2;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_C3;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_C4;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_C5;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_C5Q;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_C6;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_CLK;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_CMUX;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_CO5;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_CO6;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_CQ;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_C_CY;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_C_XOR;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_D;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_D1;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_D2;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_D3;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_D4;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_D5;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_D6;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_DMUX;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_DO5;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_DO6;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_D_CY;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_D_XOR;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_A;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_A1;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_A2;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_A3;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_A4;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_A5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_A6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_AMUX;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_AO5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_AO6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_AQ;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_AX;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_A_CY;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_A_XOR;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_B;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_B1;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_B2;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_B3;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_B4;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_B5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_B6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_BO5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_BO6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_B_CY;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_B_XOR;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_C;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_C1;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_C2;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_C3;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_C4;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_C5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_C6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_CLK;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_CO5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_CO6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_C_CY;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_C_XOR;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_D;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_D1;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_D2;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_D3;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_D4;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_D5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_D6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_DO5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_DO6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_D_CY;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_D_XOR;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_SR;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_A;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_A1;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_A2;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_A3;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_A4;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_A5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_A6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_AO5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_AO6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_AQ;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_A_CY;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_A_XOR;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_B;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_B1;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_B2;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_B3;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_B4;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_B5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_B6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_BMUX;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_BO5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_BO6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_B_CY;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_B_XOR;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_C;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_C1;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_C2;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_C3;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_C4;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_C5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_C6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_CLK;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_CO5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_CO6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_C_CY;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_C_XOR;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_D;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_D1;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_D2;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_D3;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_D4;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_D5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_D6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_DMUX;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_DO5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_DO6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_D_CY;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_D_XOR;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_A;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_A1;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_A2;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_A3;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_A4;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_A5;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_A6;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_AO5;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_AO6;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_AQ;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_A_CY;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_A_XOR;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_B;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_B1;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_B2;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_B3;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_B4;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_B5;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_B6;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_BO5;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_BO6;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_BQ;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_B_CY;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_B_XOR;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_C;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_C1;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_C2;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_C3;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_C4;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_C5;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_C6;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_CLK;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_CO5;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_CO6;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_CQ;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_C_CY;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_C_XOR;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_D;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_D1;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_D2;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_D3;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_D4;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_D5;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_D6;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_DO5;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_DO6;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_D_CY;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_D_XOR;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_A;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_A1;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_A2;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_A3;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_A4;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_A5;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_A6;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_AO5;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_AO6;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_AQ;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_A_CY;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_A_XOR;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_B;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_B1;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_B2;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_B3;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_B4;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_B5;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_B6;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_BO5;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_BO6;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_BQ;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_B_CY;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_B_XOR;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_C;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_C1;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_C2;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_C3;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_C4;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_C5;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_C6;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_CLK;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_CMUX;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_CO5;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_CO6;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_C_CY;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_C_XOR;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_D;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_D1;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_D2;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_D3;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_D4;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_D5;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_D6;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_DO5;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_DO6;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_D_CY;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_D_XOR;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_A;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_A1;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_A2;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_A3;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_A4;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_A5;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_A6;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_AO5;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_AO6;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_AQ;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_A_CY;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_A_XOR;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_B;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_B1;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_B2;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_B3;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_B4;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_B5;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_B6;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_BO5;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_BO6;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_BQ;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_B_CY;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_B_XOR;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_C;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_C1;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_C2;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_C3;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_C4;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_C5;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_C6;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_CLK;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_CO5;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_CO6;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_CQ;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_C_CY;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_C_XOR;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_D;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_D1;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_D2;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_D3;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_D4;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_D5;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_D6;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_DMUX;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_DO5;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_DO6;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_D_CY;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_D_XOR;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_A;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_A1;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_A2;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_A3;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_A4;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_A5;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_A6;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_AO5;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_AO6;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_AQ;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_A_CY;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_A_XOR;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_B;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_B1;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_B2;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_B3;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_B4;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_B5;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_B6;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_BO5;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_BO6;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_B_CY;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_B_XOR;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_C;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_C1;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_C2;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_C3;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_C4;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_C5;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_C6;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_CLK;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_CO5;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_CO6;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_C_CY;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_C_XOR;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_D;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_D1;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_D2;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_D3;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_D4;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_D5;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_D6;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_DO5;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_DO6;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_D_CY;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_D_XOR;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_A;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_A1;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_A2;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_A3;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_A4;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_A5;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_A6;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_AO5;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_AO6;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_A_CY;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_A_XOR;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_B;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_B1;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_B2;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_B3;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_B4;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_B5;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_B6;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_BO5;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_BO6;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_B_CY;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_B_XOR;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_C;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_C1;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_C2;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_C3;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_C4;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_C5;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_C6;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_CO5;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_CO6;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_C_CY;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_C_XOR;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_D;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_D1;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_D2;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_D3;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_D4;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_D5;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_D6;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_DO5;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_DO6;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_D_CY;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_D_XOR;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_A;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_A1;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_A2;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_A3;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_A4;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_A5;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_A6;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_AO5;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_AO6;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_A_CY;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_A_XOR;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_B;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_B1;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_B2;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_B3;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_B4;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_B5;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_B6;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_BO5;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_BO6;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_B_CY;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_B_XOR;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_C;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_C1;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_C2;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_C3;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_C4;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_C5;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_C6;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_CO5;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_CO6;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_C_CY;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_C_XOR;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_D;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_D1;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_D2;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_D3;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_D4;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_D5;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_D6;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_DO5;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_DO6;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_D_CY;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_D_XOR;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_A;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_A1;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_A2;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_A3;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_A4;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_A5;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_A6;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_AMUX;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_AO5;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_AO6;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_A_CY;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_A_XOR;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_B;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_B1;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_B2;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_B3;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_B4;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_B5;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_B6;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_BO5;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_BO6;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_B_CY;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_B_XOR;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_C;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_C1;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_C2;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_C3;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_C4;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_C5;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_C6;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_CO5;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_CO6;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_C_CY;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_C_XOR;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_D;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_D1;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_D2;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_D3;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_D4;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_D5;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_D6;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_DO5;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_DO6;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_D_CY;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X16Y144_D_XOR;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_A;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_A1;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_A2;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_A3;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_A4;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_A5;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_A6;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_AO5;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_AO6;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_A_CY;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_A_XOR;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_B;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_B1;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_B2;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_B3;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_B4;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_B5;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_B6;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_BO5;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_BO6;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_B_CY;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_B_XOR;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_C;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_C1;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_C2;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_C3;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_C4;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_C5;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_C6;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_CO5;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_CO6;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_C_CY;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_C_XOR;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_D;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_D1;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_D2;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_D3;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_D4;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_D5;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_D6;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_DO5;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_DO6;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_D_CY;
  wire [0:0] CLBLM_L_X12Y144_SLICE_X17Y144_D_XOR;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_A;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_A1;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_A2;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_A3;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_A4;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_A5;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_A6;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_AMUX;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_AO5;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_AO6;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_A_CY;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_A_XOR;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_B;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_B1;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_B2;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_B3;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_B4;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_B5;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_B6;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_BO5;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_BO6;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_B_CY;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_B_XOR;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_C;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_C1;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_C2;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_C3;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_C4;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_C5;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_C6;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_CO5;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_CO6;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_C_CY;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_C_XOR;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_D;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_D1;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_D2;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_D3;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_D4;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_D5;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_D6;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_DMUX;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_DO5;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_DO6;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_D_CY;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X16Y145_D_XOR;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_A;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_A1;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_A2;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_A3;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_A4;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_A5;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_A6;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_AO5;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_A_CY;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_A_XOR;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_B;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_B1;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_B2;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_B3;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_B4;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_B5;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_B6;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_BO5;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_BO6;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_B_CY;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_B_XOR;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_C;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_C1;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_C2;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_C3;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_C4;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_C5;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_C6;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_CMUX;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_CO5;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_CO6;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_C_CY;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_C_XOR;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_D;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_D1;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_D2;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_D3;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_D4;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_D5;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_D6;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_DO5;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_DO6;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_D_CY;
  wire [0:0] CLBLM_L_X12Y145_SLICE_X17Y145_D_XOR;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_A;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_A1;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_A2;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_A3;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_A4;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_A5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_A6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_AO5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_AO6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_A_CY;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_A_XOR;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_B;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_B1;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_B2;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_B3;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_B4;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_B5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_B6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_BO5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_BO6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_B_CY;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_B_XOR;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_C;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_C1;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_C2;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_C3;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_C4;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_C5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_C6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_CO5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_CO6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_C_CY;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_C_XOR;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_D;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_D1;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_D2;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_D3;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_D4;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_D5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_D6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_DO5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_DO6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_D_CY;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_D_XOR;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_A;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_A1;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_A2;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_A3;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_A4;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_A5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_A6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_AO5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_AO6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_A_CY;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_A_XOR;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_B;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_B1;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_B2;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_B3;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_B4;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_B5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_B6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_BO5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_BO6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_B_CY;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_B_XOR;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_C;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_C1;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_C2;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_C3;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_C4;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_C5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_C6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_CO5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_CO6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_C_CY;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_C_XOR;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_D;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_D1;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_D2;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_D3;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_D4;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_D5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_D6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_DO5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_DO6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_D_CY;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_D_XOR;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_A;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_A1;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_A2;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_A3;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_A4;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_A5;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_A6;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_AO5;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_AO6;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_AQ;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_A_CY;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_A_XOR;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_B;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_B1;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_B2;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_B3;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_B4;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_B5;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_B6;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_BO5;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_BO6;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_BQ;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_B_CY;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_B_XOR;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_C;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_C1;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_C2;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_C3;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_C4;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_C5;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_C6;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_CLK;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_CO5;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_CO6;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_C_CY;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_C_XOR;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_D;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_D1;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_D2;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_D3;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_D4;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_D5;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_D6;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_DMUX;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_DO5;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_DO6;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_D_CY;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_D_XOR;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_A;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_A1;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_A2;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_A3;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_A4;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_A5;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_A6;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_AO5;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_AO6;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_A_CY;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_A_XOR;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_B;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_B1;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_B2;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_B3;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_B4;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_B5;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_B6;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_BO5;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_BO6;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_B_CY;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_B_XOR;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_C;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_C1;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_C2;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_C3;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_C4;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_C5;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_C6;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_CO5;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_CO6;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_C_CY;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_C_XOR;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_D;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_D1;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_D2;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_D3;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_D4;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_D5;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_D6;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_DO5;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_DO6;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_D_CY;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_D_XOR;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_A;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_A1;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_A2;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_A3;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_A4;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_A5;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_A6;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_AO5;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_AO6;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_AQ;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_A_CY;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_A_XOR;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_B;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_B1;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_B2;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_B3;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_B4;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_B5;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_B6;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_BO5;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_BO6;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_BQ;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_B_CY;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_B_XOR;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_C;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_C1;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_C2;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_C3;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_C4;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_C5;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_C6;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_CLK;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_CMUX;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_CO5;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_CO6;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_C_CY;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_C_XOR;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_D;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_D1;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_D2;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_D3;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_D4;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_D5;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_D6;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_DO5;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_DO6;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_D_CY;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_D_XOR;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_A;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_A1;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_A2;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_A3;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_A4;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_A5;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_A6;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_AO5;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_AO6;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_A_CY;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_A_XOR;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_B;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_B1;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_B2;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_B3;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_B4;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_B5;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_B6;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_BO5;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_BO6;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_B_CY;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_B_XOR;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_C;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_C1;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_C2;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_C3;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_C4;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_C5;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_C6;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_CO5;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_CO6;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_C_CY;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_C_XOR;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_D;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_D1;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_D2;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_D3;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_D4;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_D5;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_D6;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_DO5;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_DO6;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_D_CY;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_D_XOR;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_A;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_A1;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_A2;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_A3;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_A4;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_A5;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_A5Q;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_A6;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_AMUX;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_AO5;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_AO6;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_AQ;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_A_CY;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_A_XOR;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_B;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_B1;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_B2;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_B3;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_B4;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_B5;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_B6;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_BO5;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_BO6;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_B_CY;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_B_XOR;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_C;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_C1;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_C2;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_C3;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_C4;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_C5;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_C6;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_CLK;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_CO5;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_CO6;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_C_CY;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_C_XOR;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_D;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_D1;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_D2;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_D3;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_D4;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_D5;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_D6;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_DO5;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_DO6;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_D_CY;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_D_XOR;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_SR;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_A;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_A1;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_A2;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_A3;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_A4;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_A5;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_A6;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_AO5;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_AO6;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_A_CY;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_A_XOR;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_B;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_B1;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_B2;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_B3;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_B4;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_B5;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_B6;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_BO5;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_BO6;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_B_CY;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_B_XOR;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_C;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_C1;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_C2;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_C3;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_C4;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_C5;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_C6;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_CO5;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_CO6;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_C_CY;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_C_XOR;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_D;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_D1;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_D2;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_D3;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_D4;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_D5;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_D6;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_DO5;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_DO6;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_D_CY;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_D_XOR;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_A;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_A1;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_A2;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_A3;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_A4;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_A5;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_A6;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_AO5;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_AO6;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_A_CY;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_A_XOR;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_B;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_B1;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_B2;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_B3;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_B4;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_B5;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_B6;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_BO5;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_BO6;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_BQ;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_B_CY;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_B_XOR;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_C;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_C1;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_C2;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_C3;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_C4;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_C5;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_C6;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_CLK;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_CO5;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_CO6;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_CQ;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_C_CY;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_C_XOR;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_D;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_D1;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_D2;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_D3;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_D4;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_D5;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_D6;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_DO5;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_DO6;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_D_CY;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_D_XOR;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_A;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_A1;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_A2;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_A3;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_A4;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_A5;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_A6;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_AO5;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_AO6;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_A_CY;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_A_XOR;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_B;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_B1;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_B2;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_B3;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_B4;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_B5;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_B6;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_BO5;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_BO6;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_B_CY;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_B_XOR;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_C;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_C1;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_C2;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_C3;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_C4;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_C5;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_C6;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_CO5;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_CO6;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_C_CY;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_C_XOR;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_D;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_D1;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_D2;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_D3;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_D4;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_D5;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_D6;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_DO5;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_DO6;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_D_CY;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_D_XOR;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_A;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_A1;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_A2;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_A3;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_A4;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_A5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_A5Q;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_A6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_AMUX;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_AO5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_AO6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_AQ;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_AX;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_A_CY;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_A_XOR;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_B;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_B1;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_B2;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_B3;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_B4;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_B5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_B6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_BMUX;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_BO5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_BO6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_B_CY;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_B_XOR;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_C;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_C1;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_C2;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_C3;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_C4;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_C5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_C5Q;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_C6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_CLK;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_CMUX;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_CO5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_CO6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_CQ;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_C_CY;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_C_XOR;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_D;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_D1;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_D2;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_D3;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_D4;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_D5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_D6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_DMUX;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_DO5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_DO6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_D_CY;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_D_XOR;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_SR;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_A;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_A1;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_A2;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_A3;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_A4;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_A5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_A6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_AO5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_AO6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_AQ;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_A_CY;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_A_XOR;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_B;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_B1;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_B2;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_B3;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_B4;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_B5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_B6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_BO5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_BO6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_BQ;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_B_CY;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_B_XOR;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_C;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_C1;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_C2;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_C3;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_C4;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_C5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_C5Q;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_C6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_CLK;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_CMUX;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_CO5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_CO6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_CQ;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_C_CY;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_C_XOR;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_D;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_D1;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_D2;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_D3;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_D4;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_D5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_D6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_DO5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_DO6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_D_CY;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_D_XOR;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_A;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_A1;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_A2;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_A3;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_A4;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_A5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_A6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_AO5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_AO6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_A_CY;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_A_XOR;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_B;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_B1;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_B2;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_B3;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_B4;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_B5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_B6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_BO5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_BO6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_BQ;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_B_CY;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_B_XOR;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_C;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_C1;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_C2;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_C3;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_C4;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_C5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_C6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_CLK;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_CO5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_CO6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_CQ;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_C_CY;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_C_XOR;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_D;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_D1;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_D2;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_D3;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_D4;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_D5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_D6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_DO5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_DO6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_DQ;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_D_CY;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_D_XOR;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_A;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_A1;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_A2;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_A3;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_A4;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_A5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_A5Q;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_A6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_AMUX;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_AO5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_AO6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_AQ;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_AX;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_A_CY;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_A_XOR;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_B;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_B1;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_B2;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_B3;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_B4;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_B5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_B6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_BO5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_BO6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_BQ;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_B_CY;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_B_XOR;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_C;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_C1;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_C2;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_C3;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_C4;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_C5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_C6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_CLK;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_CO5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_CO6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_CQ;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_C_CY;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_C_XOR;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_D;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_D1;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_D2;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_D3;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_D4;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_D5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_D6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_DO5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_DO6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_DQ;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_D_CY;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_D_XOR;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_A;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_A1;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_A2;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_A3;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_A4;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_A5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_A5Q;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_A6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_AMUX;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_AO5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_AO6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_AQ;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_A_CY;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_A_XOR;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_B;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_B1;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_B2;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_B3;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_B4;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_B5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_B5Q;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_B6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_BMUX;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_BO5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_BO6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_BQ;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_B_CY;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_B_XOR;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_C;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_C1;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_C2;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_C3;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_C4;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_C5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_C6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_CLK;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_CMUX;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_CO5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_CO6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_C_CY;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_C_XOR;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_D;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_D1;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_D2;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_D3;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_D4;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_D5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_D6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_DO5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_DO6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_D_CY;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_D_XOR;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_SR;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_A;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_A1;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_A2;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_A3;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_A4;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_A5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_A5Q;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_A6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_AMUX;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_AO5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_AO6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_AQ;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_A_CY;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_A_XOR;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_B;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_B1;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_B2;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_B3;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_B4;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_B5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_B6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_BO5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_BO6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_B_CY;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_B_XOR;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_C;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_C1;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_C2;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_C3;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_C4;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_C5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_C6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_CLK;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_CO5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_CO6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_C_CY;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_C_XOR;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_D;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_D1;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_D2;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_D3;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_D4;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_D5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_D6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_DO5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_DO6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_D_CY;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_D_XOR;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_SR;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_A;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_A1;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_A2;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_A3;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_A4;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_A5;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_A6;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_AMUX;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_AO5;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_AO6;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_AQ;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_AX;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_A_CY;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_A_XOR;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_B;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_B1;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_B2;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_B3;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_B4;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_B5;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_B6;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_BMUX;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_BO5;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_BO6;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_BQ;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_BX;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_B_CY;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_B_XOR;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_C;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_C1;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_C2;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_C3;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_C4;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_C5;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_C6;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_CLK;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_CMUX;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_CO5;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_CO6;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_C_CY;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_C_XOR;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_D;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_D1;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_D2;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_D3;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_D4;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_D5;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_D6;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_DO5;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_DO6;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_D_CY;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_D_XOR;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X10Y145_SR;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_A;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_A1;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_A2;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_A3;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_A4;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_A5;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_A6;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_AMUX;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_AO5;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_AO6;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_AQ;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_AX;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_A_CY;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_A_XOR;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_B;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_B1;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_B2;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_B3;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_B4;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_B5;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_B6;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_BMUX;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_BO5;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_BO6;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_B_CY;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_B_XOR;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_C;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_C1;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_C2;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_C3;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_C4;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_C5;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_C6;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_CLK;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_CO5;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_CO6;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_C_CY;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_C_XOR;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_D;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_D1;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_D2;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_D3;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_D4;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_D5;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_D6;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_DO5;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_DO6;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_D_CY;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_D_XOR;
  wire [0:0] CLBLM_L_X8Y145_SLICE_X11Y145_SR;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_A;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_A1;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_A2;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_A3;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_A4;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_A5;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_A5Q;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_A6;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_AMUX;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_AO5;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_AO6;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_AQ;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_A_CY;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_A_XOR;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_B;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_B1;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_B2;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_B3;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_B4;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_B5;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_B6;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_BO5;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_BO6;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_BQ;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_B_CY;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_B_XOR;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_C;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_C1;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_C2;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_C3;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_C4;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_C5;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_C5Q;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_C6;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_CLK;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_CMUX;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_CO5;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_CO6;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_CQ;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_C_CY;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_C_XOR;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_D;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_D1;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_D2;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_D3;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_D4;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_D5;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_D6;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_DO5;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_DO6;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_DQ;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_D_CY;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_D_XOR;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_A;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_A1;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_A2;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_A3;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_A4;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_A5;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_A5Q;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_A6;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_AMUX;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_AO5;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_AO6;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_AQ;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_A_CY;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_A_XOR;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_B;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_B1;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_B2;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_B3;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_B4;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_B5;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_B6;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_BO5;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_BO6;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_B_CY;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_B_XOR;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_C;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_C1;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_C2;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_C3;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_C4;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_C5;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_C6;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_CLK;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_CMUX;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_CO5;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_CO6;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_C_CY;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_C_XOR;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_D;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_D1;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_D2;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_D3;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_D4;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_D5;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_D6;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_DO5;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_DO6;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_D_CY;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_D_XOR;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_SR;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_A;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_A1;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_A2;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_A3;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_A4;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_A5;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_A5Q;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_A6;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_AMUX;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_AO5;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_AO6;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_AQ;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_A_CY;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_A_XOR;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_B;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_B1;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_B2;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_B3;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_B4;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_B5;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_B5Q;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_B6;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_BMUX;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_BO5;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_BO6;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_BQ;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_B_CY;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_B_XOR;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_C;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_C1;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_C2;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_C3;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_C4;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_C5;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_C6;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_CLK;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_CO5;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_CO6;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_C_CY;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_C_XOR;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_D;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_D1;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_D2;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_D3;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_D4;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_D5;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_D6;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_DO5;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_DO6;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_D_CY;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_D_XOR;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_SR;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_A;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_A1;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_A2;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_A3;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_A4;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_A5;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_A5Q;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_A6;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_AMUX;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_AO5;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_AO6;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_AQ;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_A_CY;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_A_XOR;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_B;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_B1;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_B2;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_B3;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_B4;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_B5;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_B6;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_BO5;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_BO6;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_B_CY;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_B_XOR;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_C;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_C1;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_C2;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_C3;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_C4;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_C5;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_C6;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_CLK;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_CO5;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_CO6;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_C_CY;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_C_XOR;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_D;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_D1;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_D2;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_D3;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_D4;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_D5;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_D6;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_DO5;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_DO6;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_D_CY;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_D_XOR;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_SR;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_A;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_A1;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_A2;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_A3;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_A4;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_A5;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_A5Q;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_A6;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_AMUX;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_AO5;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_AO6;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_AQ;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_A_CY;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_A_XOR;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_B;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_B1;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_B2;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_B3;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_B4;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_B5;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_B6;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_BMUX;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_BO5;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_BO6;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_BQ;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_BX;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_B_CY;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_B_XOR;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_C;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_C1;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_C2;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_C3;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_C4;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_C5;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_C6;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_CLK;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_CMUX;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_CO5;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_CO6;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_C_CY;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_C_XOR;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_D;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_D1;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_D2;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_D3;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_D4;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_D5;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_D6;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_DO5;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_DO6;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_D_CY;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_D_XOR;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_SR;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_A;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_A1;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_A2;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_A3;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_A4;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_A5;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_A6;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_AO5;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_AO6;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_AQ;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_A_CY;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_A_XOR;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_B;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_B1;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_B2;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_B3;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_B4;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_B5;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_B5Q;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_B6;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_BMUX;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_BO5;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_BO6;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_BQ;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_B_CY;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_B_XOR;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_C;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_C1;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_C2;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_C3;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_C4;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_C5;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_C5Q;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_C6;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_CLK;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_CMUX;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_CO5;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_CO6;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_CQ;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_C_CY;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_C_XOR;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_D;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_D1;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_D2;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_D3;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_D4;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_D5;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_D6;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_DO5;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_DO6;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_DQ;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_D_CY;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_D_XOR;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_A;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_A1;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_A2;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_A3;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_A4;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_A5;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_A5Q;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_A6;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_AMUX;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_AO5;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_AO6;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_AQ;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_A_CY;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_A_XOR;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_B;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_B1;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_B2;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_B3;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_B4;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_B5;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_B5Q;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_B6;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_BMUX;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_BO5;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_BO6;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_BQ;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_B_CY;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_B_XOR;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_C;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_C1;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_C2;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_C3;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_C4;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_C5;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_C6;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_CLK;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_CO5;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_CO6;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_C_CY;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_C_XOR;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_D;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_D1;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_D2;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_D3;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_D4;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_D5;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_D6;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_DO5;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_DO6;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_D_CY;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_D_XOR;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_SR;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_A;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_A1;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_A2;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_A3;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_A4;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_A5;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_A6;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_AO5;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_AO6;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_AQ;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_A_CY;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_A_XOR;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_B;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_B1;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_B2;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_B3;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_B4;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_B5;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_B5Q;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_B6;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_BMUX;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_BO5;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_BO6;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_BQ;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_B_CY;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_B_XOR;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_C;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_C1;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_C2;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_C3;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_C4;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_C5;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_C6;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_CLK;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_CO5;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_CO6;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_CQ;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_C_CY;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_C_XOR;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_D;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_D1;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_D2;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_D3;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_D4;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_D5;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_D6;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_DO5;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_DO6;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_D_CY;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_D_XOR;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_A;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_A1;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_A2;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_A3;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_A4;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_A5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_A5Q;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_A6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_AMUX;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_AO5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_AO6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_AQ;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_A_CY;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_A_XOR;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_B;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_B1;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_B2;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_B3;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_B4;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_B5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_B6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_BO5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_BO6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_B_CY;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_B_XOR;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_C;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_C1;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_C2;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_C3;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_C4;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_C5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_C6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_CLK;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_CO5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_CO6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_C_CY;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_C_XOR;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_D;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_D1;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_D2;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_D3;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_D4;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_D5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_D6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_DO5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_DO6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_D_CY;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_D_XOR;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_SR;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_A;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_A1;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_A2;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_A3;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_A4;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_A5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_A6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_AO5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_AO6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_AQ;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_A_CY;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_A_XOR;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_B;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_B1;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_B2;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_B3;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_B4;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_B5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_B5Q;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_B6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_BMUX;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_BO5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_BO6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_BQ;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_B_CY;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_B_XOR;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_C;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_C1;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_C2;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_C3;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_C4;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_C5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_C6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_CLK;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_CO5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_CO6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_CQ;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_C_CY;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_C_XOR;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_D;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_D1;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_D2;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_D3;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_D4;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_D5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_D6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_DO5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_DO6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_D_CY;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_D_XOR;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_A;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_A1;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_A2;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_A3;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_A4;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_A5;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_A6;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_AO5;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_AO6;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_AQ;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_A_CY;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_A_XOR;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_B;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_B1;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_B2;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_B3;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_B4;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_B5;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_B5Q;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_B6;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_BMUX;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_BO5;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_BO6;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_BQ;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_B_CY;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_B_XOR;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_C;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_C1;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_C2;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_C3;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_C4;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_C5;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_C6;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_CLK;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_CMUX;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_CO5;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_CO6;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_C_CY;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_C_XOR;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_D;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_D1;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_D2;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_D3;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_D4;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_D5;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_D6;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_DO5;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_DO6;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_DQ;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_D_CY;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_D_XOR;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_A;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_A1;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_A2;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_A3;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_A4;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_A5;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_A5Q;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_A6;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_AMUX;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_AO5;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_AO6;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_AQ;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_A_CY;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_A_XOR;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_B;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_B1;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_B2;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_B3;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_B4;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_B5;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_B6;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_BMUX;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_BO5;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_BO6;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_B_CY;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_B_XOR;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_C;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_C1;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_C2;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_C3;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_C4;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_C5;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_C6;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_CLK;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_CO5;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_CO6;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_C_CY;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_C_XOR;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_D;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_D1;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_D2;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_D3;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_D4;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_D5;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_D6;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_DO5;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_DO6;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_D_CY;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_D_XOR;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_SR;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_A;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_A1;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_A2;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_A3;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_A4;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_A5;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_A6;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_AO5;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_AO6;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_AQ;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_A_CY;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_A_XOR;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_B;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_B1;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_B2;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_B3;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_B4;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_B5;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_B6;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_BO5;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_BO6;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_BQ;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_B_CY;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_B_XOR;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_C;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_C1;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_C2;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_C3;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_C4;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_C5;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_C6;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_CLK;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_CO5;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_CO6;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_CQ;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_C_CY;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_C_XOR;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_D;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_D1;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_D2;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_D3;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_D4;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_D5;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_D5Q;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_D6;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_DMUX;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_DO5;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_DO6;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_DQ;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_D_CY;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_D_XOR;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_A;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_A1;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_A2;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_A3;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_A4;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_A5;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_A5Q;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_A6;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_AMUX;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_AO5;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_AO6;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_AQ;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_A_CY;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_A_XOR;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_B;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_B1;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_B2;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_B3;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_B4;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_B5;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_B5Q;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_B6;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_BMUX;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_BO5;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_BO6;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_BQ;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_B_CY;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_B_XOR;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_C;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_C1;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_C2;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_C3;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_C4;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_C5;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_C6;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_CLK;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_CO5;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_CO6;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_C_CY;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_C_XOR;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_D;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_D1;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_D2;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_D3;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_D4;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_D5;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_D6;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_DO5;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_DO6;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_D_CY;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_D_XOR;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_A;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_A1;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_A2;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_A3;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_A4;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_A5;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_A6;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_AO5;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_AO6;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_AQ;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_A_CY;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_A_XOR;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_B;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_B1;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_B2;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_B3;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_B4;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_B5;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_B6;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_BO5;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_BO6;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_BQ;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_B_CY;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_B_XOR;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_C;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_C1;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_C2;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_C3;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_C4;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_C5;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_C6;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_CLK;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_CO5;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_CO6;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_CQ;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_C_CY;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_C_XOR;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_D;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_D1;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_D2;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_D3;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_D4;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_D5;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_D6;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_DMUX;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_DO5;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_DO6;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_D_CY;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_D_XOR;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_A;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_A1;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_A2;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_A3;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_A4;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_A5;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_A6;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_AMUX;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_AO5;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_AO6;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_A_CY;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_A_XOR;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_B;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_B1;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_B2;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_B3;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_B4;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_B5;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_B6;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_BO5;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_BO6;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_BQ;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_B_CY;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_B_XOR;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_C;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_C1;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_C2;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_C3;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_C4;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_C5;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_C6;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_CLK;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_CO5;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_CO6;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_C_CY;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_C_XOR;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_D;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_D1;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_D2;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_D3;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_D4;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_D5;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_D6;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_DO5;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_DO6;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_D_CY;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_D_XOR;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_A;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_A1;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_A2;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_A3;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_A4;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_A5;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_A6;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_AO5;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_AO6;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_AQ;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_A_CY;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_A_XOR;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_B;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_B1;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_B2;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_B3;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_B4;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_B5;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_B6;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_BO5;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_BO6;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_B_CY;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_B_XOR;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_C;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_C1;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_C2;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_C3;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_C4;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_C5;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_C6;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_CLK;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_CO5;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_CO6;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_C_CY;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_C_XOR;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_D;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_D1;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_D2;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_D3;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_D4;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_D5;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_D6;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_DO5;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_DO6;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_D_CY;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_D_XOR;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_A;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_A1;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_A2;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_A3;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_A4;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_A5;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_A6;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_AO5;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_AO6;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_A_CY;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_A_XOR;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_B;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_B1;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_B2;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_B3;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_B4;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_B5;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_B6;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_BO5;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_BO6;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_B_CY;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_B_XOR;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_C;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_C1;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_C2;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_C3;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_C4;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_C5;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_C6;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_CO5;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_CO6;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_C_CY;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_C_XOR;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_D;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_D1;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_D2;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_D3;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_D4;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_D5;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_D6;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_DO5;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_DO6;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_D_CY;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_D_XOR;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_A;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_A1;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_A2;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_A3;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_A4;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_A5;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_A6;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_AO5;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_AO6;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_A_CY;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_A_XOR;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_B;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_B1;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_B2;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_B3;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_B4;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_B5;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_B6;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_BO5;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_BO6;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_B_CY;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_B_XOR;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_C;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_C1;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_C2;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_C3;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_C4;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_C5;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_C6;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_CO5;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_CO6;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_C_CY;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_C_XOR;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_D;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_D1;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_D2;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_D3;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_D4;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_D5;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_D6;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_DO5;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_DO6;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_D_CY;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_D_XOR;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_A;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_A1;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_A2;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_A3;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_A4;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_A5;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_A6;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_AO5;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_AO6;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_A_CY;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_A_XOR;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_B;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_B1;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_B2;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_B3;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_B4;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_B5;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_B6;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_BO5;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_BO6;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_B_CY;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_B_XOR;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_C;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_C1;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_C2;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_C3;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_C4;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_C5;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_C6;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_CO5;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_CO6;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_C_CY;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_C_XOR;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_D;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_D1;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_D2;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_D3;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_D4;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_D5;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_D6;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_DO5;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_DO6;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_D_CY;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_D_XOR;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_A;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_A1;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_A2;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_A3;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_A4;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_A5;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_A6;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_AO5;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_AO6;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_AQ;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_A_CY;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_A_XOR;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_B;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_B1;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_B2;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_B3;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_B4;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_B5;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_B6;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_BMUX;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_BO5;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_BO6;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_B_CY;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_B_XOR;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_C;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_C1;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_C2;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_C3;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_C4;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_C5;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_C6;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_CLK;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_CMUX;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_CO5;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_CO6;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_C_CY;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_C_XOR;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_D;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_D1;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_D2;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_D3;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_D4;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_D5;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_D6;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_DO5;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_DO6;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_D_CY;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_D_XOR;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_A;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_A1;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_A2;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_A3;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_A4;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_A5;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_A6;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_AO5;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_AO6;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_A_CY;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_A_XOR;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_B;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_B1;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_B2;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_B3;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_B4;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_B5;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_B6;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_BO5;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_BO6;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_B_CY;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_B_XOR;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_C;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_C1;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_C2;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_C3;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_C4;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_C5;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_C6;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_CO5;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_CO6;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_C_CY;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_C_XOR;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_D;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_D1;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_D2;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_D3;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_D4;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_D5;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_D6;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_DO5;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_DO6;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_D_CY;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_D_XOR;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_A;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_A1;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_A2;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_A3;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_A4;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_A5;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_A6;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_AO5;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_AO6;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_AQ;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_A_CY;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_A_XOR;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_B;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_B1;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_B2;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_B3;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_B4;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_B5;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_B6;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_BMUX;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_BO5;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_BO6;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_B_CY;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_B_XOR;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_C;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_C1;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_C2;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_C3;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_C4;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_C5;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_C6;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_CLK;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_CMUX;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_CO5;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_CO6;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_C_CY;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_C_XOR;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_D;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_D1;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_D2;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_D3;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_D4;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_D5;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_D6;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_DO5;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_DO6;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_D_CY;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X14Y143_D_XOR;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_A;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_A1;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_A2;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_A3;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_A4;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_A5;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_A6;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_AO5;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_AO6;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_A_CY;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_A_XOR;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_B;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_B1;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_B2;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_B3;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_B4;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_B5;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_B6;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_BO5;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_BO6;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_B_CY;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_B_XOR;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_C;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_C1;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_C2;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_C3;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_C4;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_C5;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_C6;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_CO5;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_CO6;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_C_CY;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_C_XOR;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_D;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_D1;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_D2;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_D3;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_D4;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_D5;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_D6;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_DO5;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_DO6;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_D_CY;
  wire [0:0] CLBLM_R_X11Y143_SLICE_X15Y143_D_XOR;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_A;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_A1;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_A2;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_A3;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_A4;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_A5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_A6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_AO5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_AO6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_AQ;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_AX;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_A_CY;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_A_XOR;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_B;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_B1;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_B2;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_B3;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_B4;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_B5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_B6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_BO5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_BO6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_B_CY;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_B_XOR;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_C;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_C1;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_C2;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_C3;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_C4;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_C5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_C6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_CE;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_CLK;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_CO5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_CO6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_C_CY;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_C_XOR;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_D;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_D1;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_D2;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_D3;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_D4;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_D5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_D6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_DO5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_DO6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_D_CY;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_D_XOR;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_A;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_A1;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_A2;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_A3;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_A4;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_A5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_A6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_AMUX;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_AO5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_AO6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_A_CY;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_A_XOR;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_B;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_B1;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_B2;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_B3;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_B4;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_B5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_B6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_BO5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_BO6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_B_CY;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_B_XOR;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_C;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_C1;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_C2;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_C3;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_C4;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_C5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_C6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_CMUX;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_CO5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_CO6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_C_CY;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_C_XOR;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_D;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_D1;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_D2;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_D3;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_D4;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_D5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_D6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_DO5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_DO6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_D_CY;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_D_XOR;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_A;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_A1;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_A2;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_A3;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_A4;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_A5;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_A6;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_AMUX;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_AO5;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_AO6;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_AQ;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_AX;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_A_CY;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_A_XOR;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_B;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_B1;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_B2;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_B3;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_B4;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_B5;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_B6;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_BMUX;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_BO5;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_BO6;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_BQ;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_BX;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_B_CY;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_B_XOR;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_C;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_C1;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_C2;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_C3;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_C4;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_C5;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_C6;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_CE;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_CLK;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_CO5;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_CO6;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_CQ;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_CX;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_C_CY;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_C_XOR;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_D;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_D1;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_D2;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_D3;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_D4;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_D5;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_D6;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_DO5;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_DO6;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_DQ;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_DX;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_D_CY;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X14Y145_D_XOR;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_A;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_A1;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_A2;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_A3;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_A4;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_A5;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_A6;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_AMUX;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_AO5;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_AO6;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_AQ;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_AX;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_A_CY;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_A_XOR;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_B;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_B1;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_B2;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_B3;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_B4;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_B5;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_B6;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_BMUX;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_BO5;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_BO6;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_B_CY;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_B_XOR;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_C;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_C1;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_C2;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_C3;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_C4;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_C5;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_C6;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_CE;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_CLK;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_CO5;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_CO6;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_C_CY;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_C_XOR;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_D;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_D1;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_D2;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_D3;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_D4;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_D5;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_D6;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_DO5;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_DO6;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_D_CY;
  wire [0:0] CLBLM_R_X11Y145_SLICE_X15Y145_D_XOR;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_A;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_A1;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_A2;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_A3;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_A4;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_A5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_A6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_AMUX;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_AO5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_AO6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_AQ;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_AX;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_A_CY;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_A_XOR;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_B;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_B1;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_B2;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_B3;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_B4;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_B5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_B6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_BO5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_BO6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_B_CY;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_B_XOR;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_C;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_C1;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_C2;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_C3;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_C4;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_C5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_C6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_CLK;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_CO5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_CO6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_C_CY;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_C_XOR;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_D;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_D1;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_D2;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_D3;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_D4;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_D5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_D6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_DO5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_DO6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_D_CY;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_D_XOR;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_SR;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_A;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_A1;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_A2;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_A3;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_A4;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_A5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_A6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_AO5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_AO6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_AQ;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_A_CY;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_A_XOR;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_B;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_B1;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_B2;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_B3;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_B4;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_B5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_B6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_BMUX;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_BO5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_BO6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_B_CY;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_B_XOR;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_C;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_C1;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_C2;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_C3;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_C4;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_C5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_C6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_CLK;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_CMUX;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_CO5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_CO6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_C_CY;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_C_XOR;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_D;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_D1;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_D2;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_D3;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_D4;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_D5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_D6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_DO5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_DO6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_D_CY;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_D_XOR;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_A;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_A1;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_A2;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_A3;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_A4;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_A5;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_A5Q;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_A6;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_AMUX;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_AO5;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_AO6;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_AQ;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_A_CY;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_A_XOR;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_B;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_B1;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_B2;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_B3;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_B4;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_B5;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_B6;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_BO5;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_BO6;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_B_CY;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_B_XOR;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_C;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_C1;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_C2;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_C3;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_C4;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_C5;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_C6;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_CLK;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_CO5;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_CO6;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_C_CY;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_C_XOR;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_D;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_D1;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_D2;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_D3;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_D4;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_D5;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_D6;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_DO5;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_DO6;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_D_CY;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_D_XOR;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_SR;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_A;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_A1;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_A2;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_A3;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_A4;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_A5;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_A6;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_AO5;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_AO6;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_AQ;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_A_CY;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_A_XOR;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_B;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_B1;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_B2;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_B3;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_B4;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_B5;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_B6;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_BO5;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_BO6;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_B_CY;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_B_XOR;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_C;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_C1;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_C2;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_C3;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_C4;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_C5;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_C6;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_CLK;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_CMUX;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_CO5;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_CO6;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_C_CY;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_C_XOR;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_D;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_D1;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_D2;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_D3;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_D4;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_D5;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_D6;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_DO5;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_DO6;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_D_CY;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_D_XOR;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_A;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_A1;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_A2;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_A3;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_A4;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_A5;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_A6;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_AO5;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_AO6;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_AQ;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_AX;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_A_CY;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_A_XOR;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_B;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_B1;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_B2;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_B3;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_B4;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_B5;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_B6;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_BO5;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_BO6;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_BQ;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_BX;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_B_CY;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_B_XOR;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_C;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_C1;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_C2;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_C3;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_C4;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_C5;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_C6;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_CE;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_CLK;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_CO5;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_CO6;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_CQ;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_CX;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_C_CY;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_C_XOR;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_D;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_D1;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_D2;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_D3;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_D4;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_D5;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_D6;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_DO5;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_DO6;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_DQ;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_DX;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_D_CY;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_D_XOR;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_A;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_A1;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_A2;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_A3;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_A4;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_A5;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_A6;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_AMUX;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_AO5;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_AO6;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_AQ;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_AX;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_A_CY;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_A_XOR;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_B;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_B1;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_B2;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_B3;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_B4;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_B5;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_B6;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_BO5;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_BO6;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_B_CY;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_B_XOR;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_C;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_C1;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_C2;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_C3;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_C4;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_C5;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_C6;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_CLK;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_CO5;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_CO6;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_C_CY;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_C_XOR;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_D;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_D1;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_D2;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_D3;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_D4;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_D5;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_D6;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_DO5;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_DO6;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_D_CY;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_D_XOR;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_SR;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_A;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_A1;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_A2;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_A3;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_A4;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_A5;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_A6;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_AMUX;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_AO5;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_AO6;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_AQ;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_AX;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_A_CY;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_A_XOR;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_B;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_B1;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_B2;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_B3;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_B4;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_B5;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_B6;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_BMUX;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_BO5;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_BO6;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_B_CY;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_B_XOR;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_C;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_C1;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_C2;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_C3;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_C4;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_C5;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_C6;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_CLK;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_CO5;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_CO6;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_C_CY;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_C_XOR;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_D;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_D1;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_D2;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_D3;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_D4;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_D5;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_D6;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_DO5;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_DO6;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_D_CY;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_D_XOR;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_SR;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_A;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_A1;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_A2;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_A3;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_A4;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_A5;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_A6;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_AO5;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_AO6;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_AQ;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_A_CY;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_A_XOR;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_B;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_B1;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_B2;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_B3;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_B4;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_B5;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_B6;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_BO5;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_BO6;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_BQ;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_B_CY;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_B_XOR;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_C;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_C1;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_C2;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_C3;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_C4;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_C5;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_C6;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_CLK;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_CO5;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_CO6;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_CQ;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_C_CY;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_C_XOR;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_D;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_D1;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_D2;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_D3;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_D4;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_D5;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_D6;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_DMUX;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_DO5;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_DO6;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_D_CY;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_D_XOR;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_A;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_A1;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_A2;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_A3;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_A4;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_A5;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_A6;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_AO5;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_AO6;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_AQ;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_A_CY;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_A_XOR;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_B;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_B1;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_B2;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_B3;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_B4;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_B5;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_B6;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_BMUX;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_BO5;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_BO6;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_B_CY;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_B_XOR;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_C;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_C1;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_C2;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_C3;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_C4;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_C5;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_C6;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_CLK;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_CO5;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_CO6;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_C_CY;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_C_XOR;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_D;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_D1;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_D2;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_D3;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_D4;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_D5;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_D6;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_DO5;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_DO6;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_D_CY;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_D_XOR;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_SR;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_A;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_A1;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_A2;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_A3;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_A4;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_A5;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_A6;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_AO5;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_AO6;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_AQ;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_A_CY;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_A_XOR;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_B;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_B1;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_B2;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_B3;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_B4;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_B5;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_B6;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_BO5;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_BO6;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_B_CY;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_B_XOR;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_C;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_C1;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_C2;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_C3;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_C4;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_C5;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_C6;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_CLK;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_CO5;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_CO6;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_C_CY;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_C_XOR;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_D;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_D1;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_D2;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_D3;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_D4;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_D5;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_D6;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_DO5;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_DO6;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_D_CY;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_D_XOR;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_A;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_A1;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_A2;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_A3;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_A4;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_A5;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_A6;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_AO5;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_AO6;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_AQ;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_A_CY;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_A_XOR;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_B;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_B1;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_B2;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_B3;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_B4;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_B5;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_B6;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_BO5;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_BO6;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_BQ;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_B_CY;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_B_XOR;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_C;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_C1;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_C2;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_C3;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_C4;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_C5;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_C6;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_CLK;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_CMUX;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_CO5;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_CO6;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_C_CY;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_C_XOR;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_D;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_D1;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_D2;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_D3;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_D4;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_D5;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_D6;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_DO5;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_DO6;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_D_CY;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_D_XOR;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_A;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_A1;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_A2;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_A3;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_A4;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_A5;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_A5Q;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_A6;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_AMUX;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_AO5;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_AO6;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_AQ;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_AX;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_A_CY;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_A_XOR;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_B;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_B1;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_B2;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_B3;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_B4;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_B5;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_B6;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_BO5;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_BO6;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_BQ;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_B_CY;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_B_XOR;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_C;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_C1;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_C2;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_C3;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_C4;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_C5;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_C6;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_CLK;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_CMUX;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_CO5;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_CO6;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_C_CY;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_C_XOR;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_D;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_D1;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_D2;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_D3;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_D4;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_D5;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_D6;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_DO5;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_DO6;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_D_CY;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_D_XOR;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_A;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_A1;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_A2;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_A3;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_A4;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_A5;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_A5Q;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_A6;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_AMUX;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_AO5;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_AO6;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_AQ;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_A_CY;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_A_XOR;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_B;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_B1;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_B2;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_B3;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_B4;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_B5;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_B6;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_BO5;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_BO6;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_B_CY;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_B_XOR;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_C;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_C1;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_C2;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_C3;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_C4;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_C5;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_C6;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_CLK;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_CO5;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_CO6;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_C_CY;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_C_XOR;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_D;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_D1;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_D2;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_D3;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_D4;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_D5;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_D6;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_DO5;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_DO6;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_D_CY;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_D_XOR;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_A;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_A1;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_A2;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_A3;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_A4;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_A5;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_A6;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_AO5;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_AO6;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_A_CY;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_A_XOR;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_B;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_B1;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_B2;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_B3;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_B4;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_B5;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_B6;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_BO5;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_BO6;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_B_CY;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_B_XOR;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_C;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_C1;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_C2;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_C3;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_C4;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_C5;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_C6;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_CO5;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_CO6;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_C_CY;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_C_XOR;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_D;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_D1;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_D2;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_D3;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_D4;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_D5;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_D6;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_DO5;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_DO6;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_D_CY;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_D_XOR;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_A;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_A1;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_A2;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_A3;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_A4;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_A5;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_A6;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_AMUX;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_AO5;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_AO6;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_A_CY;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_A_XOR;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_B;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_B1;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_B2;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_B3;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_B4;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_B5;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_B6;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_BO5;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_BO6;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_B_CY;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_B_XOR;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_C;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_C1;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_C2;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_C3;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_C4;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_C5;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_C6;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_CO5;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_CO6;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_C_CY;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_C_XOR;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_D;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_D1;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_D2;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_D3;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_D4;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_D5;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_D6;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_DO5;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_DO6;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_D_CY;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_D_XOR;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_A;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_A1;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_A2;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_A3;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_A4;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_A5;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_A6;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_AO5;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_AO6;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_A_CY;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_A_XOR;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_B;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_B1;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_B2;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_B3;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_B4;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_B5;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_B6;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_BO5;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_BO6;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_B_CY;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_B_XOR;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_C;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_C1;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_C2;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_C3;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_C4;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_C5;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_C6;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_CO5;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_CO6;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_C_CY;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_C_XOR;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_D;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_D1;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_D2;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_D3;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_D4;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_D5;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_D6;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_DO5;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_DO6;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_D_CY;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_D_XOR;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_A;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_A1;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_A2;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_A3;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_A4;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_A5;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_A6;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_AO5;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_AO6;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_A_CY;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_A_XOR;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_B;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_B1;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_B2;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_B3;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_B4;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_B5;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_B6;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_BO5;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_BO6;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_B_CY;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_B_XOR;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_C;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_C1;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_C2;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_C3;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_C4;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_C5;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_C6;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_CO5;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_CO6;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_C_CY;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_C_XOR;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_D;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_D1;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_D2;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_D3;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_D4;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_D5;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_D6;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_DO5;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_DO6;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_D_CY;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X18Y145_D_XOR;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_A;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_A1;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_A2;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_A3;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_A4;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_A5;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_A6;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_AO5;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_AO6;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_A_CY;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_A_XOR;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_B;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_B1;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_B2;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_B3;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_B4;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_B5;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_B6;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_BO5;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_BO6;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_B_CY;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_B_XOR;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_C;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_C1;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_C2;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_C3;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_C4;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_C5;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_C6;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_CO5;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_CO6;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_C_CY;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_C_XOR;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_D;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_D1;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_D2;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_D3;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_D4;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_D5;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_D6;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_DO5;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_DO6;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_D_CY;
  wire [0:0] CLBLM_R_X13Y145_SLICE_X19Y145_D_XOR;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_A;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_A1;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_A2;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_A3;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_A4;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_A5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_A6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_AMUX;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_AO5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_AO6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_A_CY;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_A_XOR;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_B;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_B1;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_B2;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_B3;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_B4;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_B5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_B6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_BO5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_BO6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_B_CY;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_B_XOR;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_C;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_C1;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_C2;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_C3;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_C4;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_C5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_C6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_CO5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_CO6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_C_CY;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_C_XOR;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_D;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_D1;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_D2;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_D3;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_D4;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_D5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_D6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_DO5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_DO6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_D_CY;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_D_XOR;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_A;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_A1;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_A2;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_A3;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_A4;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_A5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_A6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_AO5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_AO6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_A_CY;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_A_XOR;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_B;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_B1;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_B2;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_B3;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_B4;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_B5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_B6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_BO5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_BO6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_B_CY;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_B_XOR;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_C;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_C1;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_C2;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_C3;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_C4;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_C5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_C6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_CO5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_CO6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_C_CY;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_C_XOR;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_D;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_D1;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_D2;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_D3;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_D4;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_D5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_D6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_DO5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_DO6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_D_CY;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_D_XOR;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_A;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_A1;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_A2;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_A3;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_A4;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_A5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_A5Q;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_A6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_AMUX;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_AO5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_AO6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_AQ;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_AX;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_A_CY;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_A_XOR;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_B;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_B1;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_B2;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_B3;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_B4;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_B5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_B5Q;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_B6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_BMUX;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_BO5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_BO6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_BQ;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_B_CY;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_B_XOR;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_C;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_C1;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_C2;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_C3;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_C4;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_C5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_C6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_CLK;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_CMUX;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_CO5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_CO6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_C_CY;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_C_XOR;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_D;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_D1;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_D2;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_D3;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_D4;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_D5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_D6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_DO5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_DO6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_D_CY;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_D_XOR;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_A;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_A1;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_A2;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_A3;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_A4;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_A5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_A6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_AO5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_AO6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_AQ;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_A_CY;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_A_XOR;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_B;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_B1;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_B2;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_B3;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_B4;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_B5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_B6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_BO5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_BO6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_BQ;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_B_CY;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_B_XOR;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_C;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_C1;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_C2;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_C3;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_C4;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_C5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_C6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_CLK;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_CO5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_CO6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_CQ;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_C_CY;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_C_XOR;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_D;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_D1;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_D2;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_D3;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_D4;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_D5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_D6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_DMUX;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_DO5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_DO6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_D_CY;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_D_XOR;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_A;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_A1;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_A2;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_A3;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_A4;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_A5;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_A6;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_AO5;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_AO6;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_AQ;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_A_CY;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_A_XOR;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_B;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_B1;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_B2;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_B3;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_B4;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_B5;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_B6;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_BO5;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_BO6;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_BQ;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_B_CY;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_B_XOR;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_C;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_C1;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_C2;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_C3;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_C4;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_C5;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_C6;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_CLK;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_CO5;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_CO6;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_CQ;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_C_CY;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_C_XOR;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_D;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_D1;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_D2;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_D3;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_D4;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_D5;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_D6;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_DO5;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_DO6;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_DQ;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_D_CY;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X2Y143_D_XOR;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_A;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_A1;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_A2;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_A3;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_A4;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_A5;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_A6;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_AO5;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_AO6;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_AQ;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_A_CY;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_A_XOR;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_B;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_B1;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_B2;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_B3;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_B4;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_B5;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_B6;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_BMUX;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_BO5;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_BO6;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_B_CY;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_B_XOR;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_C;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_C1;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_C2;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_C3;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_C4;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_C5;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_C6;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_CLK;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_CMUX;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_CO5;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_CO6;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_C_CY;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_C_XOR;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_D;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_D1;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_D2;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_D3;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_D4;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_D5;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_D6;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_DMUX;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_DO5;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_DO6;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_D_CY;
  wire [0:0] CLBLM_R_X3Y143_SLICE_X3Y143_D_XOR;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_A;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_A1;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_A2;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_A3;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_A4;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_A5;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_A5Q;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_A6;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_AMUX;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_AO5;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_AO6;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_AQ;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_A_CY;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_A_XOR;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_B;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_B1;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_B2;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_B3;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_B4;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_B5;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_B6;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_BMUX;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_BO5;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_BO6;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_B_CY;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_B_XOR;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_C;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_C1;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_C2;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_C3;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_C4;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_C5;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_C6;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_CLK;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_CO5;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_CO6;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_C_CY;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_C_XOR;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_D;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_D1;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_D2;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_D3;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_D4;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_D5;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_D6;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_DO5;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_DO6;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_D_CY;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_D_XOR;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X2Y144_SR;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_A;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_A1;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_A2;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_A3;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_A4;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_A5;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_A5Q;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_A6;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_AMUX;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_AO5;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_AO6;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_AQ;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_A_CY;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_A_XOR;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_B;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_B1;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_B2;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_B3;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_B4;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_B5;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_B6;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_BO5;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_BO6;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_BQ;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_B_CY;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_B_XOR;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_C;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_C1;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_C2;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_C3;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_C4;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_C5;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_C6;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_CLK;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_CO5;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_CO6;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_CQ;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_C_CY;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_C_XOR;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_D;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_D1;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_D2;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_D3;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_D4;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_D5;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_D5Q;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_D6;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_DMUX;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_DO5;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_DO6;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_DQ;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_D_CY;
  wire [0:0] CLBLM_R_X3Y144_SLICE_X3Y144_D_XOR;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_A;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_A1;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_A2;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_A3;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_A4;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_A5;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_A6;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_AO5;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_AO6;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_AQ;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_A_CY;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_A_XOR;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_B;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_B1;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_B2;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_B3;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_B4;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_B5;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_B5Q;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_B6;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_BMUX;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_BO5;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_BO6;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_BQ;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_B_CY;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_B_XOR;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_C;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_C1;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_C2;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_C3;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_C4;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_C5;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_C5Q;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_C6;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_CLK;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_CMUX;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_CO5;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_CO6;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_CQ;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_C_CY;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_C_XOR;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_D;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_D1;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_D2;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_D3;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_D4;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_D5;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_D6;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_DO5;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_DO6;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_DQ;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_D_CY;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X2Y145_D_XOR;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_A;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_A1;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_A2;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_A3;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_A4;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_A5;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_A5Q;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_A6;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_AMUX;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_AO5;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_AO6;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_AQ;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_A_CY;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_A_XOR;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_B;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_B1;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_B2;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_B3;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_B4;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_B5;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_B6;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_BO5;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_BO6;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_BQ;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_B_CY;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_B_XOR;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_C;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_C1;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_C2;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_C3;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_C4;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_C5;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_C6;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_CLK;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_CO5;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_CO6;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_CQ;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_C_CY;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_C_XOR;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_D;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_D1;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_D2;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_D3;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_D4;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_D5;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_D6;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_DO5;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_DO6;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_DQ;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_D_CY;
  wire [0:0] CLBLM_R_X3Y145_SLICE_X3Y145_D_XOR;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_A;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_A1;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_A2;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_A3;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_A4;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_A5;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_A6;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_AO5;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_AO6;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_AQ;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_A_CY;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_A_XOR;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_B;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_B1;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_B2;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_B3;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_B4;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_B5;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_B5Q;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_B6;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_BMUX;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_BO5;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_BO6;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_BQ;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_B_CY;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_B_XOR;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_C;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_C1;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_C2;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_C3;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_C4;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_C5;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_C5Q;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_C6;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_CLK;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_CMUX;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_CO5;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_CO6;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_CQ;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_C_CY;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_C_XOR;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_D;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_D1;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_D2;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_D3;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_D4;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_D5;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_D6;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_DO5;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_DO6;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_D_CY;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X2Y146_D_XOR;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_A;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_A1;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_A2;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_A3;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_A4;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_A5;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_A6;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_AO5;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_AO6;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_AQ;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_A_CY;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_A_XOR;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_B;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_B1;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_B2;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_B3;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_B4;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_B5;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_B6;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_BO5;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_BO6;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_BQ;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_B_CY;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_B_XOR;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_C;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_C1;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_C2;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_C3;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_C4;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_C5;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_C5Q;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_C6;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_CLK;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_CMUX;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_CO5;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_CO6;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_CQ;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_C_CY;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_C_XOR;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_D;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_D1;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_D2;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_D3;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_D4;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_D5;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_D6;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_DO5;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_DO6;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_DQ;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_D_CY;
  wire [0:0] CLBLM_R_X3Y146_SLICE_X3Y146_D_XOR;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_A;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_A1;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_A2;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_A3;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_A4;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_A5;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_A6;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_AO5;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_AO6;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_AQ;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_A_CY;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_A_XOR;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_B;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_B1;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_B2;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_B3;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_B4;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_B5;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_B6;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_BO5;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_BO6;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_BQ;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_B_CY;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_B_XOR;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_C;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_C1;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_C2;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_C3;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_C4;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_C5;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_C5Q;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_C6;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_CLK;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_CMUX;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_CO5;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_CO6;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_CQ;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_C_CY;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_C_XOR;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_D;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_D1;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_D2;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_D3;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_D4;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_D5;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_D6;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_DMUX;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_DO5;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_DO6;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_D_CY;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X2Y147_D_XOR;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_A;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_A1;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_A2;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_A3;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_A4;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_A5;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_A5Q;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_A6;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_AMUX;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_AO5;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_AO6;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_AQ;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_AX;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_A_CY;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_A_XOR;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_B;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_B1;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_B2;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_B3;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_B4;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_B5;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_B5Q;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_B6;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_BMUX;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_BO5;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_BO6;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_BQ;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_B_CY;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_B_XOR;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_C;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_C1;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_C2;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_C3;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_C4;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_C5;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_C6;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_CLK;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_CMUX;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_CO5;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_CO6;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_C_CY;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_C_XOR;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_D;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_D1;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_D2;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_D3;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_D4;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_D5;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_D6;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_DO5;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_DO6;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_D_CY;
  wire [0:0] CLBLM_R_X3Y147_SLICE_X3Y147_D_XOR;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_A;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_A1;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_A2;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_A3;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_A4;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_A5;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_A6;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_AO5;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_AO6;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_AQ;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_A_CY;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_A_XOR;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_B;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_B1;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_B2;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_B3;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_B4;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_B5;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_B5Q;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_B6;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_BMUX;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_BO5;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_BO6;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_BQ;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_B_CY;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_B_XOR;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_C;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_C1;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_C2;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_C3;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_C4;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_C5;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_C5Q;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_C6;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_CLK;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_CMUX;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_CO5;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_CO6;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_CQ;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_C_CY;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_C_XOR;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_D;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_D1;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_D2;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_D3;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_D4;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_D5;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_D5Q;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_D6;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_DMUX;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_DO5;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_DO6;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_DQ;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_D_CY;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X2Y148_D_XOR;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_A;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_A1;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_A2;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_A3;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_A4;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_A5;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_A5Q;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_A6;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_AMUX;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_AO5;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_AO6;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_AQ;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_A_CY;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_A_XOR;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_B;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_B1;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_B2;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_B3;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_B4;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_B5;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_B6;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_BMUX;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_BO5;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_BO6;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_B_CY;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_B_XOR;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_C;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_C1;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_C2;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_C3;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_C4;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_C5;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_C6;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_CLK;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_CMUX;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_CO5;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_CO6;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_C_CY;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_C_XOR;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_D;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_D1;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_D2;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_D3;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_D4;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_D5;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_D6;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_DMUX;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_DO5;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_DO6;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_D_CY;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_D_XOR;
  wire [0:0] CLBLM_R_X3Y148_SLICE_X3Y148_SR;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_A;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_A1;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_A2;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_A3;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_A4;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_A5;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_A5Q;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_A6;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_AMUX;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_AO5;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_AO6;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_AQ;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_A_CY;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_A_XOR;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_B;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_B1;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_B2;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_B3;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_B4;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_B5;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_B6;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_BO5;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_BO6;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_BQ;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_B_CY;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_B_XOR;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_C;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_C1;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_C2;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_C3;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_C4;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_C5;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_C6;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_CLK;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_CO5;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_CO6;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_CQ;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_C_CY;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_C_XOR;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_D;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_D1;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_D2;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_D3;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_D4;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_D5;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_D6;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_DO5;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_DO6;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_D_CY;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X2Y149_D_XOR;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_A;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_A1;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_A2;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_A3;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_A4;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_A5;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_A6;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_AO5;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_AO6;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_AQ;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_A_CY;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_A_XOR;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_B;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_B1;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_B2;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_B3;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_B4;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_B5;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_B6;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_BO5;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_BO6;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_BQ;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_B_CY;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_B_XOR;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_C;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_C1;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_C2;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_C3;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_C4;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_C5;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_C6;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_CLK;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_CO5;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_CO6;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_CQ;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_C_CY;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_C_XOR;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_D;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_D1;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_D2;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_D3;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_D4;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_D5;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_D6;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_DO5;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_DO6;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_DQ;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_D_CY;
  wire [0:0] CLBLM_R_X3Y149_SLICE_X3Y149_D_XOR;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_A;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_A1;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_A2;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_A3;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_A4;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_A5;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_A6;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_AO5;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_AO6;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_AQ;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_A_CY;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_A_XOR;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_B;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_B1;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_B2;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_B3;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_B4;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_B5;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_B5Q;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_B6;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_BMUX;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_BO5;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_BO6;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_BQ;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_B_CY;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_B_XOR;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_C;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_C1;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_C2;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_C3;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_C4;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_C5;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_C6;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_CLK;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_CMUX;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_CO5;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_CO6;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_C_CY;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_C_XOR;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_D;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_D1;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_D2;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_D3;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_D4;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_D5;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_D6;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_DO5;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_DO6;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_DQ;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_D_CY;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_D_XOR;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_A;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_A1;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_A2;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_A3;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_A4;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_A5;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_A6;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_AO5;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_AQ;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_A_CY;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_A_XOR;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_B;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_B1;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_B2;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_B3;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_B4;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_B5;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_B6;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_BO5;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_BO6;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_BQ;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_B_CY;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_B_XOR;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_C;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_C1;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_C2;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_C3;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_C4;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_C5;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_C6;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_CLK;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_CO5;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_CO6;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_CQ;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_C_CY;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_C_XOR;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_D;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_D1;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_D2;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_D3;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_D4;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_D5;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_D6;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_DO5;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_DO6;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_D_CY;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_D_XOR;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_A;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_A1;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_A2;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_A3;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_A4;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_A5;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_A5Q;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_A6;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_AMUX;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_AO5;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_AO6;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_AQ;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_AX;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_A_CY;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_A_XOR;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_B;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_B1;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_B2;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_B3;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_B4;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_B5;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_B6;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_BO5;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_BO6;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_BQ;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_B_CY;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_B_XOR;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_C;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_C1;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_C2;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_C3;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_C4;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_C5;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_C6;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_CLK;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_CMUX;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_CO5;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_CO6;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_C_CY;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_C_XOR;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_D;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_D1;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_D2;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_D3;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_D4;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_D5;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_D6;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_DO5;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_DO6;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_D_CY;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_D_XOR;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_A;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_A1;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_A2;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_A3;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_A4;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_A5;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_A6;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_AO5;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_AO6;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_AQ;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_A_CY;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_A_XOR;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_B;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_B1;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_B2;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_B3;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_B4;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_B5;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_B6;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_BO5;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_BO6;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_BQ;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_B_CY;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_B_XOR;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_C;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_C1;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_C2;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_C3;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_C4;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_C5;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_C5Q;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_C6;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_CLK;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_CMUX;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_CO5;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_CO6;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_CQ;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_C_CY;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_C_XOR;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_D;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_D1;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_D2;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_D3;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_D4;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_D5;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_D5Q;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_D6;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_DMUX;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_DO5;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_DO6;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_DQ;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_D_CY;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_D_XOR;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_A;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_A1;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_A2;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_A3;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_A4;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_A5;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_A6;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_AO5;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_AO6;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_AQ;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_A_CY;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_A_XOR;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_B;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_B1;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_B2;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_B3;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_B4;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_B5;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_B6;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_BO5;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_BO6;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_BQ;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_B_CY;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_B_XOR;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_C;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_C1;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_C2;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_C3;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_C4;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_C5;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_C6;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_CLK;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_CO5;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_CO6;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_CQ;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_C_CY;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_C_XOR;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_D;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_D1;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_D2;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_D3;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_D4;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_D5;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_D6;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_DO5;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_DO6;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_D_CY;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_D_XOR;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_A;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_A1;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_A2;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_A3;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_A4;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_A5;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_A5Q;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_A6;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_AMUX;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_AO5;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_AO6;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_AQ;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_A_CY;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_A_XOR;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_B;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_B1;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_B2;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_B3;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_B4;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_B5;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_B6;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_BO5;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_BO6;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_B_CY;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_B_XOR;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_C;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_C1;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_C2;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_C3;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_C4;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_C5;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_C6;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_CLK;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_CMUX;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_CO5;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_CO6;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_C_CY;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_C_XOR;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_D;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_D1;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_D2;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_D3;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_D4;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_D5;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_D6;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_DO5;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_DO6;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_D_CY;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_D_XOR;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_A;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_A1;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_A2;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_A3;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_A4;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_A5;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_A6;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_AMUX;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_AO5;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_AO6;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_AQ;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_AX;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_A_CY;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_A_XOR;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_B;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_B1;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_B2;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_B3;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_B4;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_B5;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_B6;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_BO5;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_BO6;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_B_CY;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_B_XOR;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_C;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_C1;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_C2;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_C3;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_C4;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_C5;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_C6;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_CE;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_CLK;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_CO5;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_CO6;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_C_CY;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_C_XOR;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_D;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_D1;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_D2;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_D3;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_D4;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_D5;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_D6;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_DO5;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_DO6;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_D_CY;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_D_XOR;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_A;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_A1;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_A2;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_A3;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_A4;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_A5;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_A5Q;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_A6;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_AMUX;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_AO5;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_AO6;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_AQ;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_AX;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_A_CY;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_A_XOR;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_B;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_B1;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_B2;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_B3;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_B4;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_B5;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_B6;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_BMUX;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_BO5;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_BO6;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_BQ;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_BX;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_B_CY;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_B_XOR;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_C;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_C1;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_C2;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_C3;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_C4;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_C5;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_C6;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_CLK;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_CMUX;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_CO5;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_CO6;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_CQ;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_CX;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_C_CY;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_C_XOR;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_D;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_D1;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_D2;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_D3;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_D4;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_D5;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_D6;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_DO5;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_DO6;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_D_CY;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_D_XOR;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_A;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_A1;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_A2;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_A3;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_A4;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_A5;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_A6;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_AO5;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_AO6;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_A_CY;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_A_XOR;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_B;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_B1;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_B2;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_B3;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_B4;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_B5;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_B6;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_BO5;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_BO6;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_B_CY;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_B_XOR;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_C;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_C1;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_C2;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_C3;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_C4;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_C5;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_C6;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_CO5;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_CO6;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_C_CY;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_C_XOR;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_D;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_D1;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_D2;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_D3;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_D4;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_D5;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_D6;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_DO5;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_DO6;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_D_CY;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_D_XOR;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_A;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_A1;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_A2;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_A3;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_A4;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_A5;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_A6;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_AO5;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_AO6;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_AQ;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_A_CY;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_A_XOR;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_B;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_B1;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_B2;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_B3;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_B4;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_B5;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_B6;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_BO5;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_BO6;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_B_CY;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_B_XOR;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_C;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_C1;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_C2;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_C3;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_C4;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_C5;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_C6;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_CLK;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_CO5;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_CO6;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_C_CY;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_C_XOR;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_D;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_D1;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_D2;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_D3;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_D4;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_D5;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_D6;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_DO5;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_DO6;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_D_CY;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_D_XOR;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_A;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_A1;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_A2;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_A3;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_A4;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_A5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_A6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_AO5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_AO6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_A_CY;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_A_XOR;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_B;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_B1;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_B2;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_B3;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_B4;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_B5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_B6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_BO5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_BO6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_B_CY;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_B_XOR;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_C;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_C1;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_C2;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_C3;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_C4;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_C5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_C6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_CO5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_CO6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_C_CY;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_C_XOR;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_D;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_D1;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_D2;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_D3;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_D4;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_D5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_D6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_DO5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_DO6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_D_CY;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_D_XOR;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_A;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_A1;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_A2;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_A3;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_A4;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_A5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_A6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_AO5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_AO6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_AQ;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_A_CY;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_A_XOR;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_B;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_B1;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_B2;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_B3;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_B4;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_B5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_B5Q;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_B6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_BMUX;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_BO5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_BO6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_BQ;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_B_CY;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_B_XOR;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_C;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_C1;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_C2;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_C3;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_C4;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_C5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_C6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_CLK;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_CO5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_CO6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_C_CY;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_C_XOR;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_D;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_D1;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_D2;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_D3;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_D4;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_D5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_D6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_DO5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_DO6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_D_CY;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_D_XOR;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_A;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_A1;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_A2;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_A3;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_A4;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_A5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_A6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_AO5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_AO6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_AQ;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_A_CY;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_A_XOR;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_B;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_B1;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_B2;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_B3;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_B4;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_B5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_B6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_BO5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_BO6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_B_CY;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_B_XOR;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_C;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_C1;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_C2;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_C3;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_C4;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_C5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_C6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_CLK;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_CO5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_CO6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_C_CY;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_C_XOR;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_D;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_D1;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_D2;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_D3;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_D4;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_D5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_D6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_DO5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_DO6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_D_CY;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_D_XOR;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_A;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_A1;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_A2;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_A3;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_A4;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_A5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_A5Q;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_A6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_AMUX;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_AO5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_AO6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_AQ;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_A_CY;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_A_XOR;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_B;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_B1;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_B2;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_B3;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_B4;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_B5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_B6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_BO5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_BO6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_B_CY;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_B_XOR;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_C;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_C1;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_C2;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_C3;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_C4;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_C5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_C6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_CLK;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_CO5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_CO6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_C_CY;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_C_XOR;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_D;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_D1;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_D2;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_D3;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_D4;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_D5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_D6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_DO5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_DO6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_D_CY;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_D_XOR;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_SR;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_A;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_A1;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_A2;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_A3;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_A4;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_A5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_A6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_AO5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_AO6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_AQ;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_A_CY;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_A_XOR;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_B;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_B1;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_B2;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_B3;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_B4;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_B5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_B6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_BO5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_BO6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_BQ;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_B_CY;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_B_XOR;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_C;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_C1;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_C2;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_C3;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_C4;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_C5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_C5Q;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_C6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_CLK;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_CMUX;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_CO5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_CO6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_CQ;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_C_CY;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_C_XOR;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_D;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_D1;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_D2;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_D3;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_D4;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_D5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_D6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_DO5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_DO6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_DQ;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_D_CY;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_D_XOR;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_A;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_A1;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_A2;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_A3;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_A4;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_A5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_A6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_AMUX;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_AO5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_AO6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_A_CY;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_A_XOR;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_B;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_B1;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_B2;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_B3;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_B4;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_B5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_B5Q;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_B6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_BMUX;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_BO5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_BO6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_BQ;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_B_CY;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_B_XOR;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_C;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_C1;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_C2;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_C3;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_C4;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_C5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_C5Q;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_C6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_CLK;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_CMUX;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_CO5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_CO6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_CQ;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_C_CY;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_C_XOR;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_D;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_D1;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_D2;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_D3;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_D4;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_D5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_D6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_DO5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_DO6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_D_CY;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_D_XOR;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_SR;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_A;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_A1;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_A2;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_A3;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_A4;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_A5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_A6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_AO5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_AO6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_AQ;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_A_CY;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_A_XOR;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_B;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_B1;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_B2;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_B3;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_B4;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_B5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_B6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_BO5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_BO6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_BQ;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_B_CY;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_B_XOR;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_C;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_C1;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_C2;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_C3;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_C4;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_C5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_C6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_CLK;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_CO5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_CO6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_CQ;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_C_CY;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_C_XOR;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_D;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_D1;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_D2;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_D3;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_D4;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_D5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_D5Q;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_D6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_DMUX;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_DO5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_DO6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_DQ;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_D_CY;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_D_XOR;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_A;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_A1;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_A2;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_A3;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_A4;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_A5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_A6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_AO5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_AO6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_AQ;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_A_CY;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_A_XOR;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_B;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_B1;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_B2;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_B3;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_B4;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_B5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_B6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_BO5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_BO6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_BQ;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_B_CY;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_B_XOR;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_C;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_C1;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_C2;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_C3;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_C4;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_C5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_C6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_CLK;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_CO5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_CO6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_CQ;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_C_CY;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_C_XOR;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_D;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_D1;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_D2;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_D3;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_D4;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_D5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_D6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_DO5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_DO6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_DQ;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_D_CY;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_D_XOR;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_A;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_A1;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_A2;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_A3;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_A4;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_A5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_A6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_AO5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_AO6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_AQ;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_A_CY;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_A_XOR;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_B;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_B1;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_B2;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_B3;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_B4;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_B5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_B5Q;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_B6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_BMUX;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_BO5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_BO6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_BQ;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_B_CY;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_B_XOR;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_C;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_C1;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_C2;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_C3;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_C4;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_C5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_C5Q;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_C6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_CLK;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_CMUX;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_CO5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_CO6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_CQ;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_C_CY;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_C_XOR;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_D;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_D1;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_D2;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_D3;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_D4;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_D5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_D5Q;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_D6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_DMUX;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_DO5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_DO6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_DQ;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_D_CY;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_D_XOR;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_A;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_A1;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_A2;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_A3;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_A4;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_A5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_A6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_AO5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_AO6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_AQ;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_A_CY;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_A_XOR;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_B;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_B1;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_B2;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_B3;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_B4;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_B5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_B6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_BO5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_BO6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_BQ;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_B_CY;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_B_XOR;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_C;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_C1;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_C2;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_C3;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_C4;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_C5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_C6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_CLK;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_CO5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_CO6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_CQ;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_C_CY;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_C_XOR;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_D;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_D1;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_D2;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_D3;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_D4;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_D5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_D6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_DO5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_DO6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_DQ;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_D_CY;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_D_XOR;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_A;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_A1;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_A2;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_A3;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_A4;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_A5;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_A6;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_AO5;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_AO6;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_AQ;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_A_CY;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_A_XOR;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_B;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_B1;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_B2;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_B3;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_B4;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_B5;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_B5Q;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_B6;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_BMUX;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_BO5;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_BO6;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_BQ;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_B_CY;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_B_XOR;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_C;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_C1;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_C2;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_C3;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_C4;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_C5;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_C6;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_CLK;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_CO5;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_CO6;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_CQ;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_C_CY;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_C_XOR;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_D;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_D1;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_D2;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_D3;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_D4;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_D5;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_D6;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_DO5;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_DO6;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_DQ;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_D_CY;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X6Y145_D_XOR;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_A;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_A1;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_A2;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_A3;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_A4;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_A5;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_A5Q;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_A6;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_AMUX;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_AO5;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_AO6;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_AQ;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_A_CY;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_A_XOR;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_B;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_B1;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_B2;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_B3;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_B4;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_B5;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_B6;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_BMUX;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_BO5;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_BO6;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_B_CY;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_B_XOR;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_C;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_C1;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_C2;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_C3;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_C4;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_C5;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_C6;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_CLK;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_CO5;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_CO6;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_C_CY;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_C_XOR;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_D;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_D1;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_D2;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_D3;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_D4;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_D5;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_D6;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_DO5;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_DO6;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_D_CY;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_D_XOR;
  wire [0:0] CLBLM_R_X5Y145_SLICE_X7Y145_SR;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_A;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_A1;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_A2;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_A3;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_A4;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_A5;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_A6;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_AO5;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_AO6;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_AQ;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_A_CY;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_A_XOR;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_B;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_B1;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_B2;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_B3;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_B4;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_B5;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_B5Q;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_B6;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_BMUX;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_BO5;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_BO6;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_BQ;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_B_CY;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_B_XOR;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_C;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_C1;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_C2;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_C3;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_C4;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_C5;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_C6;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_CLK;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_CMUX;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_CO5;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_CO6;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_C_CY;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_C_XOR;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_D;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_D1;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_D2;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_D3;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_D4;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_D5;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_D6;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_DO5;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_DO6;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_D_CY;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_D_XOR;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_SR;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_A;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_A1;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_A2;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_A3;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_A4;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_A5;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_A6;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_AO5;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_AO6;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_AQ;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_A_CY;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_A_XOR;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_B;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_B1;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_B2;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_B3;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_B4;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_B5;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_B5Q;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_B6;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_BMUX;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_BO5;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_BO6;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_BQ;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_B_CY;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_B_XOR;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_C;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_C1;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_C2;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_C3;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_C4;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_C5;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_C6;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_CLK;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_CO5;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_CO6;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_CQ;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_C_CY;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_C_XOR;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_D;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_D1;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_D2;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_D3;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_D4;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_D5;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_D6;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_DO5;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_DO6;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_DQ;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_D_CY;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_D_XOR;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_A;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_A1;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_A2;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_A3;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_A4;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_A5;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_A6;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_AO5;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_AO6;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_AQ;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_A_CY;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_A_XOR;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_B;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_B1;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_B2;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_B3;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_B4;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_B5;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_B5Q;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_B6;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_BMUX;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_BO5;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_BO6;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_BQ;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_B_CY;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_B_XOR;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_C;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_C1;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_C2;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_C3;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_C4;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_C5;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_C6;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_CLK;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_CO5;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_CO6;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_CQ;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_C_CY;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_C_XOR;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_D;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_D1;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_D2;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_D3;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_D4;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_D5;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_D6;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_DO5;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_DO6;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_DQ;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_D_CY;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_D_XOR;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_A;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_A1;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_A2;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_A3;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_A4;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_A5;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_A5Q;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_A6;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_AMUX;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_AO5;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_AO6;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_AQ;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_A_CY;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_A_XOR;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_B;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_B1;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_B2;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_B3;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_B4;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_B5;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_B5Q;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_B6;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_BMUX;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_BO5;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_BO6;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_BQ;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_B_CY;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_B_XOR;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_C;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_C1;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_C2;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_C3;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_C4;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_C5;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_C5Q;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_C6;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_CLK;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_CMUX;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_CO5;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_CO6;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_CQ;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_C_CY;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_C_XOR;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_D;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_D1;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_D2;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_D3;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_D4;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_D5;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_D6;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_DO5;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_DO6;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_D_CY;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_D_XOR;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_SR;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_A;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_A1;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_A2;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_A3;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_A4;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_A5;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_A6;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_AMUX;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_AO5;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_AO6;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_AQ;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_AX;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_A_CY;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_A_XOR;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_B;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_B1;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_B2;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_B3;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_B4;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_B5;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_B5Q;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_B6;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_BMUX;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_BO5;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_BO6;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_BQ;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_B_CY;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_B_XOR;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_C;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_C1;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_C2;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_C3;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_C4;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_C5;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_C6;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_CLK;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_CMUX;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_CO5;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_CO6;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_C_CY;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_C_XOR;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_D;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_D1;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_D2;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_D3;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_D4;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_D5;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_D6;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_DO5;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_DO6;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_D_CY;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_D_XOR;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_SR;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_A;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_A1;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_A2;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_A3;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_A4;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_A5;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_A6;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_AO5;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_AO6;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_AQ;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_AX;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_A_CY;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_A_XOR;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_B;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_B1;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_B2;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_B3;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_B4;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_B5;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_B6;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_BO5;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_BO6;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_B_CY;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_B_XOR;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_C;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_C1;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_C2;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_C3;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_C4;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_C5;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_C6;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_CLK;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_CO5;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_CO6;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_C_CY;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_C_XOR;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_D;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_D1;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_D2;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_D3;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_D4;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_D5;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_D6;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_DO5;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_DO6;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_D_CY;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_D_XOR;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_SR;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_A;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_A1;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_A2;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_A3;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_A4;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_A5;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_A5Q;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_A6;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_AMUX;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_AO5;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_AO6;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_AQ;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_A_CY;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_A_XOR;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_B;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_B1;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_B2;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_B3;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_B4;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_B5;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_B6;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_BO5;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_BO6;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_BQ;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_B_CY;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_B_XOR;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_C;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_C1;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_C2;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_C3;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_C4;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_C5;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_C6;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_CLK;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_CO5;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_CO6;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_CQ;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_C_CY;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_C_XOR;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_D;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_D1;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_D2;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_D3;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_D4;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_D5;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_D5Q;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_D6;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_DMUX;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_DO5;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_DO6;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_DQ;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_D_CY;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_D_XOR;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_A;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_A1;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_A2;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_A3;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_A4;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_A5;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_A6;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_AO5;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_AO6;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_AQ;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_A_CY;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_A_XOR;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_B;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_B1;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_B2;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_B3;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_B4;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_B5;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_B5Q;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_B6;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_BMUX;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_BO5;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_BO6;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_BQ;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_B_CY;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_B_XOR;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_C;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_C1;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_C2;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_C3;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_C4;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_C5;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_C5Q;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_C6;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_CLK;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_CMUX;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_CO5;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_CO6;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_CQ;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_C_CY;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_C_XOR;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_D;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_D1;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_D2;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_D3;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_D4;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_D5;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_D5Q;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_D6;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_DMUX;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_DO5;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_DO6;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_DQ;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_D_CY;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_D_XOR;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_A;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_A1;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_A2;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_A3;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_A4;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_A5;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_A5Q;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_A6;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_AMUX;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_AO5;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_AO6;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_AQ;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_A_CY;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_A_XOR;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_B;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_B1;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_B2;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_B3;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_B4;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_B5;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_B6;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_BO5;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_BO6;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_BQ;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_B_CY;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_B_XOR;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_C;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_C1;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_C2;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_C3;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_C4;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_C5;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_C5Q;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_C6;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_CLK;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_CMUX;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_CO5;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_CO6;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_CQ;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_C_CY;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_C_XOR;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_D;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_D1;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_D2;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_D3;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_D4;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_D5;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_D6;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_DO5;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_DO6;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_DQ;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_D_CY;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_D_XOR;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_A;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_A1;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_A2;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_A3;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_A4;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_A5;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_A5Q;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_A6;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_AMUX;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_AO5;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_AO6;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_AQ;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_A_CY;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_A_XOR;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_B;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_B1;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_B2;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_B3;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_B4;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_B5;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_B6;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_BMUX;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_BO5;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_BO6;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_B_CY;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_B_XOR;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_C;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_C1;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_C2;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_C3;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_C4;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_C5;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_C6;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_CLK;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_CO5;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_CO6;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_C_CY;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_C_XOR;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_D;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_D1;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_D2;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_D3;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_D4;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_D5;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_D6;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_DO5;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_DO6;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_D_CY;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_D_XOR;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_SR;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_A;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_A1;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_A2;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_A3;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_A4;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_A5;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_A5Q;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_A6;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_AMUX;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_AO5;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_AO6;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_AQ;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_A_CY;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_A_XOR;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_B;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_B1;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_B2;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_B3;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_B4;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_B5;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_B5Q;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_B6;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_BMUX;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_BO5;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_BO6;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_BQ;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_B_CY;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_B_XOR;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_C;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_C1;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_C2;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_C3;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_C4;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_C5;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_C6;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_CLK;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_CO5;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_CO6;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_CQ;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_C_CY;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_C_XOR;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_D;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_D1;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_D2;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_D3;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_D4;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_D5;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_D5Q;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_D6;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_DMUX;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_DO5;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_DO6;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_DQ;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_D_CY;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_D_XOR;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_A;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_A1;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_A2;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_A3;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_A4;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_A5;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_A5Q;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_A6;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_AMUX;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_AO5;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_AO6;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_AQ;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_A_CY;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_A_XOR;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_B;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_B1;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_B2;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_B3;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_B4;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_B5;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_B6;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_BMUX;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_BO5;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_BO6;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_B_CY;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_B_XOR;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_C;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_C1;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_C2;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_C3;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_C4;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_C5;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_C6;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_CLK;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_CO5;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_CO6;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_C_CY;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_C_XOR;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_D;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_D1;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_D2;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_D3;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_D4;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_D5;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_D6;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_DO5;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_DO6;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_D_CY;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_D_XOR;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_SR;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_A;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_A1;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_A2;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_A3;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_A4;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_A5;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_A5Q;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_A6;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_AMUX;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_AO5;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_AO6;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_AQ;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_A_CY;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_A_XOR;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_B;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_B1;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_B2;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_B3;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_B4;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_B5;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_B5Q;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_B6;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_BMUX;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_BO5;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_BO6;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_BQ;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_B_CY;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_B_XOR;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_C;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_C1;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_C2;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_C3;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_C4;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_C5;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_C5Q;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_C6;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_CLK;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_CMUX;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_CO5;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_CO6;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_CQ;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_C_CY;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_C_XOR;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_D;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_D1;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_D2;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_D3;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_D4;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_D5;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_D6;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_DO5;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_DO6;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_DQ;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_D_CY;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_D_XOR;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_A;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_A1;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_A2;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_A3;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_A4;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_A5;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_A6;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_AO5;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_AO6;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_AQ;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_A_CY;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_A_XOR;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_B;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_B1;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_B2;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_B3;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_B4;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_B5;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_B6;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_BO5;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_BO6;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_BQ;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_B_CY;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_B_XOR;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_C;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_C1;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_C2;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_C3;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_C4;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_C5;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_C6;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_CLK;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_CO5;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_CO6;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_CQ;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_C_CY;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_C_XOR;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_D;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_D1;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_D2;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_D3;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_D4;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_D5;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_D5Q;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_D6;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_DMUX;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_DO5;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_DO6;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_DQ;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_D_CY;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_D_XOR;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_A;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_A1;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_A2;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_A3;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_A4;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_A5;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_A6;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_AO5;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_AO6;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_AQ;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_A_CY;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_A_XOR;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_B;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_B1;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_B2;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_B3;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_B4;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_B5;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_B6;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_BO5;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_BO6;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_BQ;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_B_CY;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_B_XOR;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_C;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_C1;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_C2;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_C3;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_C4;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_C5;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_C6;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_CLK;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_CO5;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_CO6;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_CQ;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_C_CY;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_C_XOR;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_D;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_D1;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_D2;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_D3;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_D4;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_D5;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_D6;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_DO5;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_DO6;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_DQ;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_D_CY;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_D_XOR;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_A;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_A1;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_A2;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_A3;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_A4;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_A5;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_A5Q;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_A6;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_AMUX;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_AO5;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_AO6;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_AQ;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_A_CY;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_A_XOR;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_B;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_B1;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_B2;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_B3;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_B4;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_B5;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_B6;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_BO5;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_BO6;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_B_CY;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_B_XOR;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_C;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_C1;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_C2;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_C3;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_C4;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_C5;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_C6;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_CLK;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_CO5;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_CO6;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_C_CY;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_C_XOR;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_D;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_D1;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_D2;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_D3;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_D4;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_D5;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_D6;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_DO5;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_DO6;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_D_CY;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_D_XOR;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_SR;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_A;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_A1;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_A2;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_A3;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_A4;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_A5;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_A6;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_AO5;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_AO6;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_AQ;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_A_CY;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_A_XOR;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_B;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_B1;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_B2;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_B3;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_B4;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_B5;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_B6;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_BO5;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_BO6;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_B_CY;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_B_XOR;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_C;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_C1;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_C2;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_C3;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_C4;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_C5;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_C6;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_CLK;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_CO5;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_CO6;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_C_CY;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_C_XOR;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_D;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_D1;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_D2;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_D3;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_D4;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_D5;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_D6;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_DO5;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_DO6;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_D_CY;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_D_XOR;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_A;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_A1;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_A2;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_A3;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_A4;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_A5;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_A6;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_AO5;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_AO6;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_AQ;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_A_CY;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_A_XOR;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_B;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_B1;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_B2;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_B3;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_B4;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_B5;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_B6;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_BO5;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_BO6;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_BQ;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_B_CY;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_B_XOR;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_C;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_C1;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_C2;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_C3;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_C4;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_C5;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_C6;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_CLK;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_CO5;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_CO6;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_CQ;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_C_CY;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_C_XOR;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_D;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_D1;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_D2;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_D3;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_D4;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_D5;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_D6;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_DO5;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_DO6;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_DQ;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_D_CY;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_D_XOR;
  wire [0:0] CLBLM_R_X5Y159_SLICE_X6Y159_A;
  wire [0:0] CLBLM_R_X5Y159_SLICE_X6Y159_A1;
  wire [0:0] CLBLM_R_X5Y159_SLICE_X6Y159_A2;
  wire [0:0] CLBLM_R_X5Y159_SLICE_X6Y159_A3;
  wire [0:0] CLBLM_R_X5Y159_SLICE_X6Y159_A4;
  wire [0:0] CLBLM_R_X5Y159_SLICE_X6Y159_A5;
  wire [0:0] CLBLM_R_X5Y159_SLICE_X6Y159_A6;
  wire [0:0] CLBLM_R_X5Y159_SLICE_X6Y159_AO5;
  wire [0:0] CLBLM_R_X5Y159_SLICE_X6Y159_AO6;
  wire [0:0] CLBLM_R_X5Y159_SLICE_X6Y159_A_CY;
  wire [0:0] CLBLM_R_X5Y159_SLICE_X6Y159_A_XOR;
  wire [0:0] CLBLM_R_X5Y159_SLICE_X6Y159_B;
  wire [0:0] CLBLM_R_X5Y159_SLICE_X6Y159_B1;
  wire [0:0] CLBLM_R_X5Y159_SLICE_X6Y159_B2;
  wire [0:0] CLBLM_R_X5Y159_SLICE_X6Y159_B3;
  wire [0:0] CLBLM_R_X5Y159_SLICE_X6Y159_B4;
  wire [0:0] CLBLM_R_X5Y159_SLICE_X6Y159_B5;
  wire [0:0] CLBLM_R_X5Y159_SLICE_X6Y159_B6;
  wire [0:0] CLBLM_R_X5Y159_SLICE_X6Y159_BO5;
  wire [0:0] CLBLM_R_X5Y159_SLICE_X6Y159_BO6;
  wire [0:0] CLBLM_R_X5Y159_SLICE_X6Y159_B_CY;
  wire [0:0] CLBLM_R_X5Y159_SLICE_X6Y159_B_XOR;
  wire [0:0] CLBLM_R_X5Y159_SLICE_X6Y159_C;
  wire [0:0] CLBLM_R_X5Y159_SLICE_X6Y159_C1;
  wire [0:0] CLBLM_R_X5Y159_SLICE_X6Y159_C2;
  wire [0:0] CLBLM_R_X5Y159_SLICE_X6Y159_C3;
  wire [0:0] CLBLM_R_X5Y159_SLICE_X6Y159_C4;
  wire [0:0] CLBLM_R_X5Y159_SLICE_X6Y159_C5;
  wire [0:0] CLBLM_R_X5Y159_SLICE_X6Y159_C6;
  wire [0:0] CLBLM_R_X5Y159_SLICE_X6Y159_CO5;
  wire [0:0] CLBLM_R_X5Y159_SLICE_X6Y159_CO6;
  wire [0:0] CLBLM_R_X5Y159_SLICE_X6Y159_C_CY;
  wire [0:0] CLBLM_R_X5Y159_SLICE_X6Y159_C_XOR;
  wire [0:0] CLBLM_R_X5Y159_SLICE_X6Y159_D;
  wire [0:0] CLBLM_R_X5Y159_SLICE_X6Y159_D1;
  wire [0:0] CLBLM_R_X5Y159_SLICE_X6Y159_D2;
  wire [0:0] CLBLM_R_X5Y159_SLICE_X6Y159_D3;
  wire [0:0] CLBLM_R_X5Y159_SLICE_X6Y159_D4;
  wire [0:0] CLBLM_R_X5Y159_SLICE_X6Y159_D5;
  wire [0:0] CLBLM_R_X5Y159_SLICE_X6Y159_D6;
  wire [0:0] CLBLM_R_X5Y159_SLICE_X6Y159_DO5;
  wire [0:0] CLBLM_R_X5Y159_SLICE_X6Y159_DO6;
  wire [0:0] CLBLM_R_X5Y159_SLICE_X6Y159_D_CY;
  wire [0:0] CLBLM_R_X5Y159_SLICE_X6Y159_D_XOR;
  wire [0:0] CLBLM_R_X5Y159_SLICE_X7Y159_A;
  wire [0:0] CLBLM_R_X5Y159_SLICE_X7Y159_A1;
  wire [0:0] CLBLM_R_X5Y159_SLICE_X7Y159_A2;
  wire [0:0] CLBLM_R_X5Y159_SLICE_X7Y159_A3;
  wire [0:0] CLBLM_R_X5Y159_SLICE_X7Y159_A4;
  wire [0:0] CLBLM_R_X5Y159_SLICE_X7Y159_A5;
  wire [0:0] CLBLM_R_X5Y159_SLICE_X7Y159_A6;
  wire [0:0] CLBLM_R_X5Y159_SLICE_X7Y159_AO5;
  wire [0:0] CLBLM_R_X5Y159_SLICE_X7Y159_AO6;
  wire [0:0] CLBLM_R_X5Y159_SLICE_X7Y159_A_CY;
  wire [0:0] CLBLM_R_X5Y159_SLICE_X7Y159_A_XOR;
  wire [0:0] CLBLM_R_X5Y159_SLICE_X7Y159_B;
  wire [0:0] CLBLM_R_X5Y159_SLICE_X7Y159_B1;
  wire [0:0] CLBLM_R_X5Y159_SLICE_X7Y159_B2;
  wire [0:0] CLBLM_R_X5Y159_SLICE_X7Y159_B3;
  wire [0:0] CLBLM_R_X5Y159_SLICE_X7Y159_B4;
  wire [0:0] CLBLM_R_X5Y159_SLICE_X7Y159_B5;
  wire [0:0] CLBLM_R_X5Y159_SLICE_X7Y159_B6;
  wire [0:0] CLBLM_R_X5Y159_SLICE_X7Y159_BO5;
  wire [0:0] CLBLM_R_X5Y159_SLICE_X7Y159_BO6;
  wire [0:0] CLBLM_R_X5Y159_SLICE_X7Y159_B_CY;
  wire [0:0] CLBLM_R_X5Y159_SLICE_X7Y159_B_XOR;
  wire [0:0] CLBLM_R_X5Y159_SLICE_X7Y159_C;
  wire [0:0] CLBLM_R_X5Y159_SLICE_X7Y159_C1;
  wire [0:0] CLBLM_R_X5Y159_SLICE_X7Y159_C2;
  wire [0:0] CLBLM_R_X5Y159_SLICE_X7Y159_C3;
  wire [0:0] CLBLM_R_X5Y159_SLICE_X7Y159_C4;
  wire [0:0] CLBLM_R_X5Y159_SLICE_X7Y159_C5;
  wire [0:0] CLBLM_R_X5Y159_SLICE_X7Y159_C6;
  wire [0:0] CLBLM_R_X5Y159_SLICE_X7Y159_CO5;
  wire [0:0] CLBLM_R_X5Y159_SLICE_X7Y159_CO6;
  wire [0:0] CLBLM_R_X5Y159_SLICE_X7Y159_C_CY;
  wire [0:0] CLBLM_R_X5Y159_SLICE_X7Y159_C_XOR;
  wire [0:0] CLBLM_R_X5Y159_SLICE_X7Y159_D;
  wire [0:0] CLBLM_R_X5Y159_SLICE_X7Y159_D1;
  wire [0:0] CLBLM_R_X5Y159_SLICE_X7Y159_D2;
  wire [0:0] CLBLM_R_X5Y159_SLICE_X7Y159_D3;
  wire [0:0] CLBLM_R_X5Y159_SLICE_X7Y159_D4;
  wire [0:0] CLBLM_R_X5Y159_SLICE_X7Y159_D5;
  wire [0:0] CLBLM_R_X5Y159_SLICE_X7Y159_D6;
  wire [0:0] CLBLM_R_X5Y159_SLICE_X7Y159_DO5;
  wire [0:0] CLBLM_R_X5Y159_SLICE_X7Y159_DO6;
  wire [0:0] CLBLM_R_X5Y159_SLICE_X7Y159_D_CY;
  wire [0:0] CLBLM_R_X5Y159_SLICE_X7Y159_D_XOR;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_A;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_A1;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_A2;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_A3;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_A4;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_A5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_A6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_AO5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_AO6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_AQ;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_A_CY;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_A_XOR;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_B;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_B1;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_B2;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_B3;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_B4;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_B5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_B6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_BO5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_BO6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_B_CY;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_B_XOR;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_C;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_C1;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_C2;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_C3;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_C4;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_C5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_C6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_CLK;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_CO5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_CO6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_C_CY;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_C_XOR;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_D;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_D1;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_D2;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_D3;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_D4;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_D5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_D6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_DO5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_DO6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_D_CY;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_D_XOR;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_A;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_A1;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_A2;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_A3;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_A4;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_A5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_A6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_AO5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_AO6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_AQ;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_A_CY;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_A_XOR;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_B;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_B1;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_B2;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_B3;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_B4;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_B5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_B6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_BO5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_BO6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_B_CY;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_B_XOR;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_C;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_C1;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_C2;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_C3;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_C4;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_C5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_C6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_CLK;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_CO5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_CO6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_C_CY;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_C_XOR;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_D;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_D1;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_D2;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_D3;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_D4;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_D5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_D6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_DO5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_DO6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_D_CY;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_D_XOR;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_A;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_A1;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_A2;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_A3;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_A4;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_A5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_A5Q;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_A6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_AMUX;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_AO5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_AO6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_AQ;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_A_CY;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_A_XOR;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_B;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_B1;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_B2;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_B3;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_B4;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_B5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_B5Q;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_B6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_BMUX;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_BO5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_BO6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_BQ;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_B_CY;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_B_XOR;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_C;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_C1;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_C2;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_C3;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_C4;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_C5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_C6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_CLK;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_CO5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_CO6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_C_CY;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_C_XOR;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_D;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_D1;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_D2;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_D3;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_D4;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_D5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_D6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_DO5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_DO6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_D_CY;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_D_XOR;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_A;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_A1;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_A2;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_A3;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_A4;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_A5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_A5Q;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_A6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_AMUX;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_AO5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_AO6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_AQ;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_AX;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_A_CY;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_A_XOR;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_B;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_B1;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_B2;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_B3;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_B4;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_B5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_B6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_BO5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_BO6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_BQ;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_B_CY;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_B_XOR;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_C;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_C1;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_C2;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_C3;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_C4;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_C5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_C6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_CLK;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_CO5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_CO6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_CQ;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_C_CY;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_C_XOR;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_D;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_D1;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_D2;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_D3;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_D4;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_D5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_D5Q;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_D6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_DMUX;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_DO5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_DO6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_DQ;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_D_CY;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_D_XOR;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_A;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_A1;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_A2;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_A3;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_A4;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_A5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_A6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_AO5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_AO6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_AQ;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_A_CY;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_A_XOR;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_B;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_B1;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_B2;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_B3;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_B4;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_B5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_B6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_BO5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_BO6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_BQ;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_B_CY;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_B_XOR;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_C;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_C1;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_C2;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_C3;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_C4;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_C5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_C6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_CLK;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_CO5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_CO6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_CQ;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_C_CY;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_C_XOR;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_D;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_D1;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_D2;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_D3;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_D4;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_D5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_D6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_DO5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_DO6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_DQ;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_D_CY;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_D_XOR;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_A;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_A1;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_A2;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_A3;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_A4;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_A5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_A6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_AO5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_AO6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_AQ;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_A_CY;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_A_XOR;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_B;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_B1;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_B2;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_B3;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_B4;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_B5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_B6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_BO5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_BO6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_BQ;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_B_CY;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_B_XOR;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_C;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_C1;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_C2;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_C3;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_C4;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_C5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_C6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_CLK;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_CO5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_CO6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_CQ;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_C_CY;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_C_XOR;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_D;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_D1;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_D2;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_D3;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_D4;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_D5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_D6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_DO5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_DO6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_DQ;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_D_CY;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_D_XOR;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_A;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_A1;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_A2;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_A3;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_A4;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_A5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_A5Q;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_A6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_AMUX;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_AO5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_AO6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_AQ;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_A_CY;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_A_XOR;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_B;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_B1;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_B2;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_B3;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_B4;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_B5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_B6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_BO5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_BO6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_BQ;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_BX;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_B_CY;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_B_XOR;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_C;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_C1;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_C2;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_C3;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_C4;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_C5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_C6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_CLK;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_CO5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_CO6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_C_CY;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_C_XOR;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_D;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_D1;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_D2;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_D3;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_D4;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_D5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_D6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_DO5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_DO6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_D_CY;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_D_XOR;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_SR;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_A;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_A1;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_A2;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_A3;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_A4;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_A5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_A5Q;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_A6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_AMUX;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_AO5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_AO6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_AQ;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_AX;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_A_CY;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_A_XOR;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_B;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_B1;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_B2;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_B3;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_B4;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_B5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_B5Q;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_B6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_BMUX;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_BO5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_BO6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_BQ;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_B_CY;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_B_XOR;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_C;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_C1;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_C2;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_C3;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_C4;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_C5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_C5Q;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_C6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_CLK;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_CMUX;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_CO5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_CO6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_CQ;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_C_CY;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_C_XOR;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_D;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_D1;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_D2;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_D3;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_D4;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_D5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_D5Q;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_D6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_DMUX;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_DO5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_DO6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_DQ;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_D_CY;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_D_XOR;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_A;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_A1;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_A2;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_A3;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_A4;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_A5;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_A6;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_AO5;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_AO6;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_AQ;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_A_CY;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_A_XOR;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_B;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_B1;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_B2;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_B3;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_B4;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_B5;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_B5Q;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_B6;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_BMUX;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_BO5;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_BO6;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_BQ;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_B_CY;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_B_XOR;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_C;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_C1;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_C2;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_C3;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_C4;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_C5;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_C5Q;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_C6;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_CLK;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_CMUX;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_CO5;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_CO6;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_CQ;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_C_CY;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_C_XOR;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_D;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_D1;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_D2;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_D3;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_D4;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_D5;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_D6;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_DO5;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_DO6;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_DQ;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_D_CY;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_D_XOR;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_A;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_A1;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_A2;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_A3;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_A4;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_A5;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_A6;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_AO5;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_AO6;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_AQ;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_A_CY;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_A_XOR;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_B;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_B1;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_B2;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_B3;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_B4;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_B5;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_B6;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_BO5;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_BO6;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_BQ;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_B_CY;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_B_XOR;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_C;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_C1;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_C2;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_C3;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_C4;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_C5;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_C6;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_CLK;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_CO5;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_CO6;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_CQ;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_C_CY;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_C_XOR;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_D;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_D1;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_D2;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_D3;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_D4;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_D5;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_D6;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_DO5;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_DO6;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_DQ;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_D_CY;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_D_XOR;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_A;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_A1;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_A2;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_A3;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_A4;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_A5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_A6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_AMUX;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_AO5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_AO6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_AX;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_A_CY;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_A_XOR;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_B;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_B1;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_B2;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_B3;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_B4;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_B5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_B6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_BO5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_BO6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_BQ;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_BX;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_B_CY;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_B_XOR;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_C;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_C1;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_C2;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_C3;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_C4;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_C5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_C6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_CE;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_CLK;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_CMUX;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_CO5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_CO6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_C_CY;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_C_XOR;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_D;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_D1;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_D2;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_D3;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_D4;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_D5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_D6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_DO5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_DO6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_D_CY;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_D_XOR;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_A;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_A1;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_A2;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_A3;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_A4;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_A5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_A6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_AMUX;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_AO5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_AO6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_A_CY;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_A_XOR;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_B;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_B1;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_B2;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_B3;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_B4;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_B5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_B5Q;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_B6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_BMUX;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_BO5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_BO6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_BQ;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_B_CY;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_B_XOR;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_C;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_C1;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_C2;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_C3;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_C4;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_C5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_C6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_CLK;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_CO5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_CO6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_C_CY;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_C_XOR;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_D;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_D1;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_D2;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_D3;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_D4;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_D5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_D6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_DO5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_DO6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_D_CY;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_D_XOR;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_SR;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_A;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_A1;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_A2;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_A3;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_A4;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_A5;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_A6;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_AO5;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_AO6;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_AQ;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_A_CY;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_A_XOR;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_B;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_B1;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_B2;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_B3;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_B4;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_B5;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_B6;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_BO5;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_BO6;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_BQ;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_B_CY;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_B_XOR;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_C;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_C1;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_C2;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_C3;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_C4;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_C5;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_C6;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_CLK;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_CO5;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_CO6;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_CQ;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_C_CY;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_C_XOR;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_D;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_D1;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_D2;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_D3;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_D4;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_D5;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_D5Q;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_D6;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_DMUX;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_DO5;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_DO6;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_DQ;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_D_CY;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_D_XOR;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_A;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_A1;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_A2;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_A3;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_A4;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_A5;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_A6;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_AO5;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_AO6;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_AQ;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_A_CY;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_A_XOR;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_B;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_B1;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_B2;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_B3;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_B4;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_B5;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_B6;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_BO5;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_BO6;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_BQ;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_B_CY;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_B_XOR;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_C;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_C1;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_C2;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_C3;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_C4;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_C5;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_C5Q;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_C6;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_CLK;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_CMUX;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_CO5;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_CO6;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_CQ;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_C_CY;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_C_XOR;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_D;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_D1;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_D2;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_D3;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_D4;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_D5;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_D6;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_DMUX;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_DO5;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_DO6;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_D_CY;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_D_XOR;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_A;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_A1;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_A2;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_A3;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_A4;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_A5;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_A6;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_AO5;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_AO6;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_AQ;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_A_CY;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_A_XOR;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_B;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_B1;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_B2;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_B3;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_B4;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_B5;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_B6;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_BMUX;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_BO5;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_BO6;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_B_CY;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_B_XOR;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_C;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_C1;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_C2;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_C3;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_C4;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_C5;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_C6;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_CLK;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_CO5;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_CO6;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_C_CY;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_C_XOR;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_D;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_D1;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_D2;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_D3;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_D4;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_D5;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_D6;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_DO5;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_DO6;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_D_CY;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_D_XOR;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_SR;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_A;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_A1;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_A2;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_A3;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_A4;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_A5;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_A6;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_AMUX;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_AO5;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_AO6;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_AQ;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_A_CY;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_A_XOR;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_B;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_B1;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_B2;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_B3;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_B4;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_B5;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_B5Q;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_B6;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_BMUX;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_BO5;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_BO6;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_BQ;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_B_CY;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_B_XOR;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_C;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_C1;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_C2;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_C3;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_C4;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_C5;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_C5Q;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_C6;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_CLK;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_CMUX;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_CO5;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_CO6;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_CQ;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_C_CY;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_C_XOR;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_D;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_D1;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_D2;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_D3;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_D4;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_D5;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_D6;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_DO5;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_DO6;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_D_CY;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_D_XOR;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_A;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_A1;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_A2;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_A3;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_A4;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_A5;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_A6;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_AO5;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_AO6;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_AQ;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_A_CY;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_A_XOR;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_B;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_B1;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_B2;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_B3;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_B4;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_B5;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_B6;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_BO5;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_BO6;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_BQ;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_B_CY;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_B_XOR;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_C;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_C1;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_C2;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_C3;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_C4;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_C5;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_C6;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_CLK;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_CO5;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_CO6;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_CQ;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_C_CY;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_C_XOR;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_D;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_D1;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_D2;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_D3;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_D4;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_D5;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_D6;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_DO5;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_DO6;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_DQ;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_D_CY;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_D_XOR;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_A;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_A1;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_A2;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_A3;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_A4;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_A5;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_A6;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_AMUX;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_AO5;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_AO6;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_AX;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_A_CY;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_A_XOR;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_B;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_B1;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_B2;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_B3;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_B4;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_B5;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_B6;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_BMUX;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_BO5;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_BO6;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_BQ;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_BX;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_B_CY;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_B_XOR;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_C;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_C1;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_C2;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_C3;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_C4;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_C5;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_C5Q;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_C6;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_CE;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_CLK;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_CMUX;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_CO5;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_CO6;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_CQ;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_CX;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_C_CY;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_C_XOR;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_D;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_D1;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_D2;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_D3;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_D4;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_D5;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_D6;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_DO5;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_DO6;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_DQ;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_DX;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_D_CY;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_D_XOR;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_A;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_A1;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_A2;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_A3;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_A4;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_A5;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_A6;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_AO5;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_AO6;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_AQ;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_A_CY;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_A_XOR;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_B;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_B1;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_B2;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_B3;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_B4;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_B5;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_B6;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_BO5;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_BO6;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_BQ;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_B_CY;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_B_XOR;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_C;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_C1;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_C2;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_C3;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_C4;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_C5;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_C5Q;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_C6;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_CLK;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_CMUX;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_CO5;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_CO6;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_CQ;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_C_CY;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_C_XOR;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_D;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_D1;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_D2;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_D3;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_D4;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_D5;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_D5Q;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_D6;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_DMUX;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_DO5;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_DO6;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_DQ;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_D_CY;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_D_XOR;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_A;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_A1;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_A2;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_A3;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_A4;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_A5;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_A6;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_AO5;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_AO6;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_AQ;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_A_CY;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_A_XOR;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_B;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_B1;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_B2;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_B3;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_B4;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_B5;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_B5Q;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_B6;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_BMUX;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_BO5;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_BO6;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_BQ;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_B_CY;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_B_XOR;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_C;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_C1;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_C2;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_C3;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_C4;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_C5;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_C5Q;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_C6;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_CLK;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_CMUX;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_CO5;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_CO6;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_CQ;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_C_CY;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_C_XOR;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_D;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_D1;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_D2;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_D3;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_D4;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_D5;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_D6;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_DO5;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_DO6;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_DQ;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_D_CY;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_D_XOR;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_A;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_A1;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_A2;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_A3;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_A4;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_A5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_A6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_AO5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_AO6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_AQ;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_A_CY;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_A_XOR;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_B;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_B1;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_B2;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_B3;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_B4;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_B5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_B6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_BO5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_BO6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_BQ;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_B_CY;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_B_XOR;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_C;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_C1;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_C2;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_C3;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_C4;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_C5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_C5Q;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_C6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_CLK;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_CMUX;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_CO5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_CO6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_CQ;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_C_CY;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_C_XOR;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_D;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_D1;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_D2;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_D3;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_D4;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_D5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_D6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_DMUX;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_DO5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_DO6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_D_CY;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_D_XOR;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_A;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_A1;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_A2;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_A3;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_A4;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_A5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_A6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_AO5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_AO6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_AQ;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_A_CY;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_A_XOR;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_B;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_B1;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_B2;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_B3;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_B4;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_B5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_B6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_BO5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_BO6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_BQ;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_B_CY;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_B_XOR;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_C;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_C1;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_C2;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_C3;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_C4;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_C5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_C6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_CLK;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_CO5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_CO6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_CQ;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_C_CY;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_C_XOR;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_D;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_D1;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_D2;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_D3;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_D4;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_D5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_D6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_DO5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_DO6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_DQ;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_D_CY;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_D_XOR;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_A;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_A1;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_A2;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_A3;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_A4;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_A5;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_A6;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_AO5;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_AO6;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_AQ;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_A_CY;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_A_XOR;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_B;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_B1;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_B2;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_B3;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_B4;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_B5;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_B6;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_BO5;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_BO6;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_BQ;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_B_CY;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_B_XOR;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_C;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_C1;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_C2;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_C3;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_C4;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_C5;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_C6;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_CLK;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_CO5;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_CO6;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_CQ;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_C_CY;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_C_XOR;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_D;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_D1;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_D2;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_D3;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_D4;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_D5;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_D6;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_DO5;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_DO6;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_D_CY;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_D_XOR;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_A;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_A1;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_A2;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_A3;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_A4;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_A5;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_A6;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_AO5;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_AO6;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_AQ;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_A_CY;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_A_XOR;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_B;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_B1;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_B2;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_B3;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_B4;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_B5;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_B6;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_BO5;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_BO6;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_BQ;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_B_CY;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_B_XOR;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_C;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_C1;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_C2;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_C3;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_C4;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_C5;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_C5Q;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_C6;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_CLK;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_CMUX;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_CO5;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_CO6;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_CQ;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_C_CY;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_C_XOR;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_D;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_D1;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_D2;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_D3;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_D4;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_D5;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_D5Q;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_D6;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_DMUX;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_DO5;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_DO6;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_DQ;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_D_CY;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_D_XOR;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_A;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_A1;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_A2;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_A3;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_A4;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_A5;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_A6;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_AO5;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_AO6;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_AQ;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_A_CY;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_A_XOR;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_B;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_B1;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_B2;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_B3;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_B4;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_B5;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_B6;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_BMUX;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_BO5;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_BO6;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_B_CY;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_B_XOR;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_C;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_C1;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_C2;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_C3;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_C4;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_C5;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_C6;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_CLK;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_CMUX;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_CO5;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_CO6;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_C_CY;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_C_XOR;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_D;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_D1;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_D2;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_D3;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_D4;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_D5;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_D6;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_DMUX;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_DO5;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_DO6;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_D_CY;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_D_XOR;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_SR;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_A;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_A1;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_A2;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_A3;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_A4;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_A5;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_A5Q;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_A6;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_AMUX;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_AO5;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_AO6;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_AQ;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_AX;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_A_CY;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_A_XOR;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_B;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_B1;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_B2;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_B3;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_B4;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_B5;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_B6;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_BO5;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_BO6;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_BQ;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_B_CY;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_B_XOR;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_C;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_C1;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_C2;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_C3;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_C4;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_C5;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_C6;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_CLK;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_CO5;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_CO6;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_CQ;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_C_CY;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_C_XOR;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_D;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_D1;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_D2;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_D3;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_D4;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_D5;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_D6;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_DMUX;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_DO5;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_DO6;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_D_CY;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_D_XOR;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_A;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_A1;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_A2;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_A3;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_A4;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_A5;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_A6;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_AO5;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_AO6;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_AQ;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_A_CY;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_A_XOR;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_B;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_B1;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_B2;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_B3;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_B4;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_B5;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_B6;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_BO5;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_BO6;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_BQ;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_B_CY;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_B_XOR;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_C;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_C1;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_C2;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_C3;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_C4;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_C5;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_C6;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_CLK;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_CO5;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_CO6;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_CQ;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_C_CY;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_C_XOR;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_D;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_D1;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_D2;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_D3;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_D4;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_D5;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_D6;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_DMUX;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_DO5;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_DO6;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_D_CY;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_D_XOR;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_A;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_A1;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_A2;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_A3;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_A4;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_A5;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_A6;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_AMUX;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_AO5;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_AO6;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_A_CY;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_A_XOR;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_B;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_B1;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_B2;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_B3;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_B4;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_B5;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_B6;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_BO5;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_BO6;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_B_CY;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_B_XOR;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_C;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_C1;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_C2;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_C3;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_C4;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_C5;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_C6;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_CO5;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_CO6;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_C_CY;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_C_XOR;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_D;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_D1;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_D2;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_D3;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_D4;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_D5;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_D6;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_DO5;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_DO6;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_D_CY;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_D_XOR;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_A;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_A1;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_A2;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_A3;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_A4;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_A5;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_A6;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_AO5;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_AO6;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_AQ;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_A_CY;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_A_XOR;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_B;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_B1;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_B2;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_B3;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_B4;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_B5;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_B6;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_BO5;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_BO6;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_BQ;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_B_CY;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_B_XOR;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_C;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_C1;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_C2;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_C3;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_C4;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_C5;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_C6;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_CLK;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_CO5;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_CO6;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_C_CY;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_C_XOR;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_D;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_D1;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_D2;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_D3;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_D4;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_D5;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_D6;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_DO5;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_DO6;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_D_CY;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_D_XOR;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_A;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_A1;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_A2;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_A3;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_A4;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_A5;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_A6;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_AMUX;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_AO5;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_AO6;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_A_CY;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_A_XOR;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_B;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_B1;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_B2;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_B3;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_B4;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_B5;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_B6;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_BO5;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_BO6;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_B_CY;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_B_XOR;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_C;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_C1;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_C2;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_C3;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_C4;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_C5;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_C6;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_CO5;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_CO6;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_C_CY;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_C_XOR;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_D;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_D1;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_D2;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_D3;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_D4;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_D5;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_D6;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_DO5;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_DO6;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_D_CY;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_D_XOR;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE1;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I1;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE1;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S1;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_CE;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_I;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  wire [0:0] CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_CE;
  wire [0:0] CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_I;
  wire [0:0] CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  wire [0:0] LIOB33_SING_X0Y100_IOB_X0Y100_O;
  wire [0:0] LIOB33_SING_X0Y149_IOB_X0Y149_O;
  wire [0:0] LIOB33_SING_X0Y150_IOB_X0Y150_O;
  wire [0:0] LIOB33_SING_X0Y199_IOB_X0Y199_O;
  wire [0:0] LIOB33_SING_X0Y50_IOB_X0Y50_I;
  wire [0:0] LIOB33_X0Y101_IOB_X0Y101_O;
  wire [0:0] LIOB33_X0Y101_IOB_X0Y102_O;
  wire [0:0] LIOB33_X0Y103_IOB_X0Y103_O;
  wire [0:0] LIOB33_X0Y103_IOB_X0Y104_O;
  wire [0:0] LIOB33_X0Y105_IOB_X0Y105_O;
  wire [0:0] LIOB33_X0Y105_IOB_X0Y106_O;
  wire [0:0] LIOB33_X0Y107_IOB_X0Y107_O;
  wire [0:0] LIOB33_X0Y107_IOB_X0Y108_O;
  wire [0:0] LIOB33_X0Y109_IOB_X0Y109_O;
  wire [0:0] LIOB33_X0Y109_IOB_X0Y110_O;
  wire [0:0] LIOB33_X0Y111_IOB_X0Y111_O;
  wire [0:0] LIOB33_X0Y111_IOB_X0Y112_O;
  wire [0:0] LIOB33_X0Y113_IOB_X0Y113_O;
  wire [0:0] LIOB33_X0Y113_IOB_X0Y114_O;
  wire [0:0] LIOB33_X0Y115_IOB_X0Y115_O;
  wire [0:0] LIOB33_X0Y115_IOB_X0Y116_O;
  wire [0:0] LIOB33_X0Y117_IOB_X0Y117_O;
  wire [0:0] LIOB33_X0Y117_IOB_X0Y118_O;
  wire [0:0] LIOB33_X0Y119_IOB_X0Y119_O;
  wire [0:0] LIOB33_X0Y119_IOB_X0Y120_O;
  wire [0:0] LIOB33_X0Y121_IOB_X0Y121_O;
  wire [0:0] LIOB33_X0Y121_IOB_X0Y122_O;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y123_O;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y124_O;
  wire [0:0] LIOB33_X0Y125_IOB_X0Y125_O;
  wire [0:0] LIOB33_X0Y125_IOB_X0Y126_O;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y127_O;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y128_O;
  wire [0:0] LIOB33_X0Y129_IOB_X0Y129_O;
  wire [0:0] LIOB33_X0Y129_IOB_X0Y130_O;
  wire [0:0] LIOB33_X0Y131_IOB_X0Y131_O;
  wire [0:0] LIOB33_X0Y131_IOB_X0Y132_O;
  wire [0:0] LIOB33_X0Y133_IOB_X0Y133_O;
  wire [0:0] LIOB33_X0Y133_IOB_X0Y134_O;
  wire [0:0] LIOB33_X0Y135_IOB_X0Y135_O;
  wire [0:0] LIOB33_X0Y135_IOB_X0Y136_O;
  wire [0:0] LIOB33_X0Y137_IOB_X0Y137_O;
  wire [0:0] LIOB33_X0Y137_IOB_X0Y138_O;
  wire [0:0] LIOB33_X0Y139_IOB_X0Y139_O;
  wire [0:0] LIOB33_X0Y139_IOB_X0Y140_O;
  wire [0:0] LIOB33_X0Y141_IOB_X0Y141_O;
  wire [0:0] LIOB33_X0Y141_IOB_X0Y142_O;
  wire [0:0] LIOB33_X0Y143_IOB_X0Y143_O;
  wire [0:0] LIOB33_X0Y145_IOB_X0Y145_O;
  wire [0:0] LIOB33_X0Y145_IOB_X0Y146_O;
  wire [0:0] LIOB33_X0Y147_IOB_X0Y147_O;
  wire [0:0] LIOB33_X0Y147_IOB_X0Y148_O;
  wire [0:0] LIOB33_X0Y151_IOB_X0Y151_O;
  wire [0:0] LIOB33_X0Y151_IOB_X0Y152_O;
  wire [0:0] LIOB33_X0Y153_IOB_X0Y153_O;
  wire [0:0] LIOB33_X0Y153_IOB_X0Y154_O;
  wire [0:0] LIOB33_X0Y155_IOB_X0Y155_O;
  wire [0:0] LIOB33_X0Y155_IOB_X0Y156_O;
  wire [0:0] LIOB33_X0Y157_IOB_X0Y157_O;
  wire [0:0] LIOB33_X0Y157_IOB_X0Y158_O;
  wire [0:0] LIOB33_X0Y159_IOB_X0Y159_O;
  wire [0:0] LIOB33_X0Y159_IOB_X0Y160_O;
  wire [0:0] LIOB33_X0Y161_IOB_X0Y161_O;
  wire [0:0] LIOB33_X0Y161_IOB_X0Y162_O;
  wire [0:0] LIOB33_X0Y163_IOB_X0Y163_O;
  wire [0:0] LIOB33_X0Y163_IOB_X0Y164_O;
  wire [0:0] LIOB33_X0Y165_IOB_X0Y165_O;
  wire [0:0] LIOB33_X0Y165_IOB_X0Y166_O;
  wire [0:0] LIOB33_X0Y167_IOB_X0Y167_O;
  wire [0:0] LIOB33_X0Y167_IOB_X0Y168_O;
  wire [0:0] LIOB33_X0Y169_IOB_X0Y169_O;
  wire [0:0] LIOB33_X0Y169_IOB_X0Y170_O;
  wire [0:0] LIOB33_X0Y171_IOB_X0Y171_O;
  wire [0:0] LIOB33_X0Y171_IOB_X0Y172_O;
  wire [0:0] LIOB33_X0Y173_IOB_X0Y173_O;
  wire [0:0] LIOB33_X0Y173_IOB_X0Y174_O;
  wire [0:0] LIOB33_X0Y175_IOB_X0Y175_O;
  wire [0:0] LIOB33_X0Y175_IOB_X0Y176_O;
  wire [0:0] LIOB33_X0Y177_IOB_X0Y177_O;
  wire [0:0] LIOB33_X0Y177_IOB_X0Y178_O;
  wire [0:0] LIOB33_X0Y179_IOB_X0Y179_O;
  wire [0:0] LIOB33_X0Y179_IOB_X0Y180_O;
  wire [0:0] LIOB33_X0Y181_IOB_X0Y181_O;
  wire [0:0] LIOB33_X0Y181_IOB_X0Y182_O;
  wire [0:0] LIOB33_X0Y183_IOB_X0Y183_O;
  wire [0:0] LIOB33_X0Y183_IOB_X0Y184_O;
  wire [0:0] LIOB33_X0Y185_IOB_X0Y185_O;
  wire [0:0] LIOB33_X0Y185_IOB_X0Y186_O;
  wire [0:0] LIOB33_X0Y187_IOB_X0Y187_O;
  wire [0:0] LIOB33_X0Y187_IOB_X0Y188_O;
  wire [0:0] LIOB33_X0Y189_IOB_X0Y189_O;
  wire [0:0] LIOB33_X0Y189_IOB_X0Y190_O;
  wire [0:0] LIOB33_X0Y191_IOB_X0Y191_O;
  wire [0:0] LIOB33_X0Y191_IOB_X0Y192_O;
  wire [0:0] LIOB33_X0Y193_IOB_X0Y193_O;
  wire [0:0] LIOB33_X0Y193_IOB_X0Y194_O;
  wire [0:0] LIOB33_X0Y195_IOB_X0Y195_O;
  wire [0:0] LIOB33_X0Y195_IOB_X0Y196_O;
  wire [0:0] LIOB33_X0Y197_IOB_X0Y197_O;
  wire [0:0] LIOB33_X0Y197_IOB_X0Y198_O;
  wire [0:0] LIOB33_X0Y51_IOB_X0Y51_I;
  wire [0:0] LIOB33_X0Y51_IOB_X0Y52_I;
  wire [0:0] LIOB33_X0Y53_IOB_X0Y53_I;
  wire [0:0] LIOB33_X0Y53_IOB_X0Y54_I;
  wire [0:0] LIOB33_X0Y55_IOB_X0Y55_I;
  wire [0:0] LIOB33_X0Y55_IOB_X0Y56_I;
  wire [0:0] LIOB33_X0Y57_IOB_X0Y57_I;
  wire [0:0] LIOB33_X0Y57_IOB_X0Y58_I;
  wire [0:0] LIOB33_X0Y59_IOB_X0Y59_I;
  wire [0:0] LIOB33_X0Y59_IOB_X0Y60_I;
  wire [0:0] LIOB33_X0Y61_IOB_X0Y61_I;
  wire [0:0] LIOB33_X0Y61_IOB_X0Y62_I;
  wire [0:0] LIOB33_X0Y63_IOB_X0Y63_I;
  wire [0:0] LIOB33_X0Y63_IOB_X0Y64_O;
  wire [0:0] LIOB33_X0Y65_IOB_X0Y65_O;
  wire [0:0] LIOB33_X0Y65_IOB_X0Y66_O;
  wire [0:0] LIOB33_X0Y77_IOB_X0Y78_I;
  wire [0:0] LIOI3_SING_X0Y100_OLOGIC_X0Y100_D1;
  wire [0:0] LIOI3_SING_X0Y100_OLOGIC_X0Y100_OQ;
  wire [0:0] LIOI3_SING_X0Y100_OLOGIC_X0Y100_T1;
  wire [0:0] LIOI3_SING_X0Y100_OLOGIC_X0Y100_TQ;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_D1;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_OQ;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_T1;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_TQ;
  wire [0:0] LIOI3_SING_X0Y150_OLOGIC_X0Y150_D1;
  wire [0:0] LIOI3_SING_X0Y150_OLOGIC_X0Y150_OQ;
  wire [0:0] LIOI3_SING_X0Y150_OLOGIC_X0Y150_T1;
  wire [0:0] LIOI3_SING_X0Y150_OLOGIC_X0Y150_TQ;
  wire [0:0] LIOI3_SING_X0Y199_OLOGIC_X0Y199_D1;
  wire [0:0] LIOI3_SING_X0Y199_OLOGIC_X0Y199_OQ;
  wire [0:0] LIOI3_SING_X0Y199_OLOGIC_X0Y199_T1;
  wire [0:0] LIOI3_SING_X0Y199_OLOGIC_X0Y199_TQ;
  wire [0:0] LIOI3_SING_X0Y50_ILOGIC_X0Y50_D;
  wire [0:0] LIOI3_SING_X0Y50_ILOGIC_X0Y50_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y57_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y57_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y58_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y58_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y63_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y63_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_OLOGIC_X0Y64_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_OLOGIC_X0Y64_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_OLOGIC_X0Y64_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_OLOGIC_X0Y64_TQ;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y101_D1;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y101_OQ;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y101_T1;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y101_TQ;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y102_D1;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y102_OQ;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y102_T1;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y102_TQ;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y103_D1;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y103_OQ;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y103_T1;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y103_TQ;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y104_D1;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y104_OQ;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y104_T1;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y104_TQ;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y105_D1;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y105_OQ;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y105_T1;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y105_TQ;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y106_D1;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y106_OQ;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y106_T1;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y106_TQ;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y109_D1;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y109_OQ;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y109_T1;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y109_TQ;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y110_D1;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y110_OQ;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y110_T1;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y110_TQ;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_D1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_OQ;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_T1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_TQ;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y112_D1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y112_OQ;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y112_T1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y112_TQ;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y115_D1;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y115_OQ;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y115_T1;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y115_TQ;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y116_D1;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y116_OQ;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y116_T1;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y116_TQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y117_D1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y117_OQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y117_T1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y117_TQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_D1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_OQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_T1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_TQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_D1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_OQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_T1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_TQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_D1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_OQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_T1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_TQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_D1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_OQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_T1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_TQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_D1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_OQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_T1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_TQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_D1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_OQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_T1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_TQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_D1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_OQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_T1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_TQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_D1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_OQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_T1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_TQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_D1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_OQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_T1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_TQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_D1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_OQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_T1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_TQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_D1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_OQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_T1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_TQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_D1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_OQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_T1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_TQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_D1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_OQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_T1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_TQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_D1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_OQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_T1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_TQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_D1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_OQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_T1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_TQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_D1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_OQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_T1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_TQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_D1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_OQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_T1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_TQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_D1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_OQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_T1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_TQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_D1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_OQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_T1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_TQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_D1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_OQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_T1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_TQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_D1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_OQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_T1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_TQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_D1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_OQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_T1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_TQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_D1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_OQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_T1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_TQ;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y151_D1;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y151_OQ;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y151_T1;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y151_TQ;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y152_D1;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y152_OQ;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y152_T1;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y152_TQ;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y153_D1;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y153_OQ;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y153_T1;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y153_TQ;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y154_D1;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y154_OQ;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y154_T1;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y154_TQ;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y155_D1;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y155_OQ;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y155_T1;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y155_TQ;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y156_D1;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y156_OQ;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y156_T1;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y156_TQ;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y159_D1;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y159_OQ;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y159_T1;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y159_TQ;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y160_D1;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y160_OQ;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y160_T1;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y160_TQ;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y161_D1;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y161_OQ;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y161_T1;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y161_TQ;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y162_D1;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y162_OQ;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y162_T1;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y162_TQ;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y165_D1;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y165_OQ;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y165_T1;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y165_TQ;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y166_D1;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y166_OQ;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y166_T1;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y166_TQ;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y167_D1;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y167_OQ;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y167_T1;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y167_TQ;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y168_D1;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y168_OQ;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y168_T1;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y168_TQ;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y171_D1;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y171_OQ;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y171_T1;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y171_TQ;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y172_D1;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y172_OQ;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y172_T1;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y172_TQ;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y173_D1;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y173_OQ;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y173_T1;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y173_TQ;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y174_D1;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y174_OQ;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y174_T1;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y174_TQ;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y175_D1;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y175_OQ;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y175_T1;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y175_TQ;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y176_D1;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y176_OQ;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y176_T1;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y176_TQ;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y177_D1;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y177_OQ;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y177_T1;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y177_TQ;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y178_D1;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y178_OQ;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y178_T1;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y178_TQ;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y179_D1;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y179_OQ;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y179_T1;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y179_TQ;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y180_D1;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y180_OQ;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y180_T1;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y180_TQ;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y183_D1;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y183_OQ;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y183_T1;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y183_TQ;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y184_D1;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y184_OQ;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y184_T1;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y184_TQ;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y185_D1;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y185_OQ;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y185_T1;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y185_TQ;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y186_D1;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y186_OQ;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y186_T1;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y186_TQ;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y189_D1;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y189_OQ;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y189_T1;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y189_TQ;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y190_D1;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y190_OQ;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y190_T1;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y190_TQ;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y191_D1;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y191_OQ;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y191_T1;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y191_TQ;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y192_D1;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y192_OQ;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y192_T1;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y192_TQ;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y195_D1;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y195_OQ;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y195_T1;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y195_TQ;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y196_D1;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y196_OQ;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y196_T1;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y196_TQ;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y197_D1;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y197_OQ;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y197_T1;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y197_TQ;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y198_D1;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y198_OQ;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y198_T1;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y198_TQ;
  wire [0:0] LIOI3_X0Y51_ILOGIC_X0Y51_D;
  wire [0:0] LIOI3_X0Y51_ILOGIC_X0Y51_O;
  wire [0:0] LIOI3_X0Y51_ILOGIC_X0Y52_D;
  wire [0:0] LIOI3_X0Y51_ILOGIC_X0Y52_O;
  wire [0:0] LIOI3_X0Y53_ILOGIC_X0Y53_D;
  wire [0:0] LIOI3_X0Y53_ILOGIC_X0Y53_O;
  wire [0:0] LIOI3_X0Y53_ILOGIC_X0Y54_D;
  wire [0:0] LIOI3_X0Y53_ILOGIC_X0Y54_O;
  wire [0:0] LIOI3_X0Y55_ILOGIC_X0Y55_D;
  wire [0:0] LIOI3_X0Y55_ILOGIC_X0Y55_O;
  wire [0:0] LIOI3_X0Y55_ILOGIC_X0Y56_D;
  wire [0:0] LIOI3_X0Y55_ILOGIC_X0Y56_O;
  wire [0:0] LIOI3_X0Y59_ILOGIC_X0Y59_D;
  wire [0:0] LIOI3_X0Y59_ILOGIC_X0Y59_O;
  wire [0:0] LIOI3_X0Y59_ILOGIC_X0Y60_D;
  wire [0:0] LIOI3_X0Y59_ILOGIC_X0Y60_O;
  wire [0:0] LIOI3_X0Y61_ILOGIC_X0Y61_D;
  wire [0:0] LIOI3_X0Y61_ILOGIC_X0Y61_O;
  wire [0:0] LIOI3_X0Y61_ILOGIC_X0Y62_D;
  wire [0:0] LIOI3_X0Y61_ILOGIC_X0Y62_O;
  wire [0:0] LIOI3_X0Y65_OLOGIC_X0Y65_D1;
  wire [0:0] LIOI3_X0Y65_OLOGIC_X0Y65_OQ;
  wire [0:0] LIOI3_X0Y65_OLOGIC_X0Y65_T1;
  wire [0:0] LIOI3_X0Y65_OLOGIC_X0Y65_TQ;
  wire [0:0] LIOI3_X0Y65_OLOGIC_X0Y66_D1;
  wire [0:0] LIOI3_X0Y65_OLOGIC_X0Y66_OQ;
  wire [0:0] LIOI3_X0Y65_OLOGIC_X0Y66_T1;
  wire [0:0] LIOI3_X0Y65_OLOGIC_X0Y66_TQ;
  wire [0:0] LIOI3_X0Y77_ILOGIC_X0Y78_D;
  wire [0:0] LIOI3_X0Y77_ILOGIC_X0Y78_O;
  wire [0:0] RIOB33_SING_X105Y100_IOB_X1Y100_I;
  wire [0:0] RIOB33_SING_X105Y149_IOB_X1Y149_I;
  wire [0:0] RIOB33_SING_X105Y150_IOB_X1Y150_O;
  wire [0:0] RIOB33_SING_X105Y199_IOB_X1Y199_O;
  wire [0:0] RIOB33_X105Y101_IOB_X1Y101_I;
  wire [0:0] RIOB33_X105Y101_IOB_X1Y102_I;
  wire [0:0] RIOB33_X105Y103_IOB_X1Y103_I;
  wire [0:0] RIOB33_X105Y103_IOB_X1Y104_I;
  wire [0:0] RIOB33_X105Y105_IOB_X1Y105_I;
  wire [0:0] RIOB33_X105Y105_IOB_X1Y106_I;
  wire [0:0] RIOB33_X105Y107_IOB_X1Y107_I;
  wire [0:0] RIOB33_X105Y107_IOB_X1Y108_I;
  wire [0:0] RIOB33_X105Y109_IOB_X1Y109_I;
  wire [0:0] RIOB33_X105Y109_IOB_X1Y110_I;
  wire [0:0] RIOB33_X105Y111_IOB_X1Y111_I;
  wire [0:0] RIOB33_X105Y111_IOB_X1Y112_I;
  wire [0:0] RIOB33_X105Y113_IOB_X1Y113_I;
  wire [0:0] RIOB33_X105Y113_IOB_X1Y114_I;
  wire [0:0] RIOB33_X105Y115_IOB_X1Y115_I;
  wire [0:0] RIOB33_X105Y115_IOB_X1Y116_I;
  wire [0:0] RIOB33_X105Y117_IOB_X1Y117_I;
  wire [0:0] RIOB33_X105Y117_IOB_X1Y118_I;
  wire [0:0] RIOB33_X105Y119_IOB_X1Y119_I;
  wire [0:0] RIOB33_X105Y119_IOB_X1Y120_I;
  wire [0:0] RIOB33_X105Y121_IOB_X1Y121_I;
  wire [0:0] RIOB33_X105Y121_IOB_X1Y122_I;
  wire [0:0] RIOB33_X105Y123_IOB_X1Y123_I;
  wire [0:0] RIOB33_X105Y123_IOB_X1Y124_I;
  wire [0:0] RIOB33_X105Y125_IOB_X1Y125_I;
  wire [0:0] RIOB33_X105Y125_IOB_X1Y126_I;
  wire [0:0] RIOB33_X105Y127_IOB_X1Y127_I;
  wire [0:0] RIOB33_X105Y127_IOB_X1Y128_I;
  wire [0:0] RIOB33_X105Y129_IOB_X1Y129_I;
  wire [0:0] RIOB33_X105Y129_IOB_X1Y130_I;
  wire [0:0] RIOB33_X105Y131_IOB_X1Y131_I;
  wire [0:0] RIOB33_X105Y131_IOB_X1Y132_I;
  wire [0:0] RIOB33_X105Y133_IOB_X1Y133_I;
  wire [0:0] RIOB33_X105Y133_IOB_X1Y134_I;
  wire [0:0] RIOB33_X105Y135_IOB_X1Y135_I;
  wire [0:0] RIOB33_X105Y135_IOB_X1Y136_I;
  wire [0:0] RIOB33_X105Y137_IOB_X1Y137_I;
  wire [0:0] RIOB33_X105Y137_IOB_X1Y138_I;
  wire [0:0] RIOB33_X105Y139_IOB_X1Y139_I;
  wire [0:0] RIOB33_X105Y139_IOB_X1Y140_I;
  wire [0:0] RIOB33_X105Y141_IOB_X1Y141_I;
  wire [0:0] RIOB33_X105Y141_IOB_X1Y142_I;
  wire [0:0] RIOB33_X105Y143_IOB_X1Y143_I;
  wire [0:0] RIOB33_X105Y143_IOB_X1Y144_I;
  wire [0:0] RIOB33_X105Y145_IOB_X1Y145_I;
  wire [0:0] RIOB33_X105Y145_IOB_X1Y146_I;
  wire [0:0] RIOB33_X105Y147_IOB_X1Y147_I;
  wire [0:0] RIOB33_X105Y147_IOB_X1Y148_I;
  wire [0:0] RIOB33_X105Y151_IOB_X1Y151_O;
  wire [0:0] RIOB33_X105Y151_IOB_X1Y152_O;
  wire [0:0] RIOB33_X105Y153_IOB_X1Y153_O;
  wire [0:0] RIOB33_X105Y153_IOB_X1Y154_O;
  wire [0:0] RIOB33_X105Y155_IOB_X1Y155_O;
  wire [0:0] RIOB33_X105Y155_IOB_X1Y156_O;
  wire [0:0] RIOB33_X105Y157_IOB_X1Y157_O;
  wire [0:0] RIOB33_X105Y157_IOB_X1Y158_O;
  wire [0:0] RIOB33_X105Y159_IOB_X1Y159_O;
  wire [0:0] RIOB33_X105Y159_IOB_X1Y160_O;
  wire [0:0] RIOB33_X105Y161_IOB_X1Y161_O;
  wire [0:0] RIOB33_X105Y161_IOB_X1Y162_O;
  wire [0:0] RIOB33_X105Y163_IOB_X1Y163_O;
  wire [0:0] RIOB33_X105Y163_IOB_X1Y164_O;
  wire [0:0] RIOB33_X105Y165_IOB_X1Y165_O;
  wire [0:0] RIOB33_X105Y165_IOB_X1Y166_O;
  wire [0:0] RIOB33_X105Y167_IOB_X1Y167_O;
  wire [0:0] RIOB33_X105Y167_IOB_X1Y168_O;
  wire [0:0] RIOB33_X105Y169_IOB_X1Y169_O;
  wire [0:0] RIOB33_X105Y169_IOB_X1Y170_O;
  wire [0:0] RIOB33_X105Y171_IOB_X1Y171_O;
  wire [0:0] RIOB33_X105Y171_IOB_X1Y172_O;
  wire [0:0] RIOB33_X105Y173_IOB_X1Y173_O;
  wire [0:0] RIOB33_X105Y173_IOB_X1Y174_O;
  wire [0:0] RIOB33_X105Y175_IOB_X1Y175_O;
  wire [0:0] RIOB33_X105Y175_IOB_X1Y176_O;
  wire [0:0] RIOB33_X105Y177_IOB_X1Y177_O;
  wire [0:0] RIOB33_X105Y177_IOB_X1Y178_O;
  wire [0:0] RIOB33_X105Y179_IOB_X1Y179_O;
  wire [0:0] RIOB33_X105Y179_IOB_X1Y180_O;
  wire [0:0] RIOB33_X105Y181_IOB_X1Y181_O;
  wire [0:0] RIOB33_X105Y181_IOB_X1Y182_O;
  wire [0:0] RIOB33_X105Y183_IOB_X1Y183_O;
  wire [0:0] RIOB33_X105Y183_IOB_X1Y184_O;
  wire [0:0] RIOB33_X105Y185_IOB_X1Y185_O;
  wire [0:0] RIOB33_X105Y185_IOB_X1Y186_O;
  wire [0:0] RIOB33_X105Y187_IOB_X1Y187_O;
  wire [0:0] RIOB33_X105Y187_IOB_X1Y188_O;
  wire [0:0] RIOB33_X105Y189_IOB_X1Y189_O;
  wire [0:0] RIOB33_X105Y189_IOB_X1Y190_O;
  wire [0:0] RIOB33_X105Y191_IOB_X1Y191_O;
  wire [0:0] RIOB33_X105Y191_IOB_X1Y192_O;
  wire [0:0] RIOB33_X105Y193_IOB_X1Y193_O;
  wire [0:0] RIOB33_X105Y193_IOB_X1Y194_O;
  wire [0:0] RIOB33_X105Y195_IOB_X1Y195_O;
  wire [0:0] RIOB33_X105Y195_IOB_X1Y196_O;
  wire [0:0] RIOB33_X105Y197_IOB_X1Y197_O;
  wire [0:0] RIOB33_X105Y197_IOB_X1Y198_O;
  wire [0:0] RIOI3_SING_X105Y100_ILOGIC_X1Y100_D;
  wire [0:0] RIOI3_SING_X105Y100_ILOGIC_X1Y100_O;
  wire [0:0] RIOI3_SING_X105Y149_ILOGIC_X1Y149_D;
  wire [0:0] RIOI3_SING_X105Y149_ILOGIC_X1Y149_O;
  wire [0:0] RIOI3_SING_X105Y150_OLOGIC_X1Y150_D1;
  wire [0:0] RIOI3_SING_X105Y150_OLOGIC_X1Y150_OQ;
  wire [0:0] RIOI3_SING_X105Y150_OLOGIC_X1Y150_T1;
  wire [0:0] RIOI3_SING_X105Y150_OLOGIC_X1Y150_TQ;
  wire [0:0] RIOI3_SING_X105Y199_OLOGIC_X1Y199_D1;
  wire [0:0] RIOI3_SING_X105Y199_OLOGIC_X1Y199_OQ;
  wire [0:0] RIOI3_SING_X105Y199_OLOGIC_X1Y199_T1;
  wire [0:0] RIOI3_SING_X105Y199_OLOGIC_X1Y199_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y120_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y120_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y131_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y131_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y132_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y132_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y143_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y143_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y144_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y144_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y137_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y137_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y138_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y138_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_TQ;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y101_D;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y101_O;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y102_D;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y102_O;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y103_D;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y103_O;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y104_D;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y104_O;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y105_D;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y105_O;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y106_D;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y106_O;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y109_D;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y109_O;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y110_D;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y110_O;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y111_D;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y111_O;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y112_D;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y112_O;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y115_D;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y115_O;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y116_D;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y116_O;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y117_D;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y117_O;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y118_D;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y118_O;
  wire [0:0] RIOI3_X105Y121_ILOGIC_X1Y121_D;
  wire [0:0] RIOI3_X105Y121_ILOGIC_X1Y121_O;
  wire [0:0] RIOI3_X105Y121_ILOGIC_X1Y122_D;
  wire [0:0] RIOI3_X105Y121_ILOGIC_X1Y122_O;
  wire [0:0] RIOI3_X105Y123_ILOGIC_X1Y123_D;
  wire [0:0] RIOI3_X105Y123_ILOGIC_X1Y123_O;
  wire [0:0] RIOI3_X105Y123_ILOGIC_X1Y124_D;
  wire [0:0] RIOI3_X105Y123_ILOGIC_X1Y124_O;
  wire [0:0] RIOI3_X105Y125_ILOGIC_X1Y125_D;
  wire [0:0] RIOI3_X105Y125_ILOGIC_X1Y125_O;
  wire [0:0] RIOI3_X105Y125_ILOGIC_X1Y126_D;
  wire [0:0] RIOI3_X105Y125_ILOGIC_X1Y126_O;
  wire [0:0] RIOI3_X105Y127_ILOGIC_X1Y127_D;
  wire [0:0] RIOI3_X105Y127_ILOGIC_X1Y127_O;
  wire [0:0] RIOI3_X105Y127_ILOGIC_X1Y128_D;
  wire [0:0] RIOI3_X105Y127_ILOGIC_X1Y128_O;
  wire [0:0] RIOI3_X105Y129_ILOGIC_X1Y129_D;
  wire [0:0] RIOI3_X105Y129_ILOGIC_X1Y129_O;
  wire [0:0] RIOI3_X105Y129_ILOGIC_X1Y130_D;
  wire [0:0] RIOI3_X105Y129_ILOGIC_X1Y130_O;
  wire [0:0] RIOI3_X105Y133_ILOGIC_X1Y133_D;
  wire [0:0] RIOI3_X105Y133_ILOGIC_X1Y133_O;
  wire [0:0] RIOI3_X105Y133_ILOGIC_X1Y134_D;
  wire [0:0] RIOI3_X105Y133_ILOGIC_X1Y134_O;
  wire [0:0] RIOI3_X105Y135_ILOGIC_X1Y135_D;
  wire [0:0] RIOI3_X105Y135_ILOGIC_X1Y135_O;
  wire [0:0] RIOI3_X105Y135_ILOGIC_X1Y136_D;
  wire [0:0] RIOI3_X105Y135_ILOGIC_X1Y136_O;
  wire [0:0] RIOI3_X105Y139_ILOGIC_X1Y139_D;
  wire [0:0] RIOI3_X105Y139_ILOGIC_X1Y139_O;
  wire [0:0] RIOI3_X105Y139_ILOGIC_X1Y140_D;
  wire [0:0] RIOI3_X105Y139_ILOGIC_X1Y140_O;
  wire [0:0] RIOI3_X105Y141_ILOGIC_X1Y141_D;
  wire [0:0] RIOI3_X105Y141_ILOGIC_X1Y141_O;
  wire [0:0] RIOI3_X105Y141_ILOGIC_X1Y142_D;
  wire [0:0] RIOI3_X105Y141_ILOGIC_X1Y142_O;
  wire [0:0] RIOI3_X105Y145_ILOGIC_X1Y145_D;
  wire [0:0] RIOI3_X105Y145_ILOGIC_X1Y145_O;
  wire [0:0] RIOI3_X105Y145_ILOGIC_X1Y146_D;
  wire [0:0] RIOI3_X105Y145_ILOGIC_X1Y146_O;
  wire [0:0] RIOI3_X105Y147_ILOGIC_X1Y147_D;
  wire [0:0] RIOI3_X105Y147_ILOGIC_X1Y147_O;
  wire [0:0] RIOI3_X105Y147_ILOGIC_X1Y148_D;
  wire [0:0] RIOI3_X105Y147_ILOGIC_X1Y148_O;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y151_D1;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y151_OQ;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y151_T1;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y151_TQ;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y152_D1;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y152_OQ;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y152_T1;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y152_TQ;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y153_D1;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y153_OQ;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y153_T1;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y153_TQ;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y154_D1;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y154_OQ;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y154_T1;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y154_TQ;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y155_D1;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y155_OQ;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y155_T1;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y155_TQ;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y156_D1;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y156_OQ;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y156_T1;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y156_TQ;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y159_D1;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y159_OQ;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y159_T1;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y159_TQ;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y160_D1;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y160_OQ;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y160_T1;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y160_TQ;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y161_D1;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y161_OQ;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y161_T1;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y161_TQ;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y162_D1;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y162_OQ;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y162_T1;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y162_TQ;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y165_D1;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y165_OQ;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y165_T1;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y165_TQ;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y166_D1;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y166_OQ;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y166_T1;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y166_TQ;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y167_D1;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y167_OQ;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y167_T1;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y167_TQ;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y168_D1;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y168_OQ;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y168_T1;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y168_TQ;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y171_D1;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y171_OQ;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y171_T1;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y171_TQ;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y172_D1;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y172_OQ;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y172_T1;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y172_TQ;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y173_D1;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y173_OQ;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y173_T1;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y173_TQ;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y174_D1;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y174_OQ;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y174_T1;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y174_TQ;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y175_D1;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y175_OQ;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y175_T1;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y175_TQ;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y176_D1;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y176_OQ;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y176_T1;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y176_TQ;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y177_D1;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y177_OQ;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y177_T1;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y177_TQ;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y178_D1;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y178_OQ;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y178_T1;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y178_TQ;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y179_D1;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y179_OQ;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y179_T1;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y179_TQ;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y180_D1;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y180_OQ;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y180_T1;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y180_TQ;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y183_D1;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y183_OQ;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y183_T1;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y183_TQ;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y184_D1;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y184_OQ;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y184_T1;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y184_TQ;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y185_D1;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y185_OQ;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y185_T1;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y185_TQ;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y186_D1;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y186_OQ;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y186_T1;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y186_TQ;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y189_D1;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y189_OQ;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y189_T1;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y189_TQ;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y190_D1;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y190_OQ;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y190_T1;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y190_TQ;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y191_D1;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y191_OQ;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y191_T1;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y191_TQ;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y192_D1;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y192_OQ;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y192_T1;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y192_TQ;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y195_D1;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y195_OQ;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y195_T1;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y195_TQ;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y196_D1;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y196_OQ;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y196_T1;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y196_TQ;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y197_D1;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y197_OQ;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y197_T1;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y197_TQ;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y198_D1;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y198_OQ;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y198_T1;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y198_TQ;


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y75_SLICE_X0Y75_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y75_SLICE_X0Y75_DO5),
.O6(CLBLL_L_X2Y75_SLICE_X0Y75_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y75_SLICE_X0Y75_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y75_SLICE_X0Y75_CO5),
.O6(CLBLL_L_X2Y75_SLICE_X0Y75_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y75_SLICE_X0Y75_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y75_SLICE_X0Y75_BO5),
.O6(CLBLL_L_X2Y75_SLICE_X0Y75_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0f0f0f0f0f)
  ) CLBLL_L_X2Y75_SLICE_X0Y75_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(LIOB33_X0Y55_IOB_X0Y56_I),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y75_SLICE_X0Y75_AO5),
.O6(CLBLL_L_X2Y75_SLICE_X0Y75_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y75_SLICE_X1Y75_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y75_SLICE_X1Y75_DO5),
.O6(CLBLL_L_X2Y75_SLICE_X1Y75_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y75_SLICE_X1Y75_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y75_SLICE_X1Y75_CO5),
.O6(CLBLL_L_X2Y75_SLICE_X1Y75_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y75_SLICE_X1Y75_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y75_SLICE_X1Y75_BO5),
.O6(CLBLL_L_X2Y75_SLICE_X1Y75_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y75_SLICE_X1Y75_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y75_SLICE_X1Y75_AO5),
.O6(CLBLL_L_X2Y75_SLICE_X1Y75_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y143_SLICE_X0Y143_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y143_SLICE_X0Y143_DO5),
.O6(CLBLL_L_X2Y143_SLICE_X0Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y143_SLICE_X0Y143_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y143_SLICE_X0Y143_CO5),
.O6(CLBLL_L_X2Y143_SLICE_X0Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y143_SLICE_X0Y143_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y143_SLICE_X0Y143_BO5),
.O6(CLBLL_L_X2Y143_SLICE_X0Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y143_SLICE_X0Y143_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y143_SLICE_X0Y143_AO5),
.O6(CLBLL_L_X2Y143_SLICE_X0Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y143_SLICE_X1Y143_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y143_SLICE_X1Y143_AO6),
.Q(CLBLL_L_X2Y143_SLICE_X1Y143_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y143_SLICE_X1Y143_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y143_SLICE_X1Y143_BO6),
.Q(CLBLL_L_X2Y143_SLICE_X1Y143_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y143_SLICE_X1Y143_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y143_SLICE_X1Y143_CO6),
.Q(CLBLL_L_X2Y143_SLICE_X1Y143_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y143_SLICE_X1Y143_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y143_SLICE_X1Y143_DO6),
.Q(CLBLL_L_X2Y143_SLICE_X1Y143_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbbbb8b88888b8b8)
  ) CLBLL_L_X2Y143_SLICE_X1Y143_DLUT (
.I0(CLBLL_L_X2Y144_SLICE_X1Y144_AQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLL_L_X2Y143_SLICE_X1Y143_DQ),
.I3(1'b1),
.I4(CLBLM_L_X10Y143_SLICE_X12Y143_BO5),
.I5(CLBLM_R_X3Y144_SLICE_X3Y144_BQ),
.O5(CLBLL_L_X2Y143_SLICE_X1Y143_DO5),
.O6(CLBLL_L_X2Y143_SLICE_X1Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf066f066f066f066)
  ) CLBLL_L_X2Y143_SLICE_X1Y143_CLUT (
.I0(LIOB33_X0Y57_IOB_X0Y58_I),
.I1(CLBLL_L_X2Y143_SLICE_X1Y143_CQ),
.I2(CLBLL_L_X2Y143_SLICE_X1Y143_DQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y143_SLICE_X1Y143_CO5),
.O6(CLBLL_L_X2Y143_SLICE_X1Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff005555aaaa)
  ) CLBLL_L_X2Y143_SLICE_X1Y143_BLUT (
.I0(CLBLM_R_X7Y152_SLICE_X8Y152_BQ),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLL_L_X4Y143_SLICE_X4Y143_DQ),
.I4(CLBLL_L_X4Y144_SLICE_X5Y144_D5Q),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLL_L_X2Y143_SLICE_X1Y143_BO5),
.O6(CLBLL_L_X2Y143_SLICE_X1Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff33fd31cc00ec20)
  ) CLBLL_L_X2Y143_SLICE_X1Y143_ALUT (
.I0(CLBLM_R_X3Y148_SLICE_X2Y148_D5Q),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLL_L_X2Y143_SLICE_X1Y143_AQ),
.I3(CLBLM_R_X3Y150_SLICE_X3Y150_BQ),
.I4(CLBLM_R_X5Y144_SLICE_X6Y144_DQ),
.I5(CLBLL_L_X4Y148_SLICE_X4Y148_A5Q),
.O5(CLBLL_L_X2Y143_SLICE_X1Y143_AO5),
.O6(CLBLL_L_X2Y143_SLICE_X1Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y144_SLICE_X0Y144_A_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y144_SLICE_X2Y144_BO6),
.Q(CLBLL_L_X2Y144_SLICE_X0Y144_AQ),
.S(CLBLM_R_X7Y144_SLICE_X8Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y144_SLICE_X0Y144_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y144_SLICE_X0Y144_DO5),
.O6(CLBLL_L_X2Y144_SLICE_X0Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y144_SLICE_X0Y144_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y144_SLICE_X0Y144_CO5),
.O6(CLBLL_L_X2Y144_SLICE_X0Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y144_SLICE_X0Y144_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y144_SLICE_X0Y144_BO5),
.O6(CLBLL_L_X2Y144_SLICE_X0Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y144_SLICE_X0Y144_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y144_SLICE_X0Y144_AO5),
.O6(CLBLL_L_X2Y144_SLICE_X0Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y144_SLICE_X1Y144_A5_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y144_SLICE_X1Y144_AO5),
.Q(CLBLL_L_X2Y144_SLICE_X1Y144_A5Q),
.S(CLBLL_L_X2Y144_SLICE_X1Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y144_SLICE_X1Y144_B5_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y144_SLICE_X1Y144_BO5),
.Q(CLBLL_L_X2Y144_SLICE_X1Y144_B5Q),
.S(CLBLL_L_X2Y144_SLICE_X1Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y144_SLICE_X1Y144_A_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y144_SLICE_X1Y144_AO6),
.Q(CLBLL_L_X2Y144_SLICE_X1Y144_AQ),
.S(CLBLL_L_X2Y144_SLICE_X1Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y144_SLICE_X1Y144_B_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y144_SLICE_X1Y144_BO6),
.Q(CLBLL_L_X2Y144_SLICE_X1Y144_BQ),
.S(CLBLL_L_X2Y144_SLICE_X1Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y144_SLICE_X1Y144_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y144_SLICE_X1Y144_DO5),
.O6(CLBLL_L_X2Y144_SLICE_X1Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000f0f0f0f0)
  ) CLBLL_L_X2Y144_SLICE_X1Y144_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X5Y144_SLICE_X7Y144_CQ),
.I3(1'b1),
.I4(1'b1),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLL_L_X2Y144_SLICE_X1Y144_CO5),
.O6(CLBLL_L_X2Y144_SLICE_X1Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000cccc0000)
  ) CLBLL_L_X2Y144_SLICE_X1Y144_BLUT (
.I0(LIOB33_X0Y63_IOB_X0Y63_I),
.I1(CLBLM_R_X3Y144_SLICE_X2Y144_AQ),
.I2(1'b1),
.I3(1'b1),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y144_SLICE_X1Y144_BO5),
.O6(CLBLL_L_X2Y144_SLICE_X1Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00ff000000)
  ) CLBLL_L_X2Y144_SLICE_X1Y144_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y142_SLICE_X7Y142_B5Q),
.I2(1'b1),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X3Y145_SLICE_X2Y145_DQ),
.I5(1'b1),
.O5(CLBLL_L_X2Y144_SLICE_X1Y144_AO5),
.O6(CLBLL_L_X2Y144_SLICE_X1Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y145_SLICE_X0Y145_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y145_SLICE_X0Y145_DO5),
.O6(CLBLL_L_X2Y145_SLICE_X0Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y145_SLICE_X0Y145_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y145_SLICE_X0Y145_CO5),
.O6(CLBLL_L_X2Y145_SLICE_X0Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y145_SLICE_X0Y145_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y145_SLICE_X0Y145_BO5),
.O6(CLBLL_L_X2Y145_SLICE_X0Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y145_SLICE_X0Y145_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y145_SLICE_X0Y145_AO5),
.O6(CLBLL_L_X2Y145_SLICE_X0Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y145_SLICE_X1Y145_A5_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y145_SLICE_X1Y145_AO5),
.Q(CLBLL_L_X2Y145_SLICE_X1Y145_A5Q),
.S(CLBLL_L_X2Y146_SLICE_X1Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y145_SLICE_X1Y145_A_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y145_SLICE_X1Y145_AO6),
.Q(CLBLL_L_X2Y145_SLICE_X1Y145_AQ),
.S(CLBLL_L_X2Y146_SLICE_X1Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y145_SLICE_X1Y145_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y145_SLICE_X1Y145_DO5),
.O6(CLBLL_L_X2Y145_SLICE_X1Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y145_SLICE_X1Y145_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y145_SLICE_X1Y145_CO5),
.O6(CLBLL_L_X2Y145_SLICE_X1Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y145_SLICE_X1Y145_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y145_SLICE_X1Y145_BO5),
.O6(CLBLL_L_X2Y145_SLICE_X1Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0000aaaa0000)
  ) CLBLL_L_X2Y145_SLICE_X1Y145_ALUT (
.I0(CLBLL_L_X2Y147_SLICE_X1Y147_A5Q),
.I1(CLBLM_R_X5Y147_SLICE_X6Y147_BQ),
.I2(1'b1),
.I3(1'b1),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y145_SLICE_X1Y145_AO5),
.O6(CLBLL_L_X2Y145_SLICE_X1Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y146_SLICE_X0Y146_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y146_SLICE_X0Y146_DO5),
.O6(CLBLL_L_X2Y146_SLICE_X0Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y146_SLICE_X0Y146_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y146_SLICE_X0Y146_CO5),
.O6(CLBLL_L_X2Y146_SLICE_X0Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y146_SLICE_X0Y146_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y146_SLICE_X0Y146_BO5),
.O6(CLBLL_L_X2Y146_SLICE_X0Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y146_SLICE_X0Y146_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y146_SLICE_X0Y146_AO5),
.O6(CLBLL_L_X2Y146_SLICE_X0Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y146_SLICE_X1Y146_A5_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y146_SLICE_X1Y146_AO5),
.Q(CLBLL_L_X2Y146_SLICE_X1Y146_A5Q),
.S(CLBLM_R_X7Y144_SLICE_X8Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y146_SLICE_X1Y146_A_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y146_SLICE_X1Y146_AO6),
.Q(CLBLL_L_X2Y146_SLICE_X1Y146_AQ),
.S(CLBLM_R_X7Y144_SLICE_X8Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y146_SLICE_X1Y146_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y146_SLICE_X1Y146_DO5),
.O6(CLBLL_L_X2Y146_SLICE_X1Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f000f000f000f00)
  ) CLBLL_L_X2Y146_SLICE_X1Y146_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X5Y149_SLICE_X7Y149_BQ),
.I3(CLBLM_R_X3Y147_SLICE_X2Y147_CQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y146_SLICE_X1Y146_CO5),
.O6(CLBLL_L_X2Y146_SLICE_X1Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555000055550000)
  ) CLBLL_L_X2Y146_SLICE_X1Y146_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X3Y151_SLICE_X3Y151_AQ),
.I5(1'b1),
.O5(CLBLL_L_X2Y146_SLICE_X1Y146_BO5),
.O6(CLBLL_L_X2Y146_SLICE_X1Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00a0a0a0a0)
  ) CLBLL_L_X2Y146_SLICE_X1Y146_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(1'b1),
.I2(CLBLM_R_X3Y154_SLICE_X3Y154_AQ),
.I3(CLBLL_L_X2Y149_SLICE_X1Y149_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y146_SLICE_X1Y146_AO5),
.O6(CLBLL_L_X2Y146_SLICE_X1Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y147_SLICE_X0Y147_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y147_SLICE_X0Y147_BO5),
.Q(CLBLL_L_X2Y147_SLICE_X0Y147_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y147_SLICE_X0Y147_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y147_SLICE_X0Y147_AO6),
.Q(CLBLL_L_X2Y147_SLICE_X0Y147_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y147_SLICE_X0Y147_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y147_SLICE_X0Y147_BO6),
.Q(CLBLL_L_X2Y147_SLICE_X0Y147_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y147_SLICE_X0Y147_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y147_SLICE_X0Y147_DO5),
.O6(CLBLL_L_X2Y147_SLICE_X0Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y147_SLICE_X0Y147_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y147_SLICE_X0Y147_CO5),
.O6(CLBLL_L_X2Y147_SLICE_X0Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5a0a08dd88dd8)
  ) CLBLL_L_X2Y147_SLICE_X0Y147_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLL_L_X4Y144_SLICE_X5Y144_D5Q),
.I2(CLBLM_L_X10Y147_SLICE_X12Y147_C5Q),
.I3(CLBLL_L_X4Y153_SLICE_X5Y153_BQ),
.I4(CLBLM_R_X3Y144_SLICE_X3Y144_A5Q),
.I5(1'b1),
.O5(CLBLL_L_X2Y147_SLICE_X0Y147_BO5),
.O6(CLBLL_L_X2Y147_SLICE_X0Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbe14be14be14be14)
  ) CLBLL_L_X2Y147_SLICE_X0Y147_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X10Y146_SLICE_X12Y146_AQ),
.I2(CLBLM_R_X7Y144_SLICE_X9Y144_AQ),
.I3(CLBLM_R_X7Y152_SLICE_X9Y152_DQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y147_SLICE_X0Y147_AO5),
.O6(CLBLL_L_X2Y147_SLICE_X0Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y147_SLICE_X1Y147_A5_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y147_SLICE_X1Y147_AO5),
.Q(CLBLL_L_X2Y147_SLICE_X1Y147_A5Q),
.S(CLBLL_L_X2Y147_SLICE_X1Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y147_SLICE_X1Y147_A_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y147_SLICE_X1Y147_AO6),
.Q(CLBLL_L_X2Y147_SLICE_X1Y147_AQ),
.S(CLBLL_L_X2Y147_SLICE_X1Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y147_SLICE_X1Y147_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y147_SLICE_X1Y147_DO5),
.O6(CLBLL_L_X2Y147_SLICE_X1Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y147_SLICE_X1Y147_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y147_SLICE_X1Y147_CO5),
.O6(CLBLL_L_X2Y147_SLICE_X1Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555555500000000)
  ) CLBLL_L_X2Y147_SLICE_X1Y147_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X3Y144_SLICE_X3Y144_CQ),
.O5(CLBLL_L_X2Y147_SLICE_X1Y147_BO5),
.O6(CLBLL_L_X2Y147_SLICE_X1Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888a0a0a0a0)
  ) CLBLL_L_X2Y147_SLICE_X1Y147_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X5Y147_SLICE_X6Y147_DQ),
.I2(CLBLM_R_X3Y146_SLICE_X3Y146_C5Q),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y147_SLICE_X1Y147_AO5),
.O6(CLBLL_L_X2Y147_SLICE_X1Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y148_SLICE_X0Y148_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y148_SLICE_X0Y148_AO5),
.Q(CLBLL_L_X2Y148_SLICE_X0Y148_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y148_SLICE_X0Y148_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y148_SLICE_X0Y148_BO5),
.Q(CLBLL_L_X2Y148_SLICE_X0Y148_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y148_SLICE_X0Y148_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y148_SLICE_X0Y148_AO6),
.Q(CLBLL_L_X2Y148_SLICE_X0Y148_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y148_SLICE_X0Y148_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y148_SLICE_X0Y148_BO6),
.Q(CLBLL_L_X2Y148_SLICE_X0Y148_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y148_SLICE_X0Y148_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y148_SLICE_X0Y148_DO5),
.O6(CLBLL_L_X2Y148_SLICE_X0Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y148_SLICE_X0Y148_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y148_SLICE_X0Y148_CO5),
.O6(CLBLL_L_X2Y148_SLICE_X0Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0aaf0aaccaaccaa)
  ) CLBLL_L_X2Y148_SLICE_X0Y148_BLUT (
.I0(CLBLM_R_X3Y150_SLICE_X2Y150_B5Q),
.I1(CLBLM_L_X10Y150_SLICE_X12Y150_AQ),
.I2(CLBLL_L_X2Y147_SLICE_X0Y147_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y148_SLICE_X0Y148_BO5),
.O6(CLBLL_L_X2Y148_SLICE_X0Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa0afa0aacacacac)
  ) CLBLL_L_X2Y148_SLICE_X0Y148_ALUT (
.I0(CLBLM_L_X8Y153_SLICE_X10Y153_AQ),
.I1(CLBLM_R_X3Y148_SLICE_X3Y148_DO6),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X3Y149_SLICE_X3Y149_DQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y148_SLICE_X0Y148_AO5),
.O6(CLBLL_L_X2Y148_SLICE_X0Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y148_SLICE_X1Y148_A5_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y148_SLICE_X1Y148_AO5),
.Q(CLBLL_L_X2Y148_SLICE_X1Y148_A5Q),
.S(CLBLL_L_X2Y146_SLICE_X1Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y148_SLICE_X1Y148_A_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y148_SLICE_X1Y148_AO6),
.Q(CLBLL_L_X2Y148_SLICE_X1Y148_AQ),
.S(CLBLL_L_X2Y146_SLICE_X1Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y148_SLICE_X1Y148_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y148_SLICE_X1Y148_DO5),
.O6(CLBLL_L_X2Y148_SLICE_X1Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y148_SLICE_X1Y148_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y148_SLICE_X1Y148_CO5),
.O6(CLBLL_L_X2Y148_SLICE_X1Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000f0f0cccc0000)
  ) CLBLL_L_X2Y148_SLICE_X1Y148_BLUT (
.I0(1'b1),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X3Y146_SLICE_X2Y146_C5Q),
.I3(1'b1),
.I4(CLBLM_R_X3Y148_SLICE_X2Y148_BQ),
.I5(1'b1),
.O5(CLBLL_L_X2Y148_SLICE_X1Y148_BO5),
.O6(CLBLL_L_X2Y148_SLICE_X1Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c088888888)
  ) CLBLL_L_X2Y148_SLICE_X1Y148_ALUT (
.I0(CLBLL_L_X4Y149_SLICE_X4Y149_C5Q),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLL_L_X4Y148_SLICE_X5Y148_BQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y148_SLICE_X1Y148_AO5),
.O6(CLBLL_L_X2Y148_SLICE_X1Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y149_SLICE_X0Y149_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y149_SLICE_X0Y149_AO6),
.Q(CLBLL_L_X2Y149_SLICE_X0Y149_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y149_SLICE_X0Y149_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y149_SLICE_X0Y149_DO5),
.O6(CLBLL_L_X2Y149_SLICE_X0Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y149_SLICE_X0Y149_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y149_SLICE_X0Y149_CO5),
.O6(CLBLL_L_X2Y149_SLICE_X0Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y149_SLICE_X0Y149_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y149_SLICE_X0Y149_BO5),
.O6(CLBLL_L_X2Y149_SLICE_X0Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00afafaaaa)
  ) CLBLL_L_X2Y149_SLICE_X0Y149_ALUT (
.I0(CLBLM_R_X3Y150_SLICE_X2Y150_B5Q),
.I1(1'b1),
.I2(CLBLM_L_X10Y150_SLICE_X12Y150_CQ),
.I3(CLBLM_R_X3Y151_SLICE_X2Y151_A5Q),
.I4(CLBLM_R_X7Y148_SLICE_X9Y148_AQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLL_L_X2Y149_SLICE_X0Y149_AO5),
.O6(CLBLL_L_X2Y149_SLICE_X0Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y149_SLICE_X1Y149_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y149_SLICE_X1Y149_AO5),
.Q(CLBLL_L_X2Y149_SLICE_X1Y149_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y149_SLICE_X1Y149_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y149_SLICE_X1Y149_AO6),
.Q(CLBLL_L_X2Y149_SLICE_X1Y149_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y149_SLICE_X1Y149_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y149_SLICE_X1Y149_BO6),
.Q(CLBLL_L_X2Y149_SLICE_X1Y149_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y149_SLICE_X1Y149_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y149_SLICE_X1Y149_CO6),
.Q(CLBLL_L_X2Y149_SLICE_X1Y149_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y149_SLICE_X1Y149_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y149_SLICE_X1Y149_DO6),
.Q(CLBLL_L_X2Y149_SLICE_X1Y149_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00de12cc00dc10)
  ) CLBLL_L_X2Y149_SLICE_X1Y149_DLUT (
.I0(CLBLL_L_X2Y149_SLICE_X1Y149_BQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLL_L_X2Y149_SLICE_X1Y149_DQ),
.I3(CLBLL_L_X2Y147_SLICE_X0Y147_B5Q),
.I4(CLBLL_L_X4Y152_SLICE_X5Y152_CQ),
.I5(CLBLL_L_X2Y149_SLICE_X1Y149_CQ),
.O5(CLBLL_L_X2Y149_SLICE_X1Y149_DO5),
.O6(CLBLL_L_X2Y149_SLICE_X1Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffec00ecffff00ff)
  ) CLBLL_L_X2Y149_SLICE_X1Y149_CLUT (
.I0(CLBLL_L_X2Y149_SLICE_X1Y149_BQ),
.I1(CLBLL_L_X4Y152_SLICE_X5Y152_CQ),
.I2(CLBLL_L_X2Y149_SLICE_X1Y149_DQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X5Y142_SLICE_X7Y142_C5Q),
.I5(CLBLL_L_X2Y149_SLICE_X1Y149_CQ),
.O5(CLBLL_L_X2Y149_SLICE_X1Y149_CO5),
.O6(CLBLL_L_X2Y149_SLICE_X1Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000010141014)
  ) CLBLL_L_X2Y149_SLICE_X1Y149_BLUT (
.I0(CLBLL_L_X4Y152_SLICE_X5Y152_CQ),
.I1(CLBLL_L_X2Y149_SLICE_X1Y149_BQ),
.I2(CLBLL_L_X2Y149_SLICE_X1Y149_CQ),
.I3(CLBLL_L_X2Y149_SLICE_X1Y149_DQ),
.I4(CLBLM_R_X3Y150_SLICE_X2Y150_DQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLL_L_X2Y149_SLICE_X1Y149_BO5),
.O6(CLBLL_L_X2Y149_SLICE_X1Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00ccf0aaffaa00)
  ) CLBLL_L_X2Y149_SLICE_X1Y149_ALUT (
.I0(CLBLM_R_X5Y149_SLICE_X7Y149_BQ),
.I1(CLBLL_L_X2Y144_SLICE_X1Y144_BQ),
.I2(CLBLM_R_X7Y148_SLICE_X9Y148_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X10Y150_SLICE_X12Y150_CQ),
.I5(1'b1),
.O5(CLBLL_L_X2Y149_SLICE_X1Y149_AO5),
.O6(CLBLL_L_X2Y149_SLICE_X1Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y150_SLICE_X0Y150_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y150_SLICE_X0Y150_DO5),
.O6(CLBLL_L_X2Y150_SLICE_X0Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y150_SLICE_X0Y150_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y150_SLICE_X0Y150_CO5),
.O6(CLBLL_L_X2Y150_SLICE_X0Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y150_SLICE_X0Y150_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y150_SLICE_X0Y150_BO5),
.O6(CLBLL_L_X2Y150_SLICE_X0Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y150_SLICE_X0Y150_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y150_SLICE_X0Y150_AO5),
.O6(CLBLL_L_X2Y150_SLICE_X0Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y150_SLICE_X1Y150_A5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X2Y150_SLICE_X1Y150_DO6),
.Q(CLBLL_L_X2Y150_SLICE_X1Y150_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y150_SLICE_X1Y150_C5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X2Y150_SLICE_X1Y150_CO5),
.Q(CLBLL_L_X2Y150_SLICE_X1Y150_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y150_SLICE_X1Y150_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X2Y150_SLICE_X1Y150_AO6),
.Q(CLBLL_L_X2Y150_SLICE_X1Y150_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y150_SLICE_X1Y150_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X2Y150_SLICE_X1Y150_CO6),
.Q(CLBLL_L_X2Y150_SLICE_X1Y150_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcdee012255aa55aa)
  ) CLBLL_L_X2Y150_SLICE_X1Y150_DLUT (
.I0(CLBLM_R_X3Y145_SLICE_X2Y145_DQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLL_L_X4Y151_SLICE_X5Y151_DQ),
.I3(CLBLM_R_X3Y143_SLICE_X2Y143_AQ),
.I4(CLBLM_R_X3Y147_SLICE_X2Y147_C5Q),
.I5(1'b1),
.O5(CLBLL_L_X2Y150_SLICE_X1Y150_DO5),
.O6(CLBLL_L_X2Y150_SLICE_X1Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff00f00fa0afa0a)
  ) CLBLL_L_X2Y150_SLICE_X1Y150_CLUT (
.I0(CLBLL_L_X2Y147_SLICE_X0Y147_BQ),
.I1(1'b1),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X3Y151_SLICE_X3Y151_CQ),
.I4(CLBLM_R_X7Y153_SLICE_X9Y153_AQ),
.I5(1'b1),
.O5(CLBLL_L_X2Y150_SLICE_X1Y150_CO5),
.O6(CLBLL_L_X2Y150_SLICE_X1Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888fffffffc)
  ) CLBLL_L_X2Y150_SLICE_X1Y150_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X3Y153_SLICE_X3Y153_CQ),
.I2(CLBLL_L_X4Y144_SLICE_X5Y144_C5Q),
.I3(CLBLM_R_X3Y151_SLICE_X3Y151_CQ),
.I4(LIOB33_X0Y61_IOB_X0Y61_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y150_SLICE_X1Y150_BO5),
.O6(CLBLL_L_X2Y150_SLICE_X1Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaf3f0c0f0)
  ) CLBLL_L_X2Y150_SLICE_X1Y150_ALUT (
.I0(CLBLM_R_X3Y152_SLICE_X2Y152_AQ),
.I1(CLBLM_L_X8Y146_SLICE_X10Y146_AQ),
.I2(CLBLL_L_X2Y150_SLICE_X1Y150_AQ),
.I3(CLBLM_R_X7Y150_SLICE_X9Y150_CQ),
.I4(CLBLM_R_X3Y148_SLICE_X2Y148_DQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLL_L_X2Y150_SLICE_X1Y150_AO5),
.O6(CLBLL_L_X2Y150_SLICE_X1Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y151_SLICE_X0Y151_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y151_SLICE_X0Y151_DO5),
.O6(CLBLL_L_X2Y151_SLICE_X0Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y151_SLICE_X0Y151_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y151_SLICE_X0Y151_CO5),
.O6(CLBLL_L_X2Y151_SLICE_X0Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y151_SLICE_X0Y151_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y151_SLICE_X0Y151_BO5),
.O6(CLBLL_L_X2Y151_SLICE_X0Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y151_SLICE_X0Y151_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y151_SLICE_X0Y151_AO5),
.O6(CLBLL_L_X2Y151_SLICE_X0Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y151_SLICE_X1Y151_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X2Y151_SLICE_X1Y151_AO6),
.Q(CLBLL_L_X2Y151_SLICE_X1Y151_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y151_SLICE_X1Y151_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X2Y151_SLICE_X1Y151_BO6),
.Q(CLBLL_L_X2Y151_SLICE_X1Y151_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y151_SLICE_X1Y151_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y151_SLICE_X1Y151_DO5),
.O6(CLBLL_L_X2Y151_SLICE_X1Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fffffff80000000)
  ) CLBLL_L_X2Y151_SLICE_X1Y151_CLUT (
.I0(CLBLM_R_X3Y151_SLICE_X2Y151_AQ),
.I1(CLBLM_R_X3Y151_SLICE_X2Y151_A5Q),
.I2(CLBLM_R_X3Y147_SLICE_X3Y147_B5Q),
.I3(CLBLM_R_X3Y151_SLICE_X3Y151_DQ),
.I4(CLBLL_L_X2Y151_SLICE_X1Y151_AQ),
.I5(LIOB33_X0Y55_IOB_X0Y55_I),
.O5(CLBLL_L_X2Y151_SLICE_X1Y151_CO5),
.O6(CLBLL_L_X2Y151_SLICE_X1Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfeffffff32333333)
  ) CLBLL_L_X2Y151_SLICE_X1Y151_BLUT (
.I0(CLBLM_R_X3Y144_SLICE_X3Y144_CQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X5Y144_SLICE_X7Y144_CQ),
.I3(CLBLM_R_X7Y144_SLICE_X9Y144_AQ),
.I4(CLBLM_R_X3Y152_SLICE_X3Y152_AQ),
.I5(CLBLL_L_X2Y149_SLICE_X1Y149_CQ),
.O5(CLBLL_L_X2Y151_SLICE_X1Y151_BO5),
.O6(CLBLL_L_X2Y151_SLICE_X1Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfeee3222dddd1111)
  ) CLBLL_L_X2Y151_SLICE_X1Y151_ALUT (
.I0(CLBLM_R_X3Y151_SLICE_X2Y151_CO6),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(LIOB33_X0Y55_IOB_X0Y55_I),
.I3(CLBLM_R_X3Y151_SLICE_X2Y151_AQ),
.I4(CLBLM_R_X5Y149_SLICE_X7Y149_CQ),
.I5(CLBLL_L_X2Y151_SLICE_X1Y151_AQ),
.O5(CLBLL_L_X2Y151_SLICE_X1Y151_AO5),
.O6(CLBLL_L_X2Y151_SLICE_X1Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y152_SLICE_X0Y152_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y152_SLICE_X0Y152_DO5),
.O6(CLBLL_L_X2Y152_SLICE_X0Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y152_SLICE_X0Y152_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y152_SLICE_X0Y152_CO5),
.O6(CLBLL_L_X2Y152_SLICE_X0Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y152_SLICE_X0Y152_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y152_SLICE_X0Y152_BO5),
.O6(CLBLL_L_X2Y152_SLICE_X0Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y152_SLICE_X0Y152_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y152_SLICE_X0Y152_AO5),
.O6(CLBLL_L_X2Y152_SLICE_X0Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y152_SLICE_X1Y152_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y152_SLICE_X1Y152_DO5),
.O6(CLBLL_L_X2Y152_SLICE_X1Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y152_SLICE_X1Y152_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y152_SLICE_X1Y152_CO5),
.O6(CLBLL_L_X2Y152_SLICE_X1Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y152_SLICE_X1Y152_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y152_SLICE_X1Y152_BO5),
.O6(CLBLL_L_X2Y152_SLICE_X1Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0ffffffff)
  ) CLBLL_L_X2Y152_SLICE_X1Y152_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLL_L_X4Y145_SLICE_X5Y145_BQ),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLL_L_X2Y150_SLICE_X1Y150_A5Q),
.O5(CLBLL_L_X2Y152_SLICE_X1Y152_AO5),
.O6(CLBLL_L_X2Y152_SLICE_X1Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y153_SLICE_X0Y153_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y153_SLICE_X0Y153_DO5),
.O6(CLBLL_L_X2Y153_SLICE_X0Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y153_SLICE_X0Y153_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y153_SLICE_X0Y153_CO5),
.O6(CLBLL_L_X2Y153_SLICE_X0Y153_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y153_SLICE_X0Y153_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y153_SLICE_X0Y153_BO5),
.O6(CLBLL_L_X2Y153_SLICE_X0Y153_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y153_SLICE_X0Y153_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y153_SLICE_X0Y153_AO5),
.O6(CLBLL_L_X2Y153_SLICE_X0Y153_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y153_SLICE_X1Y153_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X3Y153_SLICE_X2Y153_AO6),
.Q(CLBLL_L_X2Y153_SLICE_X1Y153_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y153_SLICE_X1Y153_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y153_SLICE_X1Y153_DO5),
.O6(CLBLL_L_X2Y153_SLICE_X1Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y153_SLICE_X1Y153_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y153_SLICE_X1Y153_CO5),
.O6(CLBLL_L_X2Y153_SLICE_X1Y153_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y153_SLICE_X1Y153_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y153_SLICE_X1Y153_BO5),
.O6(CLBLL_L_X2Y153_SLICE_X1Y153_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y153_SLICE_X1Y153_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y153_SLICE_X1Y153_AO5),
.O6(CLBLL_L_X2Y153_SLICE_X1Y153_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y166_SLICE_X0Y166_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y166_SLICE_X0Y166_DO5),
.O6(CLBLL_L_X2Y166_SLICE_X0Y166_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y166_SLICE_X0Y166_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y166_SLICE_X0Y166_CO5),
.O6(CLBLL_L_X2Y166_SLICE_X0Y166_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y166_SLICE_X0Y166_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y166_SLICE_X0Y166_BO5),
.O6(CLBLL_L_X2Y166_SLICE_X0Y166_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ffff0000ffff)
  ) CLBLL_L_X2Y166_SLICE_X0Y166_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X11Y143_SLICE_X14Y143_AQ),
.I5(1'b1),
.O5(CLBLL_L_X2Y166_SLICE_X0Y166_AO5),
.O6(CLBLL_L_X2Y166_SLICE_X0Y166_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y166_SLICE_X1Y166_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y166_SLICE_X1Y166_DO5),
.O6(CLBLL_L_X2Y166_SLICE_X1Y166_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y166_SLICE_X1Y166_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y166_SLICE_X1Y166_CO5),
.O6(CLBLL_L_X2Y166_SLICE_X1Y166_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y166_SLICE_X1Y166_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y166_SLICE_X1Y166_BO5),
.O6(CLBLL_L_X2Y166_SLICE_X1Y166_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y166_SLICE_X1Y166_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y166_SLICE_X1Y166_AO5),
.O6(CLBLL_L_X2Y166_SLICE_X1Y166_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y140_SLICE_X4Y140_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y140_SLICE_X4Y140_DO5),
.O6(CLBLL_L_X4Y140_SLICE_X4Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y140_SLICE_X4Y140_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y140_SLICE_X4Y140_CO5),
.O6(CLBLL_L_X4Y140_SLICE_X4Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y140_SLICE_X4Y140_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y140_SLICE_X4Y140_BO5),
.O6(CLBLL_L_X4Y140_SLICE_X4Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y140_SLICE_X4Y140_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y140_SLICE_X4Y140_AO5),
.O6(CLBLL_L_X4Y140_SLICE_X4Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y140_SLICE_X5Y140_A_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y140_SLICE_X5Y140_AO6),
.Q(CLBLL_L_X4Y140_SLICE_X5Y140_AQ),
.S(CLBLL_L_X4Y145_SLICE_X5Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y140_SLICE_X5Y140_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y140_SLICE_X5Y140_DO5),
.O6(CLBLL_L_X4Y140_SLICE_X5Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3000300000000000)
  ) CLBLL_L_X4Y140_SLICE_X5Y140_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y153_SLICE_X7Y153_CO6),
.I2(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I3(CLBLL_L_X4Y147_SLICE_X4Y147_D5Q),
.I4(1'b1),
.I5(CLBLL_L_X4Y150_SLICE_X4Y150_AQ),
.O5(CLBLL_L_X4Y140_SLICE_X5Y140_CO5),
.O6(CLBLL_L_X4Y140_SLICE_X5Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000044004400)
  ) CLBLL_L_X4Y140_SLICE_X5Y140_BLUT (
.I0(RIOB33_X105Y101_IOB_X1Y102_I),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(1'b1),
.I3(CLBLL_L_X4Y150_SLICE_X4Y150_AQ),
.I4(1'b1),
.I5(CLBLM_R_X5Y153_SLICE_X7Y153_CO6),
.O5(CLBLL_L_X4Y140_SLICE_X5Y140_BO5),
.O6(CLBLL_L_X4Y140_SLICE_X5Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000ff000000)
  ) CLBLL_L_X4Y140_SLICE_X5Y140_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X8Y150_SLICE_X11Y150_B5Q),
.I5(1'b1),
.O5(CLBLL_L_X4Y140_SLICE_X5Y140_AO5),
.O6(CLBLL_L_X4Y140_SLICE_X5Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y141_SLICE_X4Y141_A_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y141_SLICE_X2Y141_AO6),
.Q(CLBLL_L_X4Y141_SLICE_X4Y141_AQ),
.S(CLBLM_R_X11Y148_SLICE_X15Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y141_SLICE_X4Y141_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y141_SLICE_X4Y141_DO5),
.O6(CLBLL_L_X4Y141_SLICE_X4Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y141_SLICE_X4Y141_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y141_SLICE_X4Y141_CO5),
.O6(CLBLL_L_X4Y141_SLICE_X4Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y141_SLICE_X4Y141_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y141_SLICE_X4Y141_BO5),
.O6(CLBLL_L_X4Y141_SLICE_X4Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y141_SLICE_X4Y141_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y141_SLICE_X4Y141_AO5),
.O6(CLBLL_L_X4Y141_SLICE_X4Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y141_SLICE_X5Y141_A5_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y141_SLICE_X5Y141_AO5),
.Q(CLBLL_L_X4Y141_SLICE_X5Y141_A5Q),
.S(CLBLL_L_X4Y145_SLICE_X5Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y141_SLICE_X5Y141_A_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y141_SLICE_X5Y141_AO6),
.Q(CLBLL_L_X4Y141_SLICE_X5Y141_AQ),
.S(CLBLL_L_X4Y145_SLICE_X5Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y141_SLICE_X5Y141_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y141_SLICE_X5Y141_DO5),
.O6(CLBLL_L_X4Y141_SLICE_X5Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000ffff0000)
  ) CLBLL_L_X4Y141_SLICE_X5Y141_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X3Y152_SLICE_X3Y152_AQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLL_L_X4Y141_SLICE_X5Y141_CO5),
.O6(CLBLL_L_X4Y141_SLICE_X5Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h70f0f0f055ffffff)
  ) CLBLL_L_X4Y141_SLICE_X5Y141_BLUT (
.I0(LIOB33_X0Y57_IOB_X0Y58_I),
.I1(CLBLM_R_X3Y142_SLICE_X3Y142_BQ),
.I2(CLBLL_L_X4Y142_SLICE_X5Y142_AQ),
.I3(CLBLL_L_X4Y142_SLICE_X5Y142_A5Q),
.I4(CLBLL_L_X2Y143_SLICE_X1Y143_CQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y141_SLICE_X5Y141_BO5),
.O6(CLBLL_L_X4Y141_SLICE_X5Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00f000f000)
  ) CLBLL_L_X4Y141_SLICE_X5Y141_ALUT (
.I0(CLBLM_R_X5Y143_SLICE_X6Y143_D5Q),
.I1(1'b1),
.I2(CLBLL_L_X4Y140_SLICE_X5Y140_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y141_SLICE_X5Y141_AO5),
.O6(CLBLL_L_X4Y141_SLICE_X5Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y142_SLICE_X4Y142_A5_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y142_SLICE_X4Y142_CO6),
.Q(CLBLL_L_X4Y142_SLICE_X4Y142_A5Q),
.S(CLBLL_L_X4Y141_SLICE_X5Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y142_SLICE_X4Y142_A_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y142_SLICE_X4Y142_AO6),
.Q(CLBLL_L_X4Y142_SLICE_X4Y142_AQ),
.S(CLBLL_L_X4Y141_SLICE_X5Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8088800088008800)
  ) CLBLL_L_X4Y142_SLICE_X4Y142_DLUT (
.I0(CLBLL_L_X4Y142_SLICE_X5Y142_AQ),
.I1(CLBLM_R_X3Y142_SLICE_X3Y142_BQ),
.I2(CLBLL_L_X4Y141_SLICE_X5Y141_BO5),
.I3(CLBLM_L_X10Y142_SLICE_X12Y142_AQ),
.I4(CLBLL_L_X4Y142_SLICE_X5Y142_BQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y142_SLICE_X4Y142_DO5),
.O6(CLBLL_L_X4Y142_SLICE_X4Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa000030ff3030)
  ) CLBLL_L_X4Y142_SLICE_X4Y142_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X10Y143_SLICE_X12Y143_AO5),
.I2(CLBLL_L_X4Y143_SLICE_X4Y143_DQ),
.I3(CLBLM_L_X10Y143_SLICE_X12Y143_BO6),
.I4(CLBLL_L_X2Y143_SLICE_X1Y143_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y142_SLICE_X4Y142_CO5),
.O6(CLBLL_L_X4Y142_SLICE_X4Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hd1f3e2c055555555)
  ) CLBLL_L_X4Y142_SLICE_X4Y142_BLUT (
.I0(LIOB33_X0Y57_IOB_X0Y58_I),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLL_L_X4Y143_SLICE_X4Y143_AQ),
.I3(CLBLL_L_X2Y143_SLICE_X1Y143_CQ),
.I4(CLBLL_L_X4Y142_SLICE_X5Y142_A5Q),
.I5(1'b1),
.O5(CLBLL_L_X4Y142_SLICE_X4Y142_BO5),
.O6(CLBLL_L_X4Y142_SLICE_X4Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00cc00cc00)
  ) CLBLL_L_X4Y142_SLICE_X4Y142_ALUT (
.I0(1'b1),
.I1(CLBLL_L_X2Y148_SLICE_X0Y148_BQ),
.I2(1'b1),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y142_SLICE_X4Y142_AO5),
.O6(CLBLL_L_X4Y142_SLICE_X4Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y142_SLICE_X5Y142_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y142_SLICE_X4Y142_BO6),
.Q(CLBLL_L_X4Y142_SLICE_X5Y142_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y142_SLICE_X5Y142_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y142_SLICE_X5Y142_AO6),
.Q(CLBLL_L_X4Y142_SLICE_X5Y142_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y142_SLICE_X5Y142_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y142_SLICE_X5Y142_BO6),
.Q(CLBLL_L_X4Y142_SLICE_X5Y142_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y142_SLICE_X5Y142_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y142_SLICE_X5Y142_CO6),
.Q(CLBLL_L_X4Y142_SLICE_X5Y142_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0c0cff0c0c0cff0c)
  ) CLBLL_L_X4Y142_SLICE_X5Y142_DLUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y142_SLICE_X5Y142_CQ),
.I2(CLBLM_L_X10Y143_SLICE_X12Y143_AO5),
.I3(CLBLL_L_X4Y143_SLICE_X5Y143_BQ),
.I4(CLBLM_L_X10Y143_SLICE_X12Y143_BO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y142_SLICE_X5Y142_DO5),
.O6(CLBLL_L_X4Y142_SLICE_X5Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0ff00cc00)
  ) CLBLL_L_X4Y142_SLICE_X5Y142_CLUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y142_SLICE_X5Y142_CQ),
.I2(CLBLM_L_X10Y150_SLICE_X13Y150_B5Q),
.I3(CLBLM_L_X10Y143_SLICE_X12Y143_AO6),
.I4(CLBLL_L_X4Y143_SLICE_X4Y143_BQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLL_L_X4Y142_SLICE_X5Y142_CO5),
.O6(CLBLL_L_X4Y142_SLICE_X5Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'heecc2200cccc0000)
  ) CLBLL_L_X4Y142_SLICE_X5Y142_BLUT (
.I0(LIOB33_X0Y57_IOB_X0Y58_I),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(1'b1),
.I3(CLBLL_L_X2Y143_SLICE_X1Y143_CQ),
.I4(CLBLM_R_X5Y143_SLICE_X6Y143_AQ),
.I5(CLBLL_L_X4Y142_SLICE_X5Y142_A5Q),
.O5(CLBLL_L_X4Y142_SLICE_X5Y142_BO5),
.O6(CLBLL_L_X4Y142_SLICE_X5Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff000f0fff500f5)
  ) CLBLL_L_X4Y142_SLICE_X5Y142_ALUT (
.I0(CLBLM_L_X10Y142_SLICE_X12Y142_AQ),
.I1(1'b1),
.I2(CLBLL_L_X4Y141_SLICE_X5Y141_BO6),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X10Y147_SLICE_X13Y147_A5Q),
.I5(CLBLM_R_X3Y141_SLICE_X3Y141_CO6),
.O5(CLBLL_L_X4Y142_SLICE_X5Y142_AO5),
.O6(CLBLL_L_X4Y142_SLICE_X5Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y143_SLICE_X4Y143_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y143_SLICE_X4Y143_AO6),
.Q(CLBLL_L_X4Y143_SLICE_X4Y143_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y143_SLICE_X4Y143_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y143_SLICE_X4Y143_BO6),
.Q(CLBLL_L_X4Y143_SLICE_X4Y143_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y143_SLICE_X4Y143_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y143_SLICE_X4Y143_CO6),
.Q(CLBLL_L_X4Y143_SLICE_X4Y143_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y143_SLICE_X4Y143_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y143_SLICE_X4Y143_DO6),
.Q(CLBLL_L_X4Y143_SLICE_X4Y143_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000ccf0ccf0)
  ) CLBLL_L_X4Y143_SLICE_X4Y143_DLUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y143_SLICE_X4Y143_AQ),
.I2(CLBLL_L_X4Y143_SLICE_X4Y143_DQ),
.I3(CLBLM_L_X10Y143_SLICE_X12Y143_AO6),
.I4(CLBLL_L_X4Y143_SLICE_X5Y143_BQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLL_L_X4Y143_SLICE_X4Y143_DO5),
.O6(CLBLL_L_X4Y143_SLICE_X4Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f000880000)
  ) CLBLL_L_X4Y143_SLICE_X4Y143_CLUT (
.I0(CLBLL_L_X4Y142_SLICE_X5Y142_AQ),
.I1(CLBLM_L_X10Y142_SLICE_X12Y142_AQ),
.I2(CLBLL_L_X4Y147_SLICE_X4Y147_CQ),
.I3(CLBLM_R_X3Y142_SLICE_X3Y142_BQ),
.I4(CLBLM_R_X7Y150_SLICE_X9Y150_B5Q),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLL_L_X4Y143_SLICE_X4Y143_CO5),
.O6(CLBLL_L_X4Y143_SLICE_X4Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefe0e0ef0fe000e)
  ) CLBLL_L_X4Y143_SLICE_X4Y143_BLUT (
.I0(CLBLL_L_X2Y144_SLICE_X1Y144_BQ),
.I1(CLBLL_L_X4Y143_SLICE_X4Y143_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X5Y149_SLICE_X6Y149_D5Q),
.I4(CLBLL_L_X4Y150_SLICE_X4Y150_AQ),
.I5(CLBLM_L_X8Y150_SLICE_X11Y150_B5Q),
.O5(CLBLL_L_X4Y143_SLICE_X4Y143_BO5),
.O6(CLBLL_L_X4Y143_SLICE_X4Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefe5454aafe0054)
  ) CLBLL_L_X4Y143_SLICE_X4Y143_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLL_L_X2Y147_SLICE_X1Y147_AQ),
.I2(CLBLL_L_X4Y143_SLICE_X4Y143_AQ),
.I3(CLBLM_R_X5Y149_SLICE_X6Y149_D5Q),
.I4(CLBLM_L_X8Y149_SLICE_X11Y149_BQ),
.I5(CLBLM_L_X8Y150_SLICE_X11Y150_B5Q),
.O5(CLBLL_L_X4Y143_SLICE_X4Y143_AO5),
.O6(CLBLL_L_X4Y143_SLICE_X4Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y143_SLICE_X5Y143_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y143_SLICE_X5Y143_CO5),
.Q(CLBLL_L_X4Y143_SLICE_X5Y143_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y143_SLICE_X5Y143_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y143_SLICE_X5Y143_AO6),
.Q(CLBLL_L_X4Y143_SLICE_X5Y143_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y143_SLICE_X5Y143_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y143_SLICE_X5Y143_BO6),
.Q(CLBLL_L_X4Y143_SLICE_X5Y143_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y143_SLICE_X5Y143_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y143_SLICE_X5Y143_CO6),
.Q(CLBLL_L_X4Y143_SLICE_X5Y143_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y143_SLICE_X5Y143_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y143_SLICE_X5Y143_DO6),
.Q(CLBLL_L_X4Y143_SLICE_X5Y143_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffc4ffc800c400c8)
  ) CLBLL_L_X4Y143_SLICE_X5Y143_DLUT (
.I0(CLBLM_R_X5Y143_SLICE_X6Y143_D5Q),
.I1(CLBLM_L_X8Y143_SLICE_X11Y143_A5Q),
.I2(CLBLL_L_X4Y143_SLICE_X5Y143_DQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(RIOB33_X105Y109_IOB_X1Y109_I),
.I5(CLBLL_L_X2Y149_SLICE_X1Y149_BQ),
.O5(CLBLL_L_X4Y143_SLICE_X5Y143_DO5),
.O6(CLBLL_L_X4Y143_SLICE_X5Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaa00f0ccf0cc)
  ) CLBLL_L_X4Y143_SLICE_X5Y143_CLUT (
.I0(CLBLM_R_X11Y143_SLICE_X14Y143_AQ),
.I1(CLBLL_L_X2Y153_SLICE_X1Y153_AQ),
.I2(CLBLM_L_X8Y140_SLICE_X10Y140_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(RIOB33_X105Y101_IOB_X1Y101_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y143_SLICE_X5Y143_CO5),
.O6(CLBLL_L_X4Y143_SLICE_X5Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaaffca00aa00ca)
  ) CLBLL_L_X4Y143_SLICE_X5Y143_BLUT (
.I0(CLBLL_L_X2Y145_SLICE_X1Y145_AQ),
.I1(CLBLL_L_X4Y143_SLICE_X5Y143_BQ),
.I2(CLBLM_R_X3Y148_SLICE_X2Y148_D5Q),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X5Y144_SLICE_X6Y144_DQ),
.I5(CLBLM_R_X5Y150_SLICE_X7Y150_A5Q),
.O5(CLBLL_L_X4Y143_SLICE_X5Y143_BO5),
.O6(CLBLL_L_X4Y143_SLICE_X5Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaccaaf0aaccaa0f)
  ) CLBLL_L_X4Y143_SLICE_X5Y143_ALUT (
.I0(CLBLM_R_X5Y143_SLICE_X7Y143_DQ),
.I1(CLBLM_R_X5Y142_SLICE_X6Y142_CQ),
.I2(CLBLL_L_X4Y143_SLICE_X5Y143_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X8Y149_SLICE_X11Y149_BQ),
.I5(CLBLM_R_X7Y142_SLICE_X8Y142_DO6),
.O5(CLBLL_L_X4Y143_SLICE_X5Y143_AO5),
.O6(CLBLL_L_X4Y143_SLICE_X5Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y144_SLICE_X4Y144_A_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y150_SLICE_X12Y150_DO5),
.Q(CLBLL_L_X4Y144_SLICE_X4Y144_AQ),
.S(CLBLL_L_X4Y145_SLICE_X5Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0fff0fffffffffff)
  ) CLBLL_L_X4Y144_SLICE_X4Y144_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X3Y152_SLICE_X3Y152_AQ),
.I3(CLBLM_R_X7Y144_SLICE_X9Y144_AQ),
.I4(1'b1),
.I5(CLBLM_R_X7Y152_SLICE_X8Y152_BQ),
.O5(CLBLL_L_X4Y144_SLICE_X4Y144_DO5),
.O6(CLBLL_L_X4Y144_SLICE_X4Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5a5affffffff5a5a)
  ) CLBLL_L_X4Y144_SLICE_X4Y144_CLUT (
.I0(CLBLM_R_X7Y142_SLICE_X9Y142_A5Q),
.I1(1'b1),
.I2(CLBLM_R_X3Y146_SLICE_X2Y146_BQ),
.I3(1'b1),
.I4(CLBLM_R_X3Y145_SLICE_X2Y145_B5Q),
.I5(CLBLL_L_X4Y144_SLICE_X5Y144_BQ),
.O5(CLBLL_L_X4Y144_SLICE_X4Y144_CO5),
.O6(CLBLL_L_X4Y144_SLICE_X4Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000050005)
  ) CLBLL_L_X4Y144_SLICE_X4Y144_BLUT (
.I0(CLBLM_R_X3Y145_SLICE_X3Y145_AQ),
.I1(1'b1),
.I2(CLBLM_R_X7Y143_SLICE_X9Y143_DQ),
.I3(CLBLL_L_X2Y143_SLICE_X1Y143_BQ),
.I4(1'b1),
.I5(CLBLL_L_X4Y147_SLICE_X5Y147_C5Q),
.O5(CLBLL_L_X4Y144_SLICE_X4Y144_BO5),
.O6(CLBLL_L_X4Y144_SLICE_X4Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff3fcff3fc)
  ) CLBLL_L_X4Y144_SLICE_X4Y144_ALUT (
.I0(1'b1),
.I1(CLBLL_L_X2Y153_SLICE_X1Y153_AQ),
.I2(CLBLM_R_X5Y143_SLICE_X6Y143_DQ),
.I3(CLBLM_R_X3Y144_SLICE_X3Y144_DQ),
.I4(CLBLM_R_X3Y146_SLICE_X3Y146_C5Q),
.I5(CLBLL_L_X4Y144_SLICE_X4Y144_CO6),
.O5(CLBLL_L_X4Y144_SLICE_X4Y144_AO5),
.O6(CLBLL_L_X4Y144_SLICE_X4Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y144_SLICE_X5Y144_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y144_SLICE_X5Y144_BO5),
.Q(CLBLL_L_X4Y144_SLICE_X5Y144_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y144_SLICE_X5Y144_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y144_SLICE_X5Y144_CO5),
.Q(CLBLL_L_X4Y144_SLICE_X5Y144_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y144_SLICE_X5Y144_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y144_SLICE_X5Y144_DO5),
.Q(CLBLL_L_X4Y144_SLICE_X5Y144_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y144_SLICE_X5Y144_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y144_SLICE_X5Y144_AO6),
.Q(CLBLL_L_X4Y144_SLICE_X5Y144_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y144_SLICE_X5Y144_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y144_SLICE_X5Y144_BO6),
.Q(CLBLL_L_X4Y144_SLICE_X5Y144_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y144_SLICE_X5Y144_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y144_SLICE_X5Y144_CO6),
.Q(CLBLL_L_X4Y144_SLICE_X5Y144_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y144_SLICE_X5Y144_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y144_SLICE_X5Y144_DO6),
.Q(CLBLL_L_X4Y144_SLICE_X5Y144_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff33cc00bbbb8888)
  ) CLBLL_L_X4Y144_SLICE_X5Y144_DLUT (
.I0(CLBLM_R_X3Y143_SLICE_X2Y143_BQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(1'b1),
.I3(CLBLL_L_X4Y152_SLICE_X5Y152_CQ),
.I4(CLBLM_L_X8Y152_SLICE_X11Y152_A5Q),
.I5(1'b1),
.O5(CLBLL_L_X4Y144_SLICE_X5Y144_DO5),
.O6(CLBLL_L_X4Y144_SLICE_X5Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccaaccaaf0ccf0cc)
  ) CLBLL_L_X4Y144_SLICE_X5Y144_CLUT (
.I0(CLBLM_R_X5Y142_SLICE_X7Y142_CQ),
.I1(CLBLL_L_X4Y153_SLICE_X4Y153_A5Q),
.I2(CLBLL_L_X4Y146_SLICE_X5Y146_A5Q),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y144_SLICE_X5Y144_CO5),
.O6(CLBLL_L_X4Y144_SLICE_X5Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0aaf0aaaaffaa00)
  ) CLBLL_L_X4Y144_SLICE_X5Y144_BLUT (
.I0(CLBLM_R_X3Y145_SLICE_X2Y145_B5Q),
.I1(1'b1),
.I2(CLBLL_L_X4Y144_SLICE_X5Y144_CQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLL_L_X2Y149_SLICE_X1Y149_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y144_SLICE_X5Y144_BO5),
.O6(CLBLL_L_X4Y144_SLICE_X5Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000ccf0ccf0)
  ) CLBLL_L_X4Y144_SLICE_X5Y144_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y144_SLICE_X6Y144_AQ),
.I2(CLBLL_L_X4Y144_SLICE_X5Y144_AQ),
.I3(CLBLM_L_X10Y143_SLICE_X12Y143_BO6),
.I4(CLBLM_R_X7Y142_SLICE_X9Y142_A5Q),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLL_L_X4Y144_SLICE_X5Y144_AO5),
.O6(CLBLL_L_X4Y144_SLICE_X5Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y145_SLICE_X4Y145_A5_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y145_SLICE_X4Y145_AO5),
.Q(CLBLL_L_X4Y145_SLICE_X4Y145_A5Q),
.S(CLBLL_L_X4Y145_SLICE_X4Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y145_SLICE_X4Y145_A_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y145_SLICE_X4Y145_AO6),
.Q(CLBLL_L_X4Y145_SLICE_X4Y145_AQ),
.S(CLBLL_L_X4Y145_SLICE_X4Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ffff00000000)
  ) CLBLL_L_X4Y145_SLICE_X4Y145_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLL_L_X4Y153_SLICE_X5Y153_BQ),
.O5(CLBLL_L_X4Y145_SLICE_X4Y145_DO5),
.O6(CLBLL_L_X4Y145_SLICE_X4Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haffaffffffffaffa)
  ) CLBLL_L_X4Y145_SLICE_X4Y145_CLUT (
.I0(CLBLM_R_X3Y144_SLICE_X2Y144_BO5),
.I1(1'b1),
.I2(CLBLM_R_X3Y145_SLICE_X2Y145_C5Q),
.I3(CLBLM_R_X5Y145_SLICE_X6Y145_BQ),
.I4(CLBLM_R_X3Y145_SLICE_X2Y145_CQ),
.I5(CLBLL_L_X4Y147_SLICE_X5Y147_BQ),
.O5(CLBLL_L_X4Y145_SLICE_X4Y145_CO5),
.O6(CLBLL_L_X4Y145_SLICE_X4Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000054)
  ) CLBLL_L_X4Y145_SLICE_X4Y145_BLUT (
.I0(CLBLM_L_X10Y142_SLICE_X12Y142_AQ),
.I1(CLBLL_L_X4Y145_SLICE_X4Y145_CO6),
.I2(CLBLL_L_X4Y144_SLICE_X4Y144_AO6),
.I3(CLBLM_R_X3Y142_SLICE_X3Y142_BQ),
.I4(CLBLL_L_X4Y142_SLICE_X5Y142_AQ),
.I5(CLBLM_R_X3Y143_SLICE_X2Y143_CQ),
.O5(CLBLL_L_X4Y145_SLICE_X4Y145_BO5),
.O6(CLBLL_L_X4Y145_SLICE_X4Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888cc00cc00)
  ) CLBLL_L_X4Y145_SLICE_X4Y145_ALUT (
.I0(CLBLL_L_X2Y148_SLICE_X0Y148_B5Q),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(1'b1),
.I3(CLBLL_L_X2Y143_SLICE_X1Y143_CQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y145_SLICE_X4Y145_AO5),
.O6(CLBLL_L_X4Y145_SLICE_X4Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y145_SLICE_X5Y145_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLL_L_X4Y142_SLICE_X5Y142_AQ),
.Q(CLBLL_L_X4Y145_SLICE_X5Y145_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y145_SLICE_X5Y145_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_R_X5Y144_SLICE_X6Y144_CQ),
.Q(CLBLL_L_X4Y145_SLICE_X5Y145_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y145_SLICE_X5Y145_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y145_SLICE_X5Y145_DO5),
.O6(CLBLL_L_X4Y145_SLICE_X5Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000aaaaaaaa)
  ) CLBLL_L_X4Y145_SLICE_X5Y145_CLUT (
.I0(CLBLM_R_X7Y152_SLICE_X8Y152_BQ),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLL_L_X4Y145_SLICE_X5Y145_CO5),
.O6(CLBLL_L_X4Y145_SLICE_X5Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000cccc0000cccc)
  ) CLBLL_L_X4Y145_SLICE_X5Y145_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y150_SLICE_X8Y150_C5Q),
.I2(1'b1),
.I3(1'b1),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y145_SLICE_X5Y145_BO5),
.O6(CLBLL_L_X4Y145_SLICE_X5Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcccfeeefcccfeee)
  ) CLBLL_L_X4Y145_SLICE_X5Y145_ALUT (
.I0(CLBLL_L_X4Y141_SLICE_X4Y141_AQ),
.I1(CLBLM_L_X12Y149_SLICE_X16Y149_CO6),
.I2(CLBLM_L_X10Y143_SLICE_X12Y143_BO6),
.I3(CLBLM_R_X3Y145_SLICE_X2Y145_AQ),
.I4(CLBLM_R_X7Y146_SLICE_X8Y146_AO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y145_SLICE_X5Y145_AO5),
.O6(CLBLL_L_X4Y145_SLICE_X5Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y146_SLICE_X4Y146_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y146_SLICE_X4Y146_AO6),
.Q(CLBLL_L_X4Y146_SLICE_X4Y146_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y146_SLICE_X4Y146_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y146_SLICE_X4Y146_BO6),
.Q(CLBLL_L_X4Y146_SLICE_X4Y146_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y146_SLICE_X4Y146_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y146_SLICE_X4Y146_CO6),
.Q(CLBLL_L_X4Y146_SLICE_X4Y146_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y146_SLICE_X4Y146_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y146_SLICE_X4Y146_DO6),
.Q(CLBLL_L_X4Y146_SLICE_X4Y146_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefe5454aaaa0000)
  ) CLBLL_L_X4Y146_SLICE_X4Y146_DLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X3Y146_SLICE_X3Y146_BQ),
.I2(CLBLL_L_X4Y146_SLICE_X4Y146_DQ),
.I3(1'b1),
.I4(CLBLL_L_X4Y147_SLICE_X4Y147_DQ),
.I5(CLBLM_L_X10Y143_SLICE_X12Y143_AO6),
.O5(CLBLL_L_X4Y146_SLICE_X4Y146_DO5),
.O6(CLBLL_L_X4Y146_SLICE_X4Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5a0f5a0e4e4e4e4)
  ) CLBLL_L_X4Y146_SLICE_X4Y146_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLL_L_X4Y146_SLICE_X4Y146_CQ),
.I2(CLBLM_R_X3Y149_SLICE_X2Y149_CQ),
.I3(CLBLM_R_X5Y147_SLICE_X6Y147_AQ),
.I4(1'b1),
.I5(CLBLM_L_X10Y143_SLICE_X12Y143_AO6),
.O5(CLBLL_L_X4Y146_SLICE_X4Y146_CO5),
.O6(CLBLL_L_X4Y146_SLICE_X4Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f3f3f3f3f3f3c0)
  ) CLBLL_L_X4Y146_SLICE_X4Y146_BLUT (
.I0(1'b1),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X3Y142_SLICE_X2Y142_BQ),
.I3(CLBLL_L_X2Y148_SLICE_X0Y148_BQ),
.I4(CLBLM_R_X3Y144_SLICE_X3Y144_D5Q),
.I5(CLBLL_L_X4Y148_SLICE_X5Y148_CQ),
.O5(CLBLL_L_X4Y146_SLICE_X4Y146_BO5),
.O6(CLBLL_L_X4Y146_SLICE_X4Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haafcaafcaa30aa30)
  ) CLBLL_L_X4Y146_SLICE_X4Y146_ALUT (
.I0(CLBLM_L_X8Y146_SLICE_X10Y146_DQ),
.I1(CLBLM_L_X10Y143_SLICE_X12Y143_BO6),
.I2(CLBLL_L_X4Y146_SLICE_X4Y146_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(1'b1),
.I5(CLBLM_R_X3Y146_SLICE_X2Y146_AQ),
.O5(CLBLL_L_X4Y146_SLICE_X4Y146_AO5),
.O6(CLBLL_L_X4Y146_SLICE_X4Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y146_SLICE_X5Y146_A5_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y146_SLICE_X5Y146_AO5),
.Q(CLBLL_L_X4Y146_SLICE_X5Y146_A5Q),
.S(CLBLL_L_X4Y146_SLICE_X5Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y146_SLICE_X5Y146_B5_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y146_SLICE_X5Y146_BO5),
.Q(CLBLL_L_X4Y146_SLICE_X5Y146_B5Q),
.S(CLBLL_L_X4Y146_SLICE_X5Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y146_SLICE_X5Y146_A_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y146_SLICE_X5Y146_AO6),
.Q(CLBLL_L_X4Y146_SLICE_X5Y146_AQ),
.S(CLBLL_L_X4Y146_SLICE_X5Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y146_SLICE_X5Y146_B_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y146_SLICE_X5Y146_BO6),
.Q(CLBLL_L_X4Y146_SLICE_X5Y146_BQ),
.S(CLBLL_L_X4Y146_SLICE_X5Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5500550055005500)
  ) CLBLL_L_X4Y146_SLICE_X5Y146_DLUT (
.I0(CLBLM_R_X7Y142_SLICE_X8Y142_DO6),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLL_L_X4Y143_SLICE_X5Y143_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y146_SLICE_X5Y146_DO5),
.O6(CLBLL_L_X4Y146_SLICE_X5Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h4444444444444444)
  ) CLBLL_L_X4Y146_SLICE_X5Y146_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X7Y144_SLICE_X9Y144_AQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y146_SLICE_X5Y146_CO5),
.O6(CLBLL_L_X4Y146_SLICE_X5Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0000f0f00000)
  ) CLBLL_L_X4Y146_SLICE_X5Y146_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y142_SLICE_X11Y142_BQ),
.I2(CLBLL_L_X2Y146_SLICE_X1Y146_AQ),
.I3(1'b1),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y146_SLICE_X5Y146_BO5),
.O6(CLBLL_L_X4Y146_SLICE_X5Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000aa00aa00)
  ) CLBLL_L_X4Y146_SLICE_X5Y146_ALUT (
.I0(CLBLM_R_X7Y148_SLICE_X9Y148_AQ),
.I1(1'b1),
.I2(CLBLL_L_X4Y144_SLICE_X5Y144_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y146_SLICE_X5Y146_AO5),
.O6(CLBLL_L_X4Y146_SLICE_X5Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y147_SLICE_X4Y147_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y147_SLICE_X4Y147_CO5),
.Q(CLBLL_L_X4Y147_SLICE_X4Y147_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y147_SLICE_X4Y147_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y147_SLICE_X4Y147_DO5),
.Q(CLBLL_L_X4Y147_SLICE_X4Y147_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y147_SLICE_X4Y147_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y147_SLICE_X4Y147_AO6),
.Q(CLBLL_L_X4Y147_SLICE_X4Y147_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y147_SLICE_X4Y147_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y147_SLICE_X4Y147_BO6),
.Q(CLBLL_L_X4Y147_SLICE_X4Y147_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y147_SLICE_X4Y147_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y147_SLICE_X4Y147_CO6),
.Q(CLBLL_L_X4Y147_SLICE_X4Y147_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y147_SLICE_X4Y147_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y147_SLICE_X4Y147_DO6),
.Q(CLBLL_L_X4Y147_SLICE_X4Y147_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5a0a0ee44ee44)
  ) CLBLL_L_X4Y147_SLICE_X4Y147_DLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X5Y145_SLICE_X6Y145_B5Q),
.I2(CLBLL_L_X2Y148_SLICE_X1Y148_A5Q),
.I3(CLBLL_L_X2Y144_SLICE_X1Y144_B5Q),
.I4(CLBLM_R_X3Y147_SLICE_X2Y147_C5Q),
.I5(1'b1),
.O5(CLBLL_L_X4Y147_SLICE_X4Y147_DO5),
.O6(CLBLL_L_X4Y147_SLICE_X4Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hbb11ee44f5a0f5a0)
  ) CLBLL_L_X4Y147_SLICE_X4Y147_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X5Y144_SLICE_X7Y144_CQ),
.I2(CLBLL_L_X4Y143_SLICE_X5Y143_DQ),
.I3(CLBLL_L_X2Y150_SLICE_X1Y150_C5Q),
.I4(CLBLM_R_X5Y147_SLICE_X7Y147_C5Q),
.I5(1'b1),
.O5(CLBLL_L_X4Y147_SLICE_X4Y147_CO5),
.O6(CLBLL_L_X4Y147_SLICE_X4Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00000f6fc060c)
  ) CLBLL_L_X4Y147_SLICE_X4Y147_BLUT (
.I0(CLBLL_L_X4Y148_SLICE_X4Y148_CO6),
.I1(CLBLL_L_X4Y147_SLICE_X4Y147_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X3Y147_SLICE_X3Y147_AQ),
.I4(CLBLM_R_X7Y145_SLICE_X8Y145_C5Q),
.I5(CLBLM_R_X3Y146_SLICE_X3Y146_CQ),
.O5(CLBLL_L_X4Y147_SLICE_X4Y147_BO5),
.O6(CLBLL_L_X4Y147_SLICE_X4Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccf0003cccf0003)
  ) CLBLL_L_X4Y147_SLICE_X4Y147_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLL_L_X4Y148_SLICE_X4Y148_CO5),
.I3(CLBLM_R_X3Y147_SLICE_X3Y147_CO5),
.I4(CLBLM_R_X5Y144_SLICE_X7Y144_BQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y147_SLICE_X4Y147_AO5),
.O6(CLBLL_L_X4Y147_SLICE_X4Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y147_SLICE_X5Y147_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y147_SLICE_X5Y147_BO5),
.Q(CLBLL_L_X4Y147_SLICE_X5Y147_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y147_SLICE_X5Y147_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y147_SLICE_X5Y147_CO5),
.Q(CLBLL_L_X4Y147_SLICE_X5Y147_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y147_SLICE_X5Y147_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y147_SLICE_X5Y147_AO6),
.Q(CLBLL_L_X4Y147_SLICE_X5Y147_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y147_SLICE_X5Y147_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y147_SLICE_X5Y147_BO6),
.Q(CLBLL_L_X4Y147_SLICE_X5Y147_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y147_SLICE_X5Y147_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y147_SLICE_X5Y147_CO6),
.Q(CLBLL_L_X4Y147_SLICE_X5Y147_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y147_SLICE_X5Y147_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y147_SLICE_X5Y147_DO6),
.Q(CLBLL_L_X4Y147_SLICE_X5Y147_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccf0f055ff)
  ) CLBLL_L_X4Y147_SLICE_X5Y147_DLUT (
.I0(CLBLM_R_X5Y153_SLICE_X6Y153_BQ),
.I1(CLBLM_R_X3Y148_SLICE_X2Y148_CQ),
.I2(CLBLL_L_X4Y147_SLICE_X5Y147_DQ),
.I3(CLBLL_L_X4Y148_SLICE_X5Y148_CQ),
.I4(CLBLM_R_X5Y154_SLICE_X7Y154_AQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLL_L_X4Y147_SLICE_X5Y147_DO5),
.O6(CLBLL_L_X4Y147_SLICE_X5Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd88dd88bebe1414)
  ) CLBLL_L_X4Y147_SLICE_X5Y147_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X5Y146_SLICE_X6Y146_BQ),
.I2(CLBLM_R_X3Y152_SLICE_X3Y152_AQ),
.I3(CLBLM_R_X7Y148_SLICE_X9Y148_CQ),
.I4(CLBLL_L_X4Y152_SLICE_X4Y152_CQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y147_SLICE_X5Y147_CO5),
.O6(CLBLL_L_X4Y147_SLICE_X5Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hee22ee22fcfc3030)
  ) CLBLL_L_X4Y147_SLICE_X5Y147_BLUT (
.I0(CLBLM_R_X3Y145_SLICE_X2Y145_CQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X3Y147_SLICE_X3Y147_AQ),
.I3(CLBLM_L_X8Y148_SLICE_X11Y148_AQ),
.I4(CLBLL_L_X4Y147_SLICE_X5Y147_C5Q),
.I5(1'b1),
.O5(CLBLL_L_X4Y147_SLICE_X5Y147_BO5),
.O6(CLBLL_L_X4Y147_SLICE_X5Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00ccf0cc5a)
  ) CLBLL_L_X4Y147_SLICE_X5Y147_ALUT (
.I0(CLBLL_L_X4Y150_SLICE_X5Y150_BQ),
.I1(CLBLM_R_X5Y147_SLICE_X7Y147_AQ),
.I2(CLBLL_L_X4Y147_SLICE_X5Y147_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLL_L_X4Y151_SLICE_X4Y151_AO5),
.I5(CLBLM_R_X3Y146_SLICE_X3Y146_CQ),
.O5(CLBLL_L_X4Y147_SLICE_X5Y147_AO5),
.O6(CLBLL_L_X4Y147_SLICE_X5Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y148_SLICE_X4Y148_A5_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y148_SLICE_X4Y148_AO5),
.Q(CLBLL_L_X4Y148_SLICE_X4Y148_A5Q),
.S(CLBLM_R_X5Y153_SLICE_X7Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y148_SLICE_X4Y148_A_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y148_SLICE_X4Y148_AO6),
.Q(CLBLL_L_X4Y148_SLICE_X4Y148_AQ),
.S(CLBLM_R_X5Y153_SLICE_X7Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y148_SLICE_X4Y148_B_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y148_SLICE_X1Y148_BO5),
.Q(CLBLL_L_X4Y148_SLICE_X4Y148_BQ),
.S(CLBLM_R_X5Y153_SLICE_X7Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f3d1f3c0c0e2c0)
  ) CLBLL_L_X4Y148_SLICE_X4Y148_DLUT (
.I0(CLBLL_L_X4Y148_SLICE_X5Y148_AQ),
.I1(CLBLM_L_X8Y149_SLICE_X11Y149_BQ),
.I2(CLBLL_L_X4Y147_SLICE_X4Y147_DQ),
.I3(CLBLL_L_X4Y149_SLICE_X4Y149_AQ),
.I4(CLBLL_L_X4Y148_SLICE_X4Y148_BO5),
.I5(CLBLL_L_X4Y148_SLICE_X5Y148_BQ),
.O5(CLBLL_L_X4Y148_SLICE_X4Y148_DO5),
.O6(CLBLL_L_X4Y148_SLICE_X4Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h800000007fff7fff)
  ) CLBLL_L_X4Y148_SLICE_X4Y148_CLUT (
.I0(CLBLL_L_X4Y147_SLICE_X5Y147_AQ),
.I1(CLBLL_L_X4Y150_SLICE_X5Y150_BQ),
.I2(CLBLM_R_X7Y149_SLICE_X8Y149_AQ),
.I3(CLBLM_R_X7Y150_SLICE_X8Y150_AQ),
.I4(CLBLM_R_X7Y150_SLICE_X8Y150_CQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y148_SLICE_X4Y148_CO5),
.O6(CLBLL_L_X4Y148_SLICE_X4Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h20000000dfffdfff)
  ) CLBLL_L_X4Y148_SLICE_X4Y148_BLUT (
.I0(CLBLL_L_X4Y143_SLICE_X5Y143_AQ),
.I1(CLBLM_R_X7Y142_SLICE_X8Y142_DO6),
.I2(CLBLM_R_X7Y147_SLICE_X9Y147_AQ),
.I3(CLBLL_L_X2Y148_SLICE_X0Y148_A5Q),
.I4(CLBLL_L_X4Y148_SLICE_X5Y148_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y148_SLICE_X4Y148_BO5),
.O6(CLBLL_L_X4Y148_SLICE_X4Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888cc00cc00)
  ) CLBLL_L_X4Y148_SLICE_X4Y148_ALUT (
.I0(CLBLM_R_X5Y149_SLICE_X6Y149_DQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(1'b1),
.I3(CLBLM_R_X3Y149_SLICE_X3Y149_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y148_SLICE_X4Y148_AO5),
.O6(CLBLL_L_X4Y148_SLICE_X4Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y148_SLICE_X5Y148_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y148_SLICE_X5Y148_BO5),
.Q(CLBLL_L_X4Y148_SLICE_X5Y148_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y148_SLICE_X5Y148_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y148_SLICE_X5Y148_AO6),
.Q(CLBLL_L_X4Y148_SLICE_X5Y148_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y148_SLICE_X5Y148_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y148_SLICE_X5Y148_BO6),
.Q(CLBLL_L_X4Y148_SLICE_X5Y148_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y148_SLICE_X5Y148_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y148_SLICE_X5Y148_CO6),
.Q(CLBLL_L_X4Y148_SLICE_X5Y148_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y148_SLICE_X5Y148_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y148_SLICE_X5Y148_DO6),
.Q(CLBLL_L_X4Y148_SLICE_X5Y148_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5f5f5f5a0f5f5)
  ) CLBLL_L_X4Y148_SLICE_X5Y148_DLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(1'b1),
.I2(CLBLM_R_X5Y149_SLICE_X6Y149_D5Q),
.I3(CLBLM_R_X3Y143_SLICE_X2Y143_AQ),
.I4(CLBLM_R_X3Y145_SLICE_X2Y145_DQ),
.I5(CLBLM_L_X10Y147_SLICE_X13Y147_A5Q),
.O5(CLBLL_L_X4Y148_SLICE_X5Y148_DO5),
.O6(CLBLL_L_X4Y148_SLICE_X5Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888888d88dd)
  ) CLBLL_L_X4Y148_SLICE_X5Y148_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X7Y152_SLICE_X9Y152_C5Q),
.I2(CLBLL_L_X4Y146_SLICE_X4Y146_BQ),
.I3(CLBLM_R_X3Y144_SLICE_X3Y144_D5Q),
.I4(CLBLL_L_X4Y148_SLICE_X5Y148_CQ),
.I5(CLBLL_L_X2Y148_SLICE_X0Y148_BQ),
.O5(CLBLL_L_X4Y148_SLICE_X5Y148_CO5),
.O6(CLBLL_L_X4Y148_SLICE_X5Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffcc00aaf0aaf0)
  ) CLBLL_L_X4Y148_SLICE_X5Y148_BLUT (
.I0(CLBLM_R_X7Y145_SLICE_X8Y145_AQ),
.I1(CLBLM_R_X5Y145_SLICE_X6Y145_BQ),
.I2(CLBLM_R_X5Y144_SLICE_X6Y144_C5Q),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLL_L_X4Y148_SLICE_X4Y148_DO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y148_SLICE_X5Y148_BO5),
.O6(CLBLL_L_X4Y148_SLICE_X5Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccf0ccaaccf0cc55)
  ) CLBLL_L_X4Y148_SLICE_X5Y148_ALUT (
.I0(CLBLL_L_X4Y148_SLICE_X5Y148_AQ),
.I1(CLBLM_L_X10Y149_SLICE_X12Y149_B5Q),
.I2(CLBLM_R_X5Y147_SLICE_X6Y147_B5Q),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X8Y149_SLICE_X11Y149_BQ),
.I5(CLBLL_L_X4Y148_SLICE_X4Y148_BO5),
.O5(CLBLL_L_X4Y148_SLICE_X5Y148_AO5),
.O6(CLBLL_L_X4Y148_SLICE_X5Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y149_SLICE_X4Y149_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y149_SLICE_X4Y149_BO5),
.Q(CLBLL_L_X4Y149_SLICE_X4Y149_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y149_SLICE_X4Y149_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y149_SLICE_X4Y149_CO5),
.Q(CLBLL_L_X4Y149_SLICE_X4Y149_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y149_SLICE_X4Y149_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y149_SLICE_X4Y149_DO5),
.Q(CLBLL_L_X4Y149_SLICE_X4Y149_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y149_SLICE_X4Y149_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y149_SLICE_X4Y149_AO6),
.Q(CLBLL_L_X4Y149_SLICE_X4Y149_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y149_SLICE_X4Y149_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y149_SLICE_X4Y149_BO6),
.Q(CLBLL_L_X4Y149_SLICE_X4Y149_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y149_SLICE_X4Y149_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y149_SLICE_X4Y149_CO6),
.Q(CLBLL_L_X4Y149_SLICE_X4Y149_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y149_SLICE_X4Y149_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y149_SLICE_X4Y149_DO6),
.Q(CLBLL_L_X4Y149_SLICE_X4Y149_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hdddd8888a0f5f5a0)
  ) CLBLL_L_X4Y149_SLICE_X4Y149_DLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLL_L_X2Y148_SLICE_X1Y148_AQ),
.I2(CLBLM_R_X3Y148_SLICE_X2Y148_D5Q),
.I3(CLBLM_R_X5Y148_SLICE_X6Y148_CO6),
.I4(CLBLL_L_X4Y149_SLICE_X4Y149_D5Q),
.I5(1'b1),
.O5(CLBLL_L_X4Y149_SLICE_X4Y149_DO5),
.O6(CLBLL_L_X4Y149_SLICE_X4Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'he4e4e4e4fa50fa50)
  ) CLBLL_L_X4Y149_SLICE_X4Y149_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X5Y148_SLICE_X7Y148_AQ),
.I2(CLBLL_L_X4Y149_SLICE_X4Y149_DQ),
.I3(CLBLM_L_X10Y150_SLICE_X12Y150_CQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y149_SLICE_X4Y149_CO5),
.O6(CLBLL_L_X4Y149_SLICE_X4Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffcc00aa3caa3c)
  ) CLBLL_L_X4Y149_SLICE_X4Y149_BLUT (
.I0(CLBLL_L_X4Y147_SLICE_X4Y147_C5Q),
.I1(CLBLL_L_X4Y151_SLICE_X4Y151_AQ),
.I2(CLBLM_R_X3Y151_SLICE_X3Y151_BQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X10Y150_SLICE_X13Y150_B5Q),
.I5(1'b1),
.O5(CLBLL_L_X4Y149_SLICE_X4Y149_BO5),
.O6(CLBLL_L_X4Y149_SLICE_X4Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaacc0fccf0)
  ) CLBLL_L_X4Y149_SLICE_X4Y149_ALUT (
.I0(CLBLM_R_X5Y151_SLICE_X6Y151_B5Q),
.I1(CLBLL_L_X4Y149_SLICE_X4Y149_BQ),
.I2(CLBLL_L_X4Y149_SLICE_X4Y149_AQ),
.I3(CLBLM_L_X8Y149_SLICE_X11Y149_BQ),
.I4(CLBLL_L_X4Y148_SLICE_X4Y148_BO6),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLL_L_X4Y149_SLICE_X4Y149_AO5),
.O6(CLBLL_L_X4Y149_SLICE_X4Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y149_SLICE_X5Y149_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y149_SLICE_X5Y149_AO6),
.Q(CLBLL_L_X4Y149_SLICE_X5Y149_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y149_SLICE_X5Y149_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y149_SLICE_X5Y149_BO6),
.Q(CLBLL_L_X4Y149_SLICE_X5Y149_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y149_SLICE_X5Y149_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y149_SLICE_X5Y149_CO6),
.Q(CLBLL_L_X4Y149_SLICE_X5Y149_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y149_SLICE_X5Y149_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y149_SLICE_X5Y149_DO6),
.Q(CLBLL_L_X4Y149_SLICE_X5Y149_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffcf8a0000cf8a)
  ) CLBLL_L_X4Y149_SLICE_X5Y149_DLUT (
.I0(CLBLL_L_X4Y146_SLICE_X5Y146_AQ),
.I1(CLBLM_L_X8Y142_SLICE_X11Y142_CQ),
.I2(CLBLM_R_X5Y149_SLICE_X7Y149_DQ),
.I3(CLBLL_L_X4Y149_SLICE_X5Y149_DQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X5Y152_SLICE_X6Y152_CQ),
.O5(CLBLL_L_X4Y149_SLICE_X5Y149_DO5),
.O6(CLBLL_L_X4Y149_SLICE_X5Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccaaf0ccccaaaa)
  ) CLBLL_L_X4Y149_SLICE_X5Y149_CLUT (
.I0(CLBLL_L_X4Y149_SLICE_X5Y149_BQ),
.I1(CLBLM_R_X5Y149_SLICE_X6Y149_A5Q),
.I2(CLBLM_L_X10Y147_SLICE_X13Y147_AQ),
.I3(CLBLM_R_X3Y143_SLICE_X2Y143_AQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X3Y145_SLICE_X2Y145_DQ),
.O5(CLBLL_L_X4Y149_SLICE_X5Y149_CO5),
.O6(CLBLL_L_X4Y149_SLICE_X5Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'heeee2222fece3202)
  ) CLBLL_L_X4Y149_SLICE_X5Y149_BLUT (
.I0(CLBLL_L_X4Y148_SLICE_X5Y148_DQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X3Y145_SLICE_X2Y145_DQ),
.I3(CLBLM_R_X7Y150_SLICE_X8Y150_C5Q),
.I4(CLBLL_L_X4Y146_SLICE_X4Y146_AQ),
.I5(CLBLM_R_X3Y143_SLICE_X2Y143_AQ),
.O5(CLBLL_L_X4Y149_SLICE_X5Y149_BO5),
.O6(CLBLL_L_X4Y149_SLICE_X5Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00e2e2ff00f0f0)
  ) CLBLL_L_X4Y149_SLICE_X5Y149_ALUT (
.I0(CLBLM_R_X5Y149_SLICE_X6Y149_DQ),
.I1(CLBLM_L_X8Y146_SLICE_X10Y146_AQ),
.I2(CLBLL_L_X4Y149_SLICE_X5Y149_AQ),
.I3(CLBLL_L_X4Y146_SLICE_X5Y146_AQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X7Y150_SLICE_X9Y150_CQ),
.O5(CLBLL_L_X4Y149_SLICE_X5Y149_AO5),
.O6(CLBLL_L_X4Y149_SLICE_X5Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y150_SLICE_X4Y150_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLL_L_X4Y151_SLICE_X5Y151_DQ),
.Q(CLBLL_L_X4Y150_SLICE_X4Y150_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLL_L_X4Y150_SLICE_X4Y150_DLUT (
.I0(CLBLL_L_X2Y150_SLICE_X1Y150_C5Q),
.I1(CLBLL_L_X4Y147_SLICE_X4Y147_C5Q),
.I2(CLBLM_R_X3Y144_SLICE_X3Y144_A5Q),
.I3(CLBLL_L_X2Y148_SLICE_X0Y148_AQ),
.I4(CLBLM_L_X8Y153_SLICE_X10Y153_AQ),
.I5(CLBLL_L_X2Y147_SLICE_X0Y147_BQ),
.O5(CLBLL_L_X4Y150_SLICE_X4Y150_DO5),
.O6(CLBLL_L_X4Y150_SLICE_X4Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000008000000)
  ) CLBLL_L_X4Y150_SLICE_X4Y150_CLUT (
.I0(CLBLM_R_X5Y153_SLICE_X6Y153_AQ),
.I1(CLBLL_L_X4Y153_SLICE_X5Y153_BQ),
.I2(CLBLM_R_X3Y151_SLICE_X3Y151_AQ),
.I3(CLBLL_L_X4Y150_SLICE_X5Y150_CQ),
.I4(CLBLM_R_X3Y151_SLICE_X3Y151_BQ),
.I5(CLBLM_R_X5Y151_SLICE_X7Y151_BO6),
.O5(CLBLL_L_X4Y150_SLICE_X4Y150_CO5),
.O6(CLBLL_L_X4Y150_SLICE_X4Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000cccc0000cc6c)
  ) CLBLL_L_X4Y150_SLICE_X4Y150_BLUT (
.I0(CLBLM_R_X7Y152_SLICE_X8Y152_BQ),
.I1(CLBLL_L_X4Y150_SLICE_X5Y150_CQ),
.I2(CLBLM_R_X7Y144_SLICE_X9Y144_AQ),
.I3(CLBLM_R_X5Y151_SLICE_X7Y151_BO6),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLL_L_X4Y150_SLICE_X4Y150_AO5),
.O5(CLBLL_L_X4Y150_SLICE_X4Y150_BO5),
.O6(CLBLL_L_X4Y150_SLICE_X4Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h800000003f3fffff)
  ) CLBLL_L_X4Y150_SLICE_X4Y150_ALUT (
.I0(CLBLM_R_X7Y152_SLICE_X8Y152_BQ),
.I1(CLBLM_R_X5Y144_SLICE_X7Y144_CQ),
.I2(CLBLM_R_X3Y144_SLICE_X3Y144_CQ),
.I3(CLBLM_R_X7Y144_SLICE_X9Y144_AQ),
.I4(CLBLM_R_X3Y152_SLICE_X3Y152_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y150_SLICE_X4Y150_AO5),
.O6(CLBLL_L_X4Y150_SLICE_X4Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y150_SLICE_X5Y150_C5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y150_SLICE_X5Y150_CO5),
.Q(CLBLL_L_X4Y150_SLICE_X5Y150_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y150_SLICE_X5Y150_D5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y150_SLICE_X5Y150_DO5),
.Q(CLBLL_L_X4Y150_SLICE_X5Y150_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y150_SLICE_X5Y150_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y150_SLICE_X5Y150_AO6),
.Q(CLBLL_L_X4Y150_SLICE_X5Y150_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y150_SLICE_X5Y150_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y150_SLICE_X5Y150_BO6),
.Q(CLBLL_L_X4Y150_SLICE_X5Y150_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y150_SLICE_X5Y150_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y150_SLICE_X5Y150_CO6),
.Q(CLBLL_L_X4Y150_SLICE_X5Y150_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y150_SLICE_X5Y150_D_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y150_SLICE_X5Y150_DO6),
.Q(CLBLL_L_X4Y150_SLICE_X5Y150_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0aaf0aaeecceecc)
  ) CLBLL_L_X4Y150_SLICE_X5Y150_DLUT (
.I0(CLBLM_R_X5Y150_SLICE_X6Y150_C5Q),
.I1(CLBLM_R_X3Y152_SLICE_X3Y152_BO6),
.I2(CLBLM_R_X5Y144_SLICE_X7Y144_DQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y150_SLICE_X5Y150_DO5),
.O6(CLBLL_L_X4Y150_SLICE_X5Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbfbf8f8ff33cc00)
  ) CLBLL_L_X4Y150_SLICE_X5Y150_CLUT (
.I0(CLBLM_R_X5Y143_SLICE_X6Y143_DQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLL_L_X4Y150_SLICE_X4Y150_BO6),
.I3(CLBLL_L_X4Y149_SLICE_X5Y149_BQ),
.I4(CLBLL_L_X2Y148_SLICE_X0Y148_B5Q),
.I5(1'b1),
.O5(CLBLL_L_X4Y150_SLICE_X5Y150_CO5),
.O6(CLBLL_L_X4Y150_SLICE_X5Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000f0ccf033)
  ) CLBLL_L_X4Y150_SLICE_X5Y150_BLUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y150_SLICE_X5Y150_BQ),
.I2(CLBLL_L_X4Y148_SLICE_X5Y148_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLL_L_X4Y151_SLICE_X4Y151_AO5),
.I5(CLBLM_R_X3Y146_SLICE_X3Y146_CQ),
.O5(CLBLL_L_X4Y150_SLICE_X5Y150_BO5),
.O6(CLBLL_L_X4Y150_SLICE_X5Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfc0cfc0cacacfc0)
  ) CLBLL_L_X4Y150_SLICE_X5Y150_ALUT (
.I0(CLBLL_L_X4Y150_SLICE_X5Y150_AQ),
.I1(CLBLM_R_X3Y149_SLICE_X2Y149_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLL_L_X4Y148_SLICE_X4Y148_BQ),
.I4(CLBLM_R_X5Y149_SLICE_X6Y149_D5Q),
.I5(CLBLM_L_X8Y150_SLICE_X11Y150_B5Q),
.O5(CLBLL_L_X4Y150_SLICE_X5Y150_AO5),
.O6(CLBLL_L_X4Y150_SLICE_X5Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y151_SLICE_X4Y151_A_FDSE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X2Y150_SLICE_X1Y150_BO6),
.Q(CLBLL_L_X4Y151_SLICE_X4Y151_AQ),
.S(CLBLL_L_X4Y151_SLICE_X4Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y151_SLICE_X4Y151_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y151_SLICE_X4Y151_DO5),
.O6(CLBLL_L_X4Y151_SLICE_X4Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000000f0f0f0f)
  ) CLBLL_L_X4Y151_SLICE_X4Y151_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X3Y148_SLICE_X2Y148_C5Q),
.I3(1'b1),
.I4(1'b1),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLL_L_X4Y151_SLICE_X4Y151_CO5),
.O6(CLBLL_L_X4Y151_SLICE_X4Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbffffff44440000)
  ) CLBLL_L_X4Y151_SLICE_X4Y151_BLUT (
.I0(CLBLM_R_X3Y152_SLICE_X2Y152_DO6),
.I1(CLBLM_R_X5Y153_SLICE_X6Y153_AQ),
.I2(1'b1),
.I3(CLBLM_R_X3Y151_SLICE_X3Y151_AQ),
.I4(CLBLL_L_X4Y153_SLICE_X5Y153_BQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y151_SLICE_X4Y151_BO5),
.O6(CLBLL_L_X4Y151_SLICE_X4Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5a0f5a03f3fffff)
  ) CLBLL_L_X4Y151_SLICE_X4Y151_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X7Y149_SLICE_X8Y149_AQ),
.I2(CLBLM_R_X7Y150_SLICE_X8Y150_AQ),
.I3(CLBLM_R_X5Y152_SLICE_X6Y152_CQ),
.I4(CLBLM_R_X7Y150_SLICE_X8Y150_CQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y151_SLICE_X4Y151_AO5),
.O6(CLBLL_L_X4Y151_SLICE_X4Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y151_SLICE_X5Y151_A5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y151_SLICE_X4Y151_AO6),
.Q(CLBLL_L_X4Y151_SLICE_X5Y151_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y151_SLICE_X5Y151_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y151_SLICE_X5Y151_AO6),
.Q(CLBLL_L_X4Y151_SLICE_X5Y151_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y151_SLICE_X5Y151_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y151_SLICE_X5Y151_BO6),
.Q(CLBLL_L_X4Y151_SLICE_X5Y151_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y151_SLICE_X5Y151_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y151_SLICE_X5Y151_CO6),
.Q(CLBLL_L_X4Y151_SLICE_X5Y151_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y151_SLICE_X5Y151_D_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y151_SLICE_X5Y151_DO6),
.Q(CLBLL_L_X4Y151_SLICE_X5Y151_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff8cdc00008cdc)
  ) CLBLL_L_X4Y151_SLICE_X5Y151_DLUT (
.I0(CLBLM_R_X3Y143_SLICE_X2Y143_AQ),
.I1(CLBLL_L_X4Y151_SLICE_X5Y151_CQ),
.I2(CLBLM_R_X3Y145_SLICE_X2Y145_DQ),
.I3(CLBLM_L_X8Y152_SLICE_X11Y152_A5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_L_X8Y152_SLICE_X10Y152_AQ),
.O5(CLBLL_L_X4Y151_SLICE_X5Y151_DO5),
.O6(CLBLL_L_X4Y151_SLICE_X5Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccff5f0050)
  ) CLBLL_L_X4Y151_SLICE_X5Y151_CLUT (
.I0(CLBLM_L_X10Y150_SLICE_X13Y150_AQ),
.I1(CLBLM_L_X8Y151_SLICE_X10Y151_AQ),
.I2(CLBLM_R_X3Y145_SLICE_X2Y145_DQ),
.I3(CLBLM_R_X3Y143_SLICE_X2Y143_AQ),
.I4(CLBLL_L_X4Y152_SLICE_X5Y152_DQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLL_L_X4Y151_SLICE_X5Y151_CO5),
.O6(CLBLL_L_X4Y151_SLICE_X5Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafafcfc0a0a0c0c)
  ) CLBLL_L_X4Y151_SLICE_X5Y151_BLUT (
.I0(CLBLL_L_X4Y152_SLICE_X5Y152_AQ),
.I1(CLBLL_L_X4Y151_SLICE_X5Y151_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(1'b1),
.I4(CLBLM_L_X10Y143_SLICE_X12Y143_BO5),
.I5(CLBLM_L_X8Y152_SLICE_X11Y152_A5Q),
.O5(CLBLL_L_X4Y151_SLICE_X5Y151_BO5),
.O6(CLBLL_L_X4Y151_SLICE_X5Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccafccfaccafccfa)
  ) CLBLL_L_X4Y151_SLICE_X5Y151_ALUT (
.I0(CLBLL_L_X2Y148_SLICE_X0Y148_B5Q),
.I1(CLBLM_R_X5Y149_SLICE_X7Y149_B5Q),
.I2(CLBLL_L_X4Y151_SLICE_X5Y151_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLL_L_X4Y150_SLICE_X4Y150_AO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y151_SLICE_X5Y151_AO5),
.O6(CLBLL_L_X4Y151_SLICE_X5Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y152_SLICE_X4Y152_C5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y152_SLICE_X4Y152_CO5),
.Q(CLBLL_L_X4Y152_SLICE_X4Y152_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y152_SLICE_X4Y152_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y152_SLICE_X4Y152_AO6),
.Q(CLBLL_L_X4Y152_SLICE_X4Y152_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y152_SLICE_X4Y152_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y152_SLICE_X4Y152_BO6),
.Q(CLBLL_L_X4Y152_SLICE_X4Y152_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y152_SLICE_X4Y152_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y152_SLICE_X4Y152_CO6),
.Q(CLBLL_L_X4Y152_SLICE_X4Y152_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y152_SLICE_X4Y152_D_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y152_SLICE_X4Y152_DO6),
.Q(CLBLL_L_X4Y152_SLICE_X4Y152_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdccffce31003302)
  ) CLBLL_L_X4Y152_SLICE_X4Y152_DLUT (
.I0(CLBLM_R_X3Y145_SLICE_X2Y145_DQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X3Y143_SLICE_X2Y143_AQ),
.I3(CLBLM_R_X3Y151_SLICE_X2Y151_BQ),
.I4(CLBLM_L_X8Y152_SLICE_X11Y152_AQ),
.I5(CLBLM_R_X5Y154_SLICE_X7Y154_BQ),
.O5(CLBLL_L_X4Y152_SLICE_X4Y152_DO5),
.O6(CLBLL_L_X4Y152_SLICE_X4Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'heeee22228bbb8bbb)
  ) CLBLL_L_X4Y152_SLICE_X4Y152_CLUT (
.I0(CLBLM_R_X5Y151_SLICE_X6Y151_D5Q),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLL_L_X4Y152_SLICE_X4Y152_BQ),
.I3(CLBLL_L_X4Y150_SLICE_X4Y150_CO6),
.I4(CLBLM_R_X3Y153_SLICE_X3Y153_BQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y152_SLICE_X4Y152_CO5),
.O6(CLBLL_L_X4Y152_SLICE_X4Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000aabb0011)
  ) CLBLL_L_X4Y152_SLICE_X4Y152_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X7Y144_SLICE_X9Y144_AQ),
.I2(1'b1),
.I3(CLBLM_R_X7Y152_SLICE_X8Y152_BQ),
.I4(CLBLM_R_X5Y151_SLICE_X7Y151_A5Q),
.I5(CLBLL_L_X4Y150_SLICE_X4Y150_AO5),
.O5(CLBLL_L_X4Y152_SLICE_X4Y152_BO5),
.O6(CLBLL_L_X4Y152_SLICE_X4Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffa5a5a5ff000000)
  ) CLBLL_L_X4Y152_SLICE_X4Y152_ALUT (
.I0(CLBLL_L_X4Y153_SLICE_X4Y153_DO6),
.I1(1'b1),
.I2(CLBLL_L_X4Y152_SLICE_X4Y152_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLL_L_X4Y145_SLICE_X4Y145_AQ),
.I5(CLBLM_R_X5Y153_SLICE_X7Y153_BO6),
.O5(CLBLL_L_X4Y152_SLICE_X4Y152_AO5),
.O6(CLBLL_L_X4Y152_SLICE_X4Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y152_SLICE_X5Y152_B5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y152_SLICE_X5Y152_BO5),
.Q(CLBLL_L_X4Y152_SLICE_X5Y152_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y152_SLICE_X5Y152_C5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y152_SLICE_X5Y152_CO5),
.Q(CLBLL_L_X4Y152_SLICE_X5Y152_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y152_SLICE_X5Y152_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y152_SLICE_X5Y152_AO6),
.Q(CLBLL_L_X4Y152_SLICE_X5Y152_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y152_SLICE_X5Y152_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y152_SLICE_X5Y152_BO6),
.Q(CLBLL_L_X4Y152_SLICE_X5Y152_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y152_SLICE_X5Y152_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y152_SLICE_X5Y152_CO6),
.Q(CLBLL_L_X4Y152_SLICE_X5Y152_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y152_SLICE_X5Y152_D_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y152_SLICE_X5Y152_DO6),
.Q(CLBLL_L_X4Y152_SLICE_X5Y152_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff7f0f20f070002)
  ) CLBLL_L_X4Y152_SLICE_X5Y152_DLUT (
.I0(CLBLM_R_X3Y145_SLICE_X2Y145_DQ),
.I1(CLBLM_L_X10Y150_SLICE_X13Y150_A5Q),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X3Y143_SLICE_X2Y143_AQ),
.I4(CLBLL_L_X4Y152_SLICE_X4Y152_DQ),
.I5(CLBLL_L_X4Y152_SLICE_X5Y152_AQ),
.O5(CLBLL_L_X4Y152_SLICE_X5Y152_DO5),
.O6(CLBLL_L_X4Y152_SLICE_X5Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf303f303f3f30303)
  ) CLBLL_L_X4Y152_SLICE_X5Y152_CLUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y152_SLICE_X4Y152_C5Q),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X5Y141_SLICE_X6Y141_AQ),
.I4(CLBLM_L_X8Y150_SLICE_X11Y150_CQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y152_SLICE_X5Y152_CO5),
.O6(CLBLL_L_X4Y152_SLICE_X5Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5a0f5a0eeee4444)
  ) CLBLL_L_X4Y152_SLICE_X5Y152_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLL_L_X4Y150_SLICE_X4Y150_DO6),
.I2(CLBLM_R_X5Y152_SLICE_X6Y152_B5Q),
.I3(CLBLL_L_X4Y152_SLICE_X4Y152_C5Q),
.I4(CLBLL_L_X4Y152_SLICE_X5Y152_DQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y152_SLICE_X5Y152_BO5),
.O6(CLBLL_L_X4Y152_SLICE_X5Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hddd88888ddd8ddd8)
  ) CLBLL_L_X4Y152_SLICE_X5Y152_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLL_L_X4Y152_SLICE_X5Y152_BQ),
.I2(CLBLL_L_X4Y152_SLICE_X5Y152_AQ),
.I3(CLBLL_L_X4Y146_SLICE_X5Y146_BQ),
.I4(CLBLM_R_X5Y144_SLICE_X6Y144_CQ),
.I5(CLBLM_R_X3Y147_SLICE_X3Y147_BQ),
.O5(CLBLL_L_X4Y152_SLICE_X5Y152_AO5),
.O6(CLBLL_L_X4Y152_SLICE_X5Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y153_SLICE_X4Y153_A5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y154_SLICE_X4Y154_BO5),
.Q(CLBLL_L_X4Y153_SLICE_X4Y153_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y153_SLICE_X4Y153_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y153_SLICE_X4Y153_AO6),
.Q(CLBLL_L_X4Y153_SLICE_X4Y153_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y153_SLICE_X4Y153_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y153_SLICE_X4Y153_BO6),
.Q(CLBLL_L_X4Y153_SLICE_X4Y153_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y153_SLICE_X4Y153_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y153_SLICE_X4Y153_CO6),
.Q(CLBLL_L_X4Y153_SLICE_X4Y153_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fff7fff3fff3fff)
  ) CLBLL_L_X4Y153_SLICE_X4Y153_DLUT (
.I0(CLBLL_L_X4Y153_SLICE_X4Y153_BQ),
.I1(CLBLL_L_X4Y153_SLICE_X4Y153_CQ),
.I2(CLBLL_L_X4Y153_SLICE_X4Y153_AQ),
.I3(CLBLM_R_X3Y153_SLICE_X3Y153_DO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y153_SLICE_X4Y153_DO5),
.O6(CLBLL_L_X4Y153_SLICE_X4Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hb3a0b3a0eca0eca0)
  ) CLBLL_L_X4Y153_SLICE_X4Y153_CLUT (
.I0(CLBLM_R_X11Y149_SLICE_X15Y149_CQ),
.I1(CLBLL_L_X4Y153_SLICE_X4Y153_CQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X5Y153_SLICE_X7Y153_BO6),
.I4(1'b1),
.I5(CLBLM_R_X3Y153_SLICE_X3Y153_DO6),
.O5(CLBLL_L_X4Y153_SLICE_X4Y153_CO5),
.O6(CLBLL_L_X4Y153_SLICE_X4Y153_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hecb3ecb3a0a0a0a0)
  ) CLBLL_L_X4Y153_SLICE_X4Y153_BLUT (
.I0(CLBLL_L_X4Y149_SLICE_X5Y149_DQ),
.I1(CLBLL_L_X4Y153_SLICE_X4Y153_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLL_L_X4Y153_SLICE_X4Y153_DO5),
.I4(1'b1),
.I5(CLBLM_R_X5Y153_SLICE_X7Y153_BO6),
.O5(CLBLL_L_X4Y153_SLICE_X4Y153_BO5),
.O6(CLBLL_L_X4Y153_SLICE_X4Y153_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hde5acc00fcf0cc00)
  ) CLBLL_L_X4Y153_SLICE_X4Y153_ALUT (
.I0(CLBLL_L_X4Y153_SLICE_X4Y153_CQ),
.I1(CLBLM_R_X5Y154_SLICE_X6Y154_AQ),
.I2(CLBLL_L_X4Y153_SLICE_X4Y153_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X5Y153_SLICE_X7Y153_BO6),
.I5(CLBLM_R_X3Y153_SLICE_X3Y153_DO6),
.O5(CLBLL_L_X4Y153_SLICE_X4Y153_AO5),
.O6(CLBLL_L_X4Y153_SLICE_X4Y153_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y153_SLICE_X5Y153_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y153_SLICE_X5Y153_AO6),
.Q(CLBLL_L_X4Y153_SLICE_X5Y153_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y153_SLICE_X5Y153_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y153_SLICE_X5Y153_BO6),
.Q(CLBLL_L_X4Y153_SLICE_X5Y153_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffdcffffffffffff)
  ) CLBLL_L_X4Y153_SLICE_X5Y153_DLUT (
.I0(CLBLL_L_X4Y152_SLICE_X4Y152_AQ),
.I1(CLBLM_R_X7Y153_SLICE_X8Y153_CO6),
.I2(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.I3(CLBLM_R_X3Y148_SLICE_X3Y148_BO6),
.I4(CLBLM_R_X3Y149_SLICE_X3Y149_AQ),
.I5(CLBLL_L_X4Y153_SLICE_X4Y153_BQ),
.O5(CLBLL_L_X4Y153_SLICE_X5Y153_DO5),
.O6(CLBLL_L_X4Y153_SLICE_X5Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff75ff7fff)
  ) CLBLL_L_X4Y153_SLICE_X5Y153_CLUT (
.I0(CLBLL_L_X4Y153_SLICE_X4Y153_AQ),
.I1(CLBLM_R_X3Y153_SLICE_X3Y153_BQ),
.I2(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.I3(CLBLL_L_X4Y153_SLICE_X4Y153_CQ),
.I4(CLBLL_L_X4Y150_SLICE_X5Y150_D5Q),
.I5(CLBLL_L_X4Y153_SLICE_X5Y153_DO6),
.O5(CLBLL_L_X4Y153_SLICE_X5Y153_CO5),
.O6(CLBLL_L_X4Y153_SLICE_X5Y153_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffeeffbe00ee00be)
  ) CLBLL_L_X4Y153_SLICE_X5Y153_BLUT (
.I0(CLBLL_L_X2Y148_SLICE_X0Y148_B5Q),
.I1(CLBLL_L_X4Y153_SLICE_X5Y153_BQ),
.I2(CLBLM_R_X5Y153_SLICE_X6Y153_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X3Y152_SLICE_X2Y152_DO6),
.I5(CLBLM_L_X10Y152_SLICE_X13Y152_BQ),
.O5(CLBLL_L_X4Y153_SLICE_X5Y153_BO5),
.O6(CLBLL_L_X4Y153_SLICE_X5Y153_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa3faa0caa0caa3f)
  ) CLBLL_L_X4Y153_SLICE_X5Y153_ALUT (
.I0(CLBLM_R_X5Y149_SLICE_X6Y149_CQ),
.I1(CLBLM_R_X7Y153_SLICE_X8Y153_CO6),
.I2(CLBLM_R_X7Y144_SLICE_X9Y144_B5Q),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLL_L_X4Y153_SLICE_X5Y153_AQ),
.I5(CLBLL_L_X4Y153_SLICE_X5Y153_CO6),
.O5(CLBLL_L_X4Y153_SLICE_X5Y153_AO5),
.O6(CLBLL_L_X4Y153_SLICE_X5Y153_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y154_SLICE_X4Y154_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y154_SLICE_X4Y154_AO6),
.Q(CLBLL_L_X4Y154_SLICE_X4Y154_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y154_SLICE_X4Y154_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y154_SLICE_X4Y154_DO5),
.O6(CLBLL_L_X4Y154_SLICE_X4Y154_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y154_SLICE_X4Y154_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y154_SLICE_X4Y154_CO5),
.O6(CLBLL_L_X4Y154_SLICE_X4Y154_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff55ffc0c0e2c0)
  ) CLBLL_L_X4Y154_SLICE_X4Y154_BLUT (
.I0(CLBLM_R_X3Y153_SLICE_X3Y153_A5Q),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLL_L_X4Y153_SLICE_X4Y153_CQ),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(CLBLM_R_X3Y150_SLICE_X2Y150_CO5),
.I5(1'b1),
.O5(CLBLL_L_X4Y154_SLICE_X4Y154_BO5),
.O6(CLBLL_L_X4Y154_SLICE_X4Y154_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8d88888800ff00ff)
  ) CLBLL_L_X4Y154_SLICE_X4Y154_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLL_L_X4Y149_SLICE_X5Y149_AQ),
.I2(CLBLL_L_X4Y154_SLICE_X4Y154_AQ),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(CLBLM_R_X3Y151_SLICE_X3Y151_C5Q),
.I5(1'b1),
.O5(CLBLL_L_X4Y154_SLICE_X4Y154_AO5),
.O6(CLBLL_L_X4Y154_SLICE_X4Y154_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y154_SLICE_X5Y154_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y154_SLICE_X5Y154_DO5),
.O6(CLBLL_L_X4Y154_SLICE_X5Y154_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y154_SLICE_X5Y154_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y154_SLICE_X5Y154_CO5),
.O6(CLBLL_L_X4Y154_SLICE_X5Y154_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y154_SLICE_X5Y154_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y154_SLICE_X5Y154_BO5),
.O6(CLBLL_L_X4Y154_SLICE_X5Y154_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00ffffffffff)
  ) CLBLL_L_X4Y154_SLICE_X5Y154_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X5Y153_SLICE_X6Y153_BQ),
.I4(1'b1),
.I5(CLBLL_L_X4Y148_SLICE_X5Y148_CQ),
.O5(CLBLL_L_X4Y154_SLICE_X5Y154_AO5),
.O6(CLBLL_L_X4Y154_SLICE_X5Y154_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y140_SLICE_X10Y140_A5_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y140_SLICE_X10Y140_AO5),
.Q(CLBLM_L_X8Y140_SLICE_X10Y140_A5Q),
.S(CLBLM_R_X11Y148_SLICE_X15Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y140_SLICE_X10Y140_A_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y140_SLICE_X10Y140_AO6),
.Q(CLBLM_L_X8Y140_SLICE_X10Y140_AQ),
.S(CLBLM_R_X11Y148_SLICE_X15Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y140_SLICE_X10Y140_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y140_SLICE_X10Y140_DO5),
.O6(CLBLM_L_X8Y140_SLICE_X10Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y140_SLICE_X10Y140_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y140_SLICE_X10Y140_CO5),
.O6(CLBLM_L_X8Y140_SLICE_X10Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y140_SLICE_X10Y140_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y140_SLICE_X10Y140_BO5),
.O6(CLBLM_L_X8Y140_SLICE_X10Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0cc00cc00)
  ) CLBLM_L_X8Y140_SLICE_X10Y140_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X5Y142_SLICE_X6Y142_DQ),
.I3(CLBLM_R_X7Y144_SLICE_X9Y144_A5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y140_SLICE_X10Y140_AO5),
.O6(CLBLM_L_X8Y140_SLICE_X10Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y140_SLICE_X11Y140_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y140_SLICE_X11Y140_DO5),
.O6(CLBLM_L_X8Y140_SLICE_X11Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y140_SLICE_X11Y140_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y140_SLICE_X11Y140_CO5),
.O6(CLBLM_L_X8Y140_SLICE_X11Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y140_SLICE_X11Y140_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y140_SLICE_X11Y140_BO5),
.O6(CLBLM_L_X8Y140_SLICE_X11Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y140_SLICE_X11Y140_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y140_SLICE_X11Y140_AO5),
.O6(CLBLM_L_X8Y140_SLICE_X11Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y141_SLICE_X10Y141_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y141_SLICE_X10Y141_AO6),
.Q(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y141_SLICE_X10Y141_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y141_SLICE_X10Y141_BO6),
.Q(CLBLM_L_X8Y141_SLICE_X10Y141_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y141_SLICE_X10Y141_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y141_SLICE_X10Y141_CO6),
.Q(CLBLM_L_X8Y141_SLICE_X10Y141_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000aaaaaaaa)
  ) CLBLM_L_X8Y141_SLICE_X10Y141_DLUT (
.I0(CLBLM_R_X7Y143_SLICE_X9Y143_BQ),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_L_X8Y141_SLICE_X10Y141_DO5),
.O6(CLBLM_L_X8Y141_SLICE_X10Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0ffcc0000)
  ) CLBLM_L_X8Y141_SLICE_X10Y141_CLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y141_SLICE_X10Y141_CQ),
.I2(CLBLM_L_X10Y142_SLICE_X12Y142_AQ),
.I3(CLBLM_L_X8Y143_SLICE_X10Y143_BQ),
.I4(CLBLM_L_X10Y143_SLICE_X12Y143_AO6),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_L_X8Y141_SLICE_X10Y141_CO5),
.O6(CLBLM_L_X8Y141_SLICE_X10Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffcff0c00fc000c)
  ) CLBLM_L_X8Y141_SLICE_X10Y141_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y141_SLICE_X10Y141_BQ),
.I2(CLBLM_L_X10Y143_SLICE_X12Y143_AO6),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X3Y142_SLICE_X2Y142_AQ),
.I5(CLBLM_L_X8Y144_SLICE_X11Y144_A5Q),
.O5(CLBLM_L_X8Y141_SLICE_X10Y141_BO5),
.O6(CLBLM_L_X8Y141_SLICE_X10Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa003c003c)
  ) CLBLM_L_X8Y141_SLICE_X10Y141_ALUT (
.I0(CLBLM_L_X8Y142_SLICE_X10Y142_A5Q),
.I1(CLBLM_L_X8Y142_SLICE_X11Y142_BQ),
.I2(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(1'b1),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_L_X8Y141_SLICE_X10Y141_AO5),
.O6(CLBLM_L_X8Y141_SLICE_X10Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y141_SLICE_X11Y141_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y141_SLICE_X11Y141_DO5),
.O6(CLBLM_L_X8Y141_SLICE_X11Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y141_SLICE_X11Y141_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y141_SLICE_X11Y141_CO5),
.O6(CLBLM_L_X8Y141_SLICE_X11Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y141_SLICE_X11Y141_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y141_SLICE_X11Y141_BO5),
.O6(CLBLM_L_X8Y141_SLICE_X11Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y141_SLICE_X11Y141_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y141_SLICE_X11Y141_AO5),
.O6(CLBLM_L_X8Y141_SLICE_X11Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y142_SLICE_X10Y142_A5_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y142_SLICE_X7Y142_AO6),
.Q(CLBLM_L_X8Y142_SLICE_X10Y142_A5Q),
.S(CLBLM_L_X8Y141_SLICE_X10Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y142_SLICE_X10Y142_C5_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y142_SLICE_X10Y142_CO5),
.Q(CLBLM_L_X8Y142_SLICE_X10Y142_C5Q),
.S(CLBLM_L_X8Y141_SLICE_X10Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y142_SLICE_X10Y142_A_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y142_SLICE_X10Y142_AO6),
.Q(CLBLM_L_X8Y142_SLICE_X10Y142_AQ),
.S(CLBLM_L_X8Y141_SLICE_X10Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y142_SLICE_X10Y142_C_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y142_SLICE_X10Y142_CO6),
.Q(CLBLM_L_X8Y142_SLICE_X10Y142_CQ),
.S(CLBLM_L_X8Y141_SLICE_X10Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h80008000f0f00000)
  ) CLBLM_L_X8Y142_SLICE_X10Y142_DLUT (
.I0(CLBLM_L_X10Y149_SLICE_X12Y149_A5Q),
.I1(CLBLM_R_X11Y146_SLICE_X15Y146_AQ),
.I2(CLBLM_R_X5Y146_SLICE_X7Y146_AQ),
.I3(CLBLM_R_X7Y142_SLICE_X9Y142_AQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y142_SLICE_X10Y142_DO5),
.O6(CLBLM_L_X8Y142_SLICE_X10Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000aa00aa00)
  ) CLBLM_L_X8Y142_SLICE_X10Y142_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_L_X8Y148_SLICE_X11Y148_BQ),
.I4(CLBLM_R_X3Y142_SLICE_X2Y142_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y142_SLICE_X10Y142_CO5),
.O6(CLBLM_L_X8Y142_SLICE_X10Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaff007f7f7f7f)
  ) CLBLM_L_X8Y142_SLICE_X10Y142_BLUT (
.I0(CLBLM_L_X8Y150_SLICE_X10Y150_A5Q),
.I1(CLBLM_L_X8Y142_SLICE_X11Y142_DO6),
.I2(CLBLM_R_X11Y149_SLICE_X14Y149_AQ),
.I3(CLBLM_R_X3Y146_SLICE_X2Y146_BQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y142_SLICE_X10Y142_BO5),
.O6(CLBLM_L_X8Y142_SLICE_X10Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00000f0f00000)
  ) CLBLM_L_X8Y142_SLICE_X10Y142_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.I3(1'b1),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y142_SLICE_X10Y142_AO5),
.O6(CLBLM_L_X8Y142_SLICE_X10Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y142_SLICE_X11Y142_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y142_SLICE_X11Y142_CO5),
.Q(CLBLM_L_X8Y142_SLICE_X11Y142_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y142_SLICE_X11Y142_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y142_SLICE_X11Y142_AO6),
.Q(CLBLM_L_X8Y142_SLICE_X11Y142_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y142_SLICE_X11Y142_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y142_SLICE_X11Y142_BO6),
.Q(CLBLM_L_X8Y142_SLICE_X11Y142_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y142_SLICE_X11Y142_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y142_SLICE_X11Y142_CO6),
.Q(CLBLM_L_X8Y142_SLICE_X11Y142_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000004)
  ) CLBLM_L_X8Y142_SLICE_X11Y142_DLUT (
.I0(CLBLM_L_X8Y144_SLICE_X11Y144_A5Q),
.I1(CLBLM_R_X7Y146_SLICE_X9Y146_B5Q),
.I2(CLBLM_L_X8Y144_SLICE_X10Y144_B5Q),
.I3(CLBLM_R_X11Y146_SLICE_X14Y146_AQ),
.I4(CLBLM_R_X7Y144_SLICE_X8Y144_AQ),
.I5(CLBLM_R_X5Y142_SLICE_X7Y142_C5Q),
.O5(CLBLM_L_X8Y142_SLICE_X11Y142_DO5),
.O6(CLBLM_L_X8Y142_SLICE_X11Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0aaaaccccaaaa)
  ) CLBLM_L_X8Y142_SLICE_X11Y142_CLUT (
.I0(RIOB33_X105Y109_IOB_X1Y110_I),
.I1(CLBLL_L_X4Y142_SLICE_X4Y142_A5Q),
.I2(CLBLM_R_X5Y146_SLICE_X7Y146_DQ),
.I3(1'b1),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y142_SLICE_X11Y142_CO5),
.O6(CLBLM_L_X8Y142_SLICE_X11Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff11ff0100110001)
  ) CLBLM_L_X8Y142_SLICE_X11Y142_BLUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(CLBLM_L_X8Y142_SLICE_X11Y142_BQ),
.I2(CLBLM_L_X8Y142_SLICE_X11Y142_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.I5(CLBLL_L_X4Y142_SLICE_X4Y142_AQ),
.O5(CLBLM_L_X8Y142_SLICE_X11Y142_BO5),
.O6(CLBLM_L_X8Y142_SLICE_X11Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00aa3caaf0)
  ) CLBLM_L_X8Y142_SLICE_X11Y142_ALUT (
.I0(CLBLM_L_X8Y152_SLICE_X11Y152_B5Q),
.I1(CLBLM_L_X8Y142_SLICE_X11Y142_BQ),
.I2(CLBLM_L_X8Y142_SLICE_X11Y142_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.I5(RIOB33_X105Y131_IOB_X1Y131_I),
.O5(CLBLM_L_X8Y142_SLICE_X11Y142_AO5),
.O6(CLBLM_L_X8Y142_SLICE_X11Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y143_SLICE_X10Y143_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y143_SLICE_X10Y143_AO6),
.Q(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y143_SLICE_X10Y143_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y143_SLICE_X10Y143_BO6),
.Q(CLBLM_L_X8Y143_SLICE_X10Y143_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y143_SLICE_X10Y143_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y143_SLICE_X10Y143_CO6),
.Q(CLBLM_L_X8Y143_SLICE_X10Y143_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y143_SLICE_X10Y143_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y143_SLICE_X10Y143_DO6),
.Q(CLBLM_L_X8Y143_SLICE_X10Y143_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaa00aaf0aaf0)
  ) CLBLM_L_X8Y143_SLICE_X10Y143_DLUT (
.I0(CLBLM_L_X8Y146_SLICE_X11Y146_AQ),
.I1(1'b1),
.I2(CLBLM_L_X8Y143_SLICE_X10Y143_DQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X8Y143_SLICE_X11Y143_DQ),
.I5(CLBLM_R_X11Y145_SLICE_X15Y145_BO5),
.O5(CLBLM_L_X8Y143_SLICE_X10Y143_DO5),
.O6(CLBLM_L_X8Y143_SLICE_X10Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaacfccc0cc)
  ) CLBLM_L_X8Y143_SLICE_X10Y143_CLUT (
.I0(CLBLM_L_X8Y142_SLICE_X11Y142_C5Q),
.I1(CLBLM_L_X8Y143_SLICE_X10Y143_CQ),
.I2(CLBLM_L_X8Y146_SLICE_X10Y146_AQ),
.I3(CLBLM_R_X7Y150_SLICE_X9Y150_CQ),
.I4(CLBLM_R_X7Y145_SLICE_X8Y145_BQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_L_X8Y143_SLICE_X10Y143_CO5),
.O6(CLBLM_L_X8Y143_SLICE_X10Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0ccf0ccf0aaf0cc)
  ) CLBLM_L_X8Y143_SLICE_X10Y143_BLUT (
.I0(CLBLM_R_X7Y148_SLICE_X9Y148_B5Q),
.I1(CLBLM_L_X8Y143_SLICE_X10Y143_BQ),
.I2(CLBLM_R_X5Y144_SLICE_X6Y144_DQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X7Y150_SLICE_X9Y150_CQ),
.I5(CLBLM_L_X8Y146_SLICE_X10Y146_AQ),
.O5(CLBLM_L_X8Y143_SLICE_X10Y143_BO5),
.O6(CLBLM_L_X8Y143_SLICE_X10Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccfacc00ccfaccfa)
  ) CLBLM_L_X8Y143_SLICE_X10Y143_ALUT (
.I0(CLBLM_L_X8Y147_SLICE_X10Y147_BQ),
.I1(CLBLM_R_X7Y145_SLICE_X8Y145_BQ),
.I2(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X5Y144_SLICE_X6Y144_CQ),
.I5(CLBLM_R_X3Y147_SLICE_X3Y147_BQ),
.O5(CLBLM_L_X8Y143_SLICE_X10Y143_AO5),
.O6(CLBLM_L_X8Y143_SLICE_X10Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y143_SLICE_X11Y143_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y143_SLICE_X12Y143_CO5),
.Q(CLBLM_L_X8Y143_SLICE_X11Y143_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y143_SLICE_X11Y143_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y143_SLICE_X11Y143_AO6),
.Q(CLBLM_L_X8Y143_SLICE_X11Y143_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y143_SLICE_X11Y143_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y143_SLICE_X11Y143_BO6),
.Q(CLBLM_L_X8Y143_SLICE_X11Y143_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y143_SLICE_X11Y143_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y143_SLICE_X11Y143_CO6),
.Q(CLBLM_L_X8Y143_SLICE_X11Y143_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y143_SLICE_X11Y143_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y143_SLICE_X11Y143_DO6),
.Q(CLBLM_L_X8Y143_SLICE_X11Y143_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaccc0fff0)
  ) CLBLM_L_X8Y143_SLICE_X11Y143_DLUT (
.I0(CLBLM_L_X10Y150_SLICE_X12Y150_BQ),
.I1(CLBLM_L_X8Y142_SLICE_X11Y142_CQ),
.I2(CLBLM_L_X8Y143_SLICE_X11Y143_DQ),
.I3(CLBLM_L_X8Y142_SLICE_X10Y142_AQ),
.I4(CLBLM_R_X5Y149_SLICE_X7Y149_DQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_L_X8Y143_SLICE_X11Y143_DO5),
.O6(CLBLM_L_X8Y143_SLICE_X11Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdf0fef00d000e00)
  ) CLBLM_L_X8Y143_SLICE_X11Y143_CLUT (
.I0(CLBLM_L_X8Y142_SLICE_X11Y142_C5Q),
.I1(CLBLM_L_X8Y143_SLICE_X11Y143_CQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_L_X8Y143_SLICE_X11Y143_A5Q),
.I4(RIOB33_X105Y109_IOB_X1Y110_I),
.I5(CLBLM_R_X7Y146_SLICE_X8Y146_BQ),
.O5(CLBLM_L_X8Y143_SLICE_X11Y143_CO5),
.O6(CLBLM_L_X8Y143_SLICE_X11Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffc540000fc54)
  ) CLBLM_L_X8Y143_SLICE_X11Y143_BLUT (
.I0(CLBLM_R_X5Y149_SLICE_X6Y149_D5Q),
.I1(CLBLM_L_X8Y143_SLICE_X11Y143_BQ),
.I2(CLBLM_L_X8Y145_SLICE_X11Y145_AQ),
.I3(CLBLM_L_X8Y150_SLICE_X11Y150_B5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_L_X8Y141_SLICE_X10Y141_CQ),
.O5(CLBLM_L_X8Y143_SLICE_X11Y143_BO5),
.O6(CLBLM_L_X8Y143_SLICE_X11Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heefa4450eefa4450)
  ) CLBLM_L_X8Y143_SLICE_X11Y143_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X8Y143_SLICE_X11Y143_BQ),
.I2(CLBLM_L_X8Y143_SLICE_X11Y143_AQ),
.I3(CLBLM_L_X10Y143_SLICE_X12Y143_AO6),
.I4(CLBLM_L_X8Y148_SLICE_X10Y148_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y143_SLICE_X11Y143_AO5),
.O6(CLBLM_L_X8Y143_SLICE_X11Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y144_SLICE_X10Y144_A5_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y144_SLICE_X10Y144_AO5),
.Q(CLBLM_L_X8Y144_SLICE_X10Y144_A5Q),
.S(CLBLM_R_X7Y148_SLICE_X9Y148_AO5)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y144_SLICE_X10Y144_B5_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y144_SLICE_X10Y144_BO5),
.Q(CLBLM_L_X8Y144_SLICE_X10Y144_B5Q),
.S(CLBLM_R_X7Y148_SLICE_X9Y148_AO5)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y144_SLICE_X10Y144_A_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y144_SLICE_X10Y144_AO6),
.Q(CLBLM_L_X8Y144_SLICE_X10Y144_AQ),
.S(CLBLM_R_X7Y148_SLICE_X9Y148_AO5)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y144_SLICE_X10Y144_B_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y144_SLICE_X10Y144_BO6),
.Q(CLBLM_L_X8Y144_SLICE_X10Y144_BQ),
.S(CLBLM_R_X7Y148_SLICE_X9Y148_AO5)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccffcceeeeffee)
  ) CLBLM_L_X8Y144_SLICE_X10Y144_DLUT (
.I0(CLBLM_R_X5Y148_SLICE_X6Y148_BQ),
.I1(CLBLM_L_X12Y149_SLICE_X16Y149_CO6),
.I2(1'b1),
.I3(CLBLM_R_X7Y143_SLICE_X8Y143_BQ),
.I4(CLBLM_L_X10Y143_SLICE_X12Y143_DO6),
.I5(CLBLM_R_X5Y145_SLICE_X7Y145_BO6),
.O5(CLBLM_L_X8Y144_SLICE_X10Y144_DO5),
.O6(CLBLM_L_X8Y144_SLICE_X10Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0c0408000)
  ) CLBLM_L_X8Y144_SLICE_X10Y144_CLUT (
.I0(CLBLM_R_X11Y149_SLICE_X14Y149_AQ),
.I1(CLBLM_L_X10Y144_SLICE_X13Y144_CO6),
.I2(CLBLM_L_X8Y150_SLICE_X10Y150_A5Q),
.I3(CLBLM_R_X5Y142_SLICE_X7Y142_CQ),
.I4(CLBLM_R_X7Y144_SLICE_X9Y144_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X8Y144_SLICE_X10Y144_CO5),
.O6(CLBLM_L_X8Y144_SLICE_X10Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc0088888888)
  ) CLBLM_L_X8Y144_SLICE_X10Y144_BLUT (
.I0(CLBLM_R_X5Y146_SLICE_X7Y146_B5Q),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(1'b1),
.I3(CLBLL_L_X4Y152_SLICE_X5Y152_C5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y144_SLICE_X10Y144_BO5),
.O6(CLBLM_L_X8Y144_SLICE_X10Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00ff000000)
  ) CLBLM_L_X8Y144_SLICE_X10Y144_ALUT (
.I0(CLBLM_R_X5Y154_SLICE_X7Y154_DQ),
.I1(1'b1),
.I2(1'b1),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLL_L_X4Y142_SLICE_X5Y142_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X8Y144_SLICE_X10Y144_AO5),
.O6(CLBLM_L_X8Y144_SLICE_X10Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y144_SLICE_X11Y144_A5_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y144_SLICE_X11Y144_AO5),
.Q(CLBLM_L_X8Y144_SLICE_X11Y144_A5Q),
.S(CLBLL_L_X4Y145_SLICE_X5Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y144_SLICE_X11Y144_A_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y144_SLICE_X11Y144_AO6),
.Q(CLBLM_L_X8Y144_SLICE_X11Y144_AQ),
.S(CLBLL_L_X4Y145_SLICE_X5Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff22ffffff22ff22)
  ) CLBLM_L_X8Y144_SLICE_X11Y144_DLUT (
.I0(CLBLM_L_X8Y144_SLICE_X10Y144_AQ),
.I1(CLBLM_L_X8Y145_SLICE_X10Y145_CO5),
.I2(1'b1),
.I3(CLBLM_L_X8Y145_SLICE_X11Y145_AO5),
.I4(CLBLM_L_X10Y143_SLICE_X12Y143_AO5),
.I5(CLBLM_L_X8Y143_SLICE_X11Y143_AQ),
.O5(CLBLM_L_X8Y144_SLICE_X11Y144_DO5),
.O6(CLBLM_L_X8Y144_SLICE_X11Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haeaeaeaeffaeffae)
  ) CLBLM_L_X8Y144_SLICE_X11Y144_CLUT (
.I0(CLBLM_L_X12Y149_SLICE_X16Y149_CO6),
.I1(CLBLM_R_X5Y144_SLICE_X7Y144_DQ),
.I2(CLBLM_L_X8Y142_SLICE_X10Y142_BO5),
.I3(CLBLM_R_X7Y144_SLICE_X9Y144_BQ),
.I4(1'b1),
.I5(CLBLM_R_X7Y148_SLICE_X8Y148_BO5),
.O5(CLBLM_L_X8Y144_SLICE_X11Y144_CO5),
.O6(CLBLM_L_X8Y144_SLICE_X11Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h33bb00aaf3fbf0fa)
  ) CLBLM_L_X8Y144_SLICE_X11Y144_BLUT (
.I0(CLBLM_R_X5Y148_SLICE_X6Y148_B5Q),
.I1(CLBLM_R_X7Y148_SLICE_X8Y148_BO5),
.I2(CLBLM_L_X8Y141_SLICE_X10Y141_BQ),
.I3(CLBLM_L_X10Y144_SLICE_X12Y144_AO6),
.I4(CLBLL_L_X4Y143_SLICE_X5Y143_CQ),
.I5(CLBLM_L_X10Y143_SLICE_X12Y143_DO5),
.O5(CLBLM_L_X8Y144_SLICE_X11Y144_BO5),
.O6(CLBLM_L_X8Y144_SLICE_X11Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000f000f000)
  ) CLBLM_L_X8Y144_SLICE_X11Y144_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_L_X8Y142_SLICE_X10Y142_C5Q),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X5Y147_SLICE_X7Y147_C5Q),
.I5(1'b1),
.O5(CLBLM_L_X8Y144_SLICE_X11Y144_AO5),
.O6(CLBLM_L_X8Y144_SLICE_X11Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y145_SLICE_X10Y145_A_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y146_SLICE_X9Y146_AO6),
.Q(CLBLM_L_X8Y145_SLICE_X10Y145_AQ),
.S(CLBLL_L_X4Y145_SLICE_X4Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y145_SLICE_X10Y145_B_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y145_SLICE_X10Y145_AO6),
.Q(CLBLM_L_X8Y145_SLICE_X10Y145_BQ),
.S(CLBLL_L_X4Y145_SLICE_X4Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hafffafafaaffaaaa)
  ) CLBLM_L_X8Y145_SLICE_X10Y145_DLUT (
.I0(CLBLM_L_X8Y144_SLICE_X10Y144_CO5),
.I1(1'b1),
.I2(CLBLM_L_X10Y143_SLICE_X12Y143_DO6),
.I3(CLBLM_L_X10Y143_SLICE_X12Y143_DO5),
.I4(CLBLM_R_X5Y145_SLICE_X6Y145_CQ),
.I5(CLBLM_R_X7Y145_SLICE_X8Y145_DQ),
.O5(CLBLM_L_X8Y145_SLICE_X10Y145_DO5),
.O6(CLBLM_L_X8Y145_SLICE_X10Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h22800080ff77ff77)
  ) CLBLM_L_X8Y145_SLICE_X10Y145_CLUT (
.I0(CLBLM_L_X10Y143_SLICE_X13Y143_AO6),
.I1(CLBLM_L_X8Y150_SLICE_X10Y150_A5Q),
.I2(CLBLM_R_X5Y146_SLICE_X6Y146_B5Q),
.I3(CLBLM_R_X11Y149_SLICE_X14Y149_AQ),
.I4(CLBLM_R_X7Y146_SLICE_X9Y146_BQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y145_SLICE_X10Y145_CO5),
.O6(CLBLM_L_X8Y145_SLICE_X10Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5faff5facc00cc00)
  ) CLBLM_L_X8Y145_SLICE_X10Y145_BLUT (
.I0(CLBLM_R_X7Y150_SLICE_X8Y150_AQ),
.I1(CLBLM_L_X10Y142_SLICE_X12Y142_CO6),
.I2(CLBLM_R_X3Y148_SLICE_X2Y148_AQ),
.I3(CLBLM_L_X8Y140_SLICE_X10Y140_AQ),
.I4(CLBLM_L_X8Y144_SLICE_X10Y144_BQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y145_SLICE_X10Y145_BO5),
.O6(CLBLM_L_X8Y145_SLICE_X10Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c05500ddcc)
  ) CLBLM_L_X8Y145_SLICE_X10Y145_ALUT (
.I0(CLBLM_L_X8Y142_SLICE_X10Y142_BO5),
.I1(CLBLM_L_X8Y144_SLICE_X11Y144_AQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X7Y145_SLICE_X9Y145_AQ),
.I4(CLBLM_L_X8Y145_SLICE_X10Y145_CO5),
.I5(1'b1),
.O5(CLBLM_L_X8Y145_SLICE_X10Y145_AO5),
.O6(CLBLM_L_X8Y145_SLICE_X10Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y145_SLICE_X11Y145_A_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y145_SLICE_X13Y145_AO6),
.Q(CLBLM_L_X8Y145_SLICE_X11Y145_AQ),
.S(CLBLM_R_X7Y144_SLICE_X8Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffeeffcccceeee)
  ) CLBLM_L_X8Y145_SLICE_X11Y145_DLUT (
.I0(CLBLL_L_X4Y145_SLICE_X5Y145_AQ),
.I1(CLBLM_L_X8Y144_SLICE_X10Y144_DO6),
.I2(1'b1),
.I3(CLBLM_L_X10Y143_SLICE_X12Y143_AO5),
.I4(CLBLM_L_X8Y148_SLICE_X10Y148_CO6),
.I5(CLBLM_L_X10Y149_SLICE_X12Y149_DQ),
.O5(CLBLM_L_X8Y145_SLICE_X11Y145_DO5),
.O6(CLBLM_L_X8Y145_SLICE_X11Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffdfc)
  ) CLBLM_L_X8Y145_SLICE_X11Y145_CLUT (
.I0(CLBLM_L_X10Y148_SLICE_X12Y148_BO5),
.I1(CLBLM_L_X8Y145_SLICE_X10Y145_AO5),
.I2(CLBLM_L_X10Y145_SLICE_X13Y145_DO6),
.I3(CLBLL_L_X4Y141_SLICE_X5Y141_A5Q),
.I4(CLBLM_L_X8Y145_SLICE_X11Y145_DO6),
.I5(CLBLM_L_X8Y144_SLICE_X11Y144_BO6),
.O5(CLBLM_L_X8Y145_SLICE_X11Y145_CO5),
.O6(CLBLM_L_X8Y145_SLICE_X11Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffff4f4fffffff4)
  ) CLBLM_L_X8Y145_SLICE_X11Y145_BLUT (
.I0(CLBLM_L_X10Y143_SLICE_X12Y143_AO5),
.I1(CLBLM_R_X7Y143_SLICE_X8Y143_CQ),
.I2(CLBLM_R_X5Y146_SLICE_X6Y146_CO6),
.I3(CLBLM_R_X7Y142_SLICE_X9Y142_CQ),
.I4(CLBLM_L_X8Y144_SLICE_X11Y144_CO6),
.I5(CLBLM_L_X10Y143_SLICE_X12Y143_DO6),
.O5(CLBLM_L_X8Y145_SLICE_X11Y145_BO5),
.O6(CLBLM_L_X8Y145_SLICE_X11Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000f0f04444ff44)
  ) CLBLM_L_X8Y145_SLICE_X11Y145_ALUT (
.I0(CLBLM_L_X8Y148_SLICE_X10Y148_CO6),
.I1(CLBLM_R_X7Y146_SLICE_X8Y146_BQ),
.I2(CLBLM_R_X7Y148_SLICE_X8Y148_AQ),
.I3(CLBLM_L_X8Y148_SLICE_X10Y148_AQ),
.I4(CLBLM_L_X10Y144_SLICE_X12Y144_AO6),
.I5(1'b1),
.O5(CLBLM_L_X8Y145_SLICE_X11Y145_AO5),
.O6(CLBLM_L_X8Y145_SLICE_X11Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y146_SLICE_X10Y146_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y146_SLICE_X10Y146_AO5),
.Q(CLBLM_L_X8Y146_SLICE_X10Y146_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y146_SLICE_X10Y146_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y146_SLICE_X10Y146_CO5),
.Q(CLBLM_L_X8Y146_SLICE_X10Y146_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y146_SLICE_X10Y146_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y146_SLICE_X10Y146_AO6),
.Q(CLBLM_L_X8Y146_SLICE_X10Y146_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y146_SLICE_X10Y146_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y146_SLICE_X10Y146_BO6),
.Q(CLBLM_L_X8Y146_SLICE_X10Y146_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y146_SLICE_X10Y146_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y146_SLICE_X10Y146_CO6),
.Q(CLBLM_L_X8Y146_SLICE_X10Y146_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y146_SLICE_X10Y146_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y146_SLICE_X10Y146_DO6),
.Q(CLBLM_L_X8Y146_SLICE_X10Y146_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haafcaa00aafcaa00)
  ) CLBLM_L_X8Y146_SLICE_X10Y146_DLUT (
.I0(CLBLL_L_X4Y145_SLICE_X5Y145_AQ),
.I1(CLBLM_L_X8Y143_SLICE_X10Y143_CQ),
.I2(CLBLM_L_X8Y146_SLICE_X10Y146_DQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X10Y143_SLICE_X12Y143_AO6),
.I5(1'b1),
.O5(CLBLM_L_X8Y146_SLICE_X10Y146_DO5),
.O6(CLBLM_L_X8Y146_SLICE_X10Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0aaf0aaccf0ccf0)
  ) CLBLM_L_X8Y146_SLICE_X10Y146_CLUT (
.I0(CLBLL_L_X4Y144_SLICE_X5Y144_B5Q),
.I1(CLBLL_L_X4Y141_SLICE_X5Y141_A5Q),
.I2(CLBLM_L_X10Y150_SLICE_X13Y150_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y146_SLICE_X10Y146_CO5),
.O6(CLBLM_L_X8Y146_SLICE_X10Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000e0eee0ee)
  ) CLBLM_L_X8Y146_SLICE_X10Y146_BLUT (
.I0(CLBLL_L_X4Y146_SLICE_X5Y146_B5Q),
.I1(CLBLM_L_X8Y146_SLICE_X10Y146_BQ),
.I2(CLBLM_R_X5Y144_SLICE_X6Y144_DQ),
.I3(CLBLM_R_X3Y148_SLICE_X2Y148_D5Q),
.I4(CLBLM_L_X8Y141_SLICE_X10Y141_BQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_L_X8Y146_SLICE_X10Y146_BO5),
.O6(CLBLM_L_X8Y146_SLICE_X10Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'he4e4e4e4ffaa5500)
  ) CLBLM_L_X8Y146_SLICE_X10Y146_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(RIOB33_X105Y111_IOB_X1Y112_I),
.I2(CLBLM_L_X8Y143_SLICE_X10Y143_CQ),
.I3(CLBLL_L_X4Y149_SLICE_X4Y149_C5Q),
.I4(CLBLM_R_X7Y149_SLICE_X8Y149_DQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y146_SLICE_X10Y146_AO5),
.O6(CLBLM_L_X8Y146_SLICE_X10Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y146_SLICE_X11Y146_A5_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y146_SLICE_X11Y146_AO5),
.Q(CLBLM_L_X8Y146_SLICE_X11Y146_A5Q),
.S(CLBLM_R_X11Y148_SLICE_X14Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y146_SLICE_X11Y146_A_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y146_SLICE_X11Y146_AO6),
.Q(CLBLM_L_X8Y146_SLICE_X11Y146_AQ),
.S(CLBLM_R_X11Y148_SLICE_X14Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y146_SLICE_X11Y146_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y146_SLICE_X11Y146_DO5),
.O6(CLBLM_L_X8Y146_SLICE_X11Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555000055750030)
  ) CLBLM_L_X8Y146_SLICE_X11Y146_CLUT (
.I0(CLBLM_L_X10Y143_SLICE_X12Y143_DO5),
.I1(CLBLM_L_X10Y142_SLICE_X12Y142_DO6),
.I2(CLBLM_L_X8Y146_SLICE_X11Y146_AQ),
.I3(CLBLM_L_X8Y150_SLICE_X10Y150_A5Q),
.I4(CLBLM_L_X8Y146_SLICE_X10Y146_DQ),
.I5(CLBLM_R_X11Y149_SLICE_X14Y149_AQ),
.O5(CLBLM_L_X8Y146_SLICE_X11Y146_CO5),
.O6(CLBLM_L_X8Y146_SLICE_X11Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0004ffff00040004)
  ) CLBLM_L_X8Y146_SLICE_X11Y146_BLUT (
.I0(CLBLM_L_X8Y150_SLICE_X10Y150_A5Q),
.I1(CLBLM_L_X8Y140_SLICE_X10Y140_A5Q),
.I2(CLBLM_L_X10Y142_SLICE_X12Y142_DO6),
.I3(CLBLM_R_X11Y149_SLICE_X14Y149_AQ),
.I4(CLBLM_L_X10Y143_SLICE_X12Y143_DO5),
.I5(CLBLL_L_X4Y146_SLICE_X4Y146_CQ),
.O5(CLBLM_L_X8Y146_SLICE_X11Y146_BO5),
.O6(CLBLM_L_X8Y146_SLICE_X11Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00a0a0a0a0)
  ) CLBLM_L_X8Y146_SLICE_X11Y146_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(1'b1),
.I2(CLBLL_L_X4Y150_SLICE_X5Y150_C5Q),
.I3(CLBLL_L_X4Y146_SLICE_X4Y146_CQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y146_SLICE_X11Y146_AO5),
.O6(CLBLM_L_X8Y146_SLICE_X11Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y147_SLICE_X10Y147_A5_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y147_SLICE_X10Y147_AO5),
.Q(CLBLM_L_X8Y147_SLICE_X10Y147_A5Q),
.S(CLBLM_R_X7Y148_SLICE_X9Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y147_SLICE_X10Y147_B5_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y147_SLICE_X10Y147_BO5),
.Q(CLBLM_L_X8Y147_SLICE_X10Y147_B5Q),
.S(CLBLM_R_X7Y148_SLICE_X9Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y147_SLICE_X10Y147_A_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y147_SLICE_X10Y147_AO6),
.Q(CLBLM_L_X8Y147_SLICE_X10Y147_AQ),
.S(CLBLM_R_X7Y148_SLICE_X9Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y147_SLICE_X10Y147_B_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y147_SLICE_X10Y147_BO6),
.Q(CLBLM_L_X8Y147_SLICE_X10Y147_BQ),
.S(CLBLM_R_X7Y148_SLICE_X9Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff0fcf00cc)
  ) CLBLM_L_X8Y147_SLICE_X10Y147_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y148_SLICE_X10Y148_BQ),
.I2(CLBLM_R_X5Y145_SLICE_X7Y145_BO6),
.I3(CLBLM_L_X10Y148_SLICE_X12Y148_BO5),
.I4(CLBLM_L_X8Y148_SLICE_X10Y148_A5Q),
.I5(CLBLM_L_X12Y149_SLICE_X16Y149_CO6),
.O5(CLBLM_L_X8Y147_SLICE_X10Y147_DO5),
.O6(CLBLM_L_X8Y147_SLICE_X10Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff3b0a3b0a)
  ) CLBLM_L_X8Y147_SLICE_X10Y147_CLUT (
.I0(CLBLL_L_X4Y144_SLICE_X5Y144_AQ),
.I1(CLBLM_R_X5Y145_SLICE_X7Y145_BO6),
.I2(CLBLM_L_X10Y143_SLICE_X12Y143_DO6),
.I3(CLBLM_L_X8Y147_SLICE_X11Y147_AQ),
.I4(1'b1),
.I5(CLBLM_L_X12Y149_SLICE_X16Y149_CO6),
.O5(CLBLM_L_X8Y147_SLICE_X10Y147_CO5),
.O6(CLBLM_L_X8Y147_SLICE_X10Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa000088888888)
  ) CLBLM_L_X8Y147_SLICE_X10Y147_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X8Y145_SLICE_X10Y145_BQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X7Y147_SLICE_X8Y147_BQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y147_SLICE_X10Y147_BO5),
.O6(CLBLM_L_X8Y147_SLICE_X10Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0aa00aa00)
  ) CLBLM_L_X8Y147_SLICE_X10Y147_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(1'b1),
.I2(CLBLM_R_X7Y150_SLICE_X9Y150_AQ),
.I3(CLBLM_R_X5Y154_SLICE_X7Y154_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y147_SLICE_X10Y147_AO5),
.O6(CLBLM_L_X8Y147_SLICE_X10Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y147_SLICE_X11Y147_A5_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y147_SLICE_X11Y147_AO5),
.Q(CLBLM_L_X8Y147_SLICE_X11Y147_A5Q),
.S(CLBLM_R_X11Y148_SLICE_X15Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y147_SLICE_X11Y147_A_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y147_SLICE_X11Y147_AO6),
.Q(CLBLM_L_X8Y147_SLICE_X11Y147_AQ),
.S(CLBLM_R_X11Y148_SLICE_X15Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff55f500f0)
  ) CLBLM_L_X8Y147_SLICE_X11Y147_DLUT (
.I0(CLBLM_L_X10Y143_SLICE_X12Y143_AO5),
.I1(1'b1),
.I2(CLBLM_R_X7Y149_SLICE_X9Y149_DQ),
.I3(CLBLM_L_X8Y148_SLICE_X10Y148_CO6),
.I4(CLBLM_L_X10Y149_SLICE_X12Y149_CQ),
.I5(CLBLM_L_X8Y147_SLICE_X10Y147_CO6),
.O5(CLBLM_L_X8Y147_SLICE_X11Y147_DO5),
.O6(CLBLM_L_X8Y147_SLICE_X11Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h77f755f533f300f0)
  ) CLBLM_L_X8Y147_SLICE_X11Y147_CLUT (
.I0(CLBLM_L_X10Y144_SLICE_X12Y144_AO6),
.I1(CLBLM_R_X7Y148_SLICE_X8Y148_BO5),
.I2(CLBLM_R_X5Y154_SLICE_X6Y154_AQ),
.I3(CLBLM_L_X10Y143_SLICE_X12Y143_DO5),
.I4(CLBLM_L_X8Y149_SLICE_X11Y149_B5Q),
.I5(CLBLM_L_X10Y146_SLICE_X13Y146_AQ),
.O5(CLBLM_L_X8Y147_SLICE_X11Y147_CO5),
.O6(CLBLM_L_X8Y147_SLICE_X11Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffefefffe)
  ) CLBLM_L_X8Y147_SLICE_X11Y147_BLUT (
.I0(CLBLM_L_X8Y147_SLICE_X11Y147_DO6),
.I1(CLBLM_R_X7Y144_SLICE_X8Y144_CO6),
.I2(CLBLM_R_X11Y146_SLICE_X15Y146_DO6),
.I3(CLBLM_R_X7Y144_SLICE_X8Y144_A5Q),
.I4(CLBLM_L_X10Y148_SLICE_X12Y148_BO5),
.I5(CLBLM_L_X8Y147_SLICE_X11Y147_CO6),
.O5(CLBLM_L_X8Y147_SLICE_X11Y147_BO5),
.O6(CLBLM_L_X8Y147_SLICE_X11Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888aa00aa00)
  ) CLBLM_L_X8Y147_SLICE_X11Y147_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X5Y145_SLICE_X6Y145_CQ),
.I2(1'b1),
.I3(CLBLM_R_X7Y151_SLICE_X9Y151_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y147_SLICE_X11Y147_AO5),
.O6(CLBLM_L_X8Y147_SLICE_X11Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y148_SLICE_X10Y148_A5_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y148_SLICE_X10Y148_AO5),
.Q(CLBLM_L_X8Y148_SLICE_X10Y148_A5Q),
.S(CLBLM_R_X7Y148_SLICE_X9Y148_AO5)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y148_SLICE_X10Y148_A_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y148_SLICE_X10Y148_AO6),
.Q(CLBLM_L_X8Y148_SLICE_X10Y148_AQ),
.S(CLBLM_R_X7Y148_SLICE_X9Y148_AO5)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y148_SLICE_X10Y148_B_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y151_SLICE_X11Y151_BO6),
.Q(CLBLM_L_X8Y148_SLICE_X10Y148_BQ),
.S(CLBLM_R_X7Y148_SLICE_X9Y148_AO5)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffdeffde)
  ) CLBLM_L_X8Y148_SLICE_X10Y148_DLUT (
.I0(CLBLL_L_X4Y141_SLICE_X5Y141_AQ),
.I1(CLBLM_R_X3Y154_SLICE_X3Y154_AQ),
.I2(CLBLM_R_X5Y151_SLICE_X6Y151_DQ),
.I3(CLBLM_R_X7Y146_SLICE_X9Y146_AO5),
.I4(1'b1),
.I5(CLBLM_L_X8Y148_SLICE_X10Y148_BO6),
.O5(CLBLM_L_X8Y148_SLICE_X10Y148_DO5),
.O6(CLBLM_L_X8Y148_SLICE_X10Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffff3300c00088)
  ) CLBLM_L_X8Y148_SLICE_X10Y148_CLUT (
.I0(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.I1(CLBLM_L_X10Y144_SLICE_X13Y144_CO6),
.I2(CLBLL_L_X4Y149_SLICE_X4Y149_CQ),
.I3(CLBLM_L_X8Y150_SLICE_X10Y150_A5Q),
.I4(CLBLM_R_X11Y149_SLICE_X14Y149_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y148_SLICE_X10Y148_CO5),
.O6(CLBLM_L_X8Y148_SLICE_X10Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h66ffff660f000f00)
  ) CLBLM_L_X8Y148_SLICE_X10Y148_BLUT (
.I0(CLBLM_R_X5Y154_SLICE_X7Y154_DQ),
.I1(CLBLM_L_X8Y150_SLICE_X10Y150_AQ),
.I2(CLBLM_L_X10Y145_SLICE_X12Y145_AO6),
.I3(CLBLM_R_X7Y150_SLICE_X8Y150_D5Q),
.I4(CLBLM_L_X8Y151_SLICE_X10Y151_DQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y148_SLICE_X10Y148_BO5),
.O6(CLBLM_L_X8Y148_SLICE_X10Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000f0f00000)
  ) CLBLM_L_X8Y148_SLICE_X10Y148_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X7Y151_SLICE_X9Y151_AQ),
.I3(CLBLM_R_X5Y146_SLICE_X7Y146_CQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y148_SLICE_X10Y148_AO5),
.O6(CLBLM_L_X8Y148_SLICE_X10Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y148_SLICE_X11Y148_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y148_SLICE_X11Y148_BO5),
.Q(CLBLM_L_X8Y148_SLICE_X11Y148_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y148_SLICE_X11Y148_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y148_SLICE_X11Y148_CO5),
.Q(CLBLM_L_X8Y148_SLICE_X11Y148_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y148_SLICE_X11Y148_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y148_SLICE_X11Y148_AO6),
.Q(CLBLM_L_X8Y148_SLICE_X11Y148_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y148_SLICE_X11Y148_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y148_SLICE_X11Y148_BO6),
.Q(CLBLM_L_X8Y148_SLICE_X11Y148_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y148_SLICE_X11Y148_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y148_SLICE_X11Y148_CO6),
.Q(CLBLM_L_X8Y148_SLICE_X11Y148_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y148_SLICE_X11Y148_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y148_SLICE_X11Y148_DO6),
.Q(CLBLM_L_X8Y148_SLICE_X11Y148_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffc4c80000c4c8)
  ) CLBLM_L_X8Y148_SLICE_X11Y148_DLUT (
.I0(RIOB33_X105Y111_IOB_X1Y112_I),
.I1(CLBLM_L_X8Y143_SLICE_X11Y143_A5Q),
.I2(CLBLM_L_X8Y148_SLICE_X11Y148_DQ),
.I3(CLBLM_L_X8Y148_SLICE_X11Y148_BQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X7Y148_SLICE_X8Y148_AQ),
.O5(CLBLM_L_X8Y148_SLICE_X11Y148_DO5),
.O6(CLBLM_L_X8Y148_SLICE_X11Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcacacacaff0ff000)
  ) CLBLM_L_X8Y148_SLICE_X11Y148_CLUT (
.I0(CLBLL_L_X2Y149_SLICE_X0Y149_AQ),
.I1(CLBLM_L_X10Y153_SLICE_X12Y153_AQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_L_X10Y150_SLICE_X13Y150_BQ),
.I4(CLBLM_R_X7Y145_SLICE_X8Y145_C5Q),
.I5(1'b1),
.O5(CLBLM_L_X8Y148_SLICE_X11Y148_CO5),
.O6(CLBLM_L_X8Y148_SLICE_X11Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hafafa0a0cfc0cfc0)
  ) CLBLM_L_X8Y148_SLICE_X11Y148_BLUT (
.I0(CLBLM_L_X8Y151_SLICE_X10Y151_B5Q),
.I1(CLBLM_L_X8Y152_SLICE_X10Y152_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X7Y144_SLICE_X8Y144_A5Q),
.I4(RIOB33_X105Y111_IOB_X1Y112_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y148_SLICE_X11Y148_BO5),
.O6(CLBLM_L_X8Y148_SLICE_X11Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccff55f050)
  ) CLBLM_L_X8Y148_SLICE_X11Y148_ALUT (
.I0(CLBLM_R_X5Y149_SLICE_X6Y149_D5Q),
.I1(CLBLM_L_X8Y146_SLICE_X10Y146_CQ),
.I2(CLBLM_L_X8Y148_SLICE_X11Y148_AQ),
.I3(CLBLM_L_X8Y150_SLICE_X11Y150_B5Q),
.I4(CLBLM_R_X11Y148_SLICE_X15Y148_AQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_L_X8Y148_SLICE_X11Y148_AO5),
.O6(CLBLM_L_X8Y148_SLICE_X11Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y149_SLICE_X10Y149_A5_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y149_SLICE_X10Y149_AO5),
.Q(CLBLM_L_X8Y149_SLICE_X10Y149_A5Q),
.S(CLBLM_R_X11Y148_SLICE_X14Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y149_SLICE_X10Y149_B5_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y149_SLICE_X10Y149_BO5),
.Q(CLBLM_L_X8Y149_SLICE_X10Y149_B5Q),
.S(CLBLM_R_X11Y148_SLICE_X14Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y149_SLICE_X10Y149_A_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y149_SLICE_X10Y149_AO6),
.Q(CLBLM_L_X8Y149_SLICE_X10Y149_AQ),
.S(CLBLM_R_X11Y148_SLICE_X14Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y149_SLICE_X10Y149_B_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y149_SLICE_X10Y149_BO6),
.Q(CLBLM_L_X8Y149_SLICE_X10Y149_BQ),
.S(CLBLM_R_X11Y148_SLICE_X14Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3bff0aff3b3b0a0a)
  ) CLBLM_L_X8Y149_SLICE_X10Y149_DLUT (
.I0(CLBLM_L_X8Y146_SLICE_X10Y146_C5Q),
.I1(CLBLM_L_X10Y144_SLICE_X12Y144_AO6),
.I2(CLBLM_L_X10Y148_SLICE_X12Y148_BO5),
.I3(CLBLM_L_X8Y148_SLICE_X10Y148_CO6),
.I4(CLBLM_L_X8Y149_SLICE_X10Y149_B5Q),
.I5(CLBLL_L_X4Y150_SLICE_X4Y150_AQ),
.O5(CLBLM_L_X8Y149_SLICE_X10Y149_DO5),
.O6(CLBLM_L_X8Y149_SLICE_X10Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h33f3bbfb00f0aafa)
  ) CLBLM_L_X8Y149_SLICE_X10Y149_CLUT (
.I0(CLBLM_L_X8Y150_SLICE_X11Y150_BQ),
.I1(CLBLM_L_X10Y148_SLICE_X12Y148_BO5),
.I2(CLBLM_R_X7Y149_SLICE_X9Y149_CQ),
.I3(CLBLM_L_X8Y148_SLICE_X10Y148_CO6),
.I4(CLBLM_L_X10Y144_SLICE_X12Y144_AO6),
.I5(CLBLM_R_X5Y150_SLICE_X7Y150_A5Q),
.O5(CLBLM_L_X8Y149_SLICE_X10Y149_CO5),
.O6(CLBLM_L_X8Y149_SLICE_X10Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0000c0c0c0c0)
  ) CLBLM_L_X8Y149_SLICE_X10Y149_BLUT (
.I0(1'b1),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X7Y146_SLICE_X9Y146_BQ),
.I3(1'b1),
.I4(CLBLL_L_X2Y147_SLICE_X1Y147_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y149_SLICE_X10Y149_BO5),
.O6(CLBLM_L_X8Y149_SLICE_X10Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0000c0c0c0c0)
  ) CLBLM_L_X8Y149_SLICE_X10Y149_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X7Y149_SLICE_X9Y149_DQ),
.I3(1'b1),
.I4(CLBLM_R_X5Y144_SLICE_X7Y144_CQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y149_SLICE_X10Y149_AO5),
.O6(CLBLM_L_X8Y149_SLICE_X10Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y149_SLICE_X11Y149_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y149_SLICE_X11Y149_BO5),
.Q(CLBLM_L_X8Y149_SLICE_X11Y149_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y149_SLICE_X11Y149_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y149_SLICE_X11Y149_AO6),
.Q(CLBLM_L_X8Y149_SLICE_X11Y149_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y149_SLICE_X11Y149_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y149_SLICE_X11Y149_BO6),
.Q(CLBLM_L_X8Y149_SLICE_X11Y149_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y149_SLICE_X11Y149_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y149_SLICE_X11Y149_CO6),
.Q(CLBLM_L_X8Y149_SLICE_X11Y149_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffccffccffccfffc)
  ) CLBLM_L_X8Y149_SLICE_X11Y149_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y149_SLICE_X10Y149_CO6),
.I2(CLBLM_L_X8Y150_SLICE_X10Y150_AQ),
.I3(CLBLM_R_X7Y149_SLICE_X9Y149_BO6),
.I4(CLBLM_L_X10Y145_SLICE_X12Y145_AO6),
.I5(CLBLM_R_X11Y143_SLICE_X14Y143_CO5),
.O5(CLBLM_L_X8Y149_SLICE_X11Y149_DO5),
.O6(CLBLM_L_X8Y149_SLICE_X11Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0b1b1a0a0b1b1)
  ) CLBLM_L_X8Y149_SLICE_X11Y149_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLL_L_X2Y151_SLICE_X1Y151_BQ),
.I2(CLBLM_L_X8Y147_SLICE_X11Y147_AQ),
.I3(1'b1),
.I4(CLBLM_R_X7Y151_SLICE_X9Y151_CQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y149_SLICE_X11Y149_CO5),
.O6(CLBLM_L_X8Y149_SLICE_X11Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaff00f0f0cccc)
  ) CLBLM_L_X8Y149_SLICE_X11Y149_BLUT (
.I0(CLBLL_L_X4Y149_SLICE_X5Y149_CQ),
.I1(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I2(CLBLM_L_X8Y147_SLICE_X10Y147_AQ),
.I3(CLBLM_L_X8Y149_SLICE_X11Y149_CQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y149_SLICE_X11Y149_BO5),
.O6(CLBLM_L_X8Y149_SLICE_X11Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffccffe400cc00e4)
  ) CLBLM_L_X8Y149_SLICE_X11Y149_ALUT (
.I0(CLBLM_R_X3Y148_SLICE_X2Y148_D5Q),
.I1(CLBLM_L_X8Y145_SLICE_X10Y145_BQ),
.I2(CLBLM_L_X8Y149_SLICE_X11Y149_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X5Y144_SLICE_X6Y144_DQ),
.I5(CLBLM_R_X7Y151_SLICE_X9Y151_CQ),
.O5(CLBLM_L_X8Y149_SLICE_X11Y149_AO5),
.O6(CLBLM_L_X8Y149_SLICE_X11Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y150_SLICE_X10Y150_A5_FDSE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y150_SLICE_X10Y150_AO5),
.Q(CLBLM_L_X8Y150_SLICE_X10Y150_A5Q),
.S(CLBLM_R_X11Y148_SLICE_X15Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y150_SLICE_X10Y150_A_FDSE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y150_SLICE_X10Y150_AO6),
.Q(CLBLM_L_X8Y150_SLICE_X10Y150_AQ),
.S(CLBLM_R_X11Y148_SLICE_X15Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafafafafafafafa)
  ) CLBLM_L_X8Y150_SLICE_X10Y150_DLUT (
.I0(CLBLM_R_X7Y149_SLICE_X9Y149_DO6),
.I1(1'b1),
.I2(CLBLM_L_X8Y149_SLICE_X10Y149_DO6),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y150_SLICE_X10Y150_DO5),
.O6(CLBLM_L_X8Y150_SLICE_X10Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfaaafffffaaafaaa)
  ) CLBLM_L_X8Y150_SLICE_X10Y150_CLUT (
.I0(CLBLM_L_X12Y149_SLICE_X16Y149_CO6),
.I1(1'b1),
.I2(CLBLM_L_X10Y143_SLICE_X12Y143_BO6),
.I3(CLBLM_L_X8Y152_SLICE_X10Y152_CQ),
.I4(CLBLM_R_X7Y146_SLICE_X8Y146_AO6),
.I5(CLBLM_L_X8Y149_SLICE_X10Y149_BQ),
.O5(CLBLM_L_X8Y150_SLICE_X10Y150_CO5),
.O6(CLBLM_L_X8Y150_SLICE_X10Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffffec)
  ) CLBLM_L_X8Y150_SLICE_X10Y150_BLUT (
.I0(CLBLM_L_X10Y143_SLICE_X12Y143_BO5),
.I1(CLBLM_R_X7Y148_SLICE_X8Y148_CO6),
.I2(CLBLM_L_X8Y152_SLICE_X10Y152_AQ),
.I3(CLBLM_R_X5Y150_SLICE_X7Y150_DO6),
.I4(CLBLM_L_X8Y146_SLICE_X11Y146_CO6),
.I5(CLBLM_L_X8Y150_SLICE_X10Y150_CO6),
.O5(CLBLM_L_X8Y150_SLICE_X10Y150_BO5),
.O6(CLBLM_L_X8Y150_SLICE_X10Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000cc00cc00)
  ) CLBLM_L_X8Y150_SLICE_X10Y150_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y145_SLICE_X10Y145_AQ),
.I2(1'b1),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X3Y153_SLICE_X3Y153_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y150_SLICE_X10Y150_AO5),
.O6(CLBLM_L_X8Y150_SLICE_X10Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y150_SLICE_X11Y150_B5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y150_SLICE_X11Y150_BO5),
.Q(CLBLM_L_X8Y150_SLICE_X11Y150_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y150_SLICE_X11Y150_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y150_SLICE_X11Y150_AO6),
.Q(CLBLM_L_X8Y150_SLICE_X11Y150_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y150_SLICE_X11Y150_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y150_SLICE_X11Y150_BO6),
.Q(CLBLM_L_X8Y150_SLICE_X11Y150_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y150_SLICE_X11Y150_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y150_SLICE_X11Y150_CO6),
.Q(CLBLM_L_X8Y150_SLICE_X11Y150_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5fffafffff5fffa)
  ) CLBLM_L_X8Y150_SLICE_X11Y150_DLUT (
.I0(CLBLM_L_X8Y154_SLICE_X10Y154_AQ),
.I1(1'b1),
.I2(CLBLM_R_X7Y146_SLICE_X9Y146_DO6),
.I3(CLBLM_L_X10Y146_SLICE_X13Y146_AQ),
.I4(CLBLM_R_X5Y145_SLICE_X7Y145_AQ),
.I5(CLBLM_R_X7Y152_SLICE_X8Y152_CQ),
.O5(CLBLM_L_X8Y150_SLICE_X11Y150_DO5),
.O6(CLBLM_L_X8Y150_SLICE_X11Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0ffffff66)
  ) CLBLM_L_X8Y150_SLICE_X11Y150_CLUT (
.I0(CLBLM_L_X8Y149_SLICE_X10Y149_B5Q),
.I1(CLBLM_R_X3Y154_SLICE_X3Y154_AQ),
.I2(CLBLM_R_X7Y154_SLICE_X8Y154_CQ),
.I3(CLBLM_L_X8Y151_SLICE_X11Y151_CO6),
.I4(CLBLM_L_X8Y150_SLICE_X11Y150_DO6),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_L_X8Y150_SLICE_X11Y150_CO5),
.O6(CLBLM_L_X8Y150_SLICE_X11Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0aaf0aaccffcc00)
  ) CLBLM_L_X8Y150_SLICE_X11Y150_BLUT (
.I0(CLBLM_L_X8Y152_SLICE_X11Y152_A5Q),
.I1(CLBLM_R_X7Y151_SLICE_X8Y151_BQ),
.I2(CLBLM_R_X7Y153_SLICE_X9Y153_CQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(RIOB33_X105Y111_IOB_X1Y112_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y150_SLICE_X11Y150_BO5),
.O6(CLBLM_L_X8Y150_SLICE_X11Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00bbbbb0b0)
  ) CLBLM_L_X8Y150_SLICE_X11Y150_ALUT (
.I0(CLBLM_L_X8Y150_SLICE_X11Y150_B5Q),
.I1(CLBLM_R_X5Y149_SLICE_X6Y149_D5Q),
.I2(CLBLM_L_X8Y150_SLICE_X11Y150_AQ),
.I3(CLBLM_R_X5Y151_SLICE_X7Y151_AQ),
.I4(CLBLM_L_X8Y147_SLICE_X10Y147_A5Q),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_L_X8Y150_SLICE_X11Y150_AO5),
.O6(CLBLM_L_X8Y150_SLICE_X11Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y151_SLICE_X10Y151_B5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y151_SLICE_X10Y151_BO5),
.Q(CLBLM_L_X8Y151_SLICE_X10Y151_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y151_SLICE_X10Y151_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y151_SLICE_X10Y151_AO6),
.Q(CLBLM_L_X8Y151_SLICE_X10Y151_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y151_SLICE_X10Y151_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y151_SLICE_X10Y151_BO6),
.Q(CLBLM_L_X8Y151_SLICE_X10Y151_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y151_SLICE_X10Y151_D_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y151_SLICE_X10Y151_DO6),
.Q(CLBLM_L_X8Y151_SLICE_X10Y151_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccca00aa00a)
  ) CLBLM_L_X8Y151_SLICE_X10Y151_DLUT (
.I0(CLBLM_R_X3Y152_SLICE_X2Y152_BQ),
.I1(CLBLM_L_X8Y146_SLICE_X10Y146_A5Q),
.I2(CLBLM_L_X8Y151_SLICE_X10Y151_DQ),
.I3(CLBLM_L_X8Y152_SLICE_X11Y152_CO6),
.I4(1'b1),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_L_X8Y151_SLICE_X10Y151_DO5),
.O6(CLBLM_L_X8Y151_SLICE_X10Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00fffffffc)
  ) CLBLM_L_X8Y151_SLICE_X10Y151_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X5Y153_SLICE_X6Y153_AQ),
.I2(CLBLM_R_X7Y143_SLICE_X9Y143_BQ),
.I3(CLBLL_L_X4Y150_SLICE_X5Y150_CQ),
.I4(CLBLM_R_X3Y151_SLICE_X3Y151_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y151_SLICE_X10Y151_CO5),
.O6(CLBLM_L_X8Y151_SLICE_X10Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0ccf0ccfff000f0)
  ) CLBLM_L_X8Y151_SLICE_X10Y151_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y146_SLICE_X10Y146_C5Q),
.I2(CLBLM_R_X7Y148_SLICE_X9Y148_C5Q),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X11Y151_SLICE_X14Y151_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y151_SLICE_X10Y151_BO5),
.O6(CLBLM_L_X8Y151_SLICE_X10Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccaaaaf0aa)
  ) CLBLM_L_X8Y151_SLICE_X10Y151_ALUT (
.I0(CLBLL_L_X4Y148_SLICE_X4Y148_AQ),
.I1(CLBLM_L_X10Y152_SLICE_X12Y152_AQ),
.I2(CLBLM_L_X8Y151_SLICE_X10Y151_AQ),
.I3(CLBLM_R_X3Y147_SLICE_X3Y147_BQ),
.I4(CLBLM_R_X5Y144_SLICE_X6Y144_CQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_L_X8Y151_SLICE_X10Y151_AO5),
.O6(CLBLM_L_X8Y151_SLICE_X10Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y151_SLICE_X11Y151_A5_FDSE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y151_SLICE_X11Y151_AO5),
.Q(CLBLM_L_X8Y151_SLICE_X11Y151_A5Q),
.S(CLBLM_R_X11Y150_SLICE_X14Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y151_SLICE_X11Y151_A_FDSE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y151_SLICE_X11Y151_AO6),
.Q(CLBLM_L_X8Y151_SLICE_X11Y151_AQ),
.S(CLBLM_R_X11Y150_SLICE_X14Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5affff5a5affff5a)
  ) CLBLM_L_X8Y151_SLICE_X11Y151_DLUT (
.I0(CLBLM_R_X7Y148_SLICE_X8Y148_AQ),
.I1(1'b1),
.I2(CLBLM_R_X7Y154_SLICE_X8Y154_CQ),
.I3(CLBLM_R_X5Y148_SLICE_X6Y148_B5Q),
.I4(CLBLM_L_X8Y151_SLICE_X10Y151_DQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y151_SLICE_X11Y151_DO5),
.O6(CLBLM_L_X8Y151_SLICE_X11Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffdfeffffffdfe)
  ) CLBLM_L_X8Y151_SLICE_X11Y151_CLUT (
.I0(CLBLM_L_X8Y148_SLICE_X10Y148_AQ),
.I1(CLBLM_L_X8Y151_SLICE_X11Y151_DO6),
.I2(CLBLM_L_X8Y140_SLICE_X10Y140_A5Q),
.I3(CLBLM_R_X7Y151_SLICE_X9Y151_DQ),
.I4(CLBLM_L_X8Y151_SLICE_X11Y151_BO5),
.I5(CLBLM_R_X5Y151_SLICE_X6Y151_DQ),
.O5(CLBLM_L_X8Y151_SLICE_X11Y151_CO5),
.O6(CLBLM_L_X8Y151_SLICE_X11Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc00007dbe7dbe)
  ) CLBLM_L_X8Y151_SLICE_X11Y151_BLUT (
.I0(CLBLM_R_X7Y151_SLICE_X8Y151_CQ),
.I1(CLBLM_L_X8Y153_SLICE_X11Y153_BQ),
.I2(CLBLM_L_X8Y150_SLICE_X11Y150_BQ),
.I3(CLBLM_R_X5Y154_SLICE_X7Y154_DQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y151_SLICE_X11Y151_BO5),
.O6(CLBLM_L_X8Y151_SLICE_X11Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc0088888888)
  ) CLBLM_L_X8Y151_SLICE_X11Y151_ALUT (
.I0(CLBLM_R_X7Y149_SLICE_X9Y149_CQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(1'b1),
.I3(CLBLM_R_X5Y141_SLICE_X7Y141_A5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y151_SLICE_X11Y151_AO5),
.O6(CLBLM_L_X8Y151_SLICE_X11Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y152_SLICE_X10Y152_D5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y152_SLICE_X10Y152_DO5),
.Q(CLBLM_L_X8Y152_SLICE_X10Y152_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y152_SLICE_X10Y152_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y152_SLICE_X10Y152_AO6),
.Q(CLBLM_L_X8Y152_SLICE_X10Y152_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y152_SLICE_X10Y152_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y152_SLICE_X10Y152_BO6),
.Q(CLBLM_L_X8Y152_SLICE_X10Y152_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y152_SLICE_X10Y152_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y152_SLICE_X10Y152_CO6),
.Q(CLBLM_L_X8Y152_SLICE_X10Y152_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y152_SLICE_X10Y152_D_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y152_SLICE_X10Y152_DO6),
.Q(CLBLM_L_X8Y152_SLICE_X10Y152_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa50fa50e4e4e4e4)
  ) CLBLM_L_X8Y152_SLICE_X10Y152_DLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLL_L_X4Y149_SLICE_X4Y149_CQ),
.I2(CLBLM_R_X7Y152_SLICE_X9Y152_CQ),
.I3(CLBLM_L_X8Y146_SLICE_X10Y146_C5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y152_SLICE_X10Y152_DO5),
.O6(CLBLM_L_X8Y152_SLICE_X10Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hefefefaa45454500)
  ) CLBLM_L_X8Y152_SLICE_X10Y152_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X5Y144_SLICE_X6Y144_DQ),
.I2(CLBLM_R_X3Y148_SLICE_X2Y148_D5Q),
.I3(CLBLM_L_X8Y151_SLICE_X11Y151_A5Q),
.I4(CLBLM_L_X8Y152_SLICE_X10Y152_CQ),
.I5(CLBLM_R_X5Y147_SLICE_X7Y147_CQ),
.O5(CLBLM_L_X8Y152_SLICE_X10Y152_CO5),
.O6(CLBLM_L_X8Y152_SLICE_X10Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaf0aafcaaf0aa30)
  ) CLBLM_L_X8Y152_SLICE_X10Y152_BLUT (
.I0(CLBLM_L_X8Y146_SLICE_X10Y146_BQ),
.I1(CLBLM_R_X3Y147_SLICE_X3Y147_BQ),
.I2(CLBLL_L_X4Y145_SLICE_X4Y145_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X5Y144_SLICE_X6Y144_CQ),
.I5(CLBLM_L_X8Y152_SLICE_X10Y152_BQ),
.O5(CLBLM_L_X8Y152_SLICE_X10Y152_BO5),
.O6(CLBLM_L_X8Y152_SLICE_X10Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffa5550bbba1110)
  ) CLBLM_L_X8Y152_SLICE_X10Y152_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X3Y147_SLICE_X3Y147_BQ),
.I2(CLBLM_L_X8Y152_SLICE_X10Y152_AQ),
.I3(CLBLM_R_X11Y150_SLICE_X14Y150_AQ),
.I4(CLBLM_L_X10Y146_SLICE_X12Y146_AQ),
.I5(CLBLM_R_X5Y144_SLICE_X6Y144_CQ),
.O5(CLBLM_L_X8Y152_SLICE_X10Y152_AO5),
.O6(CLBLM_L_X8Y152_SLICE_X10Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y152_SLICE_X11Y152_A5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y152_SLICE_X11Y152_AO5),
.Q(CLBLM_L_X8Y152_SLICE_X11Y152_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y152_SLICE_X11Y152_B5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y152_SLICE_X11Y152_BO5),
.Q(CLBLM_L_X8Y152_SLICE_X11Y152_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y152_SLICE_X11Y152_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y152_SLICE_X11Y152_AO6),
.Q(CLBLM_L_X8Y152_SLICE_X11Y152_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y152_SLICE_X11Y152_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y152_SLICE_X11Y152_BO6),
.Q(CLBLM_L_X8Y152_SLICE_X11Y152_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h4555ffff10000000)
  ) CLBLM_L_X8Y152_SLICE_X11Y152_DLUT (
.I0(CLBLM_L_X8Y153_SLICE_X10Y153_AQ),
.I1(CLBLM_R_X3Y150_SLICE_X3Y150_BQ),
.I2(CLBLM_L_X10Y153_SLICE_X12Y153_BQ),
.I3(CLBLM_L_X8Y153_SLICE_X10Y153_BQ),
.I4(CLBLM_R_X7Y145_SLICE_X8Y145_B5Q),
.I5(CLBLM_L_X8Y152_SLICE_X11Y152_B5Q),
.O5(CLBLM_L_X8Y152_SLICE_X11Y152_DO5),
.O6(CLBLM_L_X8Y152_SLICE_X11Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fffffffffffffff)
  ) CLBLM_L_X8Y152_SLICE_X11Y152_CLUT (
.I0(CLBLM_L_X8Y154_SLICE_X10Y154_AQ),
.I1(CLBLM_R_X3Y154_SLICE_X3Y154_AQ),
.I2(CLBLM_L_X8Y153_SLICE_X11Y153_BQ),
.I3(CLBLM_R_X5Y154_SLICE_X7Y154_DQ),
.I4(CLBLM_R_X7Y154_SLICE_X8Y154_CQ),
.I5(CLBLM_R_X7Y152_SLICE_X8Y152_CQ),
.O5(CLBLM_L_X8Y152_SLICE_X11Y152_CO5),
.O6(CLBLM_L_X8Y152_SLICE_X11Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffcc00f0aaf0aa)
  ) CLBLM_L_X8Y152_SLICE_X11Y152_BLUT (
.I0(CLBLM_L_X8Y152_SLICE_X11Y152_DO6),
.I1(CLBLL_L_X2Y148_SLICE_X0Y148_A5Q),
.I2(CLBLL_L_X4Y144_SLICE_X5Y144_C5Q),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X8Y153_SLICE_X11Y153_CO6),
.I5(1'b1),
.O5(CLBLM_L_X8Y152_SLICE_X11Y152_BO5),
.O6(CLBLM_L_X8Y152_SLICE_X11Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0aaf0aaccffcc00)
  ) CLBLM_L_X8Y152_SLICE_X11Y152_ALUT (
.I0(CLBLM_L_X10Y145_SLICE_X13Y145_CO6),
.I1(CLBLM_L_X8Y140_SLICE_X10Y140_A5Q),
.I2(CLBLL_L_X4Y152_SLICE_X4Y152_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X10Y148_SLICE_X13Y148_CO6),
.I5(1'b1),
.O5(CLBLM_L_X8Y152_SLICE_X11Y152_AO5),
.O6(CLBLM_L_X8Y152_SLICE_X11Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y153_SLICE_X10Y153_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y153_SLICE_X10Y153_AO6),
.Q(CLBLM_L_X8Y153_SLICE_X10Y153_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y153_SLICE_X10Y153_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y153_SLICE_X10Y153_BO6),
.Q(CLBLM_L_X8Y153_SLICE_X10Y153_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y153_SLICE_X10Y153_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y153_SLICE_X10Y153_CO6),
.Q(CLBLM_L_X8Y153_SLICE_X10Y153_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h01000000f3f30000)
  ) CLBLM_L_X8Y153_SLICE_X10Y153_DLUT (
.I0(CLBLM_R_X11Y152_SLICE_X14Y152_DO6),
.I1(CLBLM_R_X3Y150_SLICE_X3Y150_BQ),
.I2(CLBLM_L_X8Y153_SLICE_X10Y153_AQ),
.I3(CLBLM_L_X10Y152_SLICE_X12Y152_CQ),
.I4(CLBLM_R_X7Y145_SLICE_X8Y145_B5Q),
.I5(1'b1),
.O5(CLBLM_L_X8Y153_SLICE_X10Y153_DO5),
.O6(CLBLM_L_X8Y153_SLICE_X10Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfaf3faf3faf0faf0)
  ) CLBLM_L_X8Y153_SLICE_X10Y153_CLUT (
.I0(CLBLM_L_X8Y150_SLICE_X10Y150_AQ),
.I1(CLBLM_L_X8Y153_SLICE_X10Y153_CQ),
.I2(CLBLM_R_X7Y153_SLICE_X8Y153_BO6),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(1'b1),
.I5(CLBLM_R_X7Y154_SLICE_X9Y154_BO6),
.O5(CLBLM_L_X8Y153_SLICE_X10Y153_CO5),
.O6(CLBLM_L_X8Y153_SLICE_X10Y153_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff4c004cff460046)
  ) CLBLM_L_X8Y153_SLICE_X10Y153_BLUT (
.I0(CLBLM_R_X7Y145_SLICE_X8Y145_B5Q),
.I1(CLBLM_L_X8Y153_SLICE_X10Y153_BQ),
.I2(CLBLM_L_X8Y153_SLICE_X10Y153_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X8Y147_SLICE_X10Y147_BQ),
.I5(CLBLM_R_X3Y150_SLICE_X3Y150_BQ),
.O5(CLBLM_L_X8Y153_SLICE_X10Y153_BO5),
.O6(CLBLM_L_X8Y153_SLICE_X10Y153_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff88f8000088f8)
  ) CLBLM_L_X8Y153_SLICE_X10Y153_ALUT (
.I0(CLBLM_L_X8Y153_SLICE_X10Y153_DO6),
.I1(CLBLM_L_X8Y152_SLICE_X11Y152_BQ),
.I2(CLBLM_L_X8Y153_SLICE_X10Y153_AQ),
.I3(CLBLM_L_X8Y153_SLICE_X10Y153_DO5),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X7Y143_SLICE_X9Y143_CQ),
.O5(CLBLM_L_X8Y153_SLICE_X10Y153_AO5),
.O6(CLBLM_L_X8Y153_SLICE_X10Y153_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y153_SLICE_X11Y153_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y153_SLICE_X11Y153_BO6),
.Q(CLBLM_L_X8Y153_SLICE_X11Y153_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y153_SLICE_X11Y153_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y153_SLICE_X11Y153_DO5),
.O6(CLBLM_L_X8Y153_SLICE_X11Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0fffbf00000040)
  ) CLBLM_L_X8Y153_SLICE_X11Y153_CLUT (
.I0(CLBLM_R_X11Y152_SLICE_X14Y152_DO6),
.I1(CLBLM_L_X10Y152_SLICE_X12Y152_CQ),
.I2(CLBLM_R_X7Y145_SLICE_X8Y145_B5Q),
.I3(CLBLM_R_X3Y150_SLICE_X3Y150_BQ),
.I4(CLBLM_L_X8Y153_SLICE_X10Y153_AQ),
.I5(CLBLM_L_X8Y152_SLICE_X11Y152_BQ),
.O5(CLBLM_L_X8Y153_SLICE_X11Y153_CO5),
.O6(CLBLM_L_X8Y153_SLICE_X11Y153_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf033f000f033f000)
  ) CLBLM_L_X8Y153_SLICE_X11Y153_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y153_SLICE_X11Y153_BQ),
.I2(CLBLM_L_X10Y153_SLICE_X12Y153_BQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X3Y152_SLICE_X2Y152_BQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y153_SLICE_X11Y153_BO5),
.O6(CLBLM_L_X8Y153_SLICE_X11Y153_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcecc0200a0a0a0a0)
  ) CLBLM_L_X8Y153_SLICE_X11Y153_ALUT (
.I0(CLBLM_R_X3Y150_SLICE_X2Y150_CO5),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(CLBLM_L_X12Y151_SLICE_X16Y151_BQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y153_SLICE_X11Y153_AO5),
.O6(CLBLM_L_X8Y153_SLICE_X11Y153_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y154_SLICE_X10Y154_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y154_SLICE_X10Y154_AO6),
.Q(CLBLM_L_X8Y154_SLICE_X10Y154_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y154_SLICE_X10Y154_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y154_SLICE_X10Y154_DO5),
.O6(CLBLM_L_X8Y154_SLICE_X10Y154_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y154_SLICE_X10Y154_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y154_SLICE_X10Y154_CO5),
.O6(CLBLM_L_X8Y154_SLICE_X10Y154_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0cff04ff0cff0cff)
  ) CLBLM_L_X8Y154_SLICE_X10Y154_BLUT (
.I0(CLBLM_R_X3Y151_SLICE_X3Y151_C5Q),
.I1(CLBLM_R_X7Y153_SLICE_X8Y153_DO5),
.I2(CLBLM_R_X7Y151_SLICE_X9Y151_AQ),
.I3(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I4(CLBLL_L_X4Y154_SLICE_X4Y154_AQ),
.I5(RIOB33_X105Y131_IOB_X1Y131_I),
.O5(CLBLM_L_X8Y154_SLICE_X10Y154_BO5),
.O6(CLBLM_L_X8Y154_SLICE_X10Y154_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccf0cc00cc5acc00)
  ) CLBLM_L_X8Y154_SLICE_X10Y154_ALUT (
.I0(CLBLM_R_X7Y154_SLICE_X8Y154_CQ),
.I1(CLBLM_R_X11Y151_SLICE_X15Y151_BQ),
.I2(CLBLM_L_X8Y154_SLICE_X10Y154_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X3Y152_SLICE_X2Y152_BQ),
.I5(CLBLM_R_X7Y154_SLICE_X8Y154_DO5),
.O5(CLBLM_L_X8Y154_SLICE_X10Y154_AO5),
.O6(CLBLM_L_X8Y154_SLICE_X10Y154_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y154_SLICE_X11Y154_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y154_SLICE_X11Y154_DO5),
.O6(CLBLM_L_X8Y154_SLICE_X11Y154_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y154_SLICE_X11Y154_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y154_SLICE_X11Y154_CO5),
.O6(CLBLM_L_X8Y154_SLICE_X11Y154_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y154_SLICE_X11Y154_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y154_SLICE_X11Y154_BO5),
.O6(CLBLM_L_X8Y154_SLICE_X11Y154_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y154_SLICE_X11Y154_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y154_SLICE_X11Y154_AO5),
.O6(CLBLM_L_X8Y154_SLICE_X11Y154_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y141_SLICE_X12Y141_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y141_SLICE_X12Y141_DO5),
.O6(CLBLM_L_X10Y141_SLICE_X12Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y141_SLICE_X12Y141_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y141_SLICE_X12Y141_CO5),
.O6(CLBLM_L_X10Y141_SLICE_X12Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y141_SLICE_X12Y141_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y141_SLICE_X12Y141_BO5),
.O6(CLBLM_L_X10Y141_SLICE_X12Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0200000000000000)
  ) CLBLM_L_X10Y141_SLICE_X12Y141_ALUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(RIOB33_X105Y103_IOB_X1Y103_I),
.I2(RIOB33_X105Y103_IOB_X1Y104_I),
.I3(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I4(RIOB33_X105Y101_IOB_X1Y101_I),
.I5(CLBLM_R_X5Y141_SLICE_X6Y141_AQ),
.O5(CLBLM_L_X10Y141_SLICE_X12Y141_AO5),
.O6(CLBLM_L_X10Y141_SLICE_X12Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y141_SLICE_X13Y141_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y141_SLICE_X13Y141_DO5),
.O6(CLBLM_L_X10Y141_SLICE_X13Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y141_SLICE_X13Y141_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y141_SLICE_X13Y141_CO5),
.O6(CLBLM_L_X10Y141_SLICE_X13Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y141_SLICE_X13Y141_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y141_SLICE_X13Y141_BO5),
.O6(CLBLM_L_X10Y141_SLICE_X13Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y141_SLICE_X13Y141_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y141_SLICE_X13Y141_AO5),
.O6(CLBLM_L_X10Y141_SLICE_X13Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y142_SLICE_X12Y142_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y142_SLICE_X12Y142_AO6),
.Q(CLBLM_L_X10Y142_SLICE_X12Y142_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffeffffffff)
  ) CLBLM_L_X10Y142_SLICE_X12Y142_DLUT (
.I0(CLBLM_R_X11Y146_SLICE_X14Y146_AQ),
.I1(CLBLM_R_X7Y144_SLICE_X8Y144_AQ),
.I2(CLBLM_L_X8Y144_SLICE_X10Y144_B5Q),
.I3(CLBLM_R_X7Y146_SLICE_X9Y146_B5Q),
.I4(CLBLM_L_X8Y144_SLICE_X11Y144_A5Q),
.I5(CLBLM_R_X5Y142_SLICE_X7Y142_C5Q),
.O5(CLBLM_L_X10Y142_SLICE_X12Y142_DO5),
.O6(CLBLM_L_X10Y142_SLICE_X12Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000400000000000)
  ) CLBLM_L_X10Y142_SLICE_X12Y142_CLUT (
.I0(CLBLM_R_X11Y146_SLICE_X14Y146_AQ),
.I1(CLBLM_R_X7Y146_SLICE_X9Y146_B5Q),
.I2(CLBLM_L_X8Y150_SLICE_X10Y150_A5Q),
.I3(CLBLM_L_X10Y142_SLICE_X12Y142_AO5),
.I4(CLBLM_R_X11Y149_SLICE_X14Y149_AQ),
.I5(CLBLM_R_X5Y142_SLICE_X7Y142_C5Q),
.O5(CLBLM_L_X10Y142_SLICE_X12Y142_CO5),
.O6(CLBLM_L_X10Y142_SLICE_X12Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffeffff)
  ) CLBLM_L_X10Y142_SLICE_X12Y142_BLUT (
.I0(CLBLM_L_X8Y144_SLICE_X11Y144_A5Q),
.I1(CLBLM_R_X5Y142_SLICE_X7Y142_C5Q),
.I2(CLBLM_R_X7Y146_SLICE_X9Y146_B5Q),
.I3(CLBLM_R_X7Y144_SLICE_X8Y144_AQ),
.I4(CLBLM_R_X11Y146_SLICE_X14Y146_AQ),
.I5(CLBLM_L_X8Y144_SLICE_X10Y144_B5Q),
.O5(CLBLM_L_X10Y142_SLICE_X12Y142_BO5),
.O6(CLBLM_L_X10Y142_SLICE_X12Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcfc0c000110011)
  ) CLBLM_L_X10Y142_SLICE_X12Y142_ALUT (
.I0(CLBLM_L_X8Y144_SLICE_X11Y144_A5Q),
.I1(CLBLM_R_X7Y144_SLICE_X8Y144_AQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_L_X8Y144_SLICE_X10Y144_B5Q),
.I4(CLBLM_R_X3Y141_SLICE_X3Y141_AO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y142_SLICE_X12Y142_AO5),
.O6(CLBLM_L_X10Y142_SLICE_X12Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y142_SLICE_X13Y142_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y142_SLICE_X13Y142_AO6),
.Q(CLBLM_L_X10Y142_SLICE_X13Y142_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y142_SLICE_X13Y142_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y142_SLICE_X13Y142_DO5),
.O6(CLBLM_L_X10Y142_SLICE_X13Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y142_SLICE_X13Y142_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y142_SLICE_X13Y142_CO5),
.O6(CLBLM_L_X10Y142_SLICE_X13Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0001000000110000)
  ) CLBLM_L_X10Y142_SLICE_X13Y142_BLUT (
.I0(CLBLM_L_X8Y144_SLICE_X11Y144_A5Q),
.I1(CLBLM_L_X8Y144_SLICE_X10Y144_B5Q),
.I2(CLBLM_R_X11Y146_SLICE_X14Y146_AQ),
.I3(CLBLM_R_X7Y144_SLICE_X8Y144_AQ),
.I4(CLBLM_R_X5Y142_SLICE_X7Y142_C5Q),
.I5(CLBLM_R_X7Y146_SLICE_X9Y146_B5Q),
.O5(CLBLM_L_X10Y142_SLICE_X13Y142_BO5),
.O6(CLBLM_L_X10Y142_SLICE_X13Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heeffecfc22332030)
  ) CLBLM_L_X10Y142_SLICE_X13Y142_ALUT (
.I0(CLBLM_L_X8Y142_SLICE_X11Y142_CQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_L_X10Y142_SLICE_X13Y142_AQ),
.I3(CLBLM_R_X5Y149_SLICE_X7Y149_DQ),
.I4(CLBLM_R_X3Y144_SLICE_X2Y144_A5Q),
.I5(CLBLM_L_X10Y147_SLICE_X13Y147_CQ),
.O5(CLBLM_L_X10Y142_SLICE_X13Y142_AO5),
.O6(CLBLM_L_X10Y142_SLICE_X13Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y143_SLICE_X12Y143_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_L_X8Y143_SLICE_X11Y143_AQ),
.Q(CLBLM_L_X10Y143_SLICE_X12Y143_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hafffafffffff55ff)
  ) CLBLM_L_X10Y143_SLICE_X12Y143_DLUT (
.I0(CLBLM_R_X11Y149_SLICE_X14Y149_AQ),
.I1(1'b1),
.I2(CLBLM_L_X8Y142_SLICE_X11Y142_DO6),
.I3(CLBLM_L_X8Y150_SLICE_X10Y150_A5Q),
.I4(CLBLM_L_X10Y142_SLICE_X12Y142_BO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y143_SLICE_X12Y143_DO5),
.O6(CLBLM_L_X10Y143_SLICE_X12Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffbbffbbccccf0f0)
  ) CLBLM_L_X10Y143_SLICE_X12Y143_CLUT (
.I0(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.I1(CLBLM_L_X8Y142_SLICE_X11Y142_AQ),
.I2(CLBLM_L_X10Y149_SLICE_X12Y149_B5Q),
.I3(CLBLM_L_X8Y142_SLICE_X11Y142_BQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y143_SLICE_X12Y143_CO5),
.O6(CLBLM_L_X10Y143_SLICE_X12Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefffeffefffefff)
  ) CLBLM_L_X10Y143_SLICE_X12Y143_BLUT (
.I0(CLBLM_L_X8Y150_SLICE_X10Y150_A5Q),
.I1(CLBLM_L_X12Y149_SLICE_X16Y149_CO6),
.I2(CLBLM_R_X11Y149_SLICE_X14Y149_AQ),
.I3(CLBLM_L_X8Y142_SLICE_X11Y142_DO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y143_SLICE_X12Y143_BO5),
.O6(CLBLM_L_X10Y143_SLICE_X12Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffefffefbfbfbfb)
  ) CLBLM_L_X10Y143_SLICE_X12Y143_ALUT (
.I0(CLBLM_L_X10Y142_SLICE_X12Y142_BO6),
.I1(CLBLM_L_X8Y150_SLICE_X10Y150_A5Q),
.I2(CLBLM_R_X11Y149_SLICE_X14Y149_AQ),
.I3(CLBLM_L_X12Y149_SLICE_X16Y149_CO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y143_SLICE_X12Y143_AO5),
.O6(CLBLM_L_X10Y143_SLICE_X12Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'heac0aa00c0c00000)
  ) CLBLM_L_X10Y143_SLICE_X13Y143_DLUT (
.I0(RIOB33_X105Y135_IOB_X1Y135_I),
.I1(CLBLM_R_X11Y142_SLICE_X14Y142_CO6),
.I2(LIOB33_X0Y51_IOB_X0Y51_I),
.I3(CLBLM_R_X11Y142_SLICE_X14Y142_DO6),
.I4(CLBLM_R_X11Y142_SLICE_X14Y142_BO5),
.I5(CLBLM_L_X10Y148_SLICE_X13Y148_BO6),
.O5(CLBLM_L_X10Y143_SLICE_X13Y143_DO5),
.O6(CLBLM_L_X10Y143_SLICE_X13Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffecffffffa0)
  ) CLBLM_L_X10Y143_SLICE_X13Y143_CLUT (
.I0(CLBLM_R_X5Y142_SLICE_X6Y142_DQ),
.I1(LIOB33_X0Y51_IOB_X0Y52_I),
.I2(CLBLM_R_X11Y145_SLICE_X15Y145_BO5),
.I3(CLBLM_L_X10Y146_SLICE_X13Y146_BO6),
.I4(CLBLM_L_X10Y146_SLICE_X13Y146_BO5),
.I5(CLBLM_R_X11Y142_SLICE_X14Y142_CO5),
.O5(CLBLM_L_X10Y143_SLICE_X13Y143_CO5),
.O6(CLBLM_L_X10Y143_SLICE_X13Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf888f00088880000)
  ) CLBLM_L_X10Y143_SLICE_X13Y143_BLUT (
.I0(CLBLM_R_X11Y142_SLICE_X14Y142_DO6),
.I1(CLBLM_L_X8Y144_SLICE_X10Y144_CO6),
.I2(CLBLM_R_X11Y142_SLICE_X14Y142_BO5),
.I3(LIOB33_X0Y53_IOB_X0Y53_I),
.I4(CLBLM_L_X10Y143_SLICE_X12Y143_AQ),
.I5(CLBLM_R_X11Y142_SLICE_X14Y142_CO6),
.O5(CLBLM_L_X10Y143_SLICE_X13Y143_BO5),
.O6(CLBLM_L_X10Y143_SLICE_X13Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000010000000000)
  ) CLBLM_L_X10Y143_SLICE_X13Y143_ALUT (
.I0(CLBLM_R_X5Y142_SLICE_X7Y142_C5Q),
.I1(CLBLM_R_X7Y144_SLICE_X8Y144_AQ),
.I2(CLBLM_L_X8Y144_SLICE_X10Y144_B5Q),
.I3(CLBLM_R_X11Y146_SLICE_X14Y146_AQ),
.I4(CLBLM_L_X8Y144_SLICE_X11Y144_A5Q),
.I5(CLBLM_R_X7Y146_SLICE_X9Y146_B5Q),
.O5(CLBLM_L_X10Y143_SLICE_X13Y143_AO5),
.O6(CLBLM_L_X10Y143_SLICE_X13Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ffaa0000fffe)
  ) CLBLM_L_X10Y144_SLICE_X12Y144_DLUT (
.I0(CLBLM_L_X10Y144_SLICE_X12Y144_AO5),
.I1(CLBLM_L_X10Y143_SLICE_X13Y143_CO6),
.I2(CLBLM_L_X10Y144_SLICE_X13Y144_BO6),
.I3(CLBLM_L_X10Y144_SLICE_X12Y144_CO6),
.I4(CLBLM_R_X11Y143_SLICE_X14Y143_CO5),
.I5(CLBLM_L_X10Y142_SLICE_X13Y142_BO6),
.O5(CLBLM_L_X10Y144_SLICE_X12Y144_DO5),
.O6(CLBLM_L_X10Y144_SLICE_X12Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa08000008080000)
  ) CLBLM_L_X10Y144_SLICE_X12Y144_CLUT (
.I0(CLBLM_L_X8Y150_SLICE_X10Y150_A5Q),
.I1(CLBLM_L_X10Y148_SLICE_X12Y148_AQ),
.I2(CLBLM_L_X10Y142_SLICE_X12Y142_DO6),
.I3(CLBLM_R_X3Y144_SLICE_X3Y144_DQ),
.I4(CLBLM_R_X11Y149_SLICE_X14Y149_AQ),
.I5(CLBLM_R_X11Y142_SLICE_X14Y142_BO6),
.O5(CLBLM_L_X10Y144_SLICE_X12Y144_CO5),
.O6(CLBLM_L_X10Y144_SLICE_X12Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0c0c5d0c0c0c0c0c)
  ) CLBLM_L_X10Y144_SLICE_X12Y144_BLUT (
.I0(CLBLM_L_X10Y142_SLICE_X12Y142_DO6),
.I1(CLBLM_R_X7Y142_SLICE_X9Y142_A5Q),
.I2(CLBLM_L_X10Y144_SLICE_X13Y144_AO6),
.I3(CLBLM_R_X11Y149_SLICE_X14Y149_AQ),
.I4(CLBLM_L_X8Y150_SLICE_X10Y150_A5Q),
.I5(CLBLL_L_X4Y144_SLICE_X5Y144_DQ),
.O5(CLBLM_L_X10Y144_SLICE_X12Y144_BO5),
.O6(CLBLM_L_X10Y144_SLICE_X12Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafaffff30000000)
  ) CLBLM_L_X10Y144_SLICE_X12Y144_ALUT (
.I0(CLBLM_L_X10Y142_SLICE_X12Y142_DO6),
.I1(CLBLM_L_X12Y143_SLICE_X16Y143_AO6),
.I2(CLBLM_R_X11Y149_SLICE_X14Y149_AQ),
.I3(CLBLM_R_X7Y142_SLICE_X9Y142_DQ),
.I4(CLBLM_L_X8Y150_SLICE_X10Y150_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X10Y144_SLICE_X12Y144_AO5),
.O6(CLBLM_L_X10Y144_SLICE_X12Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f5fcfcfcfd)
  ) CLBLM_L_X10Y144_SLICE_X13Y144_DLUT (
.I0(CLBLM_R_X11Y145_SLICE_X15Y145_BO5),
.I1(CLBLM_L_X8Y143_SLICE_X10Y143_DQ),
.I2(CLBLM_L_X10Y143_SLICE_X13Y143_DO6),
.I3(CLBLM_R_X11Y144_SLICE_X15Y144_AO5),
.I4(CLBLM_R_X11Y143_SLICE_X15Y143_DO6),
.I5(CLBLM_R_X11Y144_SLICE_X15Y144_CO6),
.O5(CLBLM_L_X10Y144_SLICE_X13Y144_DO5),
.O6(CLBLM_L_X10Y144_SLICE_X13Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000001)
  ) CLBLM_L_X10Y144_SLICE_X13Y144_CLUT (
.I0(CLBLM_R_X5Y142_SLICE_X7Y142_C5Q),
.I1(CLBLM_R_X11Y146_SLICE_X14Y146_AQ),
.I2(CLBLM_L_X8Y144_SLICE_X10Y144_B5Q),
.I3(CLBLM_L_X8Y144_SLICE_X11Y144_A5Q),
.I4(CLBLM_R_X7Y146_SLICE_X9Y146_B5Q),
.I5(CLBLM_R_X7Y144_SLICE_X8Y144_AQ),
.O5(CLBLM_L_X10Y144_SLICE_X13Y144_CO5),
.O6(CLBLM_L_X10Y144_SLICE_X13Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff3300ffff3705)
  ) CLBLM_L_X10Y144_SLICE_X13Y144_BLUT (
.I0(CLBLM_R_X11Y144_SLICE_X15Y144_AO5),
.I1(CLBLM_R_X11Y144_SLICE_X15Y144_CO6),
.I2(CLBLM_R_X11Y145_SLICE_X15Y145_BO5),
.I3(CLBLM_R_X5Y140_SLICE_X7Y140_AQ),
.I4(CLBLM_L_X12Y144_SLICE_X16Y144_AO5),
.I5(CLBLM_R_X11Y143_SLICE_X15Y143_DO6),
.O5(CLBLM_L_X10Y144_SLICE_X13Y144_BO5),
.O6(CLBLM_L_X10Y144_SLICE_X13Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffefffffffffff)
  ) CLBLM_L_X10Y144_SLICE_X13Y144_ALUT (
.I0(CLBLM_L_X8Y144_SLICE_X10Y144_B5Q),
.I1(CLBLM_R_X7Y144_SLICE_X8Y144_AQ),
.I2(CLBLM_R_X11Y146_SLICE_X14Y146_AQ),
.I3(CLBLM_R_X5Y142_SLICE_X7Y142_C5Q),
.I4(CLBLM_L_X8Y144_SLICE_X11Y144_A5Q),
.I5(CLBLM_L_X8Y144_SLICE_X10Y144_CO6),
.O5(CLBLM_L_X10Y144_SLICE_X13Y144_AO5),
.O6(CLBLM_L_X10Y144_SLICE_X13Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y145_SLICE_X12Y145_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_R_X7Y148_SLICE_X9Y148_BQ),
.Q(CLBLM_L_X10Y145_SLICE_X12Y145_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff5f0f5500)
  ) CLBLM_L_X10Y145_SLICE_X12Y145_DLUT (
.I0(CLBLM_L_X10Y143_SLICE_X12Y143_DO5),
.I1(1'b1),
.I2(CLBLM_L_X10Y143_SLICE_X12Y143_DO6),
.I3(CLBLM_L_X8Y141_SLICE_X10Y141_CQ),
.I4(CLBLM_R_X5Y153_SLICE_X6Y153_DQ),
.I5(CLBLM_L_X10Y148_SLICE_X12Y148_BO6),
.O5(CLBLM_L_X10Y145_SLICE_X12Y145_DO5),
.O6(CLBLM_L_X10Y145_SLICE_X12Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5fff0fff5f5f0f0)
  ) CLBLM_L_X10Y145_SLICE_X12Y145_CLUT (
.I0(CLBLM_L_X10Y143_SLICE_X12Y143_AO6),
.I1(1'b1),
.I2(CLBLM_L_X10Y146_SLICE_X12Y146_DO6),
.I3(CLBLM_L_X8Y148_SLICE_X10Y148_CO6),
.I4(CLBLM_R_X7Y145_SLICE_X9Y145_CQ),
.I5(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.O5(CLBLM_L_X10Y145_SLICE_X12Y145_CO5),
.O6(CLBLM_L_X10Y145_SLICE_X12Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_L_X10Y145_SLICE_X12Y145_BLUT (
.I0(CLBLM_L_X10Y148_SLICE_X12Y148_CO6),
.I1(CLBLM_L_X8Y145_SLICE_X11Y145_BO6),
.I2(CLBLM_L_X8Y145_SLICE_X10Y145_CO6),
.I3(CLBLM_L_X10Y144_SLICE_X12Y144_DO6),
.I4(CLBLM_L_X10Y145_SLICE_X12Y145_CO6),
.I5(CLBLM_L_X10Y145_SLICE_X12Y145_AO5),
.O5(CLBLM_L_X10Y145_SLICE_X12Y145_BO5),
.O6(CLBLM_L_X10Y145_SLICE_X12Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffffff00000050)
  ) CLBLM_L_X10Y145_SLICE_X12Y145_ALUT (
.I0(CLBLM_L_X10Y142_SLICE_X12Y142_DO6),
.I1(1'b1),
.I2(CLBLM_R_X5Y146_SLICE_X6Y146_AQ),
.I3(CLBLM_L_X8Y150_SLICE_X10Y150_A5Q),
.I4(CLBLM_R_X11Y149_SLICE_X14Y149_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y145_SLICE_X12Y145_AO5),
.O6(CLBLM_L_X10Y145_SLICE_X12Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaaffaaffaaba)
  ) CLBLM_L_X10Y145_SLICE_X13Y145_DLUT (
.I0(CLBLM_R_X7Y147_SLICE_X9Y147_DO5),
.I1(CLBLM_L_X10Y142_SLICE_X13Y142_BO6),
.I2(CLBLM_L_X10Y144_SLICE_X13Y144_DO6),
.I3(CLBLM_R_X11Y143_SLICE_X14Y143_CO5),
.I4(CLBLM_L_X10Y145_SLICE_X13Y145_BO5),
.I5(CLBLM_R_X11Y145_SLICE_X14Y145_AO5),
.O5(CLBLM_L_X10Y145_SLICE_X13Y145_DO5),
.O6(CLBLM_L_X10Y145_SLICE_X13Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffafffafe)
  ) CLBLM_L_X10Y145_SLICE_X13Y145_CLUT (
.I0(CLBLM_L_X8Y145_SLICE_X11Y145_AO6),
.I1(CLBLM_L_X10Y146_SLICE_X13Y146_CO6),
.I2(CLBLM_L_X10Y145_SLICE_X12Y145_DO6),
.I3(CLBLM_R_X11Y143_SLICE_X14Y143_CO5),
.I4(CLBLM_R_X11Y145_SLICE_X14Y145_CO6),
.I5(CLBLM_R_X7Y146_SLICE_X8Y146_BO6),
.O5(CLBLM_L_X10Y145_SLICE_X13Y145_CO5),
.O6(CLBLM_L_X10Y145_SLICE_X13Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0aff0a0a0c0c0c0c)
  ) CLBLM_L_X10Y145_SLICE_X13Y145_BLUT (
.I0(CLBLM_L_X10Y147_SLICE_X13Y147_B5Q),
.I1(CLBLL_L_X4Y141_SLICE_X5Y141_AQ),
.I2(CLBLM_L_X10Y145_SLICE_X12Y145_AO6),
.I3(CLBLM_L_X10Y144_SLICE_X13Y144_AO6),
.I4(CLBLM_R_X3Y142_SLICE_X2Y142_BQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y145_SLICE_X13Y145_BO5),
.O6(CLBLM_L_X10Y145_SLICE_X13Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c05050ff50)
  ) CLBLM_L_X10Y145_SLICE_X13Y145_ALUT (
.I0(CLBLM_R_X11Y145_SLICE_X14Y145_BO5),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_L_X8Y144_SLICE_X10Y144_BQ),
.I3(CLBLM_R_X5Y145_SLICE_X6Y145_BQ),
.I4(CLBLM_L_X10Y144_SLICE_X13Y144_AO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y145_SLICE_X13Y145_AO5),
.O6(CLBLM_L_X10Y145_SLICE_X13Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y146_SLICE_X12Y146_A_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y145_SLICE_X15Y145_AO6),
.Q(CLBLM_L_X10Y146_SLICE_X12Y146_AQ),
.S(CLBLM_R_X11Y148_SLICE_X14Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8888888f88888888)
  ) CLBLM_L_X10Y146_SLICE_X12Y146_DLUT (
.I0(CLBLM_L_X10Y142_SLICE_X12Y142_CO6),
.I1(CLBLM_L_X10Y147_SLICE_X12Y147_CQ),
.I2(CLBLM_R_X11Y143_SLICE_X14Y143_CO5),
.I3(CLBLM_R_X11Y144_SLICE_X15Y144_CO6),
.I4(CLBLM_R_X7Y146_SLICE_X9Y146_B5Q),
.I5(CLBLM_L_X10Y150_SLICE_X13Y150_A5Q),
.O5(CLBLM_L_X10Y146_SLICE_X12Y146_DO5),
.O6(CLBLM_L_X10Y146_SLICE_X12Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00f000f000aa00aa)
  ) CLBLM_L_X10Y146_SLICE_X12Y146_CLUT (
.I0(CLBLM_R_X5Y142_SLICE_X6Y142_BQ),
.I1(1'b1),
.I2(CLBLM_R_X5Y146_SLICE_X7Y146_DQ),
.I3(CLBLM_R_X11Y144_SLICE_X15Y144_CO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y146_SLICE_X12Y146_CO5),
.O6(CLBLM_L_X10Y146_SLICE_X12Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7bde7bdef0f00000)
  ) CLBLM_L_X10Y146_SLICE_X12Y146_BLUT (
.I0(CLBLL_L_X4Y147_SLICE_X4Y147_BQ),
.I1(CLBLL_L_X4Y150_SLICE_X5Y150_BQ),
.I2(CLBLM_L_X10Y148_SLICE_X13Y148_AQ),
.I3(CLBLM_L_X10Y147_SLICE_X12Y147_CQ),
.I4(CLBLM_L_X10Y142_SLICE_X12Y142_CO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y146_SLICE_X12Y146_BO5),
.O6(CLBLM_L_X10Y146_SLICE_X12Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc5cacaca55ffffff)
  ) CLBLM_L_X10Y146_SLICE_X12Y146_ALUT (
.I0(CLBLM_L_X10Y149_SLICE_X12Y149_A5Q),
.I1(CLBLM_L_X10Y147_SLICE_X12Y147_B5Q),
.I2(CLBLM_L_X8Y149_SLICE_X11Y149_BQ),
.I3(CLBLM_R_X5Y146_SLICE_X7Y146_AQ),
.I4(CLBLM_R_X11Y146_SLICE_X15Y146_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y146_SLICE_X12Y146_AO5),
.O6(CLBLM_L_X10Y146_SLICE_X12Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y146_SLICE_X13Y146_A_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y146_SLICE_X13Y146_AO6),
.Q(CLBLM_L_X10Y146_SLICE_X13Y146_AQ),
.S(CLBLM_R_X11Y148_SLICE_X15Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8888000c00000000)
  ) CLBLM_L_X10Y146_SLICE_X13Y146_DLUT (
.I0(CLBLM_R_X3Y146_SLICE_X3Y146_C5Q),
.I1(CLBLM_R_X11Y142_SLICE_X14Y142_BO6),
.I2(CLBLM_L_X8Y152_SLICE_X11Y152_AQ),
.I3(CLBLM_R_X7Y146_SLICE_X9Y146_B5Q),
.I4(CLBLM_R_X11Y149_SLICE_X14Y149_AQ),
.I5(CLBLM_L_X8Y150_SLICE_X10Y150_A5Q),
.O5(CLBLM_L_X10Y146_SLICE_X13Y146_DO5),
.O6(CLBLM_L_X10Y146_SLICE_X13Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffff5554)
  ) CLBLM_L_X10Y146_SLICE_X13Y146_CLUT (
.I0(CLBLM_L_X10Y142_SLICE_X13Y142_BO6),
.I1(CLBLM_L_X10Y146_SLICE_X12Y146_CO6),
.I2(CLBLM_R_X11Y146_SLICE_X15Y146_CO6),
.I3(CLBLM_R_X11Y144_SLICE_X14Y144_CO6),
.I4(CLBLM_R_X11Y147_SLICE_X15Y147_DO6),
.I5(CLBLM_L_X10Y146_SLICE_X13Y146_DO6),
.O5(CLBLM_L_X10Y146_SLICE_X13Y146_CO5),
.O6(CLBLM_L_X10Y146_SLICE_X13Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha000000044000000)
  ) CLBLM_L_X10Y146_SLICE_X13Y146_BLUT (
.I0(CLBLM_R_X11Y149_SLICE_X14Y149_AQ),
.I1(CLBLM_R_X5Y151_SLICE_X6Y151_BQ),
.I2(CLBLM_R_X11Y145_SLICE_X14Y145_BQ),
.I3(CLBLM_R_X11Y142_SLICE_X14Y142_DO6),
.I4(CLBLM_L_X8Y150_SLICE_X10Y150_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X10Y146_SLICE_X13Y146_BO5),
.O6(CLBLM_L_X10Y146_SLICE_X13Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00cc00cc00)
  ) CLBLM_L_X10Y146_SLICE_X13Y146_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(1'b1),
.I3(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y146_SLICE_X13Y146_AO5),
.O6(CLBLM_L_X10Y146_SLICE_X13Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y147_SLICE_X12Y147_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y147_SLICE_X12Y147_BO5),
.Q(CLBLM_L_X10Y147_SLICE_X12Y147_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y147_SLICE_X12Y147_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y147_SLICE_X12Y147_CO5),
.Q(CLBLM_L_X10Y147_SLICE_X12Y147_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y147_SLICE_X12Y147_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y147_SLICE_X12Y147_AO6),
.Q(CLBLM_L_X10Y147_SLICE_X12Y147_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y147_SLICE_X12Y147_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y147_SLICE_X12Y147_BO6),
.Q(CLBLM_L_X10Y147_SLICE_X12Y147_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y147_SLICE_X12Y147_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y147_SLICE_X12Y147_CO6),
.Q(CLBLM_L_X10Y147_SLICE_X12Y147_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0011000030303030)
  ) CLBLM_L_X10Y147_SLICE_X12Y147_DLUT (
.I0(CLBLM_R_X7Y146_SLICE_X9Y146_B5Q),
.I1(CLBLM_R_X11Y144_SLICE_X15Y144_CO6),
.I2(CLBLM_R_X7Y147_SLICE_X8Y147_BQ),
.I3(CLBLM_R_X11Y143_SLICE_X14Y143_CO5),
.I4(CLBLM_L_X10Y150_SLICE_X13Y150_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y147_SLICE_X12Y147_DO5),
.O6(CLBLM_L_X10Y147_SLICE_X12Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0aaf0aaffaa00aa)
  ) CLBLM_L_X10Y147_SLICE_X12Y147_CLUT (
.I0(CLBLM_L_X10Y150_SLICE_X13Y150_A5Q),
.I1(1'b1),
.I2(CLBLL_L_X4Y148_SLICE_X4Y148_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X11Y148_SLICE_X14Y148_DQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y147_SLICE_X12Y147_CO5),
.O6(CLBLM_L_X10Y147_SLICE_X12Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fff000ccaaccaa)
  ) CLBLM_L_X10Y147_SLICE_X12Y147_BLUT (
.I0(CLBLM_L_X10Y148_SLICE_X12Y148_A5Q),
.I1(CLBLM_L_X10Y147_SLICE_X12Y147_BQ),
.I2(CLBLM_R_X3Y151_SLICE_X3Y151_C5Q),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X8Y148_SLICE_X10Y148_BQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y147_SLICE_X12Y147_BO5),
.O6(CLBLM_L_X10Y147_SLICE_X12Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaafc30fc30)
  ) CLBLM_L_X10Y147_SLICE_X12Y147_ALUT (
.I0(CLBLM_L_X10Y147_SLICE_X12Y147_B5Q),
.I1(CLBLM_R_X11Y145_SLICE_X15Y145_BO5),
.I2(CLBLM_L_X10Y147_SLICE_X12Y147_AQ),
.I3(CLBLM_R_X7Y141_SLICE_X8Y141_AQ),
.I4(1'b1),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_L_X10Y147_SLICE_X12Y147_AO5),
.O6(CLBLM_L_X10Y147_SLICE_X12Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y147_SLICE_X13Y147_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y147_SLICE_X13Y147_AO5),
.Q(CLBLM_L_X10Y147_SLICE_X13Y147_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y147_SLICE_X13Y147_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y147_SLICE_X13Y147_BO5),
.Q(CLBLM_L_X10Y147_SLICE_X13Y147_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y147_SLICE_X13Y147_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y147_SLICE_X13Y147_AO6),
.Q(CLBLM_L_X10Y147_SLICE_X13Y147_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y147_SLICE_X13Y147_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y147_SLICE_X13Y147_BO6),
.Q(CLBLM_L_X10Y147_SLICE_X13Y147_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y147_SLICE_X13Y147_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y147_SLICE_X13Y147_CO6),
.Q(CLBLM_L_X10Y147_SLICE_X13Y147_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y147_SLICE_X13Y147_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y147_SLICE_X13Y147_DO6),
.Q(CLBLM_L_X10Y147_SLICE_X13Y147_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffddfcdc33113010)
  ) CLBLM_L_X10Y147_SLICE_X13Y147_DLUT (
.I0(CLBLM_R_X5Y149_SLICE_X7Y149_DQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_L_X10Y147_SLICE_X13Y147_DQ),
.I3(CLBLM_L_X8Y142_SLICE_X11Y142_CQ),
.I4(CLBLM_L_X8Y151_SLICE_X11Y151_AQ),
.I5(CLBLM_R_X3Y151_SLICE_X3Y151_D5Q),
.O5(CLBLM_L_X10Y147_SLICE_X13Y147_DO5),
.O6(CLBLM_L_X10Y147_SLICE_X13Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0ffcc5544)
  ) CLBLM_L_X10Y147_SLICE_X13Y147_CLUT (
.I0(CLBLM_R_X5Y149_SLICE_X7Y149_DQ),
.I1(CLBLM_L_X10Y147_SLICE_X13Y147_CQ),
.I2(CLBLM_L_X8Y151_SLICE_X11Y151_AQ),
.I3(CLBLM_L_X8Y147_SLICE_X10Y147_AQ),
.I4(CLBLM_L_X8Y142_SLICE_X11Y142_CQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_L_X10Y147_SLICE_X13Y147_CO5),
.O6(CLBLM_L_X10Y147_SLICE_X13Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f3c0c0bbbb8888)
  ) CLBLM_L_X10Y147_SLICE_X13Y147_BLUT (
.I0(CLBLM_R_X7Y147_SLICE_X8Y147_CQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLL_L_X4Y144_SLICE_X5Y144_BQ),
.I3(1'b1),
.I4(CLBLM_L_X10Y150_SLICE_X13Y150_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y147_SLICE_X13Y147_BO5),
.O6(CLBLM_L_X10Y147_SLICE_X13Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd88dd88f5f5a0a0)
  ) CLBLM_L_X10Y147_SLICE_X13Y147_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLL_L_X4Y147_SLICE_X4Y147_D5Q),
.I2(CLBLM_R_X5Y145_SLICE_X7Y145_AQ),
.I3(CLBLM_L_X8Y147_SLICE_X11Y147_BO6),
.I4(CLBLM_R_X11Y147_SLICE_X14Y147_BO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y147_SLICE_X13Y147_AO5),
.O6(CLBLM_L_X10Y147_SLICE_X13Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y148_SLICE_X12Y148_A5_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y148_SLICE_X12Y148_AO5),
.Q(CLBLM_L_X10Y148_SLICE_X12Y148_A5Q),
.S(CLBLM_R_X11Y148_SLICE_X14Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y148_SLICE_X12Y148_A_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y148_SLICE_X12Y148_AO6),
.Q(CLBLM_L_X10Y148_SLICE_X12Y148_AQ),
.S(CLBLM_R_X11Y148_SLICE_X14Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3030ff303030ff30)
  ) CLBLM_L_X10Y148_SLICE_X12Y148_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y143_SLICE_X12Y143_BO5),
.I2(CLBLM_L_X8Y152_SLICE_X10Y152_BQ),
.I3(CLBLM_L_X10Y148_SLICE_X12Y148_A5Q),
.I4(CLBLM_L_X10Y148_SLICE_X12Y148_BO5),
.I5(1'b1),
.O5(CLBLM_L_X10Y148_SLICE_X12Y148_DO5),
.O6(CLBLM_L_X10Y148_SLICE_X12Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffff5fdfffff0fc)
  ) CLBLM_L_X10Y148_SLICE_X12Y148_CLUT (
.I0(CLBLM_L_X10Y143_SLICE_X12Y143_BO6),
.I1(CLBLM_R_X7Y151_SLICE_X8Y151_CQ),
.I2(CLBLM_L_X10Y148_SLICE_X13Y148_DO6),
.I3(CLBLM_L_X10Y144_SLICE_X12Y144_AO6),
.I4(CLBLM_L_X10Y148_SLICE_X12Y148_DO6),
.I5(CLBLM_L_X8Y149_SLICE_X11Y149_AQ),
.O5(CLBLM_L_X10Y148_SLICE_X12Y148_CO5),
.O6(CLBLM_L_X10Y148_SLICE_X12Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h880080807777ffff)
  ) CLBLM_L_X10Y148_SLICE_X12Y148_BLUT (
.I0(CLBLM_L_X10Y144_SLICE_X13Y144_CO6),
.I1(CLBLM_L_X8Y150_SLICE_X10Y150_A5Q),
.I2(CLBLM_R_X7Y147_SLICE_X9Y147_C5Q),
.I3(CLBLM_R_X5Y147_SLICE_X7Y147_CQ),
.I4(CLBLM_R_X11Y149_SLICE_X14Y149_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y148_SLICE_X12Y148_BO5),
.O6(CLBLM_L_X10Y148_SLICE_X12Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa0088888888)
  ) CLBLM_L_X10Y148_SLICE_X12Y148_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X8Y148_SLICE_X10Y148_BQ),
.I2(1'b1),
.I3(CLBLM_L_X8Y147_SLICE_X10Y147_A5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y148_SLICE_X12Y148_AO5),
.O6(CLBLM_L_X10Y148_SLICE_X12Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y148_SLICE_X13Y148_A_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y150_SLICE_X13Y150_DO6),
.Q(CLBLM_L_X10Y148_SLICE_X13Y148_AQ),
.S(CLBLM_R_X11Y148_SLICE_X15Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3022002230000000)
  ) CLBLM_L_X10Y148_SLICE_X13Y148_DLUT (
.I0(CLBLM_L_X10Y147_SLICE_X12Y147_C5Q),
.I1(CLBLM_L_X8Y150_SLICE_X10Y150_A5Q),
.I2(CLBLM_L_X10Y144_SLICE_X13Y144_CO6),
.I3(CLBLM_R_X11Y149_SLICE_X14Y149_AQ),
.I4(CLBLM_L_X10Y150_SLICE_X13Y150_B5Q),
.I5(CLBLM_L_X10Y143_SLICE_X13Y143_AO6),
.O5(CLBLM_L_X10Y148_SLICE_X13Y148_DO5),
.O6(CLBLM_L_X10Y148_SLICE_X13Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_L_X10Y148_SLICE_X13Y148_CLUT (
.I0(CLBLM_L_X10Y148_SLICE_X13Y148_AO6),
.I1(CLBLM_L_X8Y149_SLICE_X11Y149_DO6),
.I2(CLBLM_L_X10Y149_SLICE_X13Y149_DO6),
.I3(CLBLM_L_X8Y145_SLICE_X10Y145_BO5),
.I4(CLBLM_R_X11Y144_SLICE_X15Y144_BO6),
.I5(CLBLM_R_X5Y148_SLICE_X7Y148_CO6),
.O5(CLBLM_L_X10Y148_SLICE_X13Y148_CO5),
.O6(CLBLM_L_X10Y148_SLICE_X13Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5500550050440000)
  ) CLBLM_L_X10Y148_SLICE_X13Y148_BLUT (
.I0(CLBLM_R_X11Y149_SLICE_X14Y149_AQ),
.I1(CLBLM_L_X10Y147_SLICE_X13Y147_BQ),
.I2(CLBLM_L_X10Y146_SLICE_X12Y146_AQ),
.I3(CLBLM_L_X8Y150_SLICE_X10Y150_A5Q),
.I4(CLBLM_L_X10Y143_SLICE_X13Y143_AO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y148_SLICE_X13Y148_BO5),
.O6(CLBLM_L_X10Y148_SLICE_X13Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000f0f00000)
  ) CLBLM_L_X10Y148_SLICE_X13Y148_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_L_X10Y143_SLICE_X12Y143_AO6),
.I3(CLBLM_R_X5Y146_SLICE_X7Y146_CQ),
.I4(CLBLM_L_X8Y148_SLICE_X11Y148_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y148_SLICE_X13Y148_AO5),
.O6(CLBLM_L_X10Y148_SLICE_X13Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y149_SLICE_X12Y149_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y149_SLICE_X12Y149_AO5),
.Q(CLBLM_L_X10Y149_SLICE_X12Y149_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y149_SLICE_X12Y149_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y149_SLICE_X12Y149_BO5),
.Q(CLBLM_L_X10Y149_SLICE_X12Y149_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y149_SLICE_X12Y149_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y149_SLICE_X12Y149_AO6),
.Q(CLBLM_L_X10Y149_SLICE_X12Y149_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y149_SLICE_X12Y149_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y149_SLICE_X12Y149_BO6),
.Q(CLBLM_L_X10Y149_SLICE_X12Y149_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y149_SLICE_X12Y149_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y149_SLICE_X12Y149_CO6),
.Q(CLBLM_L_X10Y149_SLICE_X12Y149_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y149_SLICE_X12Y149_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y149_SLICE_X12Y149_DO6),
.Q(CLBLM_L_X10Y149_SLICE_X12Y149_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaafc30fc30)
  ) CLBLM_L_X10Y149_SLICE_X12Y149_DLUT (
.I0(CLBLM_L_X8Y149_SLICE_X11Y149_AQ),
.I1(CLBLM_L_X10Y143_SLICE_X12Y143_AO6),
.I2(CLBLM_L_X10Y149_SLICE_X12Y149_DQ),
.I3(CLBLM_R_X5Y149_SLICE_X7Y149_AQ),
.I4(1'b1),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_L_X10Y149_SLICE_X12Y149_DO5),
.O6(CLBLM_L_X10Y149_SLICE_X12Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffee00eeff440044)
  ) CLBLM_L_X10Y149_SLICE_X12Y149_CLUT (
.I0(CLBLM_L_X10Y143_SLICE_X12Y143_AO6),
.I1(CLBLM_L_X10Y149_SLICE_X12Y149_CQ),
.I2(1'b1),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X10Y149_SLICE_X13Y149_A5Q),
.I5(CLBLM_L_X8Y150_SLICE_X11Y150_AQ),
.O5(CLBLM_L_X10Y149_SLICE_X12Y149_CO5),
.O6(CLBLM_L_X10Y149_SLICE_X12Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafa0a0afc0cfc0c)
  ) CLBLM_L_X10Y149_SLICE_X12Y149_BLUT (
.I0(CLBLM_R_X11Y151_SLICE_X15Y151_A5Q),
.I1(CLBLM_L_X8Y148_SLICE_X11Y148_C5Q),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_L_X10Y150_SLICE_X13Y150_CQ),
.I4(CLBLL_L_X4Y143_SLICE_X4Y143_CQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y149_SLICE_X12Y149_BO5),
.O6(CLBLM_L_X10Y149_SLICE_X12Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccaaccaaaaf0aaf0)
  ) CLBLM_L_X10Y149_SLICE_X12Y149_ALUT (
.I0(CLBLM_L_X10Y150_SLICE_X13Y150_C5Q),
.I1(CLBLM_L_X10Y148_SLICE_X12Y148_A5Q),
.I2(CLBLM_L_X10Y146_SLICE_X12Y146_AO6),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y149_SLICE_X12Y149_AO5),
.O6(CLBLM_L_X10Y149_SLICE_X12Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y149_SLICE_X13Y149_A5_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y149_SLICE_X9Y149_AO6),
.Q(CLBLM_L_X10Y149_SLICE_X13Y149_A5Q),
.S(CLBLM_R_X11Y148_SLICE_X15Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y149_SLICE_X13Y149_A_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y149_SLICE_X13Y149_AO6),
.Q(CLBLM_L_X10Y149_SLICE_X13Y149_AQ),
.S(CLBLM_R_X11Y148_SLICE_X15Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000f0a05000)
  ) CLBLM_L_X10Y149_SLICE_X13Y149_DLUT (
.I0(CLBLM_L_X8Y150_SLICE_X10Y150_A5Q),
.I1(1'b1),
.I2(CLBLM_L_X10Y143_SLICE_X13Y143_AO6),
.I3(CLBLM_L_X10Y149_SLICE_X13Y149_A5Q),
.I4(CLBLM_L_X10Y149_SLICE_X13Y149_AQ),
.I5(CLBLM_R_X11Y149_SLICE_X14Y149_AQ),
.O5(CLBLM_L_X10Y149_SLICE_X13Y149_DO5),
.O6(CLBLM_L_X10Y149_SLICE_X13Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_L_X10Y149_SLICE_X13Y149_CLUT (
.I0(CLBLM_L_X8Y150_SLICE_X10Y150_BO6),
.I1(CLBLM_L_X10Y148_SLICE_X13Y148_AO5),
.I2(CLBLM_L_X10Y147_SLICE_X12Y147_DO6),
.I3(CLBLM_L_X8Y150_SLICE_X10Y150_DO6),
.I4(CLBLM_L_X10Y148_SLICE_X13Y148_BO5),
.I5(CLBLM_R_X11Y144_SLICE_X14Y144_BO6),
.O5(CLBLM_L_X10Y149_SLICE_X13Y149_CO5),
.O6(CLBLM_L_X10Y149_SLICE_X13Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0000bb88bb88)
  ) CLBLM_L_X10Y149_SLICE_X13Y149_BLUT (
.I0(CLBLM_R_X7Y148_SLICE_X9Y148_B5Q),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(1'b1),
.I3(CLBLM_R_X11Y149_SLICE_X15Y149_AQ),
.I4(CLBLM_R_X3Y152_SLICE_X3Y152_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X10Y149_SLICE_X13Y149_BO5),
.O6(CLBLM_L_X10Y149_SLICE_X13Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0c0c0c0c0)
  ) CLBLM_L_X10Y149_SLICE_X13Y149_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_L_X8Y152_SLICE_X11Y152_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y149_SLICE_X13Y149_AO5),
.O6(CLBLM_L_X10Y149_SLICE_X13Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y150_SLICE_X12Y150_A5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y150_SLICE_X12Y150_AO5),
.Q(CLBLM_L_X10Y150_SLICE_X12Y150_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y150_SLICE_X12Y150_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y150_SLICE_X12Y150_AO6),
.Q(CLBLM_L_X10Y150_SLICE_X12Y150_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y150_SLICE_X12Y150_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y150_SLICE_X12Y150_BO6),
.Q(CLBLM_L_X10Y150_SLICE_X12Y150_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y150_SLICE_X12Y150_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y150_SLICE_X12Y150_CO6),
.Q(CLBLM_L_X10Y150_SLICE_X12Y150_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h55ffffff88888888)
  ) CLBLM_L_X10Y150_SLICE_X12Y150_DLUT (
.I0(CLBLM_R_X11Y150_SLICE_X15Y150_AQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(1'b1),
.I3(CLBLM_L_X8Y146_SLICE_X10Y146_A5Q),
.I4(CLBLM_L_X10Y150_SLICE_X13Y150_BQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y150_SLICE_X12Y150_DO5),
.O6(CLBLM_L_X10Y150_SLICE_X12Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaf0aac0aaf0aac0)
  ) CLBLM_L_X10Y150_SLICE_X12Y150_CLUT (
.I0(CLBLM_L_X8Y150_SLICE_X11Y150_AQ),
.I1(CLBLM_L_X10Y150_SLICE_X12Y150_CQ),
.I2(CLBLM_L_X10Y143_SLICE_X12Y143_CO6),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X10Y151_SLICE_X12Y151_CO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y150_SLICE_X12Y150_CO5),
.O6(CLBLM_L_X10Y150_SLICE_X12Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haeabaeab04010401)
  ) CLBLM_L_X10Y150_SLICE_X12Y150_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X10Y150_SLICE_X12Y150_BQ),
.I2(CLBLM_R_X3Y148_SLICE_X2Y148_B5Q),
.I3(CLBLM_L_X10Y150_SLICE_X12Y150_DO6),
.I4(1'b1),
.I5(CLBLM_R_X11Y152_SLICE_X14Y152_A5Q),
.O5(CLBLM_L_X10Y150_SLICE_X12Y150_BO5),
.O6(CLBLM_L_X10Y150_SLICE_X12Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafa5050ee44ee44)
  ) CLBLM_L_X10Y150_SLICE_X12Y150_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X10Y151_SLICE_X12Y151_BO6),
.I2(CLBLM_R_X11Y151_SLICE_X14Y151_CO6),
.I3(CLBLL_L_X4Y150_SLICE_X5Y150_BQ),
.I4(CLBLM_L_X8Y145_SLICE_X11Y145_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y150_SLICE_X12Y150_AO5),
.O6(CLBLM_L_X10Y150_SLICE_X12Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y150_SLICE_X13Y150_A5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y150_SLICE_X13Y150_AO5),
.Q(CLBLM_L_X10Y150_SLICE_X13Y150_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y150_SLICE_X13Y150_B5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y151_SLICE_X13Y151_BO6),
.Q(CLBLM_L_X10Y150_SLICE_X13Y150_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y150_SLICE_X13Y150_C5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y150_SLICE_X13Y150_CO5),
.Q(CLBLM_L_X10Y150_SLICE_X13Y150_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y150_SLICE_X13Y150_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y150_SLICE_X13Y150_AO6),
.Q(CLBLM_L_X10Y150_SLICE_X13Y150_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y150_SLICE_X13Y150_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y150_SLICE_X13Y150_BO6),
.Q(CLBLM_L_X10Y150_SLICE_X13Y150_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y150_SLICE_X13Y150_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y150_SLICE_X13Y150_CO6),
.Q(CLBLM_L_X10Y150_SLICE_X13Y150_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a077ddbbee)
  ) CLBLM_L_X10Y150_SLICE_X13Y150_DLUT (
.I0(CLBLM_L_X8Y154_SLICE_X10Y154_AQ),
.I1(CLBLM_L_X10Y147_SLICE_X13Y147_B5Q),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X7Y154_SLICE_X8Y154_CQ),
.I4(CLBLM_L_X10Y148_SLICE_X12Y148_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y150_SLICE_X13Y150_DO5),
.O6(CLBLM_L_X10Y150_SLICE_X13Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf505fa0acfc0cfc0)
  ) CLBLM_L_X10Y150_SLICE_X13Y150_CLUT (
.I0(CLBLM_L_X10Y149_SLICE_X13Y149_A5Q),
.I1(CLBLM_R_X11Y151_SLICE_X14Y151_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_L_X10Y149_SLICE_X12Y149_BQ),
.I4(CLBLL_L_X4Y150_SLICE_X5Y150_CQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y150_SLICE_X13Y150_CO5),
.O6(CLBLM_L_X10Y150_SLICE_X13Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00be14aa00ee44)
  ) CLBLM_L_X10Y150_SLICE_X13Y150_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X10Y150_SLICE_X13Y150_BQ),
.I2(CLBLM_R_X11Y150_SLICE_X15Y150_AQ),
.I3(CLBLM_R_X11Y152_SLICE_X14Y152_AQ),
.I4(CLBLM_R_X3Y148_SLICE_X2Y148_B5Q),
.I5(CLBLM_L_X8Y146_SLICE_X10Y146_A5Q),
.O5(CLBLM_L_X10Y150_SLICE_X13Y150_BO5),
.O6(CLBLM_L_X10Y150_SLICE_X13Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5a0f5a0eeee4444)
  ) CLBLM_L_X10Y150_SLICE_X13Y150_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X10Y145_SLICE_X12Y145_BO6),
.I2(CLBLM_L_X10Y149_SLICE_X12Y149_DQ),
.I3(CLBLM_L_X10Y149_SLICE_X13Y149_CO6),
.I4(CLBLM_L_X8Y152_SLICE_X10Y152_D5Q),
.I5(1'b1),
.O5(CLBLM_L_X10Y150_SLICE_X13Y150_AO5),
.O6(CLBLM_L_X10Y150_SLICE_X13Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y151_SLICE_X12Y151_A_FDSE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y151_SLICE_X10Y151_CO6),
.Q(CLBLM_L_X10Y151_SLICE_X12Y151_AQ),
.S(CLBLM_R_X11Y148_SLICE_X14Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00f000f000f000f0)
  ) CLBLM_L_X10Y151_SLICE_X12Y151_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X7Y145_SLICE_X8Y145_B5Q),
.I3(CLBLM_R_X3Y150_SLICE_X3Y150_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y151_SLICE_X12Y151_DO5),
.O6(CLBLM_L_X10Y151_SLICE_X12Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccffffdcccffff)
  ) CLBLM_L_X10Y151_SLICE_X12Y151_CLUT (
.I0(RIOB33_X105Y101_IOB_X1Y102_I),
.I1(CLBLM_L_X10Y141_SLICE_X12Y141_AO6),
.I2(CLBLM_R_X7Y151_SLICE_X9Y151_BQ),
.I3(CLBLM_R_X5Y149_SLICE_X7Y149_D5Q),
.I4(CLBLM_R_X7Y153_SLICE_X8Y153_DO5),
.I5(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.O5(CLBLM_L_X10Y151_SLICE_X12Y151_CO5),
.O6(CLBLM_L_X10Y151_SLICE_X12Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hbeeeeeeeeeeeeeee)
  ) CLBLM_L_X10Y151_SLICE_X12Y151_BLUT (
.I0(CLBLM_R_X3Y148_SLICE_X2Y148_B5Q),
.I1(CLBLM_L_X10Y150_SLICE_X12Y150_A5Q),
.I2(CLBLM_R_X11Y150_SLICE_X15Y150_AQ),
.I3(CLBLM_L_X10Y150_SLICE_X12Y150_BQ),
.I4(CLBLM_L_X10Y150_SLICE_X13Y150_BQ),
.I5(CLBLM_L_X8Y146_SLICE_X10Y146_A5Q),
.O5(CLBLM_L_X10Y151_SLICE_X12Y151_BO5),
.O6(CLBLM_L_X10Y151_SLICE_X12Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h80000000c0000000)
  ) CLBLM_L_X10Y151_SLICE_X12Y151_ALUT (
.I0(CLBLM_L_X8Y146_SLICE_X10Y146_A5Q),
.I1(CLBLM_L_X10Y150_SLICE_X12Y150_A5Q),
.I2(CLBLM_R_X11Y150_SLICE_X15Y150_AQ),
.I3(CLBLM_L_X10Y150_SLICE_X12Y150_BQ),
.I4(CLBLM_L_X10Y150_SLICE_X13Y150_BQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y151_SLICE_X12Y151_AO5),
.O6(CLBLM_L_X10Y151_SLICE_X12Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y151_SLICE_X13Y151_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y151_SLICE_X13Y151_AO6),
.Q(CLBLM_L_X10Y151_SLICE_X13Y151_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_L_X10Y151_SLICE_X13Y151_DLUT (
.I0(CLBLM_R_X11Y151_SLICE_X14Y151_BQ),
.I1(CLBLM_L_X10Y151_SLICE_X12Y151_AO6),
.I2(CLBLM_R_X7Y152_SLICE_X9Y152_AQ),
.I3(CLBLM_L_X10Y151_SLICE_X13Y151_CO6),
.I4(CLBLM_L_X10Y151_SLICE_X13Y151_AQ),
.I5(CLBLM_L_X10Y152_SLICE_X13Y152_BQ),
.O5(CLBLM_L_X10Y151_SLICE_X13Y151_DO5),
.O6(CLBLM_L_X10Y151_SLICE_X13Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fffffffffffffff)
  ) CLBLM_L_X10Y151_SLICE_X13Y151_CLUT (
.I0(CLBLM_R_X11Y151_SLICE_X15Y151_AQ),
.I1(CLBLM_L_X10Y151_SLICE_X12Y151_AO5),
.I2(CLBLM_R_X11Y151_SLICE_X14Y151_BQ),
.I3(CLBLM_L_X10Y151_SLICE_X13Y151_AQ),
.I4(CLBLM_R_X7Y152_SLICE_X9Y152_AQ),
.I5(CLBLM_L_X10Y152_SLICE_X13Y152_BQ),
.O5(CLBLM_L_X10Y151_SLICE_X13Y151_CO5),
.O6(CLBLM_L_X10Y151_SLICE_X13Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f3c0c05fff5fff)
  ) CLBLM_L_X10Y151_SLICE_X13Y151_BLUT (
.I0(CLBLM_R_X7Y152_SLICE_X9Y152_AQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_L_X10Y151_SLICE_X13Y151_AQ),
.I3(CLBLM_L_X10Y151_SLICE_X12Y151_AO6),
.I4(CLBLM_L_X10Y151_SLICE_X12Y151_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y151_SLICE_X13Y151_BO5),
.O6(CLBLM_L_X10Y151_SLICE_X13Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccafffccccfaaa)
  ) CLBLM_L_X10Y151_SLICE_X13Y151_ALUT (
.I0(CLBLM_R_X3Y148_SLICE_X2Y148_B5Q),
.I1(CLBLM_R_X3Y142_SLICE_X2Y142_A5Q),
.I2(CLBLM_L_X10Y151_SLICE_X12Y151_AO6),
.I3(CLBLM_R_X7Y152_SLICE_X9Y152_AQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_L_X10Y151_SLICE_X13Y151_AQ),
.O5(CLBLM_L_X10Y151_SLICE_X13Y151_AO5),
.O6(CLBLM_L_X10Y151_SLICE_X13Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y152_SLICE_X12Y152_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y152_SLICE_X12Y152_AO6),
.Q(CLBLM_L_X10Y152_SLICE_X12Y152_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y152_SLICE_X12Y152_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y152_SLICE_X12Y152_BO6),
.Q(CLBLM_L_X10Y152_SLICE_X12Y152_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y152_SLICE_X12Y152_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y152_SLICE_X12Y152_CO6),
.Q(CLBLM_L_X10Y152_SLICE_X12Y152_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fffffffffffffff)
  ) CLBLM_L_X10Y152_SLICE_X12Y152_DLUT (
.I0(CLBLM_R_X11Y151_SLICE_X14Y151_AQ),
.I1(CLBLM_R_X11Y152_SLICE_X14Y152_A5Q),
.I2(CLBLM_L_X10Y153_SLICE_X12Y153_BQ),
.I3(CLBLM_L_X10Y153_SLICE_X12Y153_AQ),
.I4(CLBLM_L_X8Y152_SLICE_X11Y152_B5Q),
.I5(CLBLM_L_X8Y153_SLICE_X10Y153_BQ),
.O5(CLBLM_L_X10Y152_SLICE_X12Y152_DO5),
.O6(CLBLM_L_X10Y152_SLICE_X12Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaa00aaff0c0c0c)
  ) CLBLM_L_X10Y152_SLICE_X12Y152_CLUT (
.I0(CLBLM_R_X11Y152_SLICE_X15Y152_BO6),
.I1(CLBLM_L_X10Y152_SLICE_X13Y152_CO6),
.I2(CLBLM_R_X11Y152_SLICE_X14Y152_DO6),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X7Y144_SLICE_X8Y144_A5Q),
.I5(CLBLM_L_X10Y152_SLICE_X12Y152_CQ),
.O5(CLBLM_L_X10Y152_SLICE_X12Y152_CO5),
.O6(CLBLM_L_X10Y152_SLICE_X12Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff90c0000090c0)
  ) CLBLM_L_X10Y152_SLICE_X12Y152_BLUT (
.I0(CLBLM_R_X11Y152_SLICE_X14Y152_CO6),
.I1(CLBLM_L_X10Y152_SLICE_X12Y152_BQ),
.I2(CLBLM_L_X10Y152_SLICE_X13Y152_CO5),
.I3(CLBLM_L_X10Y151_SLICE_X12Y151_DO6),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X7Y155_SLICE_X8Y155_AQ),
.O5(CLBLM_L_X10Y152_SLICE_X12Y152_BO5),
.O6(CLBLM_L_X10Y152_SLICE_X12Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccca050ccccf000)
  ) CLBLM_L_X10Y152_SLICE_X12Y152_ALUT (
.I0(CLBLM_L_X10Y152_SLICE_X12Y152_DO6),
.I1(CLBLM_R_X5Y149_SLICE_X7Y149_D5Q),
.I2(CLBLM_L_X10Y152_SLICE_X13Y152_CO5),
.I3(CLBLM_L_X10Y152_SLICE_X12Y152_AQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_L_X10Y151_SLICE_X12Y151_DO6),
.O5(CLBLM_L_X10Y152_SLICE_X12Y152_AO5),
.O6(CLBLM_L_X10Y152_SLICE_X12Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y152_SLICE_X13Y152_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y152_SLICE_X13Y152_AO6),
.Q(CLBLM_L_X10Y152_SLICE_X13Y152_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y152_SLICE_X13Y152_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y152_SLICE_X13Y152_BO6),
.Q(CLBLM_L_X10Y152_SLICE_X13Y152_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000000000cc00)
  ) CLBLM_L_X10Y152_SLICE_X13Y152_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X12Y151_SLICE_X16Y151_BQ),
.I2(1'b1),
.I3(CLBLM_L_X10Y152_SLICE_X13Y152_CO6),
.I4(CLBLM_L_X10Y152_SLICE_X13Y152_AQ),
.I5(CLBLM_L_X12Y151_SLICE_X16Y151_DO6),
.O5(CLBLM_L_X10Y152_SLICE_X13Y152_DO5),
.O6(CLBLM_L_X10Y152_SLICE_X13Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h001000100fff0fff)
  ) CLBLM_L_X10Y152_SLICE_X13Y152_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X3Y150_SLICE_X3Y150_BQ),
.I2(CLBLM_R_X7Y145_SLICE_X8Y145_B5Q),
.I3(CLBLM_L_X8Y153_SLICE_X10Y153_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y152_SLICE_X13Y152_CO5),
.O6(CLBLM_L_X10Y152_SLICE_X13Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff00ffff9c009c)
  ) CLBLM_L_X10Y152_SLICE_X13Y152_BLUT (
.I0(CLBLM_L_X10Y151_SLICE_X13Y151_BO5),
.I1(CLBLM_L_X10Y152_SLICE_X13Y152_BQ),
.I2(CLBLM_R_X11Y151_SLICE_X14Y151_BQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X10Y152_SLICE_X12Y152_CQ),
.I5(CLBLM_R_X3Y148_SLICE_X2Y148_B5Q),
.O5(CLBLM_L_X10Y152_SLICE_X13Y152_BO5),
.O6(CLBLM_L_X10Y152_SLICE_X13Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffaaaaaaafaaa)
  ) CLBLM_L_X10Y152_SLICE_X13Y152_ALUT (
.I0(CLBLM_L_X10Y152_SLICE_X13Y152_DO6),
.I1(1'b1),
.I2(CLBLM_L_X10Y152_SLICE_X13Y152_AQ),
.I3(CLBLM_R_X11Y152_SLICE_X15Y152_BO6),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_L_X10Y150_SLICE_X12Y150_A5Q),
.O5(CLBLM_L_X10Y152_SLICE_X13Y152_AO5),
.O6(CLBLM_L_X10Y152_SLICE_X13Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y153_SLICE_X12Y153_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y153_SLICE_X12Y153_AO6),
.Q(CLBLM_L_X10Y153_SLICE_X12Y153_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y153_SLICE_X12Y153_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y153_SLICE_X12Y153_BO6),
.Q(CLBLM_L_X10Y153_SLICE_X12Y153_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y153_SLICE_X12Y153_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y153_SLICE_X12Y153_CO6),
.Q(CLBLM_L_X10Y153_SLICE_X12Y153_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7f7fffff5f5fffff)
  ) CLBLM_L_X10Y153_SLICE_X12Y153_DLUT (
.I0(CLBLM_L_X10Y153_SLICE_X12Y153_BQ),
.I1(CLBLM_L_X10Y153_SLICE_X12Y153_AQ),
.I2(CLBLM_L_X8Y153_SLICE_X10Y153_BQ),
.I3(1'b1),
.I4(CLBLM_L_X8Y152_SLICE_X11Y152_B5Q),
.I5(1'b1),
.O5(CLBLM_L_X10Y153_SLICE_X12Y153_DO5),
.O6(CLBLM_L_X10Y153_SLICE_X12Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafafcf30a0a0c03)
  ) CLBLM_L_X10Y153_SLICE_X12Y153_CLUT (
.I0(CLBLM_L_X8Y152_SLICE_X10Y152_D5Q),
.I1(CLBLM_L_X10Y153_SLICE_X12Y153_CQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X5Y148_SLICE_X6Y148_AO5),
.I4(CLBLM_L_X8Y149_SLICE_X11Y149_BQ),
.I5(CLBLL_L_X4Y151_SLICE_X5Y151_A5Q),
.O5(CLBLM_L_X10Y153_SLICE_X12Y153_CO5),
.O6(CLBLM_L_X10Y153_SLICE_X12Y153_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa3caa00aaccaa00)
  ) CLBLM_L_X10Y153_SLICE_X12Y153_BLUT (
.I0(CLBLM_L_X10Y153_SLICE_X12Y153_CQ),
.I1(CLBLM_L_X10Y153_SLICE_X12Y153_BQ),
.I2(CLBLM_L_X10Y151_SLICE_X12Y151_DO6),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X10Y152_SLICE_X13Y152_CO5),
.I5(CLBLM_L_X8Y153_SLICE_X10Y153_BQ),
.O5(CLBLM_L_X10Y153_SLICE_X12Y153_BO5),
.O6(CLBLM_L_X10Y153_SLICE_X12Y153_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaf03c0000)
  ) CLBLM_L_X10Y153_SLICE_X12Y153_ALUT (
.I0(CLBLM_R_X7Y147_SLICE_X9Y147_C5Q),
.I1(CLBLM_L_X10Y151_SLICE_X12Y151_DO6),
.I2(CLBLM_L_X10Y153_SLICE_X12Y153_AQ),
.I3(CLBLM_L_X10Y153_SLICE_X12Y153_DO5),
.I4(CLBLM_L_X10Y152_SLICE_X13Y152_CO5),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_L_X10Y153_SLICE_X12Y153_AO5),
.O6(CLBLM_L_X10Y153_SLICE_X12Y153_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y153_SLICE_X13Y153_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y153_SLICE_X13Y153_AO6),
.Q(CLBLM_L_X10Y153_SLICE_X13Y153_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y153_SLICE_X13Y153_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y153_SLICE_X13Y153_DO5),
.O6(CLBLM_L_X10Y153_SLICE_X13Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y153_SLICE_X13Y153_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y153_SLICE_X13Y153_CO5),
.O6(CLBLM_L_X10Y153_SLICE_X13Y153_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y153_SLICE_X13Y153_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y153_SLICE_X13Y153_BO5),
.O6(CLBLM_L_X10Y153_SLICE_X13Y153_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00ccf5cc00ccf0)
  ) CLBLM_L_X10Y153_SLICE_X13Y153_ALUT (
.I0(CLBLM_R_X5Y148_SLICE_X6Y148_AO5),
.I1(CLBLM_R_X11Y149_SLICE_X15Y149_AQ),
.I2(CLBLM_L_X10Y153_SLICE_X13Y153_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X8Y149_SLICE_X11Y149_BQ),
.I5(CLBLM_L_X10Y153_SLICE_X12Y153_CQ),
.O5(CLBLM_L_X10Y153_SLICE_X13Y153_AO5),
.O6(CLBLM_L_X10Y153_SLICE_X13Y153_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y143_SLICE_X16Y143_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y143_SLICE_X16Y143_DO5),
.O6(CLBLM_L_X12Y143_SLICE_X16Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y143_SLICE_X16Y143_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y143_SLICE_X16Y143_CO5),
.O6(CLBLM_L_X12Y143_SLICE_X16Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y143_SLICE_X16Y143_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y143_SLICE_X16Y143_BO5),
.O6(CLBLM_L_X12Y143_SLICE_X16Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffefffff)
  ) CLBLM_L_X12Y143_SLICE_X16Y143_ALUT (
.I0(CLBLM_L_X8Y144_SLICE_X11Y144_A5Q),
.I1(CLBLM_R_X11Y146_SLICE_X14Y146_AQ),
.I2(CLBLM_R_X7Y146_SLICE_X9Y146_B5Q),
.I3(CLBLM_R_X7Y144_SLICE_X8Y144_AQ),
.I4(CLBLM_R_X5Y142_SLICE_X7Y142_C5Q),
.I5(CLBLM_L_X8Y144_SLICE_X10Y144_B5Q),
.O5(CLBLM_L_X12Y143_SLICE_X16Y143_AO5),
.O6(CLBLM_L_X12Y143_SLICE_X16Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y143_SLICE_X17Y143_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y143_SLICE_X17Y143_DO5),
.O6(CLBLM_L_X12Y143_SLICE_X17Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y143_SLICE_X17Y143_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y143_SLICE_X17Y143_CO5),
.O6(CLBLM_L_X12Y143_SLICE_X17Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y143_SLICE_X17Y143_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y143_SLICE_X17Y143_BO5),
.O6(CLBLM_L_X12Y143_SLICE_X17Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y143_SLICE_X17Y143_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y143_SLICE_X17Y143_AO5),
.O6(CLBLM_L_X12Y143_SLICE_X17Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbbbaaaabbbfaaaf)
  ) CLBLM_L_X12Y144_SLICE_X16Y144_DLUT (
.I0(CLBLM_L_X12Y146_SLICE_X16Y146_AO6),
.I1(CLBLM_L_X12Y144_SLICE_X16Y144_AO6),
.I2(CLBLM_R_X11Y144_SLICE_X15Y144_AO5),
.I3(CLBLM_R_X11Y145_SLICE_X15Y145_BO5),
.I4(RIOB33_X105Y143_IOB_X1Y143_I),
.I5(CLBLM_R_X11Y143_SLICE_X15Y143_DO6),
.O5(CLBLM_L_X12Y144_SLICE_X16Y144_DO5),
.O6(CLBLM_L_X12Y144_SLICE_X16Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hddccddccddccdfcf)
  ) CLBLM_L_X12Y144_SLICE_X16Y144_CLUT (
.I0(CLBLM_L_X12Y144_SLICE_X16Y144_AO6),
.I1(CLBLM_L_X12Y145_SLICE_X16Y145_BO6),
.I2(CLBLM_R_X11Y145_SLICE_X15Y145_BO5),
.I3(RIOB33_X105Y141_IOB_X1Y142_I),
.I4(CLBLM_R_X11Y144_SLICE_X15Y144_AO5),
.I5(CLBLM_R_X11Y143_SLICE_X15Y143_DO6),
.O5(CLBLM_L_X12Y144_SLICE_X16Y144_CO5),
.O6(CLBLM_L_X12Y144_SLICE_X16Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffefffcfefefcfc)
  ) CLBLM_L_X12Y144_SLICE_X16Y144_BLUT (
.I0(RIOB33_X105Y137_IOB_X1Y137_I),
.I1(CLBLM_L_X12Y145_SLICE_X17Y145_BO6),
.I2(CLBLM_L_X12Y145_SLICE_X17Y145_AO6),
.I3(RIOB33_X105Y135_IOB_X1Y136_I),
.I4(CLBLM_R_X7Y149_SLICE_X9Y149_BQ),
.I5(CLBLM_R_X11Y144_SLICE_X14Y144_AQ),
.O5(CLBLM_L_X12Y144_SLICE_X16Y144_BO5),
.O6(CLBLM_L_X12Y144_SLICE_X16Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff5fff500a80008)
  ) CLBLM_L_X12Y144_SLICE_X16Y144_ALUT (
.I0(CLBLM_R_X11Y142_SLICE_X14Y142_DO6),
.I1(RIOB33_X105Y143_IOB_X1Y144_I),
.I2(CLBLM_R_X11Y149_SLICE_X14Y149_AQ),
.I3(CLBLM_L_X8Y150_SLICE_X10Y150_A5Q),
.I4(CLBLM_R_X11Y148_SLICE_X14Y148_DQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y144_SLICE_X16Y144_AO5),
.O6(CLBLM_L_X12Y144_SLICE_X16Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y144_SLICE_X17Y144_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y144_SLICE_X17Y144_DO5),
.O6(CLBLM_L_X12Y144_SLICE_X17Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y144_SLICE_X17Y144_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y144_SLICE_X17Y144_CO5),
.O6(CLBLM_L_X12Y144_SLICE_X17Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y144_SLICE_X17Y144_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y144_SLICE_X17Y144_BO5),
.O6(CLBLM_L_X12Y144_SLICE_X17Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y144_SLICE_X17Y144_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y144_SLICE_X17Y144_AO5),
.O6(CLBLM_L_X12Y144_SLICE_X17Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hba30ba30ba30ba30)
  ) CLBLM_L_X12Y145_SLICE_X16Y145_DLUT (
.I0(CLBLM_R_X11Y145_SLICE_X15Y145_BO5),
.I1(CLBLM_L_X12Y145_SLICE_X16Y145_AO6),
.I2(RIOB33_X105Y137_IOB_X1Y138_I),
.I3(CLBLM_R_X3Y145_SLICE_X3Y145_DQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y145_SLICE_X16Y145_DO5),
.O6(CLBLM_L_X12Y145_SLICE_X16Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha202a00000000000)
  ) CLBLM_L_X12Y145_SLICE_X16Y145_CLUT (
.I0(CLBLM_R_X11Y142_SLICE_X14Y142_BO6),
.I1(CLBLM_R_X7Y146_SLICE_X9Y146_B5Q),
.I2(CLBLM_R_X11Y149_SLICE_X14Y149_AQ),
.I3(CLBLL_L_X4Y144_SLICE_X5Y144_BQ),
.I4(CLBLM_L_X10Y147_SLICE_X13Y147_AQ),
.I5(CLBLM_L_X8Y150_SLICE_X10Y150_A5Q),
.O5(CLBLM_L_X12Y145_SLICE_X16Y145_CO5),
.O6(CLBLM_L_X12Y145_SLICE_X16Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5088008850000000)
  ) CLBLM_L_X12Y145_SLICE_X16Y145_BLUT (
.I0(CLBLM_R_X11Y149_SLICE_X14Y149_AQ),
.I1(CLBLM_R_X11Y145_SLICE_X14Y145_CQ),
.I2(CLBLM_R_X11Y142_SLICE_X14Y142_BO6),
.I3(CLBLM_L_X8Y150_SLICE_X10Y150_A5Q),
.I4(CLBLM_L_X10Y147_SLICE_X12Y147_AQ),
.I5(CLBLM_R_X11Y142_SLICE_X14Y142_DO6),
.O5(CLBLM_L_X12Y145_SLICE_X16Y145_BO5),
.O6(CLBLM_L_X12Y145_SLICE_X16Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff33ff22003000)
  ) CLBLM_L_X12Y145_SLICE_X16Y145_ALUT (
.I0(CLBLM_R_X11Y145_SLICE_X14Y145_DQ),
.I1(CLBLM_L_X8Y150_SLICE_X10Y150_A5Q),
.I2(RIOB33_X105Y145_IOB_X1Y146_I),
.I3(CLBLM_R_X11Y142_SLICE_X14Y142_DO6),
.I4(CLBLM_R_X11Y149_SLICE_X14Y149_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y145_SLICE_X16Y145_AO5),
.O6(CLBLM_L_X12Y145_SLICE_X16Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y145_SLICE_X17Y145_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y145_SLICE_X17Y145_DO5),
.O6(CLBLM_L_X12Y145_SLICE_X17Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaffaa0000ff00)
  ) CLBLM_L_X12Y145_SLICE_X17Y145_CLUT (
.I0(CLBLM_R_X11Y145_SLICE_X15Y145_BO5),
.I1(1'b1),
.I2(1'b1),
.I3(RIOB33_X105Y137_IOB_X1Y137_I),
.I4(CLBLM_L_X12Y145_SLICE_X16Y145_AO6),
.I5(CLBLM_R_X7Y145_SLICE_X9Y145_BQ),
.O5(CLBLM_L_X12Y145_SLICE_X17Y145_CO5),
.O6(CLBLM_L_X12Y145_SLICE_X17Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefafefaeeaaeeaa)
  ) CLBLM_L_X12Y145_SLICE_X17Y145_BLUT (
.I0(CLBLM_R_X11Y146_SLICE_X15Y146_BO5),
.I1(RIOB33_X105Y135_IOB_X1Y135_I),
.I2(CLBLM_L_X10Y145_SLICE_X12Y145_AQ),
.I3(CLBLM_R_X11Y145_SLICE_X15Y145_AQ),
.I4(1'b1),
.I5(RIOB33_X105Y137_IOB_X1Y138_I),
.O5(CLBLM_L_X12Y145_SLICE_X17Y145_BO5),
.O6(CLBLM_L_X12Y145_SLICE_X17Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffcccfcccfccc)
  ) CLBLM_L_X12Y145_SLICE_X17Y145_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X13Y145_SLICE_X18Y145_AO6),
.I2(RIOB33_X105Y141_IOB_X1Y142_I),
.I3(CLBLM_R_X11Y145_SLICE_X14Y145_CQ),
.I4(RIOB33_X105Y145_IOB_X1Y146_I),
.I5(CLBLM_R_X11Y145_SLICE_X14Y145_DQ),
.O5(CLBLM_L_X12Y145_SLICE_X17Y145_AO5),
.O6(CLBLM_L_X12Y145_SLICE_X17Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y146_SLICE_X16Y146_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y146_SLICE_X16Y146_DO5),
.O6(CLBLM_L_X12Y146_SLICE_X16Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y146_SLICE_X16Y146_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y146_SLICE_X16Y146_CO5),
.O6(CLBLM_L_X12Y146_SLICE_X16Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fc00ccf0fc00cc)
  ) CLBLM_L_X12Y146_SLICE_X16Y146_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y149_SLICE_X9Y149_BQ),
.I2(RIOB33_X105Y147_IOB_X1Y148_I),
.I3(CLBLM_R_X11Y146_SLICE_X15Y146_CO5),
.I4(CLBLM_R_X11Y142_SLICE_X14Y142_CO5),
.I5(1'b1),
.O5(CLBLM_L_X12Y146_SLICE_X16Y146_BO5),
.O6(CLBLM_L_X12Y146_SLICE_X16Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5000888850000000)
  ) CLBLM_L_X12Y146_SLICE_X16Y146_ALUT (
.I0(CLBLM_R_X11Y149_SLICE_X14Y149_AQ),
.I1(CLBLM_R_X11Y148_SLICE_X14Y148_BQ),
.I2(CLBLM_R_X11Y142_SLICE_X14Y142_BO6),
.I3(CLBLM_L_X12Y149_SLICE_X16Y149_BQ),
.I4(CLBLM_L_X8Y150_SLICE_X10Y150_A5Q),
.I5(CLBLM_R_X11Y142_SLICE_X14Y142_DO6),
.O5(CLBLM_L_X12Y146_SLICE_X16Y146_AO5),
.O6(CLBLM_L_X12Y146_SLICE_X16Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y146_SLICE_X17Y146_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y146_SLICE_X17Y146_DO5),
.O6(CLBLM_L_X12Y146_SLICE_X17Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y146_SLICE_X17Y146_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y146_SLICE_X17Y146_CO5),
.O6(CLBLM_L_X12Y146_SLICE_X17Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y146_SLICE_X17Y146_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y146_SLICE_X17Y146_BO5),
.O6(CLBLM_L_X12Y146_SLICE_X17Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y146_SLICE_X17Y146_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y146_SLICE_X17Y146_AO5),
.O6(CLBLM_L_X12Y146_SLICE_X17Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y149_SLICE_X16Y149_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y149_SLICE_X16Y149_AO6),
.Q(CLBLM_L_X12Y149_SLICE_X16Y149_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y149_SLICE_X16Y149_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y149_SLICE_X16Y149_BO6),
.Q(CLBLM_L_X12Y149_SLICE_X16Y149_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0a0a05050a0a0505)
  ) CLBLM_L_X12Y149_SLICE_X16Y149_DLUT (
.I0(CLBLM_R_X11Y149_SLICE_X15Y149_BQ),
.I1(1'b1),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(1'b1),
.I4(CLBLM_R_X11Y148_SLICE_X14Y148_AO6),
.I5(1'b1),
.O5(CLBLM_L_X12Y149_SLICE_X16Y149_DO5),
.O6(CLBLM_L_X12Y149_SLICE_X16Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffeeffff)
  ) CLBLM_L_X12Y149_SLICE_X16Y149_CLUT (
.I0(RIOB33_X105Y133_IOB_X1Y133_I),
.I1(CLBLM_L_X12Y149_SLICE_X16Y149_AQ),
.I2(1'b1),
.I3(RIOB33_X105Y129_IOB_X1Y130_I),
.I4(RIOB33_X105Y131_IOB_X1Y132_I),
.I5(RIOB33_X105Y129_IOB_X1Y129_I),
.O5(CLBLM_L_X12Y149_SLICE_X16Y149_CO5),
.O6(CLBLM_L_X12Y149_SLICE_X16Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000e4e4e4e4)
  ) CLBLM_L_X12Y149_SLICE_X16Y149_BLUT (
.I0(CLBLM_R_X11Y145_SLICE_X15Y145_BO5),
.I1(CLBLM_L_X12Y149_SLICE_X16Y149_BQ),
.I2(CLBLL_L_X4Y149_SLICE_X5Y149_DQ),
.I3(1'b1),
.I4(CLBLM_L_X10Y149_SLICE_X12Y149_AQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_L_X12Y149_SLICE_X16Y149_BO5),
.O6(CLBLM_L_X12Y149_SLICE_X16Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00a5a56565)
  ) CLBLM_L_X12Y149_SLICE_X16Y149_ALUT (
.I0(CLBLM_R_X11Y148_SLICE_X14Y148_AO6),
.I1(RIOB33_X105Y131_IOB_X1Y132_I),
.I2(CLBLM_R_X11Y149_SLICE_X15Y149_BQ),
.I3(CLBLM_L_X10Y147_SLICE_X13Y147_AQ),
.I4(RIOB33_X105Y133_IOB_X1Y133_I),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_L_X12Y149_SLICE_X16Y149_AO5),
.O6(CLBLM_L_X12Y149_SLICE_X16Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y149_SLICE_X17Y149_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y149_SLICE_X17Y149_DO5),
.O6(CLBLM_L_X12Y149_SLICE_X17Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y149_SLICE_X17Y149_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y149_SLICE_X17Y149_CO5),
.O6(CLBLM_L_X12Y149_SLICE_X17Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y149_SLICE_X17Y149_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y149_SLICE_X17Y149_BO5),
.O6(CLBLM_L_X12Y149_SLICE_X17Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y149_SLICE_X17Y149_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y149_SLICE_X17Y149_AO5),
.O6(CLBLM_L_X12Y149_SLICE_X17Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y151_SLICE_X16Y151_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X12Y151_SLICE_X16Y151_AO6),
.Q(CLBLM_L_X12Y151_SLICE_X16Y151_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y151_SLICE_X16Y151_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X12Y151_SLICE_X16Y151_BO6),
.Q(CLBLM_L_X12Y151_SLICE_X16Y151_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff7f7f7f7f)
  ) CLBLM_L_X12Y151_SLICE_X16Y151_DLUT (
.I0(CLBLM_R_X11Y152_SLICE_X14Y152_AQ),
.I1(CLBLM_L_X10Y152_SLICE_X12Y152_BQ),
.I2(CLBLM_L_X12Y151_SLICE_X16Y151_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X11Y151_SLICE_X14Y151_DO6),
.O5(CLBLM_L_X12Y151_SLICE_X16Y151_DO5),
.O6(CLBLM_L_X12Y151_SLICE_X16Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffccffaaffaaff)
  ) CLBLM_L_X12Y151_SLICE_X16Y151_CLUT (
.I0(CLBLM_R_X11Y146_SLICE_X14Y146_BO6),
.I1(CLBLM_L_X10Y145_SLICE_X12Y145_BO6),
.I2(1'b1),
.I3(CLBLM_R_X3Y151_SLICE_X3Y151_D5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y151_SLICE_X16Y151_CO5),
.O6(CLBLM_L_X12Y151_SLICE_X16Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f09900cc00)
  ) CLBLM_L_X12Y151_SLICE_X16Y151_BLUT (
.I0(CLBLM_L_X12Y151_SLICE_X16Y151_DO6),
.I1(CLBLM_L_X12Y151_SLICE_X16Y151_BQ),
.I2(CLBLM_R_X11Y148_SLICE_X15Y148_AQ),
.I3(CLBLM_L_X10Y152_SLICE_X13Y152_CO5),
.I4(CLBLM_L_X10Y151_SLICE_X12Y151_DO6),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_L_X12Y151_SLICE_X16Y151_BO5),
.O6(CLBLM_L_X12Y151_SLICE_X16Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heecc2200decc1200)
  ) CLBLM_L_X12Y151_SLICE_X16Y151_ALUT (
.I0(CLBLM_L_X12Y151_SLICE_X16Y151_AQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_L_X10Y151_SLICE_X12Y151_DO6),
.I3(CLBLM_L_X10Y152_SLICE_X13Y152_CO5),
.I4(CLBLM_L_X10Y151_SLICE_X12Y151_AQ),
.I5(CLBLM_R_X11Y151_SLICE_X14Y151_DO6),
.O5(CLBLM_L_X12Y151_SLICE_X16Y151_AO5),
.O6(CLBLM_L_X12Y151_SLICE_X16Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y151_SLICE_X17Y151_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y151_SLICE_X17Y151_DO5),
.O6(CLBLM_L_X12Y151_SLICE_X17Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y151_SLICE_X17Y151_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y151_SLICE_X17Y151_CO5),
.O6(CLBLM_L_X12Y151_SLICE_X17Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y151_SLICE_X17Y151_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y151_SLICE_X17Y151_BO5),
.O6(CLBLM_L_X12Y151_SLICE_X17Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y151_SLICE_X17Y151_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y151_SLICE_X17Y151_AO5),
.O6(CLBLM_L_X12Y151_SLICE_X17Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y141_SLICE_X2Y141_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y141_SLICE_X2Y141_DO5),
.O6(CLBLM_R_X3Y141_SLICE_X2Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y141_SLICE_X2Y141_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y141_SLICE_X2Y141_CO5),
.O6(CLBLM_R_X3Y141_SLICE_X2Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffc)
  ) CLBLM_R_X3Y141_SLICE_X2Y141_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y146_SLICE_X2Y146_BQ),
.I2(CLBLL_L_X4Y143_SLICE_X5Y143_C5Q),
.I3(CLBLM_R_X3Y145_SLICE_X2Y145_CQ),
.I4(CLBLM_R_X3Y145_SLICE_X2Y145_B5Q),
.I5(CLBLM_R_X3Y141_SLICE_X2Y141_AO5),
.O5(CLBLM_R_X3Y141_SLICE_X2Y141_BO5),
.O6(CLBLM_R_X3Y141_SLICE_X2Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000fffffffc)
  ) CLBLM_R_X3Y141_SLICE_X2Y141_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLL_L_X2Y153_SLICE_X1Y153_AQ),
.I2(CLBLM_R_X3Y145_SLICE_X2Y145_C5Q),
.I3(CLBLM_R_X5Y143_SLICE_X6Y143_DQ),
.I4(CLBLM_R_X3Y146_SLICE_X2Y146_CQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y141_SLICE_X2Y141_AO5),
.O6(CLBLM_R_X3Y141_SLICE_X2Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000303000cc0000)
  ) CLBLM_R_X3Y141_SLICE_X3Y141_DLUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y142_SLICE_X5Y142_AQ),
.I2(CLBLM_R_X5Y142_SLICE_X6Y142_C5Q),
.I3(CLBLL_L_X4Y143_SLICE_X4Y143_CQ),
.I4(CLBLM_L_X10Y142_SLICE_X12Y142_AQ),
.I5(CLBLM_R_X3Y142_SLICE_X3Y142_BQ),
.O5(CLBLM_R_X3Y141_SLICE_X3Y141_DO5),
.O6(CLBLM_R_X3Y141_SLICE_X3Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000333300331333)
  ) CLBLM_R_X3Y141_SLICE_X3Y141_CLUT (
.I0(CLBLM_R_X3Y141_SLICE_X2Y141_BO6),
.I1(CLBLL_L_X4Y142_SLICE_X5Y142_AQ),
.I2(CLBLM_R_X5Y142_SLICE_X6Y142_C5Q),
.I3(CLBLL_L_X4Y141_SLICE_X5Y141_BO5),
.I4(CLBLM_R_X5Y144_SLICE_X6Y144_D5Q),
.I5(CLBLM_R_X3Y142_SLICE_X3Y142_BQ),
.O5(CLBLM_R_X3Y141_SLICE_X3Y141_CO5),
.O6(CLBLM_R_X3Y141_SLICE_X3Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffcdcfcdcd)
  ) CLBLM_R_X3Y141_SLICE_X3Y141_BLUT (
.I0(CLBLL_L_X4Y141_SLICE_X5Y141_BO5),
.I1(CLBLL_L_X4Y142_SLICE_X5Y142_AQ),
.I2(CLBLM_R_X3Y142_SLICE_X3Y142_BQ),
.I3(CLBLM_R_X5Y142_SLICE_X6Y142_C5Q),
.I4(CLBLM_R_X3Y141_SLICE_X2Y141_BO6),
.I5(CLBLM_L_X10Y142_SLICE_X12Y142_AQ),
.O5(CLBLM_R_X3Y141_SLICE_X3Y141_BO5),
.O6(CLBLM_R_X3Y141_SLICE_X3Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heeaaaaaeaaaaaaae)
  ) CLBLM_R_X3Y141_SLICE_X3Y141_ALUT (
.I0(CLBLM_R_X3Y141_SLICE_X3Y141_DO6),
.I1(CLBLL_L_X4Y142_SLICE_X5Y142_AQ),
.I2(CLBLM_R_X7Y150_SLICE_X9Y150_B5Q),
.I3(CLBLM_R_X3Y142_SLICE_X3Y142_BQ),
.I4(CLBLM_L_X10Y142_SLICE_X12Y142_AQ),
.I5(CLBLL_L_X4Y141_SLICE_X5Y141_BO5),
.O5(CLBLM_R_X3Y141_SLICE_X3Y141_AO5),
.O6(CLBLM_R_X3Y141_SLICE_X3Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y142_SLICE_X2Y142_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y142_SLICE_X2Y142_CO6),
.Q(CLBLM_R_X3Y142_SLICE_X2Y142_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y142_SLICE_X2Y142_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y142_SLICE_X2Y142_BO5),
.Q(CLBLM_R_X3Y142_SLICE_X2Y142_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y142_SLICE_X2Y142_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y142_SLICE_X2Y142_AO6),
.Q(CLBLM_R_X3Y142_SLICE_X2Y142_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y142_SLICE_X2Y142_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y142_SLICE_X2Y142_BO6),
.Q(CLBLM_R_X3Y142_SLICE_X2Y142_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y142_SLICE_X2Y142_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y142_SLICE_X2Y142_DO5),
.O6(CLBLM_R_X3Y142_SLICE_X2Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha3acafa033333333)
  ) CLBLM_R_X3Y142_SLICE_X2Y142_CLUT (
.I0(CLBLM_R_X5Y145_SLICE_X7Y145_A5Q),
.I1(LIOB33_X0Y59_IOB_X0Y60_I),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X3Y142_SLICE_X2Y142_A5Q),
.I4(CLBLM_R_X3Y143_SLICE_X2Y143_DQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y142_SLICE_X2Y142_CO5),
.O6(CLBLM_R_X3Y142_SLICE_X2Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'heeee4444f5a0f5a0)
  ) CLBLM_R_X3Y142_SLICE_X2Y142_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLL_L_X4Y143_SLICE_X5Y143_C5Q),
.I2(CLBLM_R_X5Y153_SLICE_X6Y153_DQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_R_X3Y142_SLICE_X3Y142_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y142_SLICE_X2Y142_BO5),
.O6(CLBLM_R_X3Y142_SLICE_X2Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfaeefafa50445050)
  ) CLBLM_R_X3Y142_SLICE_X2Y142_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X3Y145_SLICE_X3Y145_A5Q),
.I2(CLBLM_R_X3Y142_SLICE_X2Y142_AQ),
.I3(CLBLM_L_X8Y146_SLICE_X10Y146_AQ),
.I4(CLBLM_R_X7Y150_SLICE_X9Y150_CQ),
.I5(CLBLM_R_X3Y142_SLICE_X3Y142_CQ),
.O5(CLBLM_R_X3Y142_SLICE_X2Y142_AO5),
.O6(CLBLM_R_X3Y142_SLICE_X2Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y142_SLICE_X3Y142_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y142_SLICE_X3Y142_AO6),
.Q(CLBLM_R_X3Y142_SLICE_X3Y142_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y142_SLICE_X3Y142_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y142_SLICE_X3Y142_BO6),
.Q(CLBLM_R_X3Y142_SLICE_X3Y142_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y142_SLICE_X3Y142_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y142_SLICE_X3Y142_CO6),
.Q(CLBLM_R_X3Y142_SLICE_X3Y142_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000020000)
  ) CLBLM_R_X3Y142_SLICE_X3Y142_DLUT (
.I0(CLBLL_L_X4Y142_SLICE_X5Y142_AQ),
.I1(CLBLM_R_X5Y144_SLICE_X6Y144_D5Q),
.I2(CLBLM_R_X3Y142_SLICE_X3Y142_BQ),
.I3(CLBLL_L_X4Y143_SLICE_X4Y143_CQ),
.I4(CLBLM_L_X10Y142_SLICE_X12Y142_AQ),
.I5(CLBLM_R_X5Y142_SLICE_X6Y142_C5Q),
.O5(CLBLM_R_X3Y142_SLICE_X3Y142_DO5),
.O6(CLBLM_R_X3Y142_SLICE_X3Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0cc33f0f00000)
  ) CLBLM_R_X3Y142_SLICE_X3Y142_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y142_SLICE_X3Y142_CQ),
.I2(CLBLM_R_X3Y145_SLICE_X3Y145_CQ),
.I3(CLBLM_R_X3Y143_SLICE_X3Y143_CO6),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(LIOB33_X0Y53_IOB_X0Y54_I),
.O5(CLBLM_R_X3Y142_SLICE_X3Y142_CO5),
.O6(CLBLM_R_X3Y142_SLICE_X3Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff5555ffab5501)
  ) CLBLM_R_X3Y142_SLICE_X3Y142_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X5Y144_SLICE_X6Y144_D5Q),
.I2(CLBLM_R_X3Y141_SLICE_X3Y141_BO6),
.I3(CLBLM_R_X3Y142_SLICE_X3Y142_DO6),
.I4(CLBLM_L_X8Y148_SLICE_X11Y148_CQ),
.I5(CLBLL_L_X4Y142_SLICE_X4Y142_DO6),
.O5(CLBLM_R_X3Y142_SLICE_X3Y142_BO5),
.O6(CLBLM_R_X3Y142_SLICE_X3Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbffbfff51551555)
  ) CLBLM_R_X3Y142_SLICE_X3Y142_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(LIOB33_X0Y53_IOB_X0Y54_I),
.I2(CLBLM_R_X3Y142_SLICE_X3Y142_AQ),
.I3(CLBLM_R_X3Y143_SLICE_X3Y143_DO6),
.I4(CLBLM_R_X3Y143_SLICE_X3Y143_CO5),
.I5(CLBLL_L_X4Y142_SLICE_X5Y142_CQ),
.O5(CLBLM_R_X3Y142_SLICE_X3Y142_AO5),
.O6(CLBLM_R_X3Y142_SLICE_X3Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y143_SLICE_X2Y143_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y143_SLICE_X2Y143_AO6),
.Q(CLBLM_R_X3Y143_SLICE_X2Y143_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y143_SLICE_X2Y143_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y143_SLICE_X2Y143_BO6),
.Q(CLBLM_R_X3Y143_SLICE_X2Y143_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y143_SLICE_X2Y143_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y143_SLICE_X2Y143_CO6),
.Q(CLBLM_R_X3Y143_SLICE_X2Y143_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y143_SLICE_X2Y143_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y143_SLICE_X2Y143_DO6),
.Q(CLBLM_R_X3Y143_SLICE_X2Y143_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0f0faaaaf0f0)
  ) CLBLM_R_X3Y143_SLICE_X2Y143_DLUT (
.I0(CLBLL_L_X4Y141_SLICE_X5Y141_AQ),
.I1(1'b1),
.I2(CLBLM_R_X3Y143_SLICE_X2Y143_DQ),
.I3(1'b1),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(LIOB33_X0Y59_IOB_X0Y60_I),
.O5(CLBLM_R_X3Y143_SLICE_X2Y143_DO5),
.O6(CLBLM_R_X3Y143_SLICE_X2Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ccccf0f066cc)
  ) CLBLM_R_X3Y143_SLICE_X2Y143_CLUT (
.I0(CLBLM_R_X3Y143_SLICE_X2Y143_BQ),
.I1(CLBLM_R_X3Y143_SLICE_X2Y143_CQ),
.I2(CLBLL_L_X4Y154_SLICE_X4Y154_AQ),
.I3(CLBLM_R_X3Y142_SLICE_X3Y142_CQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X3Y143_SLICE_X3Y143_CO6),
.O5(CLBLM_R_X3Y143_SLICE_X2Y143_CO5),
.O6(CLBLM_R_X3Y143_SLICE_X2Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hec20ce02ee22cc00)
  ) CLBLM_R_X3Y143_SLICE_X2Y143_BLUT (
.I0(LIOB33_X0Y53_IOB_X0Y54_I),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X3Y143_SLICE_X3Y143_CO6),
.I3(CLBLM_L_X8Y143_SLICE_X11Y143_DQ),
.I4(CLBLM_R_X3Y143_SLICE_X2Y143_BQ),
.I5(CLBLM_R_X3Y142_SLICE_X3Y142_CQ),
.O5(CLBLM_R_X3Y143_SLICE_X2Y143_BO5),
.O6(CLBLM_R_X3Y143_SLICE_X2Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbfaa1500ffaa5500)
  ) CLBLM_R_X3Y143_SLICE_X2Y143_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X3Y143_SLICE_X2Y143_DQ),
.I2(CLBLM_R_X3Y142_SLICE_X2Y142_A5Q),
.I3(CLBLL_L_X2Y150_SLICE_X1Y150_DO5),
.I4(CLBLM_R_X5Y149_SLICE_X6Y149_BQ),
.I5(LIOB33_X0Y59_IOB_X0Y60_I),
.O5(CLBLM_R_X3Y143_SLICE_X2Y143_AO5),
.O6(CLBLM_R_X3Y143_SLICE_X2Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y143_SLICE_X3Y143_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y143_SLICE_X3Y143_AO6),
.Q(CLBLM_R_X3Y143_SLICE_X3Y143_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fffffffffffffff)
  ) CLBLM_R_X3Y143_SLICE_X3Y143_DLUT (
.I0(CLBLM_R_X3Y142_SLICE_X3Y142_AQ),
.I1(CLBLM_R_X3Y142_SLICE_X3Y142_CQ),
.I2(CLBLM_R_X3Y145_SLICE_X3Y145_BQ),
.I3(CLBLM_R_X3Y145_SLICE_X3Y145_CQ),
.I4(CLBLM_R_X3Y143_SLICE_X3Y143_AQ),
.I5(CLBLM_R_X3Y143_SLICE_X2Y143_BQ),
.O5(CLBLM_R_X3Y143_SLICE_X3Y143_DO5),
.O6(CLBLM_R_X3Y143_SLICE_X3Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h77ffffff33ffffff)
  ) CLBLM_R_X3Y143_SLICE_X3Y143_CLUT (
.I0(CLBLM_R_X3Y142_SLICE_X3Y142_AQ),
.I1(CLBLM_R_X3Y145_SLICE_X3Y145_BQ),
.I2(1'b1),
.I3(CLBLM_R_X3Y145_SLICE_X3Y145_CQ),
.I4(CLBLM_R_X3Y143_SLICE_X3Y143_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y143_SLICE_X3Y143_CO5),
.O6(CLBLM_R_X3Y143_SLICE_X3Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00008aaa75557555)
  ) CLBLM_R_X3Y143_SLICE_X3Y143_BLUT (
.I0(LIOB33_X0Y53_IOB_X0Y54_I),
.I1(CLBLM_R_X3Y143_SLICE_X3Y143_CO6),
.I2(CLBLM_R_X3Y142_SLICE_X3Y142_CQ),
.I3(CLBLM_R_X3Y143_SLICE_X2Y143_BQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y143_SLICE_X3Y143_BO5),
.O6(CLBLM_R_X3Y143_SLICE_X3Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffbe00befffa00fa)
  ) CLBLM_R_X3Y143_SLICE_X3Y143_ALUT (
.I0(CLBLM_R_X3Y143_SLICE_X3Y143_BO5),
.I1(CLBLM_R_X3Y145_SLICE_X3Y145_BQ),
.I2(CLBLM_R_X3Y143_SLICE_X3Y143_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLL_L_X2Y143_SLICE_X1Y143_BQ),
.I5(CLBLM_R_X3Y145_SLICE_X3Y145_CQ),
.O5(CLBLM_R_X3Y143_SLICE_X3Y143_AO5),
.O6(CLBLM_R_X3Y143_SLICE_X3Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y144_SLICE_X2Y144_A5_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y144_SLICE_X2Y144_AO5),
.Q(CLBLM_R_X3Y144_SLICE_X2Y144_A5Q),
.S(CLBLM_R_X3Y146_SLICE_X2Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y144_SLICE_X2Y144_A_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y144_SLICE_X2Y144_AO6),
.Q(CLBLM_R_X3Y144_SLICE_X2Y144_AQ),
.S(CLBLM_R_X3Y146_SLICE_X2Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y144_SLICE_X2Y144_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y144_SLICE_X2Y144_DO5),
.O6(CLBLM_R_X3Y144_SLICE_X2Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000020000000200)
  ) CLBLM_R_X3Y144_SLICE_X2Y144_CLUT (
.I0(CLBLM_R_X5Y148_SLICE_X7Y148_AO6),
.I1(CLBLM_R_X7Y144_SLICE_X9Y144_CQ),
.I2(CLBLL_L_X2Y147_SLICE_X0Y147_B5Q),
.I3(CLBLM_R_X5Y142_SLICE_X7Y142_AO5),
.I4(CLBLL_L_X2Y147_SLICE_X0Y147_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y144_SLICE_X2Y144_CO5),
.O6(CLBLM_R_X3Y144_SLICE_X2Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f00077bbddee)
  ) CLBLM_R_X3Y144_SLICE_X2Y144_BLUT (
.I0(CLBLM_R_X3Y146_SLICE_X2Y146_CQ),
.I1(CLBLM_R_X3Y142_SLICE_X2Y142_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X3Y145_SLICE_X2Y145_BQ),
.I4(CLBLL_L_X4Y143_SLICE_X5Y143_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X3Y144_SLICE_X2Y144_BO5),
.O6(CLBLM_R_X3Y144_SLICE_X2Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0000cc00cc00)
  ) CLBLM_R_X3Y144_SLICE_X2Y144_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(1'b1),
.I3(CLBLM_R_X3Y144_SLICE_X3Y144_BQ),
.I4(CLBLM_L_X8Y142_SLICE_X11Y142_CQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y144_SLICE_X2Y144_AO5),
.O6(CLBLM_R_X3Y144_SLICE_X2Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y144_SLICE_X3Y144_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y144_SLICE_X3Y144_AO5),
.Q(CLBLM_R_X3Y144_SLICE_X3Y144_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y144_SLICE_X3Y144_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y144_SLICE_X3Y144_DO5),
.Q(CLBLM_R_X3Y144_SLICE_X3Y144_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y144_SLICE_X3Y144_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y144_SLICE_X3Y144_AO6),
.Q(CLBLM_R_X3Y144_SLICE_X3Y144_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y144_SLICE_X3Y144_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y144_SLICE_X3Y144_BO6),
.Q(CLBLM_R_X3Y144_SLICE_X3Y144_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y144_SLICE_X3Y144_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y144_SLICE_X3Y144_CO6),
.Q(CLBLM_R_X3Y144_SLICE_X3Y144_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y144_SLICE_X3Y144_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y144_SLICE_X3Y144_DO6),
.Q(CLBLM_R_X3Y144_SLICE_X3Y144_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd88dd88f5f5a0a0)
  ) CLBLM_R_X3Y144_SLICE_X3Y144_DLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X3Y143_SLICE_X3Y143_AQ),
.I2(CLBLM_R_X3Y144_SLICE_X3Y144_DQ),
.I3(CLBLL_L_X2Y153_SLICE_X1Y153_AQ),
.I4(CLBLL_L_X4Y152_SLICE_X5Y152_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X3Y144_SLICE_X3Y144_DO5),
.O6(CLBLM_R_X3Y144_SLICE_X3Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hafafaca3afafacac)
  ) CLBLM_R_X3Y144_SLICE_X3Y144_CLUT (
.I0(CLBLM_R_X3Y145_SLICE_X3Y145_AQ),
.I1(CLBLM_R_X3Y144_SLICE_X3Y144_CQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLL_L_X4Y144_SLICE_X4Y144_DO6),
.I4(CLBLL_L_X2Y148_SLICE_X0Y148_B5Q),
.I5(CLBLM_R_X5Y144_SLICE_X7Y144_CQ),
.O5(CLBLM_R_X3Y144_SLICE_X3Y144_CO5),
.O6(CLBLM_R_X3Y144_SLICE_X3Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hafa0aca0afafacac)
  ) CLBLM_R_X3Y144_SLICE_X3Y144_BLUT (
.I0(CLBLM_R_X7Y144_SLICE_X9Y144_D5Q),
.I1(CLBLM_R_X3Y144_SLICE_X3Y144_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X5Y144_SLICE_X6Y144_CQ),
.I4(CLBLL_L_X2Y146_SLICE_X1Y146_AQ),
.I5(CLBLM_R_X3Y147_SLICE_X3Y147_BQ),
.O5(CLBLM_R_X3Y144_SLICE_X3Y144_BO5),
.O6(CLBLM_R_X3Y144_SLICE_X3Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heeaaeeaaf3f3c0c0)
  ) CLBLM_R_X3Y144_SLICE_X3Y144_ALUT (
.I0(CLBLM_R_X3Y147_SLICE_X3Y147_DO6),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X3Y145_SLICE_X3Y145_DQ),
.I3(CLBLM_R_X5Y144_SLICE_X6Y144_AQ),
.I4(CLBLL_L_X2Y148_SLICE_X0Y148_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y144_SLICE_X3Y144_AO5),
.O6(CLBLM_R_X3Y144_SLICE_X3Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y145_SLICE_X2Y145_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y145_SLICE_X2Y145_BO5),
.Q(CLBLM_R_X3Y145_SLICE_X2Y145_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y145_SLICE_X2Y145_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y145_SLICE_X2Y145_CO5),
.Q(CLBLM_R_X3Y145_SLICE_X2Y145_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y145_SLICE_X2Y145_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y145_SLICE_X2Y145_AO6),
.Q(CLBLM_R_X3Y145_SLICE_X2Y145_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y145_SLICE_X2Y145_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y145_SLICE_X2Y145_BO6),
.Q(CLBLM_R_X3Y145_SLICE_X2Y145_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y145_SLICE_X2Y145_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y145_SLICE_X2Y145_CO6),
.Q(CLBLM_R_X3Y145_SLICE_X2Y145_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y145_SLICE_X2Y145_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y145_SLICE_X2Y145_DO6),
.Q(CLBLM_R_X3Y145_SLICE_X2Y145_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff5ff0000f50000)
  ) CLBLM_R_X3Y145_SLICE_X2Y145_DLUT (
.I0(CLBLM_R_X3Y143_SLICE_X2Y143_AQ),
.I1(1'b1),
.I2(CLBLM_R_X3Y145_SLICE_X2Y145_DQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X3Y146_SLICE_X2Y146_B5Q),
.I5(CLBLL_L_X2Y153_SLICE_X1Y153_AQ),
.O5(CLBLM_R_X3Y145_SLICE_X2Y145_DO5),
.O6(CLBLM_R_X3Y145_SLICE_X2Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'heeee4444f5a0f5a0)
  ) CLBLM_R_X3Y145_SLICE_X2Y145_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X3Y145_SLICE_X2Y145_B5Q),
.I2(CLBLM_R_X5Y146_SLICE_X6Y146_AQ),
.I3(CLBLM_R_X5Y144_SLICE_X6Y144_D5Q),
.I4(CLBLL_L_X2Y145_SLICE_X1Y145_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X3Y145_SLICE_X2Y145_CO5),
.O6(CLBLM_R_X3Y145_SLICE_X2Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccaaaaff00aaaa)
  ) CLBLM_R_X3Y145_SLICE_X2Y145_BLUT (
.I0(CLBLM_R_X3Y146_SLICE_X2Y146_CQ),
.I1(CLBLL_L_X4Y148_SLICE_X4Y148_A5Q),
.I2(1'b1),
.I3(CLBLL_L_X4Y148_SLICE_X5Y148_CQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y145_SLICE_X2Y145_BO5),
.O6(CLBLM_R_X3Y145_SLICE_X2Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaf3aaf3aaf3aa00)
  ) CLBLM_R_X3Y145_SLICE_X2Y145_ALUT (
.I0(CLBLM_R_X3Y146_SLICE_X2Y146_B5Q),
.I1(CLBLM_R_X3Y148_SLICE_X2Y148_D5Q),
.I2(CLBLM_R_X5Y144_SLICE_X6Y144_DQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X3Y144_SLICE_X2Y144_AQ),
.I5(CLBLM_R_X3Y145_SLICE_X2Y145_AQ),
.O5(CLBLM_R_X3Y145_SLICE_X2Y145_AO5),
.O6(CLBLM_R_X3Y145_SLICE_X2Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y145_SLICE_X3Y145_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y145_SLICE_X3Y145_AO5),
.Q(CLBLM_R_X3Y145_SLICE_X3Y145_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y145_SLICE_X3Y145_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y145_SLICE_X3Y145_AO6),
.Q(CLBLM_R_X3Y145_SLICE_X3Y145_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y145_SLICE_X3Y145_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y145_SLICE_X3Y145_BO6),
.Q(CLBLM_R_X3Y145_SLICE_X3Y145_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y145_SLICE_X3Y145_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y145_SLICE_X3Y145_CO6),
.Q(CLBLM_R_X3Y145_SLICE_X3Y145_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y145_SLICE_X3Y145_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y145_SLICE_X3Y145_DO6),
.Q(CLBLM_R_X3Y145_SLICE_X3Y145_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbbbb8b888bb88b8)
  ) CLBLM_R_X3Y145_SLICE_X3Y145_DLUT (
.I0(CLBLM_R_X3Y147_SLICE_X2Y147_AQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X3Y145_SLICE_X3Y145_DQ),
.I3(CLBLM_R_X5Y149_SLICE_X7Y149_DQ),
.I4(CLBLL_L_X2Y145_SLICE_X1Y145_A5Q),
.I5(CLBLM_L_X8Y142_SLICE_X11Y142_CQ),
.O5(CLBLM_R_X3Y145_SLICE_X3Y145_DO5),
.O6(CLBLM_R_X3Y145_SLICE_X3Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccceeee0000aaaa)
  ) CLBLM_R_X3Y145_SLICE_X3Y145_CLUT (
.I0(CLBLM_R_X3Y143_SLICE_X3Y143_BO6),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X3Y145_SLICE_X3Y145_CQ),
.I5(CLBLM_R_X3Y151_SLICE_X2Y151_BQ),
.O5(CLBLM_R_X3Y145_SLICE_X3Y145_CO5),
.O6(CLBLM_R_X3Y145_SLICE_X3Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hddcc5500eeccaa00)
  ) CLBLM_R_X3Y145_SLICE_X3Y145_BLUT (
.I0(CLBLM_R_X3Y145_SLICE_X3Y145_CQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(1'b1),
.I3(CLBLM_R_X3Y143_SLICE_X3Y143_BO6),
.I4(CLBLM_R_X11Y147_SLICE_X14Y147_AQ),
.I5(CLBLM_R_X3Y145_SLICE_X3Y145_BQ),
.O5(CLBLM_R_X3Y145_SLICE_X3Y145_BO5),
.O6(CLBLM_R_X3Y145_SLICE_X3Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88bbbb88fcfc3030)
  ) CLBLM_R_X3Y145_SLICE_X3Y145_ALUT (
.I0(CLBLM_R_X3Y146_SLICE_X3Y146_BQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X3Y146_SLICE_X3Y146_AQ),
.I3(CLBLL_L_X4Y150_SLICE_X5Y150_CQ),
.I4(CLBLL_L_X4Y141_SLICE_X4Y141_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y145_SLICE_X3Y145_AO5),
.O6(CLBLM_R_X3Y145_SLICE_X3Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y146_SLICE_X2Y146_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y146_SLICE_X2Y146_BO5),
.Q(CLBLM_R_X3Y146_SLICE_X2Y146_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y146_SLICE_X2Y146_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y146_SLICE_X2Y146_CO5),
.Q(CLBLM_R_X3Y146_SLICE_X2Y146_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y146_SLICE_X2Y146_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y146_SLICE_X2Y146_AO6),
.Q(CLBLM_R_X3Y146_SLICE_X2Y146_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y146_SLICE_X2Y146_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y146_SLICE_X2Y146_BO6),
.Q(CLBLM_R_X3Y146_SLICE_X2Y146_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y146_SLICE_X2Y146_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y146_SLICE_X2Y146_CO6),
.Q(CLBLM_R_X3Y146_SLICE_X2Y146_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00aa00aa00aa00aa)
  ) CLBLM_R_X3Y146_SLICE_X2Y146_DLUT (
.I0(CLBLL_L_X4Y150_SLICE_X5Y150_CQ),
.I1(1'b1),
.I2(1'b1),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y146_SLICE_X2Y146_DO5),
.O6(CLBLM_R_X3Y146_SLICE_X2Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0aaf0aaccffcc00)
  ) CLBLM_R_X3Y146_SLICE_X2Y146_CLUT (
.I0(CLBLM_R_X3Y145_SLICE_X2Y145_C5Q),
.I1(CLBLM_R_X3Y145_SLICE_X3Y145_A5Q),
.I2(CLBLM_R_X3Y150_SLICE_X2Y150_B5Q),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(RIOB33_X105Y121_IOB_X1Y122_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y146_SLICE_X2Y146_CO5),
.O6(CLBLM_R_X3Y146_SLICE_X2Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff33cc00e2e2e2e2)
  ) CLBLM_R_X3Y146_SLICE_X2Y146_BLUT (
.I0(LIOB33_X0Y59_IOB_X0Y59_I),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X3Y146_SLICE_X2Y146_AQ),
.I3(CLBLM_R_X3Y147_SLICE_X2Y147_BQ),
.I4(CLBLL_L_X4Y143_SLICE_X5Y143_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X3Y146_SLICE_X2Y146_BO5),
.O6(CLBLM_R_X3Y146_SLICE_X2Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heeffeafa44554050)
  ) CLBLM_R_X3Y146_SLICE_X2Y146_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X5Y144_SLICE_X6Y144_DQ),
.I2(CLBLM_R_X3Y146_SLICE_X2Y146_AQ),
.I3(CLBLM_R_X3Y148_SLICE_X2Y148_D5Q),
.I4(CLBLL_L_X2Y144_SLICE_X0Y144_AQ),
.I5(CLBLM_R_X3Y151_SLICE_X3Y151_AQ),
.O5(CLBLM_R_X3Y146_SLICE_X2Y146_AO5),
.O6(CLBLM_R_X3Y146_SLICE_X2Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y146_SLICE_X3Y146_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y146_SLICE_X3Y146_CO5),
.Q(CLBLM_R_X3Y146_SLICE_X3Y146_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y146_SLICE_X3Y146_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y146_SLICE_X3Y146_AO6),
.Q(CLBLM_R_X3Y146_SLICE_X3Y146_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y146_SLICE_X3Y146_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y146_SLICE_X3Y146_BO6),
.Q(CLBLM_R_X3Y146_SLICE_X3Y146_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y146_SLICE_X3Y146_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y146_SLICE_X3Y146_CO6),
.Q(CLBLM_R_X3Y146_SLICE_X3Y146_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y146_SLICE_X3Y146_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y146_SLICE_X3Y146_DO6),
.Q(CLBLM_R_X3Y146_SLICE_X3Y146_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000c8fac8fa)
  ) CLBLM_R_X3Y146_SLICE_X3Y146_DLUT (
.I0(CLBLL_L_X2Y144_SLICE_X1Y144_A5Q),
.I1(CLBLM_L_X8Y142_SLICE_X11Y142_CQ),
.I2(CLBLM_R_X3Y146_SLICE_X3Y146_DQ),
.I3(CLBLM_R_X5Y149_SLICE_X7Y149_DQ),
.I4(CLBLM_R_X3Y147_SLICE_X2Y147_CQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X3Y146_SLICE_X3Y146_DO5),
.O6(CLBLM_R_X3Y146_SLICE_X3Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcc00ccf0aaf0aa)
  ) CLBLM_R_X3Y146_SLICE_X3Y146_CLUT (
.I0(CLBLM_R_X5Y143_SLICE_X6Y143_DQ),
.I1(CLBLM_R_X5Y149_SLICE_X6Y149_AQ),
.I2(CLBLM_R_X3Y145_SLICE_X3Y145_BQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLL_L_X4Y143_SLICE_X5Y143_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X3Y146_SLICE_X3Y146_CO5),
.O6(CLBLM_R_X3Y146_SLICE_X3Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0cceef0f0cc44)
  ) CLBLM_R_X3Y146_SLICE_X3Y146_BLUT (
.I0(CLBLM_R_X7Y150_SLICE_X9Y150_CQ),
.I1(CLBLM_R_X3Y146_SLICE_X3Y146_BQ),
.I2(CLBLL_L_X2Y144_SLICE_X0Y144_AQ),
.I3(CLBLM_L_X8Y146_SLICE_X10Y146_AQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X3Y148_SLICE_X2Y148_CQ),
.O5(CLBLM_R_X3Y146_SLICE_X3Y146_BO5),
.O6(CLBLM_R_X3Y146_SLICE_X3Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff005050ff000505)
  ) CLBLM_R_X3Y146_SLICE_X3Y146_ALUT (
.I0(CLBLM_R_X3Y146_SLICE_X3Y146_CQ),
.I1(1'b1),
.I2(CLBLM_R_X3Y146_SLICE_X3Y146_AQ),
.I3(CLBLM_R_X7Y142_SLICE_X9Y142_D5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X3Y147_SLICE_X3Y147_CO6),
.O5(CLBLM_R_X3Y146_SLICE_X3Y146_AO5),
.O6(CLBLM_R_X3Y146_SLICE_X3Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y147_SLICE_X2Y147_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y147_SLICE_X2Y147_CO5),
.Q(CLBLM_R_X3Y147_SLICE_X2Y147_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y147_SLICE_X2Y147_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y147_SLICE_X2Y147_AO6),
.Q(CLBLM_R_X3Y147_SLICE_X2Y147_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y147_SLICE_X2Y147_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y147_SLICE_X2Y147_BO6),
.Q(CLBLM_R_X3Y147_SLICE_X2Y147_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y147_SLICE_X2Y147_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y147_SLICE_X2Y147_CO6),
.Q(CLBLM_R_X3Y147_SLICE_X2Y147_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f3f3f3ebc3aa00)
  ) CLBLM_R_X3Y147_SLICE_X2Y147_DLUT (
.I0(CLBLM_R_X11Y147_SLICE_X15Y147_AQ),
.I1(CLBLM_R_X3Y147_SLICE_X3Y147_A5Q),
.I2(CLBLM_R_X3Y150_SLICE_X3Y150_BQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X5Y153_SLICE_X7Y153_BO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y147_SLICE_X2Y147_DO5),
.O6(CLBLM_R_X3Y147_SLICE_X2Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hb8b8b8b8ffcc3300)
  ) CLBLM_R_X3Y147_SLICE_X2Y147_CLUT (
.I0(CLBLM_R_X3Y151_SLICE_X2Y151_AQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLM_R_X5Y147_SLICE_X7Y147_AQ),
.I4(CLBLM_R_X3Y146_SLICE_X3Y146_DQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y147_SLICE_X2Y147_CO5),
.O6(CLBLM_R_X3Y147_SLICE_X2Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcf6cc66f0f00000)
  ) CLBLM_R_X3Y147_SLICE_X2Y147_BLUT (
.I0(CLBLM_R_X3Y147_SLICE_X3Y147_A5Q),
.I1(CLBLM_R_X3Y147_SLICE_X2Y147_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X3Y150_SLICE_X3Y150_BQ),
.I4(CLBLM_R_X3Y146_SLICE_X2Y146_C5Q),
.I5(CLBLM_R_X5Y153_SLICE_X7Y153_BO6),
.O5(CLBLM_R_X3Y147_SLICE_X2Y147_BO5),
.O6(CLBLM_R_X3Y147_SLICE_X2Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffb400b400b400)
  ) CLBLM_R_X3Y147_SLICE_X2Y147_ALUT (
.I0(CLBLM_R_X3Y147_SLICE_X2Y147_DO6),
.I1(CLBLM_R_X3Y147_SLICE_X2Y147_BQ),
.I2(CLBLM_R_X3Y147_SLICE_X2Y147_AQ),
.I3(CLBLM_R_X5Y153_SLICE_X7Y153_BO6),
.I4(CLBLM_R_X7Y144_SLICE_X8Y144_BQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X3Y147_SLICE_X2Y147_AO5),
.O6(CLBLM_R_X3Y147_SLICE_X2Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y147_SLICE_X3Y147_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y147_SLICE_X2Y147_DO5),
.Q(CLBLM_R_X3Y147_SLICE_X3Y147_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y147_SLICE_X3Y147_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y147_SLICE_X3Y147_BO5),
.Q(CLBLM_R_X3Y147_SLICE_X3Y147_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y147_SLICE_X3Y147_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y147_SLICE_X3Y147_AO6),
.Q(CLBLM_R_X3Y147_SLICE_X3Y147_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y147_SLICE_X3Y147_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y147_SLICE_X3Y147_BO6),
.Q(CLBLM_R_X3Y147_SLICE_X3Y147_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff7f008000000000)
  ) CLBLM_R_X3Y147_SLICE_X3Y147_DLUT (
.I0(CLBLM_R_X3Y147_SLICE_X2Y147_AQ),
.I1(CLBLM_R_X3Y147_SLICE_X2Y147_BQ),
.I2(CLBLM_R_X3Y147_SLICE_X3Y147_A5Q),
.I3(CLBLM_R_X3Y150_SLICE_X3Y150_BQ),
.I4(CLBLM_R_X3Y144_SLICE_X3Y144_AQ),
.I5(CLBLM_R_X5Y153_SLICE_X7Y153_BO6),
.O5(CLBLM_R_X3Y147_SLICE_X3Y147_DO5),
.O6(CLBLM_R_X3Y147_SLICE_X3Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3fff3fff77ffffff)
  ) CLBLM_R_X3Y147_SLICE_X3Y147_CLUT (
.I0(CLBLM_R_X3Y148_SLICE_X2Y148_AQ),
.I1(CLBLL_L_X4Y147_SLICE_X4Y147_BQ),
.I2(CLBLL_L_X4Y148_SLICE_X4Y148_CO6),
.I3(CLBLM_R_X3Y147_SLICE_X3Y147_AQ),
.I4(CLBLM_R_X3Y146_SLICE_X3Y146_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y147_SLICE_X3Y147_CO5),
.O6(CLBLM_R_X3Y147_SLICE_X3Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcc00ccf055f055)
  ) CLBLM_R_X3Y147_SLICE_X3Y147_BLUT (
.I0(CLBLM_R_X3Y147_SLICE_X3Y147_B5Q),
.I1(CLBLM_R_X5Y144_SLICE_X6Y144_CQ),
.I2(CLBLM_L_X10Y147_SLICE_X13Y147_DQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X5Y147_SLICE_X6Y147_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y147_SLICE_X3Y147_BO5),
.O6(CLBLM_R_X3Y147_SLICE_X3Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaf3aaffaafcaaff)
  ) CLBLM_R_X3Y147_SLICE_X3Y147_ALUT (
.I0(CLBLL_L_X2Y147_SLICE_X0Y147_BQ),
.I1(CLBLL_L_X4Y148_SLICE_X4Y148_CO6),
.I2(CLBLM_R_X3Y146_SLICE_X3Y146_CQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X3Y147_SLICE_X3Y147_CO5),
.I5(CLBLM_R_X3Y147_SLICE_X3Y147_AQ),
.O5(CLBLM_R_X3Y147_SLICE_X3Y147_AO5),
.O6(CLBLM_R_X3Y147_SLICE_X3Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y148_SLICE_X2Y148_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y148_SLICE_X2Y148_BO5),
.Q(CLBLM_R_X3Y148_SLICE_X2Y148_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y148_SLICE_X2Y148_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y148_SLICE_X2Y148_CO5),
.Q(CLBLM_R_X3Y148_SLICE_X2Y148_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y148_SLICE_X2Y148_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y148_SLICE_X2Y148_DO5),
.Q(CLBLM_R_X3Y148_SLICE_X2Y148_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y148_SLICE_X2Y148_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y148_SLICE_X2Y148_AO6),
.Q(CLBLM_R_X3Y148_SLICE_X2Y148_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y148_SLICE_X2Y148_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y148_SLICE_X2Y148_BO6),
.Q(CLBLM_R_X3Y148_SLICE_X2Y148_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y148_SLICE_X2Y148_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y148_SLICE_X2Y148_CO6),
.Q(CLBLM_R_X3Y148_SLICE_X2Y148_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y148_SLICE_X2Y148_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y148_SLICE_X2Y148_DO6),
.Q(CLBLM_R_X3Y148_SLICE_X2Y148_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaccaaccccffcc00)
  ) CLBLM_R_X3Y148_SLICE_X2Y148_DLUT (
.I0(CLBLM_R_X3Y144_SLICE_X3Y144_D5Q),
.I1(CLBLL_L_X4Y147_SLICE_X4Y147_BQ),
.I2(1'b1),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X5Y144_SLICE_X6Y144_DQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y148_SLICE_X2Y148_DO5),
.O6(CLBLM_R_X3Y148_SLICE_X2Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaccccccccff00)
  ) CLBLM_R_X3Y148_SLICE_X2Y148_CLUT (
.I0(CLBLM_R_X3Y150_SLICE_X3Y150_AQ),
.I1(CLBLM_R_X3Y148_SLICE_X2Y148_AQ),
.I2(1'b1),
.I3(CLBLM_R_X11Y146_SLICE_X14Y146_BO6),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y148_SLICE_X2Y148_CO5),
.O6(CLBLM_R_X3Y148_SLICE_X2Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaa5500e4e4e4e4)
  ) CLBLM_R_X3Y148_SLICE_X2Y148_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLL_L_X4Y152_SLICE_X4Y152_CQ),
.I2(CLBLM_R_X3Y147_SLICE_X3Y147_A5Q),
.I3(CLBLM_R_X3Y149_SLICE_X2Y149_A5Q),
.I4(CLBLM_R_X3Y142_SLICE_X2Y142_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X3Y148_SLICE_X2Y148_BO5),
.O6(CLBLM_R_X3Y148_SLICE_X2Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0000eded2121)
  ) CLBLM_R_X3Y148_SLICE_X2Y148_ALUT (
.I0(CLBLM_R_X3Y148_SLICE_X3Y148_CO6),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X3Y148_SLICE_X2Y148_AQ),
.I3(1'b1),
.I4(CLBLL_L_X2Y149_SLICE_X1Y149_DQ),
.I5(CLBLM_R_X3Y146_SLICE_X3Y146_CQ),
.O5(CLBLM_R_X3Y148_SLICE_X2Y148_AO5),
.O6(CLBLM_R_X3Y148_SLICE_X2Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y148_SLICE_X3Y148_A5_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y148_SLICE_X3Y148_AO5),
.Q(CLBLM_R_X3Y148_SLICE_X3Y148_A5Q),
.S(CLBLM_R_X3Y146_SLICE_X2Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y148_SLICE_X3Y148_A_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y148_SLICE_X3Y148_AO6),
.Q(CLBLM_R_X3Y148_SLICE_X3Y148_AQ),
.S(CLBLM_R_X3Y146_SLICE_X2Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3d1c0e2f3f3c0c0)
  ) CLBLM_R_X3Y148_SLICE_X3Y148_DLUT (
.I0(CLBLM_R_X7Y147_SLICE_X9Y147_AQ),
.I1(CLBLM_L_X8Y149_SLICE_X11Y149_BQ),
.I2(CLBLL_L_X4Y147_SLICE_X5Y147_CQ),
.I3(CLBLM_R_X7Y142_SLICE_X8Y142_DO6),
.I4(CLBLL_L_X2Y148_SLICE_X0Y148_A5Q),
.I5(CLBLL_L_X4Y143_SLICE_X5Y143_AQ),
.O5(CLBLM_R_X3Y148_SLICE_X3Y148_DO5),
.O6(CLBLM_R_X3Y148_SLICE_X3Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7f7fffff006600aa)
  ) CLBLM_R_X3Y148_SLICE_X3Y148_CLUT (
.I0(CLBLL_L_X4Y147_SLICE_X4Y147_BQ),
.I1(CLBLM_R_X3Y147_SLICE_X3Y147_AQ),
.I2(CLBLM_R_X3Y146_SLICE_X3Y146_AQ),
.I3(CLBLM_R_X3Y146_SLICE_X3Y146_CQ),
.I4(CLBLL_L_X4Y148_SLICE_X4Y148_CO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y148_SLICE_X3Y148_CO5),
.O6(CLBLM_R_X3Y148_SLICE_X3Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hdfffffff5fffffff)
  ) CLBLM_R_X3Y148_SLICE_X3Y148_BLUT (
.I0(CLBLM_R_X3Y144_SLICE_X3Y144_AQ),
.I1(CLBLM_R_X3Y150_SLICE_X3Y150_BQ),
.I2(CLBLM_R_X3Y147_SLICE_X2Y147_AQ),
.I3(CLBLM_R_X3Y147_SLICE_X2Y147_BQ),
.I4(CLBLM_R_X3Y147_SLICE_X3Y147_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X3Y148_SLICE_X3Y148_BO5),
.O6(CLBLM_R_X3Y148_SLICE_X3Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00000cccc0000)
  ) CLBLM_R_X3Y148_SLICE_X3Y148_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y150_SLICE_X6Y150_BQ),
.I2(CLBLM_R_X5Y144_SLICE_X6Y144_C5Q),
.I3(1'b1),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y148_SLICE_X3Y148_AO5),
.O6(CLBLM_R_X3Y148_SLICE_X3Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y149_SLICE_X2Y149_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y149_SLICE_X2Y149_AO5),
.Q(CLBLM_R_X3Y149_SLICE_X2Y149_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y149_SLICE_X2Y149_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y149_SLICE_X2Y149_AO6),
.Q(CLBLM_R_X3Y149_SLICE_X2Y149_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y149_SLICE_X2Y149_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y149_SLICE_X2Y149_BO6),
.Q(CLBLM_R_X3Y149_SLICE_X2Y149_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y149_SLICE_X2Y149_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y149_SLICE_X2Y149_CO6),
.Q(CLBLM_R_X3Y149_SLICE_X2Y149_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f000f000f000f00)
  ) CLBLM_R_X3Y149_SLICE_X2Y149_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X5Y149_SLICE_X6Y149_A5Q),
.I3(CLBLM_R_X5Y151_SLICE_X6Y151_B5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y149_SLICE_X2Y149_DO5),
.O6(CLBLM_R_X3Y149_SLICE_X2Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h888888d8888888d8)
  ) CLBLM_R_X3Y149_SLICE_X2Y149_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X3Y147_SLICE_X3Y147_B5Q),
.I2(CLBLL_L_X2Y149_SLICE_X1Y149_BQ),
.I3(CLBLL_L_X2Y149_SLICE_X1Y149_DQ),
.I4(CLBLL_L_X2Y149_SLICE_X1Y149_CQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y149_SLICE_X2Y149_CO5),
.O6(CLBLM_R_X3Y149_SLICE_X2Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0cacac0c0c0c0)
  ) CLBLM_R_X3Y149_SLICE_X2Y149_BLUT (
.I0(CLBLL_L_X2Y149_SLICE_X1Y149_CQ),
.I1(CLBLM_R_X7Y150_SLICE_X8Y150_D5Q),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(1'b1),
.I4(CLBLL_L_X2Y149_SLICE_X1Y149_BQ),
.I5(CLBLL_L_X2Y149_SLICE_X1Y149_DQ),
.O5(CLBLM_R_X3Y149_SLICE_X2Y149_BO5),
.O6(CLBLM_R_X3Y149_SLICE_X2Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heeee4444f5a0f5a0)
  ) CLBLM_R_X3Y149_SLICE_X2Y149_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X5Y150_SLICE_X6Y150_A5Q),
.I2(CLBLM_R_X3Y149_SLICE_X2Y149_AQ),
.I3(CLBLM_L_X8Y152_SLICE_X10Y152_DQ),
.I4(CLBLM_R_X7Y153_SLICE_X9Y153_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X3Y149_SLICE_X2Y149_AO5),
.O6(CLBLM_R_X3Y149_SLICE_X2Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y149_SLICE_X3Y149_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y149_SLICE_X3Y149_AO6),
.Q(CLBLM_R_X3Y149_SLICE_X3Y149_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y149_SLICE_X3Y149_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y149_SLICE_X3Y149_BO6),
.Q(CLBLM_R_X3Y149_SLICE_X3Y149_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y149_SLICE_X3Y149_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y149_SLICE_X3Y149_CO6),
.Q(CLBLM_R_X3Y149_SLICE_X3Y149_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y149_SLICE_X3Y149_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y149_SLICE_X3Y149_DO6),
.Q(CLBLM_R_X3Y149_SLICE_X3Y149_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000077777777)
  ) CLBLM_R_X3Y149_SLICE_X3Y149_DLUT (
.I0(CLBLL_L_X4Y147_SLICE_X4Y147_AQ),
.I1(CLBLM_R_X3Y150_SLICE_X3Y150_DO6),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X7Y143_SLICE_X8Y143_DQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X3Y149_SLICE_X3Y149_DO5),
.O6(CLBLM_R_X3Y149_SLICE_X3Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffefaaea55450040)
  ) CLBLM_R_X3Y149_SLICE_X3Y149_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLL_L_X4Y147_SLICE_X5Y147_B5Q),
.I2(CLBLM_R_X7Y150_SLICE_X9Y150_CQ),
.I3(CLBLM_L_X8Y146_SLICE_X10Y146_AQ),
.I4(CLBLM_R_X3Y149_SLICE_X3Y149_CQ),
.I5(CLBLM_R_X3Y149_SLICE_X3Y149_AQ),
.O5(CLBLM_R_X3Y149_SLICE_X3Y149_CO5),
.O6(CLBLM_R_X3Y149_SLICE_X3Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00a8a8fcfc)
  ) CLBLM_R_X3Y149_SLICE_X3Y149_BLUT (
.I0(CLBLM_R_X5Y144_SLICE_X6Y144_CQ),
.I1(CLBLM_R_X3Y149_SLICE_X3Y149_BQ),
.I2(CLBLM_R_X3Y148_SLICE_X3Y148_AQ),
.I3(CLBLM_R_X5Y148_SLICE_X7Y148_AQ),
.I4(CLBLM_R_X3Y147_SLICE_X3Y147_BQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X3Y149_SLICE_X3Y149_BO5),
.O6(CLBLM_R_X3Y149_SLICE_X3Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff848484ff848484)
  ) CLBLM_R_X3Y149_SLICE_X3Y149_ALUT (
.I0(CLBLM_R_X3Y152_SLICE_X3Y152_DO6),
.I1(CLBLM_R_X5Y153_SLICE_X7Y153_BO6),
.I2(CLBLM_R_X3Y149_SLICE_X3Y149_AQ),
.I3(CLBLL_L_X4Y147_SLICE_X4Y147_AQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y149_SLICE_X3Y149_AO5),
.O6(CLBLM_R_X3Y149_SLICE_X3Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y150_SLICE_X2Y150_B5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X3Y150_SLICE_X2Y150_BO5),
.Q(CLBLM_R_X3Y150_SLICE_X2Y150_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y150_SLICE_X2Y150_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X3Y150_SLICE_X2Y150_AO6),
.Q(CLBLM_R_X3Y150_SLICE_X2Y150_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y150_SLICE_X2Y150_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X3Y150_SLICE_X2Y150_BO6),
.Q(CLBLM_R_X3Y150_SLICE_X2Y150_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y150_SLICE_X2Y150_D_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X3Y150_SLICE_X2Y150_DO6),
.Q(CLBLM_R_X3Y150_SLICE_X2Y150_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00a5a5ff000000)
  ) CLBLM_R_X3Y150_SLICE_X2Y150_DLUT (
.I0(CLBLM_R_X5Y150_SLICE_X7Y150_BO6),
.I1(1'b1),
.I2(CLBLM_R_X3Y150_SLICE_X2Y150_DQ),
.I3(CLBLM_R_X3Y144_SLICE_X3Y144_A5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X3Y152_SLICE_X2Y152_BQ),
.O5(CLBLM_R_X3Y150_SLICE_X2Y150_DO5),
.O6(CLBLM_R_X3Y150_SLICE_X2Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00000ffffffee)
  ) CLBLM_R_X3Y150_SLICE_X2Y150_CLUT (
.I0(CLBLM_R_X3Y150_SLICE_X2Y150_BQ),
.I1(CLBLL_L_X4Y153_SLICE_X4Y153_A5Q),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLL_L_X2Y150_SLICE_X1Y150_BO5),
.I4(CLBLL_L_X2Y150_SLICE_X1Y150_CQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y150_SLICE_X2Y150_CO5),
.O6(CLBLM_R_X3Y150_SLICE_X2Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcc00ccf0aaf0aa)
  ) CLBLM_R_X3Y150_SLICE_X2Y150_BLUT (
.I0(CLBLM_R_X5Y152_SLICE_X6Y152_CQ),
.I1(CLBLL_L_X4Y154_SLICE_X4Y154_AQ),
.I2(CLBLM_R_X3Y150_SLICE_X2Y150_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X3Y148_SLICE_X3Y148_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y150_SLICE_X2Y150_BO5),
.O6(CLBLM_R_X3Y150_SLICE_X2Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccfffafffa)
  ) CLBLM_R_X3Y150_SLICE_X2Y150_ALUT (
.I0(CLBLM_L_X8Y153_SLICE_X11Y153_BQ),
.I1(CLBLM_R_X3Y150_SLICE_X2Y150_BQ),
.I2(CLBLM_R_X11Y150_SLICE_X14Y150_CO6),
.I3(CLBLM_L_X8Y148_SLICE_X10Y148_DO6),
.I4(1'b1),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X3Y150_SLICE_X2Y150_AO5),
.O6(CLBLM_R_X3Y150_SLICE_X2Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y150_SLICE_X3Y150_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.Q(CLBLM_R_X3Y150_SLICE_X3Y150_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y150_SLICE_X3Y150_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X3Y150_SLICE_X3Y150_BO6),
.Q(CLBLM_R_X3Y150_SLICE_X3Y150_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y150_SLICE_X3Y150_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X3Y150_SLICE_X3Y150_CO6),
.Q(CLBLM_R_X3Y150_SLICE_X3Y150_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hee00ee00ffffffff)
  ) CLBLM_R_X3Y150_SLICE_X3Y150_DLUT (
.I0(CLBLM_R_X3Y152_SLICE_X2Y152_AQ),
.I1(CLBLM_R_X3Y150_SLICE_X3Y150_CQ),
.I2(1'b1),
.I3(CLBLL_L_X4Y150_SLICE_X4Y150_CO6),
.I4(1'b1),
.I5(CLBLM_R_X3Y152_SLICE_X2Y152_BQ),
.O5(CLBLM_R_X3Y150_SLICE_X3Y150_DO5),
.O6(CLBLM_R_X3Y150_SLICE_X3Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0a0aca0ac)
  ) CLBLM_R_X3Y150_SLICE_X3Y150_CLUT (
.I0(CLBLM_R_X5Y148_SLICE_X6Y148_BQ),
.I1(CLBLM_R_X7Y152_SLICE_X8Y152_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X7Y144_SLICE_X9Y144_AQ),
.I4(1'b1),
.I5(CLBLL_L_X4Y150_SLICE_X4Y150_AO5),
.O5(CLBLM_R_X3Y150_SLICE_X3Y150_CO5),
.O6(CLBLM_R_X3Y150_SLICE_X3Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0044444c4c)
  ) CLBLM_R_X3Y150_SLICE_X3Y150_BLUT (
.I0(CLBLL_L_X4Y150_SLICE_X4Y150_CO6),
.I1(CLBLM_R_X3Y152_SLICE_X2Y152_BQ),
.I2(CLBLM_R_X3Y150_SLICE_X3Y150_CQ),
.I3(CLBLM_L_X10Y148_SLICE_X12Y148_AQ),
.I4(CLBLM_R_X3Y152_SLICE_X2Y152_AQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X3Y150_SLICE_X3Y150_BO5),
.O6(CLBLM_R_X3Y150_SLICE_X3Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff005f5f5f5f)
  ) CLBLM_R_X3Y150_SLICE_X3Y150_ALUT (
.I0(CLBLL_L_X4Y150_SLICE_X4Y150_CO6),
.I1(1'b1),
.I2(CLBLM_R_X3Y150_SLICE_X3Y150_CQ),
.I3(CLBLL_L_X4Y149_SLICE_X4Y149_BQ),
.I4(1'b1),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X3Y150_SLICE_X3Y150_AO5),
.O6(CLBLM_R_X3Y150_SLICE_X3Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y151_SLICE_X2Y151_A5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X3Y151_SLICE_X2Y151_CO5),
.Q(CLBLM_R_X3Y151_SLICE_X2Y151_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y151_SLICE_X2Y151_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X3Y151_SLICE_X2Y151_AO6),
.Q(CLBLM_R_X3Y151_SLICE_X2Y151_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y151_SLICE_X2Y151_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X3Y151_SLICE_X2Y151_BO6),
.Q(CLBLM_R_X3Y151_SLICE_X2Y151_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8ffff0000ffff000)
  ) CLBLM_R_X3Y151_SLICE_X2Y151_DLUT (
.I0(LIOB33_X0Y55_IOB_X0Y55_I),
.I1(CLBLM_R_X3Y151_SLICE_X2Y151_AQ),
.I2(CLBLM_R_X3Y147_SLICE_X3Y147_B5Q),
.I3(CLBLM_R_X3Y151_SLICE_X2Y151_A5Q),
.I4(CLBLM_R_X3Y151_SLICE_X3Y151_DQ),
.I5(CLBLL_L_X2Y151_SLICE_X1Y151_AQ),
.O5(CLBLM_R_X3Y151_SLICE_X2Y151_DO5),
.O6(CLBLM_R_X3Y151_SLICE_X2Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0fffffff8bb88bb8)
  ) CLBLM_R_X3Y151_SLICE_X2Y151_CLUT (
.I0(CLBLM_R_X7Y152_SLICE_X8Y152_AQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X3Y147_SLICE_X3Y147_B5Q),
.I3(CLBLM_R_X3Y151_SLICE_X2Y151_A5Q),
.I4(CLBLM_R_X3Y151_SLICE_X3Y151_DQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y151_SLICE_X2Y151_CO5),
.O6(CLBLM_R_X3Y151_SLICE_X2Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff008c8cdcdc)
  ) CLBLM_R_X3Y151_SLICE_X2Y151_BLUT (
.I0(CLBLM_R_X3Y143_SLICE_X2Y143_AQ),
.I1(CLBLL_L_X4Y149_SLICE_X5Y149_CQ),
.I2(CLBLM_R_X3Y145_SLICE_X2Y145_DQ),
.I3(CLBLM_R_X7Y152_SLICE_X9Y152_BQ),
.I4(CLBLM_R_X3Y148_SLICE_X2Y148_C5Q),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X3Y151_SLICE_X2Y151_BO5),
.O6(CLBLM_R_X3Y151_SLICE_X2Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccf0f0cccc0ff0)
  ) CLBLM_R_X3Y151_SLICE_X2Y151_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y150_SLICE_X6Y150_A5Q),
.I2(CLBLM_R_X3Y151_SLICE_X2Y151_AQ),
.I3(CLBLL_L_X2Y151_SLICE_X1Y151_AQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X3Y151_SLICE_X2Y151_CO6),
.O5(CLBLM_R_X3Y151_SLICE_X2Y151_AO5),
.O6(CLBLM_R_X3Y151_SLICE_X2Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y151_SLICE_X3Y151_C5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X3Y151_SLICE_X3Y151_CO5),
.Q(CLBLM_R_X3Y151_SLICE_X3Y151_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y151_SLICE_X3Y151_D5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X3Y151_SLICE_X3Y151_DO5),
.Q(CLBLM_R_X3Y151_SLICE_X3Y151_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y151_SLICE_X3Y151_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X3Y151_SLICE_X3Y151_AO6),
.Q(CLBLM_R_X3Y151_SLICE_X3Y151_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y151_SLICE_X3Y151_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X3Y151_SLICE_X3Y151_BO6),
.Q(CLBLM_R_X3Y151_SLICE_X3Y151_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y151_SLICE_X3Y151_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X3Y151_SLICE_X3Y151_CO6),
.Q(CLBLM_R_X3Y151_SLICE_X3Y151_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y151_SLICE_X3Y151_D_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X3Y151_SLICE_X3Y151_DO6),
.Q(CLBLM_R_X3Y151_SLICE_X3Y151_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccf0f0aaaa00ff)
  ) CLBLM_R_X3Y151_SLICE_X3Y151_DLUT (
.I0(CLBLM_R_X3Y147_SLICE_X3Y147_BQ),
.I1(CLBLL_L_X4Y147_SLICE_X5Y147_B5Q),
.I2(CLBLM_R_X3Y151_SLICE_X2Y151_DO6),
.I3(CLBLM_L_X12Y149_SLICE_X16Y149_CO6),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y151_SLICE_X3Y151_DO5),
.O6(CLBLM_R_X3Y151_SLICE_X3Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h88dd88dda0a0a0f5)
  ) CLBLM_R_X3Y151_SLICE_X3Y151_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X7Y144_SLICE_X9Y144_AQ),
.I2(CLBLM_R_X5Y145_SLICE_X6Y145_B5Q),
.I3(CLBLM_R_X7Y153_SLICE_X8Y153_DO5),
.I4(CLBLL_L_X4Y154_SLICE_X4Y154_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y151_SLICE_X3Y151_CO5),
.O6(CLBLM_R_X3Y151_SLICE_X3Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00f9f9f0f0)
  ) CLBLM_R_X3Y151_SLICE_X3Y151_BLUT (
.I0(CLBLL_L_X4Y151_SLICE_X4Y151_BO6),
.I1(CLBLM_R_X3Y151_SLICE_X3Y151_BQ),
.I2(CLBLL_L_X2Y148_SLICE_X0Y148_B5Q),
.I3(CLBLL_L_X4Y143_SLICE_X5Y143_AQ),
.I4(CLBLM_R_X3Y150_SLICE_X3Y150_AQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X3Y151_SLICE_X3Y151_BO5),
.O6(CLBLM_R_X3Y151_SLICE_X3Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc5acc00cc00)
  ) CLBLM_R_X3Y151_SLICE_X3Y151_ALUT (
.I0(CLBLL_L_X4Y151_SLICE_X4Y151_BO5),
.I1(CLBLM_R_X5Y148_SLICE_X6Y148_B5Q),
.I2(CLBLM_R_X3Y151_SLICE_X3Y151_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLL_L_X2Y148_SLICE_X0Y148_B5Q),
.I5(CLBLM_R_X3Y150_SLICE_X3Y150_AQ),
.O5(CLBLM_R_X3Y151_SLICE_X3Y151_AO5),
.O6(CLBLM_R_X3Y151_SLICE_X3Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y152_SLICE_X2Y152_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X3Y152_SLICE_X2Y152_AO6),
.Q(CLBLM_R_X3Y152_SLICE_X2Y152_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y152_SLICE_X2Y152_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X3Y152_SLICE_X2Y152_BO6),
.Q(CLBLM_R_X3Y152_SLICE_X2Y152_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y152_SLICE_X2Y152_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X3Y152_SLICE_X2Y152_CO6),
.Q(CLBLM_R_X3Y152_SLICE_X2Y152_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hefffefffffffffff)
  ) CLBLM_R_X3Y152_SLICE_X2Y152_DLUT (
.I0(CLBLM_R_X5Y151_SLICE_X7Y151_BO6),
.I1(CLBLL_L_X4Y150_SLICE_X4Y150_AO5),
.I2(CLBLM_R_X7Y152_SLICE_X8Y152_BQ),
.I3(CLBLL_L_X4Y150_SLICE_X5Y150_CQ),
.I4(1'b1),
.I5(CLBLM_R_X7Y144_SLICE_X9Y144_AQ),
.O5(CLBLM_R_X3Y152_SLICE_X2Y152_DO5),
.O6(CLBLM_R_X3Y152_SLICE_X2Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fff055f0ccf044)
  ) CLBLM_R_X3Y152_SLICE_X2Y152_CLUT (
.I0(CLBLM_R_X3Y148_SLICE_X2Y148_D5Q),
.I1(CLBLM_R_X3Y152_SLICE_X2Y152_CQ),
.I2(CLBLM_R_X7Y152_SLICE_X8Y152_BQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X5Y144_SLICE_X6Y144_DQ),
.I5(CLBLL_L_X2Y144_SLICE_X1Y144_B5Q),
.O5(CLBLM_R_X3Y152_SLICE_X2Y152_CO5),
.O6(CLBLM_R_X3Y152_SLICE_X2Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8bbb8bbb8bbb8bbb)
  ) CLBLM_R_X3Y152_SLICE_X2Y152_BLUT (
.I0(CLBLM_R_X5Y152_SLICE_X7Y152_DQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X3Y152_SLICE_X2Y152_AQ),
.I3(CLBLL_L_X4Y150_SLICE_X4Y150_CO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y152_SLICE_X2Y152_BO5),
.O6(CLBLM_R_X3Y152_SLICE_X2Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c5c0c5c0c0c0c0)
  ) CLBLM_R_X3Y152_SLICE_X2Y152_ALUT (
.I0(CLBLM_R_X7Y152_SLICE_X8Y152_BQ),
.I1(CLBLL_L_X4Y152_SLICE_X4Y152_DQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLL_L_X4Y150_SLICE_X4Y150_AO5),
.I4(1'b1),
.I5(CLBLM_R_X7Y144_SLICE_X9Y144_AQ),
.O5(CLBLM_R_X3Y152_SLICE_X2Y152_AO5),
.O6(CLBLM_R_X3Y152_SLICE_X2Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y152_SLICE_X3Y152_A5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X3Y152_SLICE_X3Y152_AO5),
.Q(CLBLM_R_X3Y152_SLICE_X3Y152_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y152_SLICE_X3Y152_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X3Y152_SLICE_X3Y152_AO6),
.Q(CLBLM_R_X3Y152_SLICE_X3Y152_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffdfffdfff)
  ) CLBLM_R_X3Y152_SLICE_X3Y152_DLUT (
.I0(CLBLM_R_X3Y153_SLICE_X3Y153_AQ),
.I1(CLBLM_R_X3Y148_SLICE_X3Y148_BO5),
.I2(CLBLM_R_X3Y153_SLICE_X3Y153_BQ),
.I3(CLBLL_L_X4Y150_SLICE_X5Y150_D5Q),
.I4(1'b1),
.I5(CLBLM_R_X3Y150_SLICE_X3Y150_BQ),
.O5(CLBLM_R_X3Y152_SLICE_X3Y152_DO5),
.O6(CLBLM_R_X3Y152_SLICE_X3Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000002a80)
  ) CLBLM_R_X3Y152_SLICE_X3Y152_CLUT (
.I0(CLBLM_R_X3Y150_SLICE_X3Y150_AQ),
.I1(CLBLM_R_X7Y144_SLICE_X9Y144_AQ),
.I2(CLBLM_R_X7Y152_SLICE_X8Y152_BQ),
.I3(CLBLM_R_X3Y152_SLICE_X3Y152_AQ),
.I4(CLBLL_L_X2Y148_SLICE_X0Y148_B5Q),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X3Y152_SLICE_X3Y152_CO5),
.O6(CLBLM_R_X3Y152_SLICE_X3Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha082a0a0a0a0a0a0)
  ) CLBLM_R_X3Y152_SLICE_X3Y152_BLUT (
.I0(CLBLM_R_X5Y153_SLICE_X7Y153_BO6),
.I1(CLBLM_R_X3Y148_SLICE_X3Y148_BO5),
.I2(CLBLL_L_X4Y150_SLICE_X5Y150_D5Q),
.I3(CLBLM_R_X3Y150_SLICE_X3Y150_BQ),
.I4(CLBLM_R_X3Y153_SLICE_X3Y153_AQ),
.I5(CLBLM_R_X3Y153_SLICE_X3Y153_BQ),
.O5(CLBLM_R_X3Y152_SLICE_X3Y152_BO5),
.O6(CLBLM_R_X3Y152_SLICE_X3Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffff000afa3afa3)
  ) CLBLM_R_X3Y152_SLICE_X3Y152_ALUT (
.I0(CLBLL_L_X4Y149_SLICE_X4Y149_B5Q),
.I1(CLBLL_L_X2Y150_SLICE_X1Y150_A5Q),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLL_L_X4Y145_SLICE_X5Y145_BQ),
.I4(CLBLM_R_X3Y152_SLICE_X3Y152_CO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y152_SLICE_X3Y152_AO5),
.O6(CLBLM_R_X3Y152_SLICE_X3Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y153_SLICE_X2Y153_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_R_X3Y152_SLICE_X2Y152_CQ),
.Q(CLBLM_R_X3Y153_SLICE_X2Y153_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y153_SLICE_X2Y153_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y153_SLICE_X2Y153_DO5),
.O6(CLBLM_R_X3Y153_SLICE_X2Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y153_SLICE_X2Y153_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y153_SLICE_X2Y153_CO5),
.O6(CLBLM_R_X3Y153_SLICE_X2Y153_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y153_SLICE_X2Y153_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y153_SLICE_X2Y153_BO5),
.O6(CLBLM_R_X3Y153_SLICE_X2Y153_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5a0a0cccfcccf)
  ) CLBLM_R_X3Y153_SLICE_X2Y153_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(RIOB33_X105Y133_IOB_X1Y133_I),
.I2(CLBLM_R_X3Y153_SLICE_X2Y153_AQ),
.I3(CLBLM_R_X3Y151_SLICE_X3Y151_D5Q),
.I4(CLBLM_R_X5Y143_SLICE_X6Y143_DQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y153_SLICE_X2Y153_AO5),
.O6(CLBLM_R_X3Y153_SLICE_X2Y153_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y153_SLICE_X3Y153_A5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X3Y153_SLICE_X3Y153_BO6),
.Q(CLBLM_R_X3Y153_SLICE_X3Y153_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y153_SLICE_X3Y153_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X3Y153_SLICE_X3Y153_AO6),
.Q(CLBLM_R_X3Y153_SLICE_X3Y153_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y153_SLICE_X3Y153_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X3Y153_SLICE_X3Y153_CO5),
.Q(CLBLM_R_X3Y153_SLICE_X3Y153_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y153_SLICE_X3Y153_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y153_SLICE_X8Y153_BO5),
.Q(CLBLM_R_X3Y153_SLICE_X3Y153_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0200000000000000)
  ) CLBLM_R_X3Y153_SLICE_X3Y153_DLUT (
.I0(CLBLM_R_X3Y153_SLICE_X3Y153_BQ),
.I1(CLBLM_R_X3Y148_SLICE_X3Y148_BO5),
.I2(CLBLM_R_X3Y150_SLICE_X3Y150_BQ),
.I3(CLBLM_R_X3Y149_SLICE_X3Y149_AQ),
.I4(CLBLM_R_X3Y153_SLICE_X3Y153_AQ),
.I5(CLBLL_L_X4Y150_SLICE_X5Y150_D5Q),
.O5(CLBLM_R_X3Y153_SLICE_X3Y153_DO5),
.O6(CLBLM_R_X3Y153_SLICE_X3Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ffffff909090)
  ) CLBLM_R_X3Y153_SLICE_X3Y153_CLUT (
.I0(CLBLM_R_X3Y153_SLICE_X3Y153_BQ),
.I1(CLBLM_R_X3Y148_SLICE_X3Y148_BO6),
.I2(CLBLM_R_X5Y153_SLICE_X7Y153_BO6),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLL_L_X4Y153_SLICE_X5Y153_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y153_SLICE_X3Y153_CO5),
.O6(CLBLM_R_X3Y153_SLICE_X3Y153_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haca0a0a000ff0000)
  ) CLBLM_R_X3Y153_SLICE_X3Y153_BLUT (
.I0(CLBLM_R_X3Y143_SLICE_X2Y143_AQ),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I4(CLBLM_R_X3Y150_SLICE_X2Y150_CO5),
.I5(1'b1),
.O5(CLBLM_R_X3Y153_SLICE_X3Y153_BO5),
.O6(CLBLM_R_X3Y153_SLICE_X3Y153_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hebaafaaac300f000)
  ) CLBLM_R_X3Y153_SLICE_X3Y153_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X3Y148_SLICE_X3Y148_BO6),
.I2(CLBLM_R_X3Y153_SLICE_X3Y153_AQ),
.I3(CLBLM_R_X5Y153_SLICE_X7Y153_BO6),
.I4(CLBLM_R_X3Y153_SLICE_X3Y153_BQ),
.I5(CLBLM_L_X8Y151_SLICE_X10Y151_BQ),
.O5(CLBLM_R_X3Y153_SLICE_X3Y153_AO5),
.O6(CLBLM_R_X3Y153_SLICE_X3Y153_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y154_SLICE_X2Y154_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y154_SLICE_X2Y154_DO5),
.O6(CLBLM_R_X3Y154_SLICE_X2Y154_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y154_SLICE_X2Y154_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y154_SLICE_X2Y154_CO5),
.O6(CLBLM_R_X3Y154_SLICE_X2Y154_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y154_SLICE_X2Y154_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y154_SLICE_X2Y154_BO5),
.O6(CLBLM_R_X3Y154_SLICE_X2Y154_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y154_SLICE_X2Y154_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y154_SLICE_X2Y154_AO5),
.O6(CLBLM_R_X3Y154_SLICE_X2Y154_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y154_SLICE_X3Y154_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X3Y154_SLICE_X3Y154_AO6),
.Q(CLBLM_R_X3Y154_SLICE_X3Y154_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y154_SLICE_X3Y154_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y154_SLICE_X3Y154_DO5),
.O6(CLBLM_R_X3Y154_SLICE_X3Y154_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y154_SLICE_X3Y154_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y154_SLICE_X3Y154_CO5),
.O6(CLBLM_R_X3Y154_SLICE_X3Y154_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y154_SLICE_X3Y154_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y154_SLICE_X3Y154_BO5),
.O6(CLBLM_R_X3Y154_SLICE_X3Y154_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff00003c003c00)
  ) CLBLM_R_X3Y154_SLICE_X3Y154_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y153_SLICE_X11Y153_BQ),
.I2(CLBLM_R_X3Y154_SLICE_X3Y154_AQ),
.I3(CLBLM_R_X3Y152_SLICE_X2Y152_BQ),
.I4(CLBLL_L_X2Y151_SLICE_X1Y151_AQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X3Y154_SLICE_X3Y154_AO5),
.O6(CLBLM_R_X3Y154_SLICE_X3Y154_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y140_SLICE_X6Y140_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y140_SLICE_X6Y140_DO5),
.O6(CLBLM_R_X5Y140_SLICE_X6Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y140_SLICE_X6Y140_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y140_SLICE_X6Y140_CO5),
.O6(CLBLM_R_X5Y140_SLICE_X6Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y140_SLICE_X6Y140_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y140_SLICE_X6Y140_BO5),
.O6(CLBLM_R_X5Y140_SLICE_X6Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y140_SLICE_X6Y140_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y140_SLICE_X6Y140_AO5),
.O6(CLBLM_R_X5Y140_SLICE_X6Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y140_SLICE_X7Y140_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y140_SLICE_X7Y140_BO5),
.Q(CLBLM_R_X5Y140_SLICE_X7Y140_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y140_SLICE_X7Y140_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y140_SLICE_X7Y140_AO6),
.Q(CLBLM_R_X5Y140_SLICE_X7Y140_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y140_SLICE_X7Y140_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y140_SLICE_X7Y140_BO6),
.Q(CLBLM_R_X5Y140_SLICE_X7Y140_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y140_SLICE_X7Y140_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y140_SLICE_X7Y140_DO5),
.O6(CLBLM_R_X5Y140_SLICE_X7Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y140_SLICE_X7Y140_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y140_SLICE_X7Y140_CO5),
.O6(CLBLM_R_X5Y140_SLICE_X7Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbbb8888f3c0f3c0)
  ) CLBLM_R_X5Y140_SLICE_X7Y140_BLUT (
.I0(CLBLM_R_X7Y143_SLICE_X9Y143_DQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X5Y140_SLICE_X7Y140_AQ),
.I3(RIOB33_X105Y123_IOB_X1Y123_I),
.I4(RIOB33_X105Y107_IOB_X1Y108_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y140_SLICE_X7Y140_BO5),
.O6(CLBLM_R_X5Y140_SLICE_X7Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccaaf0ccccaaf0)
  ) CLBLM_R_X5Y140_SLICE_X7Y140_ALUT (
.I0(CLBLM_R_X5Y143_SLICE_X7Y143_DQ),
.I1(CLBLM_R_X5Y140_SLICE_X7Y140_BQ),
.I2(CLBLM_R_X5Y140_SLICE_X7Y140_AQ),
.I3(CLBLM_R_X11Y145_SLICE_X15Y145_BO5),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y140_SLICE_X7Y140_AO5),
.O6(CLBLM_R_X5Y140_SLICE_X7Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y141_SLICE_X6Y141_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y141_SLICE_X6Y141_AO6),
.Q(CLBLM_R_X5Y141_SLICE_X6Y141_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y141_SLICE_X6Y141_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y141_SLICE_X6Y141_DO5),
.O6(CLBLM_R_X5Y141_SLICE_X6Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y141_SLICE_X6Y141_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y141_SLICE_X6Y141_CO5),
.O6(CLBLM_R_X5Y141_SLICE_X6Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000080000000000)
  ) CLBLM_R_X5Y141_SLICE_X6Y141_BLUT (
.I0(CLBLL_L_X4Y147_SLICE_X4Y147_D5Q),
.I1(RIOB33_X105Y101_IOB_X1Y101_I),
.I2(CLBLL_L_X4Y150_SLICE_X4Y150_AQ),
.I3(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(RIOB33_X105Y131_IOB_X1Y131_I),
.O5(CLBLM_R_X5Y141_SLICE_X6Y141_BO5),
.O6(CLBLM_R_X5Y141_SLICE_X6Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0ffa0ffa0)
  ) CLBLM_R_X5Y141_SLICE_X6Y141_ALUT (
.I0(CLBLM_R_X5Y143_SLICE_X7Y143_CQ),
.I1(1'b1),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X5Y141_SLICE_X6Y141_BO6),
.I4(1'b1),
.I5(CLBLM_R_X5Y153_SLICE_X7Y153_CO6),
.O5(CLBLM_R_X5Y141_SLICE_X6Y141_AO5),
.O6(CLBLM_R_X5Y141_SLICE_X6Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y141_SLICE_X7Y141_A5_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y141_SLICE_X7Y141_AO5),
.Q(CLBLM_R_X5Y141_SLICE_X7Y141_A5Q),
.S(CLBLL_L_X4Y141_SLICE_X5Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y141_SLICE_X7Y141_A_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y141_SLICE_X7Y141_AO6),
.Q(CLBLM_R_X5Y141_SLICE_X7Y141_AQ),
.S(CLBLL_L_X4Y141_SLICE_X5Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y141_SLICE_X7Y141_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y141_SLICE_X7Y141_DO5),
.O6(CLBLM_R_X5Y141_SLICE_X7Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y141_SLICE_X7Y141_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y141_SLICE_X7Y141_CO5),
.O6(CLBLM_R_X5Y141_SLICE_X7Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y141_SLICE_X7Y141_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y141_SLICE_X7Y141_BO5),
.O6(CLBLM_R_X5Y141_SLICE_X7Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000cccc0000)
  ) CLBLM_R_X5Y141_SLICE_X7Y141_ALUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y153_SLICE_X4Y153_AQ),
.I2(1'b1),
.I3(CLBLM_R_X7Y141_SLICE_X9Y141_AQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y141_SLICE_X7Y141_AO5),
.O6(CLBLM_R_X5Y141_SLICE_X7Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y142_SLICE_X6Y142_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y142_SLICE_X6Y142_CO5),
.Q(CLBLM_R_X5Y142_SLICE_X6Y142_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y142_SLICE_X6Y142_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y142_SLICE_X6Y142_AO6),
.Q(CLBLM_R_X5Y142_SLICE_X6Y142_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y142_SLICE_X6Y142_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y142_SLICE_X6Y142_BO6),
.Q(CLBLM_R_X5Y142_SLICE_X6Y142_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y142_SLICE_X6Y142_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y142_SLICE_X6Y142_CO6),
.Q(CLBLM_R_X5Y142_SLICE_X6Y142_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y142_SLICE_X6Y142_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y142_SLICE_X6Y142_DO6),
.Q(CLBLM_R_X5Y142_SLICE_X6Y142_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0bbbbbb00)
  ) CLBLM_R_X5Y142_SLICE_X6Y142_DLUT (
.I0(CLBLM_L_X8Y142_SLICE_X11Y142_CQ),
.I1(CLBLM_R_X5Y149_SLICE_X7Y149_DQ),
.I2(CLBLM_R_X7Y144_SLICE_X9Y144_C5Q),
.I3(CLBLM_R_X5Y142_SLICE_X6Y142_DQ),
.I4(CLBLL_L_X4Y145_SLICE_X4Y145_A5Q),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X5Y142_SLICE_X6Y142_DO5),
.O6(CLBLM_R_X5Y142_SLICE_X6Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5a0f5a0baba1010)
  ) CLBLM_R_X5Y142_SLICE_X6Y142_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X7Y150_SLICE_X9Y150_B5Q),
.I2(CLBLL_L_X4Y142_SLICE_X5Y142_BQ),
.I3(CLBLL_L_X4Y141_SLICE_X5Y141_A5Q),
.I4(CLBLL_L_X4Y143_SLICE_X4Y143_BQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y142_SLICE_X6Y142_CO5),
.O6(CLBLM_R_X5Y142_SLICE_X6Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaafc0cfc0c)
  ) CLBLM_R_X5Y142_SLICE_X6Y142_BLUT (
.I0(CLBLM_R_X5Y144_SLICE_X6Y144_B5Q),
.I1(CLBLM_R_X5Y142_SLICE_X6Y142_BQ),
.I2(CLBLM_R_X11Y145_SLICE_X15Y145_BO5),
.I3(CLBLM_R_X5Y143_SLICE_X6Y143_AQ),
.I4(1'b1),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X5Y142_SLICE_X6Y142_BO5),
.O6(CLBLM_R_X5Y142_SLICE_X6Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccff5acccc005a)
  ) CLBLM_R_X5Y142_SLICE_X6Y142_ALUT (
.I0(CLBLM_L_X8Y142_SLICE_X10Y142_DO6),
.I1(CLBLM_R_X7Y143_SLICE_X9Y143_BQ),
.I2(CLBLM_R_X5Y142_SLICE_X6Y142_AQ),
.I3(CLBLM_L_X8Y149_SLICE_X11Y149_BQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLL_L_X4Y144_SLICE_X5Y144_CQ),
.O5(CLBLM_R_X5Y142_SLICE_X6Y142_AO5),
.O6(CLBLM_R_X5Y142_SLICE_X6Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y142_SLICE_X7Y142_B5_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y142_SLICE_X7Y142_BO5),
.Q(CLBLM_R_X5Y142_SLICE_X7Y142_B5Q),
.S(CLBLL_L_X4Y151_SLICE_X4Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y142_SLICE_X7Y142_C5_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y142_SLICE_X7Y142_CO5),
.Q(CLBLM_R_X5Y142_SLICE_X7Y142_C5Q),
.S(CLBLL_L_X4Y151_SLICE_X4Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y142_SLICE_X7Y142_B_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y142_SLICE_X7Y142_BO6),
.Q(CLBLM_R_X5Y142_SLICE_X7Y142_BQ),
.S(CLBLL_L_X4Y151_SLICE_X4Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y142_SLICE_X7Y142_C_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y142_SLICE_X7Y142_CO6),
.Q(CLBLM_R_X5Y142_SLICE_X7Y142_CQ),
.S(CLBLL_L_X4Y151_SLICE_X4Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y142_SLICE_X7Y142_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y142_SLICE_X7Y142_DO5),
.O6(CLBLM_R_X5Y142_SLICE_X7Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888c0c0c0c0)
  ) CLBLM_R_X5Y142_SLICE_X7Y142_CLUT (
.I0(CLBLM_R_X5Y141_SLICE_X7Y141_AQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X3Y144_SLICE_X3Y144_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y142_SLICE_X7Y142_CO5),
.O6(CLBLM_R_X5Y142_SLICE_X7Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888cccc0000)
  ) CLBLM_R_X5Y142_SLICE_X7Y142_BLUT (
.I0(CLBLM_R_X5Y142_SLICE_X7Y142_CQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X5Y142_SLICE_X6Y142_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y142_SLICE_X7Y142_BO5),
.O6(CLBLM_R_X5Y142_SLICE_X7Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa000000010001)
  ) CLBLM_R_X5Y142_SLICE_X7Y142_ALUT (
.I0(CLBLM_R_X5Y143_SLICE_X7Y143_BQ),
.I1(CLBLM_R_X5Y149_SLICE_X7Y149_CQ),
.I2(CLBLM_R_X5Y143_SLICE_X7Y143_CQ),
.I3(CLBLM_R_X7Y147_SLICE_X8Y147_DQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y142_SLICE_X7Y142_AO5),
.O6(CLBLM_R_X5Y142_SLICE_X7Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y143_SLICE_X6Y143_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y143_SLICE_X6Y143_DO5),
.Q(CLBLM_R_X5Y143_SLICE_X6Y143_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y143_SLICE_X6Y143_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y143_SLICE_X6Y143_AO6),
.Q(CLBLM_R_X5Y143_SLICE_X6Y143_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y143_SLICE_X6Y143_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y143_SLICE_X6Y143_BO6),
.Q(CLBLM_R_X5Y143_SLICE_X6Y143_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y143_SLICE_X6Y143_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y143_SLICE_X6Y143_CO6),
.Q(CLBLM_R_X5Y143_SLICE_X6Y143_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y143_SLICE_X6Y143_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y143_SLICE_X6Y143_DO6),
.Q(CLBLM_R_X5Y143_SLICE_X6Y143_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hd8d8d8d8ffaa5500)
  ) CLBLM_R_X5Y143_SLICE_X6Y143_DLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLL_L_X4Y144_SLICE_X4Y144_AQ),
.I2(CLBLM_R_X3Y145_SLICE_X2Y145_CQ),
.I3(RIOB33_X105Y109_IOB_X1Y109_I),
.I4(CLBLM_R_X7Y147_SLICE_X8Y147_DQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y143_SLICE_X6Y143_DO5),
.O6(CLBLM_R_X5Y143_SLICE_X6Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfeaa5400fefe5454)
  ) CLBLM_R_X5Y143_SLICE_X6Y143_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X5Y143_SLICE_X6Y143_CQ),
.I2(CLBLL_L_X4Y144_SLICE_X4Y144_AQ),
.I3(CLBLM_R_X5Y144_SLICE_X6Y144_CQ),
.I4(CLBLL_L_X4Y143_SLICE_X5Y143_CQ),
.I5(CLBLM_R_X3Y147_SLICE_X3Y147_BQ),
.O5(CLBLM_R_X5Y143_SLICE_X6Y143_CO5),
.O6(CLBLM_R_X5Y143_SLICE_X6Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haafcaa00aafcaafc)
  ) CLBLM_R_X5Y143_SLICE_X6Y143_BLUT (
.I0(CLBLL_L_X4Y148_SLICE_X5Y148_B5Q),
.I1(CLBLM_R_X5Y143_SLICE_X6Y143_BQ),
.I2(CLBLL_L_X4Y142_SLICE_X4Y142_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X8Y150_SLICE_X11Y150_B5Q),
.I5(CLBLM_R_X5Y149_SLICE_X6Y149_D5Q),
.O5(CLBLM_R_X5Y143_SLICE_X6Y143_BO5),
.O6(CLBLM_R_X5Y143_SLICE_X6Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00c8c8ff00fafa)
  ) CLBLM_R_X5Y143_SLICE_X6Y143_ALUT (
.I0(CLBLM_R_X5Y153_SLICE_X7Y153_A5Q),
.I1(CLBLM_L_X8Y142_SLICE_X11Y142_CQ),
.I2(CLBLM_R_X5Y143_SLICE_X6Y143_AQ),
.I3(CLBLM_R_X5Y151_SLICE_X6Y151_DQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X5Y149_SLICE_X7Y149_DQ),
.O5(CLBLM_R_X5Y143_SLICE_X6Y143_AO5),
.O6(CLBLM_R_X5Y143_SLICE_X6Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y143_SLICE_X7Y143_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y143_SLICE_X7Y143_AO6),
.Q(CLBLM_R_X5Y143_SLICE_X7Y143_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y143_SLICE_X7Y143_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y143_SLICE_X7Y143_BO6),
.Q(CLBLM_R_X5Y143_SLICE_X7Y143_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y143_SLICE_X7Y143_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y143_SLICE_X7Y143_CO6),
.Q(CLBLM_R_X5Y143_SLICE_X7Y143_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y143_SLICE_X7Y143_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y143_SLICE_X7Y143_DO6),
.Q(CLBLM_R_X5Y143_SLICE_X7Y143_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffabbba55501110)
  ) CLBLM_R_X5Y143_SLICE_X7Y143_DLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X5Y149_SLICE_X7Y149_DQ),
.I2(CLBLM_R_X5Y143_SLICE_X7Y143_DQ),
.I3(CLBLM_R_X5Y141_SLICE_X7Y141_AQ),
.I4(CLBLM_L_X8Y142_SLICE_X11Y142_CQ),
.I5(CLBLL_L_X4Y153_SLICE_X5Y153_BQ),
.O5(CLBLM_R_X5Y143_SLICE_X7Y143_DO5),
.O6(CLBLM_R_X5Y143_SLICE_X7Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hb1b1e4e4b1b1e4e4)
  ) CLBLM_R_X5Y143_SLICE_X7Y143_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X8Y144_SLICE_X10Y144_AQ),
.I2(CLBLM_R_X3Y143_SLICE_X2Y143_DQ),
.I3(1'b1),
.I4(CLBLM_R_X7Y143_SLICE_X9Y143_CQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y143_SLICE_X7Y143_CO5),
.O6(CLBLM_R_X5Y143_SLICE_X7Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff33cc000033cc)
  ) CLBLM_R_X5Y143_SLICE_X7Y143_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y143_SLICE_X9Y143_BQ),
.I2(1'b1),
.I3(CLBLM_L_X8Y144_SLICE_X11Y144_AQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLL_L_X2Y145_SLICE_X1Y145_AQ),
.O5(CLBLM_R_X5Y143_SLICE_X7Y143_BO5),
.O6(CLBLM_R_X5Y143_SLICE_X7Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff003333ff00cccc)
  ) CLBLM_R_X5Y143_SLICE_X7Y143_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y144_SLICE_X3Y144_CQ),
.I2(1'b1),
.I3(CLBLM_R_X5Y143_SLICE_X6Y143_BQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X5Y145_SLICE_X7Y145_A5Q),
.O5(CLBLM_R_X5Y143_SLICE_X7Y143_AO5),
.O6(CLBLM_R_X5Y143_SLICE_X7Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y144_SLICE_X6Y144_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y144_SLICE_X6Y144_BO5),
.Q(CLBLM_R_X5Y144_SLICE_X6Y144_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y144_SLICE_X6Y144_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y144_SLICE_X6Y144_CO5),
.Q(CLBLM_R_X5Y144_SLICE_X6Y144_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y144_SLICE_X6Y144_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y144_SLICE_X6Y144_DO5),
.Q(CLBLM_R_X5Y144_SLICE_X6Y144_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y144_SLICE_X6Y144_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y144_SLICE_X6Y144_AO6),
.Q(CLBLM_R_X5Y144_SLICE_X6Y144_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y144_SLICE_X6Y144_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y144_SLICE_X6Y144_BO6),
.Q(CLBLM_R_X5Y144_SLICE_X6Y144_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y144_SLICE_X6Y144_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y144_SLICE_X6Y144_CO6),
.Q(CLBLM_R_X5Y144_SLICE_X6Y144_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y144_SLICE_X6Y144_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y144_SLICE_X6Y144_DO6),
.Q(CLBLM_R_X5Y144_SLICE_X6Y144_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0aaf0aaffcc00cc)
  ) CLBLM_R_X5Y144_SLICE_X6Y144_DLUT (
.I0(RIOB33_X105Y107_IOB_X1Y107_I),
.I1(CLBLM_R_X7Y150_SLICE_X9Y150_B5Q),
.I2(CLBLM_L_X10Y150_SLICE_X13Y150_A5Q),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X5Y153_SLICE_X7Y153_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X5Y144_SLICE_X6Y144_DO5),
.O6(CLBLM_R_X5Y144_SLICE_X6Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccf0f0aaaaff00)
  ) CLBLM_R_X5Y144_SLICE_X6Y144_CLUT (
.I0(CLBLM_R_X7Y152_SLICE_X9Y152_AQ),
.I1(CLBLM_R_X5Y144_SLICE_X6Y144_D5Q),
.I2(RIOB33_X105Y109_IOB_X1Y109_I),
.I3(CLBLM_L_X8Y148_SLICE_X11Y148_CQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y144_SLICE_X6Y144_CO5),
.O6(CLBLM_R_X5Y144_SLICE_X6Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcfc0c0fa0afa0a)
  ) CLBLM_R_X5Y144_SLICE_X6Y144_BLUT (
.I0(CLBLL_L_X4Y150_SLICE_X5Y150_C5Q),
.I1(CLBLM_L_X8Y147_SLICE_X10Y147_B5Q),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_L_X8Y143_SLICE_X11Y143_BQ),
.I4(RIOB33_X105Y119_IOB_X1Y119_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y144_SLICE_X6Y144_BO5),
.O6(CLBLM_R_X5Y144_SLICE_X6Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffddd00000ddd0)
  ) CLBLM_R_X5Y144_SLICE_X6Y144_ALUT (
.I0(CLBLM_R_X3Y148_SLICE_X2Y148_D5Q),
.I1(CLBLM_R_X5Y144_SLICE_X6Y144_DQ),
.I2(CLBLM_R_X5Y144_SLICE_X6Y144_AQ),
.I3(CLBLM_L_X8Y147_SLICE_X10Y147_B5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X3Y146_SLICE_X3Y146_CQ),
.O5(CLBLM_R_X5Y144_SLICE_X6Y144_AO5),
.O6(CLBLM_R_X5Y144_SLICE_X6Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y144_SLICE_X7Y144_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y144_SLICE_X7Y144_AO6),
.Q(CLBLM_R_X5Y144_SLICE_X7Y144_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y144_SLICE_X7Y144_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y144_SLICE_X7Y144_BO6),
.Q(CLBLM_R_X5Y144_SLICE_X7Y144_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y144_SLICE_X7Y144_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y144_SLICE_X7Y144_CO6),
.Q(CLBLM_R_X5Y144_SLICE_X7Y144_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y144_SLICE_X7Y144_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y144_SLICE_X7Y144_DO6),
.Q(CLBLM_R_X5Y144_SLICE_X7Y144_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hddddd8d88888d8d8)
  ) CLBLM_R_X5Y144_SLICE_X7Y144_DLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X5Y144_SLICE_X7Y144_AQ),
.I2(CLBLM_R_X5Y144_SLICE_X7Y144_DQ),
.I3(1'b1),
.I4(CLBLM_L_X10Y143_SLICE_X12Y143_BO5),
.I5(CLBLM_R_X7Y143_SLICE_X9Y143_AQ),
.O5(CLBLM_R_X5Y144_SLICE_X7Y144_DO5),
.O6(CLBLM_R_X5Y144_SLICE_X7Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefb5451fefb5451)
  ) CLBLM_R_X5Y144_SLICE_X7Y144_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X5Y144_SLICE_X7Y144_CQ),
.I2(CLBLL_L_X2Y148_SLICE_X0Y148_B5Q),
.I3(CLBLL_L_X4Y144_SLICE_X4Y144_DO6),
.I4(CLBLM_L_X8Y149_SLICE_X10Y149_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X5Y144_SLICE_X7Y144_CO5),
.O6(CLBLM_R_X5Y144_SLICE_X7Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ececff002020)
  ) CLBLM_R_X5Y144_SLICE_X7Y144_BLUT (
.I0(CLBLM_R_X7Y142_SLICE_X8Y142_CO6),
.I1(CLBLM_L_X8Y149_SLICE_X11Y149_BQ),
.I2(CLBLM_R_X7Y142_SLICE_X8Y142_DO6),
.I3(CLBLM_R_X3Y149_SLICE_X2Y149_A5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_L_X8Y148_SLICE_X11Y148_B5Q),
.O5(CLBLM_R_X5Y144_SLICE_X7Y144_BO5),
.O6(CLBLM_R_X5Y144_SLICE_X7Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ddddf0f0dd00)
  ) CLBLM_R_X5Y144_SLICE_X7Y144_ALUT (
.I0(CLBLM_R_X5Y149_SLICE_X6Y149_D5Q),
.I1(CLBLM_L_X8Y150_SLICE_X11Y150_B5Q),
.I2(CLBLM_L_X10Y143_SLICE_X12Y143_AQ),
.I3(CLBLM_R_X5Y144_SLICE_X7Y144_AQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLL_L_X4Y146_SLICE_X5Y146_A5Q),
.O5(CLBLM_R_X5Y144_SLICE_X7Y144_AO5),
.O6(CLBLM_R_X5Y144_SLICE_X7Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y145_SLICE_X6Y145_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y145_SLICE_X6Y145_BO5),
.Q(CLBLM_R_X5Y145_SLICE_X6Y145_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y145_SLICE_X6Y145_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y145_SLICE_X6Y145_AO6),
.Q(CLBLM_R_X5Y145_SLICE_X6Y145_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y145_SLICE_X6Y145_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y145_SLICE_X6Y145_BO6),
.Q(CLBLM_R_X5Y145_SLICE_X6Y145_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y145_SLICE_X6Y145_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y145_SLICE_X6Y145_CO6),
.Q(CLBLM_R_X5Y145_SLICE_X6Y145_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y145_SLICE_X6Y145_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y145_SLICE_X6Y145_DO6),
.Q(CLBLM_R_X5Y145_SLICE_X6Y145_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffa5550aafa0050)
  ) CLBLM_R_X5Y145_SLICE_X6Y145_DLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(1'b1),
.I2(CLBLM_R_X5Y145_SLICE_X6Y145_DQ),
.I3(CLBLM_L_X10Y143_SLICE_X12Y143_BO5),
.I4(CLBLL_L_X4Y145_SLICE_X4Y145_A5Q),
.I5(CLBLM_R_X5Y145_SLICE_X6Y145_AQ),
.O5(CLBLM_R_X5Y145_SLICE_X6Y145_DO5),
.O6(CLBLM_R_X5Y145_SLICE_X6Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfe54fe54aa00aa00)
  ) CLBLM_R_X5Y145_SLICE_X6Y145_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X5Y145_SLICE_X6Y145_CQ),
.I2(CLBLM_R_X3Y149_SLICE_X3Y149_CQ),
.I3(CLBLM_R_X5Y142_SLICE_X6Y142_CQ),
.I4(1'b1),
.I5(CLBLM_L_X10Y143_SLICE_X12Y143_AO6),
.O5(CLBLM_R_X5Y145_SLICE_X6Y145_CO5),
.O6(CLBLM_R_X5Y145_SLICE_X6Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff00f00fa0afa0a)
  ) CLBLM_R_X5Y145_SLICE_X6Y145_BLUT (
.I0(CLBLM_R_X5Y146_SLICE_X7Y146_B5Q),
.I1(1'b1),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X3Y145_SLICE_X2Y145_C5Q),
.I4(CLBLM_R_X11Y146_SLICE_X14Y146_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y145_SLICE_X6Y145_BO5),
.O6(CLBLM_R_X5Y145_SLICE_X6Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00fcfcff005454)
  ) CLBLM_R_X5Y145_SLICE_X6Y145_ALUT (
.I0(CLBLM_R_X3Y147_SLICE_X3Y147_BQ),
.I1(CLBLL_L_X2Y147_SLICE_X1Y147_A5Q),
.I2(CLBLM_R_X5Y145_SLICE_X6Y145_AQ),
.I3(CLBLM_R_X5Y153_SLICE_X6Y153_BQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X5Y144_SLICE_X6Y144_CQ),
.O5(CLBLM_R_X5Y145_SLICE_X6Y145_AO5),
.O6(CLBLM_R_X5Y145_SLICE_X6Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y145_SLICE_X7Y145_A5_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y145_SLICE_X7Y145_AO5),
.Q(CLBLM_R_X5Y145_SLICE_X7Y145_A5Q),
.S(CLBLL_L_X4Y151_SLICE_X4Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y145_SLICE_X7Y145_A_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y145_SLICE_X7Y145_AO6),
.Q(CLBLM_R_X5Y145_SLICE_X7Y145_AQ),
.S(CLBLL_L_X4Y151_SLICE_X4Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff2f22ffff2f22)
  ) CLBLM_R_X5Y145_SLICE_X7Y145_DLUT (
.I0(CLBLM_R_X5Y145_SLICE_X6Y145_DQ),
.I1(CLBLM_L_X8Y142_SLICE_X10Y142_BO5),
.I2(CLBLM_L_X8Y145_SLICE_X10Y145_CO5),
.I3(CLBLM_R_X5Y145_SLICE_X7Y145_A5Q),
.I4(CLBLM_R_X5Y145_SLICE_X7Y145_BO5),
.I5(1'b1),
.O5(CLBLM_R_X5Y145_SLICE_X7Y145_DO5),
.O6(CLBLM_R_X5Y145_SLICE_X7Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffffae)
  ) CLBLM_R_X5Y145_SLICE_X7Y145_CLUT (
.I0(CLBLM_L_X8Y148_SLICE_X10Y148_CO5),
.I1(CLBLM_R_X5Y142_SLICE_X7Y142_B5Q),
.I2(CLBLM_R_X5Y145_SLICE_X7Y145_BO6),
.I3(CLBLL_L_X4Y142_SLICE_X4Y142_CO5),
.I4(CLBLM_R_X5Y145_SLICE_X7Y145_DO6),
.I5(CLBLM_R_X5Y151_SLICE_X7Y151_DO6),
.O5(CLBLM_R_X5Y145_SLICE_X7Y145_CO5),
.O6(CLBLM_R_X5Y145_SLICE_X7Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h55ffffff44500000)
  ) CLBLM_R_X5Y145_SLICE_X7Y145_BLUT (
.I0(CLBLM_L_X8Y150_SLICE_X10Y150_A5Q),
.I1(CLBLL_L_X4Y151_SLICE_X4Y151_AQ),
.I2(CLBLM_R_X5Y142_SLICE_X7Y142_BQ),
.I3(CLBLM_R_X11Y149_SLICE_X14Y149_AQ),
.I4(CLBLM_L_X10Y143_SLICE_X13Y143_AO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y145_SLICE_X7Y145_BO5),
.O6(CLBLM_R_X5Y145_SLICE_X7Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0f000f000)
  ) CLBLM_R_X5Y145_SLICE_X7Y145_ALUT (
.I0(CLBLM_R_X5Y145_SLICE_X6Y145_DQ),
.I1(1'b1),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLL_L_X2Y144_SLICE_X1Y144_A5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y145_SLICE_X7Y145_AO5),
.O6(CLBLM_R_X5Y145_SLICE_X7Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y146_SLICE_X6Y146_B5_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y146_SLICE_X6Y146_BO5),
.Q(CLBLM_R_X5Y146_SLICE_X6Y146_B5Q),
.S(CLBLM_R_X11Y148_SLICE_X14Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y146_SLICE_X6Y146_A_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y146_SLICE_X6Y146_AO6),
.Q(CLBLM_R_X5Y146_SLICE_X6Y146_AQ),
.S(CLBLM_R_X11Y148_SLICE_X14Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y146_SLICE_X6Y146_B_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y146_SLICE_X6Y146_BO6),
.Q(CLBLM_R_X5Y146_SLICE_X6Y146_BQ),
.S(CLBLM_R_X11Y148_SLICE_X14Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y146_SLICE_X6Y146_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y146_SLICE_X6Y146_DO5),
.O6(CLBLM_R_X5Y146_SLICE_X6Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h50ff505050ff5050)
  ) CLBLM_R_X5Y146_SLICE_X6Y146_CLUT (
.I0(CLBLM_R_X5Y145_SLICE_X7Y145_BO6),
.I1(1'b1),
.I2(CLBLM_R_X5Y146_SLICE_X6Y146_BQ),
.I3(CLBLM_L_X10Y143_SLICE_X12Y143_DO5),
.I4(CLBLM_R_X5Y147_SLICE_X6Y147_CQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y146_SLICE_X6Y146_CO5),
.O6(CLBLM_R_X5Y146_SLICE_X6Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00000aaaa0000)
  ) CLBLM_R_X5Y146_SLICE_X6Y146_BLUT (
.I0(CLBLM_L_X10Y153_SLICE_X13Y153_AQ),
.I1(1'b1),
.I2(CLBLL_L_X4Y146_SLICE_X5Y146_BQ),
.I3(1'b1),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y146_SLICE_X6Y146_BO5),
.O6(CLBLM_R_X5Y146_SLICE_X6Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0c0c0c0c0)
  ) CLBLM_R_X5Y146_SLICE_X6Y146_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y145_SLICE_X2Y145_CQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y146_SLICE_X6Y146_AO5),
.O6(CLBLM_R_X5Y146_SLICE_X6Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y146_SLICE_X7Y146_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y146_SLICE_X7Y146_BO5),
.Q(CLBLM_R_X5Y146_SLICE_X7Y146_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y146_SLICE_X7Y146_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y146_SLICE_X7Y146_AO6),
.Q(CLBLM_R_X5Y146_SLICE_X7Y146_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y146_SLICE_X7Y146_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y146_SLICE_X7Y146_BO6),
.Q(CLBLM_R_X5Y146_SLICE_X7Y146_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y146_SLICE_X7Y146_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y146_SLICE_X7Y146_CO6),
.Q(CLBLM_R_X5Y146_SLICE_X7Y146_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y146_SLICE_X7Y146_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y146_SLICE_X7Y146_DO6),
.Q(CLBLM_R_X5Y146_SLICE_X7Y146_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccfacc50ccfacc50)
  ) CLBLM_R_X5Y146_SLICE_X7Y146_DLUT (
.I0(CLBLM_R_X11Y145_SLICE_X15Y145_BO5),
.I1(CLBLL_L_X4Y146_SLICE_X4Y146_DQ),
.I2(CLBLM_R_X5Y146_SLICE_X7Y146_DQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X3Y146_SLICE_X3Y146_DQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y146_SLICE_X7Y146_DO5),
.O6(CLBLM_R_X5Y146_SLICE_X7Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfe54fe54aa00fe54)
  ) CLBLM_R_X5Y146_SLICE_X7Y146_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X5Y146_SLICE_X7Y146_CQ),
.I2(CLBLM_R_X3Y148_SLICE_X3Y148_A5Q),
.I3(CLBLM_R_X3Y142_SLICE_X3Y142_BQ),
.I4(CLBLM_R_X5Y149_SLICE_X6Y149_D5Q),
.I5(CLBLM_L_X8Y150_SLICE_X11Y150_B5Q),
.O5(CLBLM_R_X5Y146_SLICE_X7Y146_CO5),
.O6(CLBLM_R_X5Y146_SLICE_X7Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc5cac5caff0ff000)
  ) CLBLM_R_X5Y146_SLICE_X7Y146_BLUT (
.I0(CLBLM_R_X3Y152_SLICE_X3Y152_AQ),
.I1(CLBLM_R_X5Y147_SLICE_X7Y147_A5Q),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X5Y146_SLICE_X6Y146_B5Q),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y146_SLICE_X7Y146_BO5),
.O6(CLBLM_R_X5Y146_SLICE_X7Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccff00cccc0f0f)
  ) CLBLM_R_X5Y146_SLICE_X7Y146_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y143_SLICE_X11Y143_A5Q),
.I2(CLBLM_R_X5Y146_SLICE_X7Y146_AQ),
.I3(CLBLM_R_X5Y147_SLICE_X6Y147_BQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_L_X8Y149_SLICE_X11Y149_BQ),
.O5(CLBLM_R_X5Y146_SLICE_X7Y146_AO5),
.O6(CLBLM_R_X5Y146_SLICE_X7Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y147_SLICE_X6Y147_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y147_SLICE_X6Y147_BO5),
.Q(CLBLM_R_X5Y147_SLICE_X6Y147_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y147_SLICE_X6Y147_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y147_SLICE_X6Y147_AO6),
.Q(CLBLM_R_X5Y147_SLICE_X6Y147_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y147_SLICE_X6Y147_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y147_SLICE_X6Y147_BO6),
.Q(CLBLM_R_X5Y147_SLICE_X6Y147_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y147_SLICE_X6Y147_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y147_SLICE_X6Y147_CO6),
.Q(CLBLM_R_X5Y147_SLICE_X6Y147_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y147_SLICE_X6Y147_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y147_SLICE_X6Y147_DO6),
.Q(CLBLM_R_X5Y147_SLICE_X6Y147_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccaaccffcca0ccf0)
  ) CLBLM_R_X5Y147_SLICE_X6Y147_DLUT (
.I0(CLBLM_L_X8Y142_SLICE_X11Y142_CQ),
.I1(CLBLL_L_X4Y144_SLICE_X5Y144_DQ),
.I2(CLBLM_R_X5Y147_SLICE_X6Y147_DQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X5Y149_SLICE_X7Y149_DQ),
.I5(CLBLL_L_X2Y146_SLICE_X1Y146_A5Q),
.O5(CLBLM_R_X5Y147_SLICE_X6Y147_DO5),
.O6(CLBLM_R_X5Y147_SLICE_X6Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hafa0afa0aca0aca0)
  ) CLBLM_R_X5Y147_SLICE_X6Y147_CLUT (
.I0(CLBLM_R_X5Y142_SLICE_X6Y142_BQ),
.I1(CLBLM_R_X5Y147_SLICE_X6Y147_CQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_L_X10Y143_SLICE_X12Y143_AO6),
.I4(1'b1),
.I5(CLBLL_L_X4Y149_SLICE_X5Y149_AQ),
.O5(CLBLM_R_X5Y147_SLICE_X6Y147_CO5),
.O6(CLBLM_R_X5Y147_SLICE_X6Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hafa0afa0fafa0a0a)
  ) CLBLM_R_X5Y147_SLICE_X6Y147_BLUT (
.I0(CLBLM_R_X5Y149_SLICE_X7Y149_C5Q),
.I1(1'b1),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X5Y150_SLICE_X7Y150_A5Q),
.I4(CLBLM_R_X5Y147_SLICE_X6Y147_CQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y147_SLICE_X6Y147_BO5),
.O6(CLBLM_R_X5Y147_SLICE_X6Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00f0f0d8d8)
  ) CLBLM_R_X5Y147_SLICE_X6Y147_ALUT (
.I0(CLBLM_R_X7Y150_SLICE_X9Y150_CQ),
.I1(CLBLM_R_X5Y151_SLICE_X6Y151_AQ),
.I2(CLBLM_R_X5Y147_SLICE_X6Y147_AQ),
.I3(CLBLM_R_X11Y144_SLICE_X14Y144_AQ),
.I4(CLBLM_L_X8Y146_SLICE_X10Y146_AQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X5Y147_SLICE_X6Y147_AO5),
.O6(CLBLM_R_X5Y147_SLICE_X6Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y147_SLICE_X7Y147_A5_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y147_SLICE_X7Y147_AO5),
.Q(CLBLM_R_X5Y147_SLICE_X7Y147_A5Q),
.S(CLBLM_R_X11Y148_SLICE_X15Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y147_SLICE_X7Y147_B5_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y147_SLICE_X7Y147_BO5),
.Q(CLBLM_R_X5Y147_SLICE_X7Y147_B5Q),
.S(CLBLM_R_X11Y148_SLICE_X15Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y147_SLICE_X7Y147_C5_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y147_SLICE_X7Y147_CO5),
.Q(CLBLM_R_X5Y147_SLICE_X7Y147_C5Q),
.S(CLBLM_R_X11Y148_SLICE_X15Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y147_SLICE_X7Y147_A_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y147_SLICE_X7Y147_AO6),
.Q(CLBLM_R_X5Y147_SLICE_X7Y147_AQ),
.S(CLBLM_R_X11Y148_SLICE_X15Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y147_SLICE_X7Y147_B_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y147_SLICE_X7Y147_BO6),
.Q(CLBLM_R_X5Y147_SLICE_X7Y147_BQ),
.S(CLBLM_R_X11Y148_SLICE_X15Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y147_SLICE_X7Y147_C_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y147_SLICE_X7Y147_CO6),
.Q(CLBLM_R_X5Y147_SLICE_X7Y147_CQ),
.S(CLBLM_R_X11Y148_SLICE_X15Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3030303030303030)
  ) CLBLM_R_X5Y147_SLICE_X7Y147_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y151_SLICE_X10Y151_B5Q),
.I2(CLBLM_R_X5Y140_SLICE_X7Y140_B5Q),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y147_SLICE_X7Y147_DO5),
.O6(CLBLM_R_X5Y147_SLICE_X7Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a088888888)
  ) CLBLM_R_X5Y147_SLICE_X7Y147_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X3Y148_SLICE_X3Y148_A5Q),
.I2(CLBLM_R_X7Y148_SLICE_X9Y148_CQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y147_SLICE_X7Y147_CO5),
.O6(CLBLM_R_X5Y147_SLICE_X7Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0000f0f00000)
  ) CLBLM_R_X5Y147_SLICE_X7Y147_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y147_SLICE_X6Y147_B5Q),
.I2(CLBLM_R_X5Y149_SLICE_X6Y149_AQ),
.I3(1'b1),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y147_SLICE_X7Y147_BO5),
.O6(CLBLM_R_X5Y147_SLICE_X7Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00000cccc0000)
  ) CLBLM_R_X5Y147_SLICE_X7Y147_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y151_SLICE_X9Y151_DQ),
.I2(CLBLM_R_X5Y143_SLICE_X7Y143_AQ),
.I3(1'b1),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y147_SLICE_X7Y147_AO5),
.O6(CLBLM_R_X5Y147_SLICE_X7Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y148_SLICE_X6Y148_B5_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y148_SLICE_X6Y148_BO5),
.Q(CLBLM_R_X5Y148_SLICE_X6Y148_B5Q),
.S(CLBLL_L_X4Y145_SLICE_X5Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y148_SLICE_X6Y148_A_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y150_SLICE_X2Y150_CO6),
.Q(CLBLM_R_X5Y148_SLICE_X6Y148_AQ),
.S(CLBLL_L_X4Y145_SLICE_X5Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y148_SLICE_X6Y148_B_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y148_SLICE_X6Y148_BO6),
.Q(CLBLM_R_X5Y148_SLICE_X6Y148_BQ),
.S(CLBLL_L_X4Y145_SLICE_X5Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y148_SLICE_X6Y148_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y148_SLICE_X6Y148_DO5),
.O6(CLBLM_R_X5Y148_SLICE_X6Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff808080c0c0c0c0)
  ) CLBLM_R_X5Y148_SLICE_X6Y148_CLUT (
.I0(CLBLL_L_X4Y147_SLICE_X4Y147_C5Q),
.I1(CLBLM_R_X7Y145_SLICE_X8Y145_B5Q),
.I2(CLBLM_R_X5Y151_SLICE_X6Y151_BQ),
.I3(CLBLM_L_X10Y150_SLICE_X12Y150_AQ),
.I4(CLBLL_L_X4Y149_SLICE_X4Y149_D5Q),
.I5(1'b1),
.O5(CLBLM_R_X5Y148_SLICE_X6Y148_CO5),
.O6(CLBLM_R_X5Y148_SLICE_X6Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000f0f00000)
  ) CLBLM_R_X5Y148_SLICE_X6Y148_BLUT (
.I0(CLBLL_L_X2Y150_SLICE_X1Y150_AQ),
.I1(1'b1),
.I2(CLBLL_L_X4Y147_SLICE_X5Y147_DQ),
.I3(1'b1),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y148_SLICE_X6Y148_BO5),
.O6(CLBLM_R_X5Y148_SLICE_X6Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0afffffff)
  ) CLBLM_R_X5Y148_SLICE_X6Y148_ALUT (
.I0(CLBLL_L_X4Y148_SLICE_X4Y148_BO5),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLL_L_X4Y149_SLICE_X4Y149_AQ),
.I3(CLBLL_L_X4Y148_SLICE_X5Y148_AQ),
.I4(CLBLL_L_X4Y148_SLICE_X5Y148_BQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y148_SLICE_X6Y148_AO5),
.O6(CLBLM_R_X5Y148_SLICE_X6Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y148_SLICE_X7Y148_A_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y148_SLICE_X6Y148_AO6),
.Q(CLBLM_R_X5Y148_SLICE_X7Y148_AQ),
.S(CLBLL_L_X4Y151_SLICE_X4Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ff00f0f0fff0)
  ) CLBLM_R_X5Y148_SLICE_X7Y148_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X7Y149_SLICE_X8Y149_BQ),
.I3(CLBLM_R_X5Y149_SLICE_X6Y149_CQ),
.I4(CLBLM_L_X8Y142_SLICE_X10Y142_BO5),
.I5(CLBLM_L_X10Y143_SLICE_X12Y143_AO5),
.O5(CLBLM_R_X5Y148_SLICE_X7Y148_DO5),
.O6(CLBLM_R_X5Y148_SLICE_X7Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffeee)
  ) CLBLM_R_X5Y148_SLICE_X7Y148_CLUT (
.I0(CLBLL_L_X4Y145_SLICE_X5Y145_AO6),
.I1(CLBLM_L_X8Y146_SLICE_X11Y146_BO6),
.I2(CLBLM_L_X10Y143_SLICE_X12Y143_BO5),
.I3(CLBLM_R_X3Y149_SLICE_X3Y149_BQ),
.I4(CLBLM_R_X5Y148_SLICE_X7Y148_DO6),
.I5(CLBLM_R_X5Y148_SLICE_X7Y148_BO6),
.O5(CLBLM_R_X5Y148_SLICE_X7Y148_CO5),
.O6(CLBLM_R_X5Y148_SLICE_X7Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h2f220f000f000f00)
  ) CLBLM_R_X5Y148_SLICE_X7Y148_BLUT (
.I0(CLBLM_R_X11Y149_SLICE_X14Y149_AQ),
.I1(CLBLM_L_X8Y150_SLICE_X10Y150_A5Q),
.I2(CLBLM_R_X5Y145_SLICE_X7Y145_BO6),
.I3(CLBLL_L_X4Y144_SLICE_X5Y144_D5Q),
.I4(CLBLM_L_X10Y144_SLICE_X13Y144_CO6),
.I5(CLBLM_R_X7Y148_SLICE_X9Y148_CQ),
.O5(CLBLM_R_X5Y148_SLICE_X7Y148_BO5),
.O6(CLBLM_R_X5Y148_SLICE_X7Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000001)
  ) CLBLM_R_X5Y148_SLICE_X7Y148_ALUT (
.I0(CLBLM_L_X10Y150_SLICE_X13Y150_CQ),
.I1(CLBLM_R_X7Y149_SLICE_X8Y149_CQ),
.I2(CLBLM_R_X5Y150_SLICE_X6Y150_AQ),
.I3(CLBLM_R_X5Y146_SLICE_X7Y146_BQ),
.I4(CLBLM_R_X5Y143_SLICE_X7Y143_AQ),
.I5(CLBLM_R_X7Y147_SLICE_X9Y147_BQ),
.O5(CLBLM_R_X5Y148_SLICE_X7Y148_AO5),
.O6(CLBLM_R_X5Y148_SLICE_X7Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y149_SLICE_X6Y149_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y149_SLICE_X6Y149_AO5),
.Q(CLBLM_R_X5Y149_SLICE_X6Y149_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y149_SLICE_X6Y149_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y149_SLICE_X6Y149_DO5),
.Q(CLBLM_R_X5Y149_SLICE_X6Y149_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y149_SLICE_X6Y149_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y149_SLICE_X6Y149_AO6),
.Q(CLBLM_R_X5Y149_SLICE_X6Y149_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y149_SLICE_X6Y149_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y149_SLICE_X6Y149_BO6),
.Q(CLBLM_R_X5Y149_SLICE_X6Y149_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y149_SLICE_X6Y149_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y149_SLICE_X6Y149_CO6),
.Q(CLBLM_R_X5Y149_SLICE_X6Y149_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y149_SLICE_X6Y149_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y149_SLICE_X6Y149_DO6),
.Q(CLBLM_R_X5Y149_SLICE_X6Y149_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccaaccaaf0fff000)
  ) CLBLM_R_X5Y149_SLICE_X6Y149_DLUT (
.I0(CLBLL_L_X4Y150_SLICE_X5Y150_BQ),
.I1(CLBLM_R_X5Y152_SLICE_X6Y152_DQ),
.I2(CLBLL_L_X4Y146_SLICE_X5Y146_B5Q),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X8Y150_SLICE_X11Y150_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X5Y149_SLICE_X6Y149_DO5),
.O6(CLBLM_R_X5Y149_SLICE_X6Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaffccaaaa00cc)
  ) CLBLM_R_X5Y149_SLICE_X6Y149_CLUT (
.I0(CLBLL_L_X4Y147_SLICE_X5Y147_BQ),
.I1(CLBLM_R_X5Y149_SLICE_X6Y149_CQ),
.I2(1'b1),
.I3(CLBLM_L_X10Y143_SLICE_X12Y143_BO5),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X5Y143_SLICE_X6Y143_CQ),
.O5(CLBLM_R_X5Y149_SLICE_X6Y149_CO5),
.O6(CLBLM_R_X5Y149_SLICE_X6Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffcca0cca0cca0)
  ) CLBLM_R_X5Y149_SLICE_X6Y149_BLUT (
.I0(CLBLM_L_X10Y150_SLICE_X12Y150_AQ),
.I1(CLBLM_L_X8Y148_SLICE_X11Y148_DQ),
.I2(CLBLL_L_X4Y149_SLICE_X4Y149_D5Q),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X5Y148_SLICE_X6Y148_CO5),
.I5(CLBLL_L_X4Y152_SLICE_X5Y152_B5Q),
.O5(CLBLM_R_X5Y149_SLICE_X6Y149_BO5),
.O6(CLBLM_R_X5Y149_SLICE_X6Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa0afa0acfcfc0c0)
  ) CLBLM_R_X5Y149_SLICE_X6Y149_ALUT (
.I0(CLBLL_L_X4Y148_SLICE_X5Y148_B5Q),
.I1(CLBLM_R_X7Y147_SLICE_X8Y147_D5Q),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_L_X8Y149_SLICE_X11Y149_CQ),
.I4(CLBLM_R_X5Y150_SLICE_X6Y150_CQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y149_SLICE_X6Y149_AO5),
.O6(CLBLM_R_X5Y149_SLICE_X6Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y149_SLICE_X7Y149_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y149_SLICE_X7Y149_BO5),
.Q(CLBLM_R_X5Y149_SLICE_X7Y149_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y149_SLICE_X7Y149_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y149_SLICE_X7Y149_CO5),
.Q(CLBLM_R_X5Y149_SLICE_X7Y149_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y149_SLICE_X7Y149_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y149_SLICE_X7Y149_DO5),
.Q(CLBLM_R_X5Y149_SLICE_X7Y149_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y149_SLICE_X7Y149_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y149_SLICE_X7Y149_AO6),
.Q(CLBLM_R_X5Y149_SLICE_X7Y149_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y149_SLICE_X7Y149_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y149_SLICE_X7Y149_BO6),
.Q(CLBLM_R_X5Y149_SLICE_X7Y149_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y149_SLICE_X7Y149_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y149_SLICE_X7Y149_CO6),
.Q(CLBLM_R_X5Y149_SLICE_X7Y149_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y149_SLICE_X7Y149_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y149_SLICE_X7Y149_DO6),
.Q(CLBLM_R_X5Y149_SLICE_X7Y149_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'he2e2e2e2ffcc3300)
  ) CLBLM_R_X5Y149_SLICE_X7Y149_DLUT (
.I0(CLBLM_L_X8Y142_SLICE_X11Y142_CQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X5Y140_SLICE_X7Y140_B5Q),
.I3(CLBLM_R_X7Y152_SLICE_X9Y152_C5Q),
.I4(CLBLM_R_X5Y149_SLICE_X7Y149_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y149_SLICE_X7Y149_DO5),
.O6(CLBLM_R_X5Y149_SLICE_X7Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa33aaccf0aaf0aa)
  ) CLBLM_R_X5Y149_SLICE_X7Y149_CLUT (
.I0(CLBLM_L_X8Y149_SLICE_X10Y149_AQ),
.I1(CLBLM_R_X5Y147_SLICE_X7Y147_A5Q),
.I2(CLBLL_L_X4Y151_SLICE_X5Y151_CQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X3Y151_SLICE_X3Y151_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y149_SLICE_X7Y149_CO5),
.O6(CLBLM_R_X5Y149_SLICE_X7Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcfc0c0fa0afa0a)
  ) CLBLM_R_X5Y149_SLICE_X7Y149_BLUT (
.I0(CLBLM_R_X7Y145_SLICE_X8Y145_CQ),
.I1(CLBLM_R_X5Y152_SLICE_X6Y152_A5Q),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X7Y150_SLICE_X8Y150_CQ),
.I4(CLBLM_R_X7Y144_SLICE_X9Y144_DQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y149_SLICE_X7Y149_BO5),
.O6(CLBLM_R_X5Y149_SLICE_X7Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00fafaff003232)
  ) CLBLM_R_X5Y149_SLICE_X7Y149_ALUT (
.I0(CLBLM_L_X8Y142_SLICE_X10Y142_C5Q),
.I1(CLBLM_R_X5Y149_SLICE_X6Y149_D5Q),
.I2(CLBLM_R_X5Y149_SLICE_X7Y149_AQ),
.I3(CLBLM_R_X3Y150_SLICE_X3Y150_CQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_L_X8Y150_SLICE_X11Y150_B5Q),
.O5(CLBLM_R_X5Y149_SLICE_X7Y149_AO5),
.O6(CLBLM_R_X5Y149_SLICE_X7Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y150_SLICE_X6Y150_A5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y150_SLICE_X6Y150_AO5),
.Q(CLBLM_R_X5Y150_SLICE_X6Y150_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y150_SLICE_X6Y150_C5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y150_SLICE_X6Y150_CO5),
.Q(CLBLM_R_X5Y150_SLICE_X6Y150_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y150_SLICE_X6Y150_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y150_SLICE_X6Y150_AO6),
.Q(CLBLM_R_X5Y150_SLICE_X6Y150_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y150_SLICE_X6Y150_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y150_SLICE_X6Y150_BO6),
.Q(CLBLM_R_X5Y150_SLICE_X6Y150_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y150_SLICE_X6Y150_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y150_SLICE_X6Y150_CO6),
.Q(CLBLM_R_X5Y150_SLICE_X6Y150_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y150_SLICE_X6Y150_D_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y150_SLICE_X6Y150_DO6),
.Q(CLBLM_R_X5Y150_SLICE_X6Y150_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccf00fcccc0000)
  ) CLBLM_R_X5Y150_SLICE_X6Y150_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y145_SLICE_X8Y145_CQ),
.I2(CLBLM_R_X5Y150_SLICE_X7Y150_BO5),
.I3(CLBLM_R_X5Y150_SLICE_X6Y150_DQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X3Y152_SLICE_X2Y152_BQ),
.O5(CLBLM_R_X5Y150_SLICE_X6Y150_DO5),
.O6(CLBLM_R_X5Y150_SLICE_X6Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefe5454ff55aa00)
  ) CLBLM_R_X5Y150_SLICE_X6Y150_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X7Y145_SLICE_X9Y145_DQ),
.I2(CLBLM_L_X8Y152_SLICE_X10Y152_DQ),
.I3(CLBLL_L_X4Y150_SLICE_X5Y150_AQ),
.I4(CLBLM_R_X5Y144_SLICE_X6Y144_BQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y150_SLICE_X6Y150_CO5),
.O6(CLBLM_R_X5Y150_SLICE_X6Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf6f6f6f606060606)
  ) CLBLM_R_X5Y150_SLICE_X6Y150_BLUT (
.I0(CLBLL_L_X4Y153_SLICE_X5Y153_BQ),
.I1(CLBLM_R_X7Y146_SLICE_X9Y146_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X5Y154_SLICE_X7Y154_CQ),
.O5(CLBLM_R_X5Y150_SLICE_X6Y150_BO5),
.O6(CLBLM_R_X5Y150_SLICE_X6Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf6f60606afa0afa0)
  ) CLBLM_R_X5Y150_SLICE_X6Y150_ALUT (
.I0(CLBLM_L_X10Y147_SLICE_X13Y147_BQ),
.I1(CLBLM_R_X5Y153_SLICE_X6Y153_AQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X5Y152_SLICE_X6Y152_A5Q),
.I4(CLBLL_L_X2Y148_SLICE_X0Y148_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y150_SLICE_X6Y150_AO5),
.O6(CLBLM_R_X5Y150_SLICE_X6Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y150_SLICE_X7Y150_A5_FDSE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y150_SLICE_X7Y150_AO5),
.Q(CLBLM_R_X5Y150_SLICE_X7Y150_A5Q),
.S(CLBLM_R_X11Y148_SLICE_X15Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y150_SLICE_X7Y150_A_FDSE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y150_SLICE_X7Y150_AO6),
.Q(CLBLM_R_X5Y150_SLICE_X7Y150_AQ),
.S(CLBLM_R_X11Y148_SLICE_X15Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h44ff44ff44444444)
  ) CLBLM_R_X5Y150_SLICE_X7Y150_DLUT (
.I0(CLBLM_L_X10Y143_SLICE_X12Y143_AO5),
.I1(CLBLM_R_X5Y154_SLICE_X7Y154_CQ),
.I2(1'b1),
.I3(CLBLM_L_X8Y142_SLICE_X10Y142_BO5),
.I4(1'b1),
.I5(CLBLL_L_X4Y151_SLICE_X5Y151_BQ),
.O5(CLBLM_R_X5Y150_SLICE_X7Y150_DO5),
.O6(CLBLM_R_X5Y150_SLICE_X7Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000001)
  ) CLBLM_R_X5Y150_SLICE_X7Y150_CLUT (
.I0(CLBLM_R_X5Y152_SLICE_X7Y152_AQ),
.I1(CLBLM_R_X7Y150_SLICE_X8Y150_BQ),
.I2(CLBLM_R_X7Y148_SLICE_X9Y148_BQ),
.I3(CLBLL_L_X4Y147_SLICE_X4Y147_CQ),
.I4(CLBLL_L_X4Y149_SLICE_X4Y149_B5Q),
.I5(CLBLM_R_X5Y150_SLICE_X6Y150_BQ),
.O5(CLBLM_R_X5Y150_SLICE_X7Y150_CO5),
.O6(CLBLM_R_X5Y150_SLICE_X7Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff7fffffff3fffff)
  ) CLBLM_R_X5Y150_SLICE_X7Y150_BLUT (
.I0(CLBLM_R_X5Y150_SLICE_X6Y150_DQ),
.I1(CLBLM_R_X7Y151_SLICE_X9Y151_DQ),
.I2(CLBLM_L_X8Y151_SLICE_X10Y151_DQ),
.I3(CLBLM_L_X8Y152_SLICE_X11Y152_CO6),
.I4(CLBLM_R_X5Y151_SLICE_X6Y151_DQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y150_SLICE_X7Y150_BO5),
.O6(CLBLM_R_X5Y150_SLICE_X7Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00000aaaa0000)
  ) CLBLM_R_X5Y150_SLICE_X7Y150_ALUT (
.I0(CLBLM_R_X5Y152_SLICE_X7Y152_CQ),
.I1(1'b1),
.I2(CLBLL_L_X4Y150_SLICE_X5Y150_DQ),
.I3(1'b1),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y150_SLICE_X7Y150_AO5),
.O6(CLBLM_R_X5Y150_SLICE_X7Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y151_SLICE_X6Y151_A5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y151_SLICE_X6Y151_AO5),
.Q(CLBLM_R_X5Y151_SLICE_X6Y151_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y151_SLICE_X6Y151_B5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y151_SLICE_X6Y151_BO5),
.Q(CLBLM_R_X5Y151_SLICE_X6Y151_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y151_SLICE_X6Y151_D5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y151_SLICE_X6Y151_DO5),
.Q(CLBLM_R_X5Y151_SLICE_X6Y151_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y151_SLICE_X6Y151_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y151_SLICE_X6Y151_AO6),
.Q(CLBLM_R_X5Y151_SLICE_X6Y151_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y151_SLICE_X6Y151_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y151_SLICE_X6Y151_BO6),
.Q(CLBLM_R_X5Y151_SLICE_X6Y151_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y151_SLICE_X6Y151_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y151_SLICE_X6Y151_CO6),
.Q(CLBLM_R_X5Y151_SLICE_X6Y151_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y151_SLICE_X6Y151_D_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y151_SLICE_X6Y151_DO6),
.Q(CLBLM_R_X5Y151_SLICE_X6Y151_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'heecceeccf5a0f5a0)
  ) CLBLM_R_X5Y151_SLICE_X6Y151_DLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X5Y151_SLICE_X7Y151_CO6),
.I2(CLBLM_L_X8Y151_SLICE_X10Y151_DQ),
.I3(CLBLM_R_X5Y151_SLICE_X6Y151_A5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y151_SLICE_X6Y151_DO5),
.O6(CLBLM_R_X5Y151_SLICE_X6Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf8f0f8f088008800)
  ) CLBLM_R_X5Y151_SLICE_X6Y151_CLUT (
.I0(CLBLL_L_X4Y144_SLICE_X4Y144_BO6),
.I1(CLBLM_R_X5Y150_SLICE_X7Y150_CO6),
.I2(CLBLM_R_X7Y145_SLICE_X9Y145_DQ),
.I3(CLBLM_R_X7Y151_SLICE_X8Y151_DO5),
.I4(1'b1),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X5Y151_SLICE_X6Y151_CO5),
.O6(CLBLM_R_X5Y151_SLICE_X6Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'heeee2222fc30fc30)
  ) CLBLM_R_X5Y151_SLICE_X6Y151_BLUT (
.I0(CLBLM_R_X7Y152_SLICE_X9Y152_D5Q),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(RIOB33_X105Y123_IOB_X1Y124_I),
.I3(CLBLM_R_X11Y151_SLICE_X15Y151_AQ),
.I4(CLBLM_R_X5Y153_SLICE_X7Y153_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y151_SLICE_X6Y151_BO5),
.O6(CLBLM_R_X5Y151_SLICE_X6Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbbb8888f3c0f3c0)
  ) CLBLM_R_X5Y151_SLICE_X6Y151_ALUT (
.I0(CLBLM_R_X3Y148_SLICE_X2Y148_B5Q),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X5Y151_SLICE_X6Y151_AQ),
.I3(CLBLM_R_X5Y149_SLICE_X6Y149_BQ),
.I4(CLBLM_R_X7Y150_SLICE_X8Y150_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y151_SLICE_X6Y151_AO5),
.O6(CLBLM_R_X5Y151_SLICE_X6Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y151_SLICE_X7Y151_A5_FDSE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y151_SLICE_X7Y151_AO5),
.Q(CLBLM_R_X5Y151_SLICE_X7Y151_A5Q),
.S(CLBLL_L_X4Y145_SLICE_X5Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y151_SLICE_X7Y151_A_FDSE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y151_SLICE_X7Y151_AO6),
.Q(CLBLM_R_X5Y151_SLICE_X7Y151_AQ),
.S(CLBLL_L_X4Y145_SLICE_X5Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff5f0fffff5500)
  ) CLBLM_R_X5Y151_SLICE_X7Y151_DLUT (
.I0(CLBLM_L_X10Y143_SLICE_X12Y143_AO6),
.I1(1'b1),
.I2(CLBLM_L_X10Y143_SLICE_X12Y143_BO5),
.I3(CLBLL_L_X4Y150_SLICE_X5Y150_AQ),
.I4(CLBLM_L_X12Y149_SLICE_X16Y149_CO6),
.I5(CLBLM_L_X8Y151_SLICE_X10Y151_AQ),
.O5(CLBLM_R_X5Y151_SLICE_X7Y151_DO5),
.O6(CLBLM_R_X5Y151_SLICE_X7Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h4555100000000000)
  ) CLBLM_R_X5Y151_SLICE_X7Y151_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X8Y152_SLICE_X11Y152_CO6),
.I2(CLBLM_R_X7Y151_SLICE_X9Y151_DQ),
.I3(CLBLM_L_X8Y151_SLICE_X10Y151_DQ),
.I4(CLBLM_R_X5Y151_SLICE_X6Y151_DQ),
.I5(CLBLM_R_X3Y152_SLICE_X2Y152_BQ),
.O5(CLBLM_R_X5Y151_SLICE_X7Y151_CO5),
.O6(CLBLM_R_X5Y151_SLICE_X7Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h55fffffffffefffe)
  ) CLBLM_R_X5Y151_SLICE_X7Y151_BLUT (
.I0(CLBLM_R_X7Y143_SLICE_X9Y143_CQ),
.I1(CLBLM_R_X3Y151_SLICE_X3Y151_BQ),
.I2(CLBLL_L_X4Y153_SLICE_X5Y153_BQ),
.I3(CLBLL_L_X4Y151_SLICE_X5Y151_AQ),
.I4(CLBLM_R_X7Y143_SLICE_X9Y143_BQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y151_SLICE_X7Y151_BO5),
.O6(CLBLM_R_X5Y151_SLICE_X7Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000cc00cc00)
  ) CLBLM_R_X5Y151_SLICE_X7Y151_ALUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y148_SLICE_X4Y148_BQ),
.I2(CLBLM_R_X5Y152_SLICE_X6Y152_C5Q),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y151_SLICE_X7Y151_AO5),
.O6(CLBLM_R_X5Y151_SLICE_X7Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y152_SLICE_X6Y152_A5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y152_SLICE_X6Y152_AO5),
.Q(CLBLM_R_X5Y152_SLICE_X6Y152_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y152_SLICE_X6Y152_B5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y152_SLICE_X6Y152_BO5),
.Q(CLBLM_R_X5Y152_SLICE_X6Y152_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y152_SLICE_X6Y152_C5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y152_SLICE_X6Y152_CO5),
.Q(CLBLM_R_X5Y152_SLICE_X6Y152_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y152_SLICE_X6Y152_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y152_SLICE_X6Y152_AO6),
.Q(CLBLM_R_X5Y152_SLICE_X6Y152_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y152_SLICE_X6Y152_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y152_SLICE_X6Y152_BO6),
.Q(CLBLM_R_X5Y152_SLICE_X6Y152_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y152_SLICE_X6Y152_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y152_SLICE_X6Y152_CO6),
.Q(CLBLM_R_X5Y152_SLICE_X6Y152_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y152_SLICE_X6Y152_D_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y152_SLICE_X6Y152_DO6),
.Q(CLBLM_R_X5Y152_SLICE_X6Y152_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfb51fe54aa00aa00)
  ) CLBLM_R_X5Y152_SLICE_X6Y152_DLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(RIOB33_X105Y107_IOB_X1Y107_I),
.I2(CLBLM_R_X5Y152_SLICE_X6Y152_DQ),
.I3(CLBLM_R_X7Y153_SLICE_X8Y153_AQ),
.I4(CLBLM_R_X5Y152_SLICE_X6Y152_BQ),
.I5(CLBLM_L_X8Y143_SLICE_X11Y143_A5Q),
.O5(CLBLM_R_X5Y152_SLICE_X6Y152_DO5),
.O6(CLBLM_R_X5Y152_SLICE_X6Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccf0ccf0ff550055)
  ) CLBLM_R_X5Y152_SLICE_X6Y152_CLUT (
.I0(CLBLL_L_X4Y152_SLICE_X5Y152_BQ),
.I1(CLBLM_R_X7Y149_SLICE_X9Y149_C5Q),
.I2(RIOB33_X105Y113_IOB_X1Y113_I),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLL_L_X4Y153_SLICE_X4Y153_BQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y152_SLICE_X6Y152_CO5),
.O6(CLBLM_R_X5Y152_SLICE_X6Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0aaf0aaccffcc00)
  ) CLBLM_R_X5Y152_SLICE_X6Y152_BLUT (
.I0(RIOB33_X105Y107_IOB_X1Y107_I),
.I1(CLBLM_R_X5Y152_SLICE_X6Y152_BQ),
.I2(CLBLL_L_X2Y150_SLICE_X1Y150_A5Q),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLL_L_X4Y151_SLICE_X5Y151_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X5Y152_SLICE_X6Y152_BO5),
.O6(CLBLM_R_X5Y152_SLICE_X6Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0ff000cacacaca)
  ) CLBLM_R_X5Y152_SLICE_X6Y152_ALUT (
.I0(RIOB33_X105Y117_IOB_X1Y117_I),
.I1(CLBLM_R_X7Y152_SLICE_X8Y152_CQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLL_L_X4Y150_SLICE_X5Y150_D5Q),
.I4(CLBLM_R_X3Y150_SLICE_X2Y150_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y152_SLICE_X6Y152_AO5),
.O6(CLBLM_R_X5Y152_SLICE_X6Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y152_SLICE_X7Y152_D5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y152_SLICE_X7Y152_DO5),
.Q(CLBLM_R_X5Y152_SLICE_X7Y152_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y152_SLICE_X7Y152_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y152_SLICE_X7Y152_AO6),
.Q(CLBLM_R_X5Y152_SLICE_X7Y152_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y152_SLICE_X7Y152_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y152_SLICE_X7Y152_BO6),
.Q(CLBLM_R_X5Y152_SLICE_X7Y152_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y152_SLICE_X7Y152_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y152_SLICE_X7Y152_CO6),
.Q(CLBLM_R_X5Y152_SLICE_X7Y152_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y152_SLICE_X7Y152_D_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y152_SLICE_X7Y152_DO6),
.Q(CLBLM_R_X5Y152_SLICE_X7Y152_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccff00338b8bb8b8)
  ) CLBLM_R_X5Y152_SLICE_X7Y152_DLUT (
.I0(CLBLM_R_X3Y147_SLICE_X3Y147_AQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X7Y143_SLICE_X9Y143_CQ),
.I3(CLBLL_L_X4Y152_SLICE_X5Y152_BQ),
.I4(CLBLM_L_X8Y148_SLICE_X10Y148_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X5Y152_SLICE_X7Y152_DO5),
.O6(CLBLM_R_X5Y152_SLICE_X7Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafa5050eeee4444)
  ) CLBLM_R_X5Y152_SLICE_X7Y152_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X5Y152_SLICE_X7Y152_CQ),
.I2(CLBLM_R_X5Y152_SLICE_X7Y152_BQ),
.I3(1'b1),
.I4(CLBLM_L_X8Y152_SLICE_X10Y152_DQ),
.I5(CLBLM_L_X10Y143_SLICE_X12Y143_BO6),
.O5(CLBLM_R_X5Y152_SLICE_X7Y152_CO5),
.O6(CLBLM_R_X5Y152_SLICE_X7Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0aa88ffcc)
  ) CLBLM_R_X5Y152_SLICE_X7Y152_BLUT (
.I0(CLBLM_R_X5Y144_SLICE_X6Y144_DQ),
.I1(CLBLM_R_X5Y152_SLICE_X7Y152_BQ),
.I2(CLBLM_R_X7Y150_SLICE_X9Y150_C5Q),
.I3(CLBLM_R_X5Y151_SLICE_X7Y151_A5Q),
.I4(CLBLM_R_X3Y148_SLICE_X2Y148_D5Q),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X5Y152_SLICE_X7Y152_BO5),
.O6(CLBLM_R_X5Y152_SLICE_X7Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa0ff00ff0)
  ) CLBLM_R_X5Y152_SLICE_X7Y152_ALUT (
.I0(CLBLL_L_X4Y152_SLICE_X5Y152_B5Q),
.I1(1'b1),
.I2(CLBLM_R_X5Y153_SLICE_X6Y153_AQ),
.I3(CLBLM_L_X8Y149_SLICE_X10Y149_BQ),
.I4(1'b1),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X5Y152_SLICE_X7Y152_AO5),
.O6(CLBLM_R_X5Y152_SLICE_X7Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y153_SLICE_X6Y153_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y153_SLICE_X6Y153_AO6),
.Q(CLBLM_R_X5Y153_SLICE_X6Y153_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y153_SLICE_X6Y153_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y153_SLICE_X6Y153_BO6),
.Q(CLBLM_R_X5Y153_SLICE_X6Y153_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y153_SLICE_X6Y153_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y153_SLICE_X6Y153_CO6),
.Q(CLBLM_R_X5Y153_SLICE_X6Y153_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y153_SLICE_X6Y153_D_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y153_SLICE_X6Y153_DO6),
.Q(CLBLM_R_X5Y153_SLICE_X6Y153_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hee44ee44ea40ea40)
  ) CLBLM_R_X5Y153_SLICE_X6Y153_DLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X10Y143_SLICE_X12Y143_BO6),
.I2(CLBLM_R_X5Y153_SLICE_X6Y153_DQ),
.I3(CLBLM_R_X7Y154_SLICE_X8Y154_AQ),
.I4(1'b1),
.I5(CLBLM_R_X3Y152_SLICE_X2Y152_CQ),
.O5(CLBLM_R_X5Y153_SLICE_X6Y153_DO5),
.O6(CLBLM_R_X5Y153_SLICE_X6Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffee33333322)
  ) CLBLM_R_X5Y153_SLICE_X6Y153_CLUT (
.I0(CLBLM_R_X5Y153_SLICE_X6Y153_BQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(1'b1),
.I3(CLBLM_R_X5Y152_SLICE_X6Y152_B5Q),
.I4(CLBLM_R_X5Y152_SLICE_X7Y152_DQ),
.I5(CLBLM_L_X8Y150_SLICE_X11Y150_BQ),
.O5(CLBLM_R_X5Y153_SLICE_X6Y153_CO5),
.O6(CLBLM_R_X5Y153_SLICE_X6Y153_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000ff001515)
  ) CLBLM_R_X5Y153_SLICE_X6Y153_BLUT (
.I0(CLBLM_R_X5Y152_SLICE_X7Y152_DQ),
.I1(CLBLM_R_X5Y153_SLICE_X6Y153_BQ),
.I2(CLBLM_R_X5Y153_SLICE_X6Y153_CQ),
.I3(CLBLM_R_X7Y152_SLICE_X9Y152_D5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X5Y152_SLICE_X6Y152_B5Q),
.O5(CLBLM_R_X5Y153_SLICE_X6Y153_BO5),
.O6(CLBLM_R_X5Y153_SLICE_X6Y153_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaafccffccf)
  ) CLBLM_R_X5Y153_SLICE_X6Y153_ALUT (
.I0(CLBLM_R_X5Y153_SLICE_X6Y153_CQ),
.I1(CLBLL_L_X2Y148_SLICE_X0Y148_B5Q),
.I2(CLBLM_R_X5Y153_SLICE_X6Y153_AQ),
.I3(CLBLM_R_X3Y152_SLICE_X2Y152_DO6),
.I4(1'b1),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X5Y153_SLICE_X6Y153_AO5),
.O6(CLBLM_R_X5Y153_SLICE_X6Y153_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y153_SLICE_X7Y153_A5_FDSE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y153_SLICE_X7Y153_AO5),
.Q(CLBLM_R_X5Y153_SLICE_X7Y153_A5Q),
.S(CLBLL_L_X2Y147_SLICE_X1Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y153_SLICE_X7Y153_A_FDSE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y153_SLICE_X7Y153_AO6),
.Q(CLBLM_R_X5Y153_SLICE_X7Y153_AQ),
.S(CLBLL_L_X2Y147_SLICE_X1Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333333300000000)
  ) CLBLM_R_X5Y153_SLICE_X7Y153_DLUT (
.I0(1'b1),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X3Y151_SLICE_X3Y151_BQ),
.O5(CLBLM_R_X5Y153_SLICE_X7Y153_DO5),
.O6(CLBLM_R_X5Y153_SLICE_X7Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffeffffffffff)
  ) CLBLM_R_X5Y153_SLICE_X7Y153_CLUT (
.I0(CLBLM_R_X3Y150_SLICE_X2Y150_CO5),
.I1(CLBLM_L_X10Y150_SLICE_X12Y150_CQ),
.I2(CLBLL_L_X4Y154_SLICE_X4Y154_AQ),
.I3(CLBLM_R_X7Y153_SLICE_X8Y153_DO5),
.I4(CLBLM_R_X7Y154_SLICE_X9Y154_AO6),
.I5(CLBLL_L_X4Y154_SLICE_X4Y154_BO6),
.O5(CLBLM_R_X5Y153_SLICE_X7Y153_CO5),
.O6(CLBLM_R_X5Y153_SLICE_X7Y153_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000cc8ccc4c)
  ) CLBLM_R_X5Y153_SLICE_X7Y153_BLUT (
.I0(CLBLM_R_X7Y150_SLICE_X9Y150_C5Q),
.I1(CLBLL_L_X4Y153_SLICE_X5Y153_CO6),
.I2(CLBLM_R_X7Y149_SLICE_X9Y149_DQ),
.I3(CLBLM_L_X10Y150_SLICE_X12Y150_CQ),
.I4(CLBLM_R_X7Y144_SLICE_X9Y144_B5Q),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X5Y153_SLICE_X7Y153_BO5),
.O6(CLBLM_R_X5Y153_SLICE_X7Y153_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00aaaa0000)
  ) CLBLM_R_X5Y153_SLICE_X7Y153_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_L_X8Y151_SLICE_X11Y151_A5Q),
.I4(CLBLM_R_X7Y155_SLICE_X8Y155_BQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y153_SLICE_X7Y153_AO5),
.O6(CLBLM_R_X5Y153_SLICE_X7Y153_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y154_SLICE_X6Y154_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y154_SLICE_X6Y154_AO6),
.Q(CLBLM_R_X5Y154_SLICE_X6Y154_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y154_SLICE_X6Y154_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y154_SLICE_X6Y154_DO5),
.O6(CLBLM_R_X5Y154_SLICE_X6Y154_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y154_SLICE_X6Y154_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y154_SLICE_X6Y154_CO5),
.O6(CLBLM_R_X5Y154_SLICE_X6Y154_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y154_SLICE_X6Y154_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y154_SLICE_X6Y154_BO5),
.O6(CLBLM_R_X5Y154_SLICE_X6Y154_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccaaaaccccf0f0)
  ) CLBLM_R_X5Y154_SLICE_X6Y154_ALUT (
.I0(CLBLL_L_X2Y150_SLICE_X1Y150_AQ),
.I1(CLBLM_L_X8Y153_SLICE_X10Y153_CQ),
.I2(CLBLM_R_X5Y154_SLICE_X6Y154_AQ),
.I3(1'b1),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_L_X10Y143_SLICE_X12Y143_AO6),
.O5(CLBLM_R_X5Y154_SLICE_X6Y154_AO5),
.O6(CLBLM_R_X5Y154_SLICE_X6Y154_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y154_SLICE_X7Y154_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y154_SLICE_X7Y154_AO6),
.Q(CLBLM_R_X5Y154_SLICE_X7Y154_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y154_SLICE_X7Y154_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y154_SLICE_X7Y154_BO6),
.Q(CLBLM_R_X5Y154_SLICE_X7Y154_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y154_SLICE_X7Y154_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y154_SLICE_X7Y154_CO6),
.Q(CLBLM_R_X5Y154_SLICE_X7Y154_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y154_SLICE_X7Y154_D_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y154_SLICE_X7Y154_DO6),
.Q(CLBLM_R_X5Y154_SLICE_X7Y154_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff780078ff000000)
  ) CLBLM_R_X5Y154_SLICE_X7Y154_DLUT (
.I0(CLBLM_R_X3Y154_SLICE_X3Y154_AQ),
.I1(CLBLM_L_X8Y153_SLICE_X11Y153_BQ),
.I2(CLBLM_R_X5Y154_SLICE_X7Y154_DQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLL_L_X4Y146_SLICE_X4Y146_BQ),
.I5(CLBLM_R_X3Y152_SLICE_X2Y152_BQ),
.O5(CLBLM_R_X5Y154_SLICE_X7Y154_DO5),
.O6(CLBLM_R_X5Y154_SLICE_X7Y154_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaa00aaccaacc)
  ) CLBLM_R_X5Y154_SLICE_X7Y154_CLUT (
.I0(CLBLM_L_X8Y152_SLICE_X11Y152_BQ),
.I1(CLBLM_R_X5Y154_SLICE_X7Y154_CQ),
.I2(1'b1),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X5Y144_SLICE_X7Y144_AQ),
.I5(CLBLM_L_X10Y143_SLICE_X12Y143_AO6),
.O5(CLBLM_R_X5Y154_SLICE_X7Y154_CO5),
.O6(CLBLM_R_X5Y154_SLICE_X7Y154_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa00003030)
  ) CLBLM_R_X5Y154_SLICE_X7Y154_BLUT (
.I0(CLBLM_R_X7Y153_SLICE_X9Y153_BQ),
.I1(CLBLM_R_X5Y154_SLICE_X7Y154_BQ),
.I2(CLBLM_R_X5Y154_SLICE_X7Y154_AQ),
.I3(1'b1),
.I4(CLBLL_L_X4Y152_SLICE_X5Y152_C5Q),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X5Y154_SLICE_X7Y154_BO5),
.O6(CLBLM_R_X5Y154_SLICE_X7Y154_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00ffff0303)
  ) CLBLM_R_X5Y154_SLICE_X7Y154_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y154_SLICE_X7Y154_BQ),
.I2(CLBLM_R_X5Y154_SLICE_X7Y154_AQ),
.I3(CLBLM_R_X7Y149_SLICE_X8Y149_BQ),
.I4(CLBLL_L_X4Y152_SLICE_X5Y152_C5Q),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X5Y154_SLICE_X7Y154_AO5),
.O6(CLBLM_R_X5Y154_SLICE_X7Y154_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y159_SLICE_X6Y159_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y159_SLICE_X6Y159_DO5),
.O6(CLBLM_R_X5Y159_SLICE_X6Y159_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y159_SLICE_X6Y159_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y159_SLICE_X6Y159_CO5),
.O6(CLBLM_R_X5Y159_SLICE_X6Y159_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y159_SLICE_X6Y159_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y159_SLICE_X6Y159_BO5),
.O6(CLBLM_R_X5Y159_SLICE_X6Y159_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaaffaaffaaffaa)
  ) CLBLM_R_X5Y159_SLICE_X6Y159_ALUT (
.I0(CLBLM_R_X7Y145_SLICE_X9Y145_DQ),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_L_X8Y152_SLICE_X10Y152_DQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y159_SLICE_X6Y159_AO5),
.O6(CLBLM_R_X5Y159_SLICE_X6Y159_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y159_SLICE_X7Y159_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y159_SLICE_X7Y159_DO5),
.O6(CLBLM_R_X5Y159_SLICE_X7Y159_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y159_SLICE_X7Y159_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y159_SLICE_X7Y159_CO5),
.O6(CLBLM_R_X5Y159_SLICE_X7Y159_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y159_SLICE_X7Y159_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y159_SLICE_X7Y159_BO5),
.O6(CLBLM_R_X5Y159_SLICE_X7Y159_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y159_SLICE_X7Y159_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y159_SLICE_X7Y159_AO5),
.O6(CLBLM_R_X5Y159_SLICE_X7Y159_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y141_SLICE_X8Y141_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y141_SLICE_X8Y141_AO6),
.Q(CLBLM_R_X7Y141_SLICE_X8Y141_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y141_SLICE_X8Y141_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y141_SLICE_X8Y141_DO5),
.O6(CLBLM_R_X7Y141_SLICE_X8Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y141_SLICE_X8Y141_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y141_SLICE_X8Y141_CO5),
.O6(CLBLM_R_X7Y141_SLICE_X8Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y141_SLICE_X8Y141_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y141_SLICE_X8Y141_BO5),
.O6(CLBLM_R_X7Y141_SLICE_X8Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffddd00000ddd0)
  ) CLBLM_R_X7Y141_SLICE_X8Y141_ALUT (
.I0(CLBLM_R_X5Y149_SLICE_X7Y149_DQ),
.I1(CLBLM_L_X8Y142_SLICE_X11Y142_CQ),
.I2(CLBLM_R_X7Y141_SLICE_X8Y141_AQ),
.I3(CLBLL_L_X4Y140_SLICE_X5Y140_AQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X7Y143_SLICE_X8Y143_BQ),
.O5(CLBLM_R_X7Y141_SLICE_X8Y141_AO5),
.O6(CLBLM_R_X7Y141_SLICE_X8Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y141_SLICE_X9Y141_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y141_SLICE_X9Y141_AO6),
.Q(CLBLM_R_X7Y141_SLICE_X9Y141_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y141_SLICE_X9Y141_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y141_SLICE_X9Y141_DO5),
.O6(CLBLM_R_X7Y141_SLICE_X9Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y141_SLICE_X9Y141_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y141_SLICE_X9Y141_CO5),
.O6(CLBLM_R_X7Y141_SLICE_X9Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y141_SLICE_X9Y141_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y141_SLICE_X9Y141_BO5),
.O6(CLBLM_R_X7Y141_SLICE_X9Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfe32cc00fe32fe32)
  ) CLBLM_R_X7Y141_SLICE_X9Y141_ALUT (
.I0(CLBLM_L_X8Y142_SLICE_X10Y142_A5Q),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X7Y141_SLICE_X9Y141_AQ),
.I3(CLBLM_L_X8Y148_SLICE_X11Y148_C5Q),
.I4(CLBLM_R_X5Y144_SLICE_X6Y144_DQ),
.I5(CLBLM_R_X3Y148_SLICE_X2Y148_D5Q),
.O5(CLBLM_R_X7Y141_SLICE_X9Y141_AO5),
.O6(CLBLM_R_X7Y141_SLICE_X9Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y142_SLICE_X8Y142_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y142_SLICE_X8Y142_AO5),
.Q(CLBLM_R_X7Y142_SLICE_X8Y142_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y142_SLICE_X8Y142_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y142_SLICE_X8Y142_BO5),
.Q(CLBLM_R_X7Y142_SLICE_X8Y142_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y142_SLICE_X8Y142_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y142_SLICE_X8Y142_AO6),
.Q(CLBLM_R_X7Y142_SLICE_X8Y142_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y142_SLICE_X8Y142_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y142_SLICE_X8Y142_BO6),
.Q(CLBLM_R_X7Y142_SLICE_X8Y142_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fffffffffffffff)
  ) CLBLM_R_X7Y142_SLICE_X8Y142_DLUT (
.I0(CLBLM_L_X10Y149_SLICE_X12Y149_A5Q),
.I1(CLBLM_R_X5Y142_SLICE_X6Y142_AQ),
.I2(CLBLM_R_X7Y142_SLICE_X9Y142_AQ),
.I3(CLBLM_R_X11Y146_SLICE_X15Y146_AQ),
.I4(CLBLM_R_X5Y146_SLICE_X7Y146_AQ),
.I5(CLBLM_R_X5Y144_SLICE_X7Y144_BQ),
.O5(CLBLM_R_X7Y142_SLICE_X8Y142_DO5),
.O6(CLBLM_R_X7Y142_SLICE_X8Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff80000000)
  ) CLBLM_R_X7Y142_SLICE_X8Y142_CLUT (
.I0(CLBLM_R_X7Y142_SLICE_X9Y142_AQ),
.I1(CLBLM_R_X5Y142_SLICE_X6Y142_AQ),
.I2(CLBLM_L_X10Y149_SLICE_X12Y149_A5Q),
.I3(CLBLM_R_X11Y146_SLICE_X15Y146_AQ),
.I4(CLBLM_R_X5Y146_SLICE_X7Y146_AQ),
.I5(CLBLM_R_X5Y144_SLICE_X7Y144_BQ),
.O5(CLBLM_R_X7Y142_SLICE_X8Y142_CO5),
.O6(CLBLM_R_X7Y142_SLICE_X8Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccc3c3a9a9aaaa)
  ) CLBLM_R_X7Y142_SLICE_X8Y142_BLUT (
.I0(CLBLM_R_X7Y142_SLICE_X8Y142_B5Q),
.I1(CLBLM_R_X7Y142_SLICE_X8Y142_BQ),
.I2(CLBLM_R_X7Y148_SLICE_X8Y148_DO6),
.I3(1'b1),
.I4(CLBLM_R_X7Y142_SLICE_X8Y142_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X7Y142_SLICE_X8Y142_BO5),
.O6(CLBLM_R_X7Y142_SLICE_X8Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h111100000f0ff0f0)
  ) CLBLM_R_X7Y142_SLICE_X8Y142_ALUT (
.I0(CLBLM_R_X7Y142_SLICE_X8Y142_B5Q),
.I1(CLBLM_R_X7Y142_SLICE_X8Y142_BQ),
.I2(CLBLM_R_X7Y148_SLICE_X8Y148_DO6),
.I3(1'b1),
.I4(CLBLM_R_X7Y142_SLICE_X8Y142_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X7Y142_SLICE_X8Y142_AO5),
.O6(CLBLM_R_X7Y142_SLICE_X8Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y142_SLICE_X9Y142_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y142_SLICE_X10Y142_BO6),
.Q(CLBLM_R_X7Y142_SLICE_X9Y142_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y142_SLICE_X9Y142_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y142_SLICE_X9Y142_DO5),
.Q(CLBLM_R_X7Y142_SLICE_X9Y142_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y142_SLICE_X9Y142_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y142_SLICE_X9Y142_AO6),
.Q(CLBLM_R_X7Y142_SLICE_X9Y142_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y142_SLICE_X9Y142_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y142_SLICE_X9Y142_BO6),
.Q(CLBLM_R_X7Y142_SLICE_X9Y142_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y142_SLICE_X9Y142_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y142_SLICE_X9Y142_CO6),
.Q(CLBLM_R_X7Y142_SLICE_X9Y142_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y142_SLICE_X9Y142_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y142_SLICE_X9Y142_DO6),
.Q(CLBLM_R_X7Y142_SLICE_X9Y142_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfe32fe32bbbb8888)
  ) CLBLM_R_X7Y142_SLICE_X9Y142_DLUT (
.I0(CLBLM_R_X5Y142_SLICE_X6Y142_C5Q),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X7Y142_SLICE_X9Y142_DQ),
.I3(CLBLM_R_X7Y142_SLICE_X9Y142_AQ),
.I4(RIOB33_X105Y111_IOB_X1Y111_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y142_SLICE_X9Y142_DO5),
.O6(CLBLM_R_X7Y142_SLICE_X9Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5a0e4e4f5a0e4e4)
  ) CLBLM_R_X7Y142_SLICE_X9Y142_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X7Y142_SLICE_X9Y142_CQ),
.I2(CLBLM_R_X7Y150_SLICE_X9Y150_B5Q),
.I3(CLBLM_R_X7Y142_SLICE_X9Y142_BQ),
.I4(CLBLM_L_X10Y143_SLICE_X12Y143_BO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y142_SLICE_X9Y142_CO5),
.O6(CLBLM_R_X7Y142_SLICE_X9Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaf0c0aaaaffcc)
  ) CLBLM_R_X7Y142_SLICE_X9Y142_BLUT (
.I0(CLBLM_L_X10Y152_SLICE_X12Y152_BQ),
.I1(CLBLM_R_X7Y142_SLICE_X9Y142_BQ),
.I2(CLBLM_R_X5Y144_SLICE_X6Y144_DQ),
.I3(CLBLL_L_X4Y142_SLICE_X4Y142_A5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X3Y148_SLICE_X2Y148_D5Q),
.O5(CLBLM_R_X7Y142_SLICE_X9Y142_BO5),
.O6(CLBLM_R_X7Y142_SLICE_X9Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaffc3aaaa00c3)
  ) CLBLM_R_X7Y142_SLICE_X9Y142_ALUT (
.I0(CLBLM_R_X7Y150_SLICE_X9Y150_CQ),
.I1(CLBLM_L_X10Y146_SLICE_X12Y146_AO5),
.I2(CLBLM_R_X7Y142_SLICE_X9Y142_AQ),
.I3(CLBLM_L_X8Y149_SLICE_X11Y149_BQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X7Y147_SLICE_X9Y147_CQ),
.O5(CLBLM_R_X7Y142_SLICE_X9Y142_AO5),
.O6(CLBLM_R_X7Y142_SLICE_X9Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y143_SLICE_X8Y143_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y143_SLICE_X8Y143_AO6),
.Q(CLBLM_R_X7Y143_SLICE_X8Y143_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y143_SLICE_X8Y143_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y143_SLICE_X8Y143_BO6),
.Q(CLBLM_R_X7Y143_SLICE_X8Y143_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y143_SLICE_X8Y143_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y143_SLICE_X8Y143_CO6),
.Q(CLBLM_R_X7Y143_SLICE_X8Y143_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y143_SLICE_X8Y143_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y143_SLICE_X8Y143_DO6),
.Q(CLBLM_R_X7Y143_SLICE_X8Y143_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ccccff00f0f0)
  ) CLBLM_R_X7Y143_SLICE_X8Y143_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.I2(CLBLM_R_X7Y143_SLICE_X8Y143_DQ),
.I3(CLBLM_R_X3Y144_SLICE_X2Y144_A5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_L_X10Y143_SLICE_X12Y143_BO5),
.O5(CLBLM_R_X7Y143_SLICE_X8Y143_DO5),
.O6(CLBLM_R_X7Y143_SLICE_X8Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0aaaaf0f08888)
  ) CLBLM_R_X7Y143_SLICE_X8Y143_CLUT (
.I0(CLBLM_L_X10Y143_SLICE_X12Y143_AO6),
.I1(CLBLM_R_X7Y143_SLICE_X8Y143_CQ),
.I2(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.I3(1'b1),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X5Y143_SLICE_X6Y143_BQ),
.O5(CLBLM_R_X7Y143_SLICE_X8Y143_CO5),
.O6(CLBLM_R_X7Y143_SLICE_X8Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haf05fa50fe54fe54)
  ) CLBLM_R_X7Y143_SLICE_X8Y143_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X7Y143_SLICE_X8Y143_BQ),
.I2(CLBLM_R_X7Y142_SLICE_X8Y142_AQ),
.I3(CLBLM_R_X7Y150_SLICE_X8Y150_C5Q),
.I4(CLBLM_R_X7Y141_SLICE_X9Y141_AQ),
.I5(CLBLM_L_X10Y143_SLICE_X12Y143_BO6),
.O5(CLBLM_R_X7Y143_SLICE_X8Y143_BO5),
.O6(CLBLM_R_X7Y143_SLICE_X8Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hddd88888ddd8ddd8)
  ) CLBLM_R_X7Y143_SLICE_X8Y143_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X7Y142_SLICE_X9Y142_BQ),
.I2(CLBLM_R_X7Y143_SLICE_X8Y143_AQ),
.I3(CLBLL_L_X2Y144_SLICE_X1Y144_AQ),
.I4(CLBLM_R_X5Y144_SLICE_X6Y144_CQ),
.I5(CLBLM_R_X3Y147_SLICE_X3Y147_BQ),
.O5(CLBLM_R_X7Y143_SLICE_X8Y143_AO5),
.O6(CLBLM_R_X7Y143_SLICE_X8Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y143_SLICE_X9Y143_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y143_SLICE_X9Y143_AO6),
.Q(CLBLM_R_X7Y143_SLICE_X9Y143_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y143_SLICE_X9Y143_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y143_SLICE_X9Y143_BO6),
.Q(CLBLM_R_X7Y143_SLICE_X9Y143_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y143_SLICE_X9Y143_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y143_SLICE_X9Y143_CO6),
.Q(CLBLM_R_X7Y143_SLICE_X9Y143_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y143_SLICE_X9Y143_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y143_SLICE_X9Y143_DO6),
.Q(CLBLM_R_X7Y143_SLICE_X9Y143_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0afa0afafa0afa0)
  ) CLBLM_R_X7Y143_SLICE_X9Y143_DLUT (
.I0(CLBLM_L_X10Y142_SLICE_X13Y142_AQ),
.I1(1'b1),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X7Y143_SLICE_X9Y143_BQ),
.I4(1'b1),
.I5(CLBLM_R_X5Y148_SLICE_X6Y148_BQ),
.O5(CLBLM_R_X7Y143_SLICE_X9Y143_DO5),
.O6(CLBLM_R_X7Y143_SLICE_X9Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5f5f5e4e4b1e4)
  ) CLBLM_R_X7Y143_SLICE_X9Y143_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X7Y143_SLICE_X9Y143_CQ),
.I2(CLBLL_L_X4Y144_SLICE_X5Y144_B5Q),
.I3(CLBLM_R_X7Y143_SLICE_X9Y143_BQ),
.I4(CLBLM_R_X7Y144_SLICE_X8Y144_BO6),
.I5(CLBLL_L_X2Y148_SLICE_X0Y148_B5Q),
.O5(CLBLM_R_X7Y143_SLICE_X9Y143_CO5),
.O6(CLBLM_R_X7Y143_SLICE_X9Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff9fff90f090f09)
  ) CLBLM_R_X7Y143_SLICE_X9Y143_BLUT (
.I0(CLBLM_R_X7Y144_SLICE_X8Y144_BO6),
.I1(CLBLM_R_X7Y143_SLICE_X9Y143_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLL_L_X2Y148_SLICE_X0Y148_B5Q),
.I4(1'b1),
.I5(CLBLM_L_X8Y143_SLICE_X10Y143_BQ),
.O5(CLBLM_R_X7Y143_SLICE_X9Y143_BO5),
.O6(CLBLM_R_X7Y143_SLICE_X9Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaff33aaaaf030)
  ) CLBLM_R_X7Y143_SLICE_X9Y143_ALUT (
.I0(CLBLM_L_X8Y142_SLICE_X10Y142_CQ),
.I1(CLBLM_R_X3Y147_SLICE_X3Y147_BQ),
.I2(CLBLM_R_X7Y143_SLICE_X9Y143_AQ),
.I3(CLBLM_R_X5Y144_SLICE_X6Y144_CQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X5Y141_SLICE_X7Y141_A5Q),
.O5(CLBLM_R_X7Y143_SLICE_X9Y143_AO5),
.O6(CLBLM_R_X7Y143_SLICE_X9Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y144_SLICE_X8Y144_A5_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y144_SLICE_X8Y144_AO5),
.Q(CLBLM_R_X7Y144_SLICE_X8Y144_A5Q),
.S(CLBLM_R_X11Y148_SLICE_X15Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y144_SLICE_X8Y144_A_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y144_SLICE_X8Y144_AO6),
.Q(CLBLM_R_X7Y144_SLICE_X8Y144_AQ),
.S(CLBLM_R_X11Y148_SLICE_X15Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y144_SLICE_X8Y144_B_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y142_SLICE_X10Y142_DO5),
.Q(CLBLM_R_X7Y144_SLICE_X8Y144_BQ),
.S(CLBLM_R_X11Y148_SLICE_X15Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000ff00ff00)
  ) CLBLM_R_X7Y144_SLICE_X8Y144_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X7Y143_SLICE_X9Y143_CQ),
.I4(1'b1),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X7Y144_SLICE_X8Y144_DO5),
.O6(CLBLM_R_X7Y144_SLICE_X8Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00aaf0fa00aaf0fa)
  ) CLBLM_R_X7Y144_SLICE_X8Y144_CLUT (
.I0(CLBLM_R_X7Y144_SLICE_X8Y144_BQ),
.I1(1'b1),
.I2(CLBLM_R_X7Y143_SLICE_X8Y143_DQ),
.I3(CLBLM_L_X8Y145_SLICE_X10Y145_CO5),
.I4(CLBLM_L_X8Y142_SLICE_X10Y142_BO5),
.I5(1'b1),
.O5(CLBLM_R_X7Y144_SLICE_X8Y144_CO5),
.O6(CLBLM_R_X7Y144_SLICE_X8Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fffffffffffffff)
  ) CLBLM_R_X7Y144_SLICE_X8Y144_BLUT (
.I0(CLBLM_R_X3Y152_SLICE_X3Y152_AQ),
.I1(CLBLM_R_X7Y152_SLICE_X8Y152_BQ),
.I2(CLBLM_R_X3Y144_SLICE_X3Y144_CQ),
.I3(CLBLL_L_X4Y151_SLICE_X5Y151_AQ),
.I4(CLBLM_R_X7Y144_SLICE_X9Y144_AQ),
.I5(CLBLM_R_X5Y144_SLICE_X7Y144_CQ),
.O5(CLBLM_R_X7Y144_SLICE_X8Y144_BO5),
.O6(CLBLM_R_X7Y144_SLICE_X8Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888cc00cc00)
  ) CLBLM_R_X7Y144_SLICE_X8Y144_ALUT (
.I0(CLBLM_R_X5Y150_SLICE_X6Y150_CQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(1'b1),
.I3(CLBLM_L_X8Y144_SLICE_X10Y144_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y144_SLICE_X8Y144_AO5),
.O6(CLBLM_R_X7Y144_SLICE_X8Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y144_SLICE_X9Y144_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y151_SLICE_X8Y151_DO6),
.Q(CLBLM_R_X7Y144_SLICE_X9Y144_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y144_SLICE_X9Y144_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y144_SLICE_X9Y144_BO5),
.Q(CLBLM_R_X7Y144_SLICE_X9Y144_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y144_SLICE_X9Y144_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y144_SLICE_X9Y144_CO5),
.Q(CLBLM_R_X7Y144_SLICE_X9Y144_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y144_SLICE_X9Y144_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y144_SLICE_X9Y144_DO5),
.Q(CLBLM_R_X7Y144_SLICE_X9Y144_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y144_SLICE_X9Y144_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y144_SLICE_X9Y144_AO6),
.Q(CLBLM_R_X7Y144_SLICE_X9Y144_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y144_SLICE_X9Y144_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y144_SLICE_X9Y144_BO6),
.Q(CLBLM_R_X7Y144_SLICE_X9Y144_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y144_SLICE_X9Y144_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y144_SLICE_X9Y144_CO6),
.Q(CLBLM_R_X7Y144_SLICE_X9Y144_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y144_SLICE_X9Y144_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y144_SLICE_X9Y144_DO6),
.Q(CLBLM_R_X7Y144_SLICE_X9Y144_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaa00aaf0ccf0cc)
  ) CLBLM_R_X7Y144_SLICE_X9Y144_DLUT (
.I0(CLBLM_R_X3Y150_SLICE_X3Y150_BQ),
.I1(CLBLM_R_X11Y147_SLICE_X15Y147_AQ),
.I2(CLBLM_R_X7Y146_SLICE_X9Y146_B5Q),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X8Y143_SLICE_X10Y143_DQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y144_SLICE_X9Y144_DO5),
.O6(CLBLM_R_X7Y144_SLICE_X9Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcf03fc30e2e2e2e2)
  ) CLBLM_R_X7Y144_SLICE_X9Y144_CLUT (
.I0(CLBLM_R_X7Y142_SLICE_X9Y142_D5Q),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_L_X10Y149_SLICE_X13Y149_AQ),
.I3(CLBLM_L_X10Y147_SLICE_X12Y147_CQ),
.I4(CLBLM_R_X7Y152_SLICE_X8Y152_BQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y144_SLICE_X9Y144_CO5),
.O6(CLBLM_R_X7Y144_SLICE_X9Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00aaaaccccf0f0)
  ) CLBLM_R_X7Y144_SLICE_X9Y144_BLUT (
.I0(CLBLM_L_X8Y143_SLICE_X11Y143_CQ),
.I1(CLBLM_R_X7Y144_SLICE_X9Y144_BQ),
.I2(RIOB33_X105Y127_IOB_X1Y128_I),
.I3(CLBLM_L_X8Y148_SLICE_X11Y148_B5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y144_SLICE_X9Y144_BO5),
.O6(CLBLM_R_X7Y144_SLICE_X9Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaacffccffc)
  ) CLBLM_R_X7Y144_SLICE_X9Y144_ALUT (
.I0(CLBLM_R_X7Y142_SLICE_X9Y142_DQ),
.I1(CLBLL_L_X2Y148_SLICE_X0Y148_B5Q),
.I2(CLBLM_R_X7Y144_SLICE_X9Y144_AQ),
.I3(CLBLM_R_X7Y152_SLICE_X8Y152_BQ),
.I4(1'b1),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X7Y144_SLICE_X9Y144_AO5),
.O6(CLBLM_R_X7Y144_SLICE_X9Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y145_SLICE_X8Y145_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y145_SLICE_X8Y145_BO5),
.Q(CLBLM_R_X7Y145_SLICE_X8Y145_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y145_SLICE_X8Y145_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y145_SLICE_X8Y145_CO5),
.Q(CLBLM_R_X7Y145_SLICE_X8Y145_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y145_SLICE_X8Y145_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y145_SLICE_X8Y145_AO6),
.Q(CLBLM_R_X7Y145_SLICE_X8Y145_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y145_SLICE_X8Y145_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y145_SLICE_X8Y145_BO6),
.Q(CLBLM_R_X7Y145_SLICE_X8Y145_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y145_SLICE_X8Y145_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y145_SLICE_X8Y145_CO6),
.Q(CLBLM_R_X7Y145_SLICE_X8Y145_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y145_SLICE_X8Y145_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y145_SLICE_X8Y145_DO6),
.Q(CLBLM_R_X7Y145_SLICE_X8Y145_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hbb88bb88b888b888)
  ) CLBLM_R_X7Y145_SLICE_X8Y145_DLUT (
.I0(CLBLM_R_X7Y143_SLICE_X8Y143_AQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X7Y145_SLICE_X8Y145_DQ),
.I3(CLBLM_L_X10Y143_SLICE_X12Y143_BO6),
.I4(1'b1),
.I5(CLBLM_R_X7Y151_SLICE_X8Y151_BQ),
.O5(CLBLM_R_X7Y145_SLICE_X8Y145_DO5),
.O6(CLBLM_R_X7Y145_SLICE_X8Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0aaaacccc00ff)
  ) CLBLM_R_X7Y145_SLICE_X8Y145_CLUT (
.I0(CLBLM_R_X7Y144_SLICE_X9Y144_D5Q),
.I1(CLBLM_R_X3Y143_SLICE_X2Y143_CQ),
.I2(CLBLM_R_X7Y145_SLICE_X8Y145_DQ),
.I3(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y145_SLICE_X8Y145_CO5),
.O6(CLBLM_R_X7Y145_SLICE_X8Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'he4e4e4e4ff55aa00)
  ) CLBLM_R_X7Y145_SLICE_X8Y145_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X7Y149_SLICE_X8Y149_AQ),
.I2(CLBLM_R_X3Y149_SLICE_X3Y149_CQ),
.I3(CLBLM_R_X7Y143_SLICE_X8Y143_CQ),
.I4(CLBLM_R_X5Y149_SLICE_X7Y149_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X7Y145_SLICE_X8Y145_BO5),
.O6(CLBLM_R_X7Y145_SLICE_X8Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaccc0aaaafff0)
  ) CLBLM_R_X7Y145_SLICE_X8Y145_ALUT (
.I0(CLBLM_R_X7Y145_SLICE_X8Y145_B5Q),
.I1(CLBLM_R_X5Y144_SLICE_X6Y144_CQ),
.I2(CLBLM_R_X7Y145_SLICE_X8Y145_AQ),
.I3(CLBLM_L_X8Y142_SLICE_X10Y142_CQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X3Y147_SLICE_X3Y147_BQ),
.O5(CLBLM_R_X7Y145_SLICE_X8Y145_AO5),
.O6(CLBLM_R_X7Y145_SLICE_X8Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y145_SLICE_X9Y145_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y145_SLICE_X9Y145_AO6),
.Q(CLBLM_R_X7Y145_SLICE_X9Y145_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y145_SLICE_X9Y145_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y145_SLICE_X9Y145_BO6),
.Q(CLBLM_R_X7Y145_SLICE_X9Y145_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y145_SLICE_X9Y145_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y145_SLICE_X9Y145_CO6),
.Q(CLBLM_R_X7Y145_SLICE_X9Y145_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y145_SLICE_X9Y145_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y145_SLICE_X9Y145_DO6),
.Q(CLBLM_R_X7Y145_SLICE_X9Y145_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hafafafafafafafac)
  ) CLBLM_R_X7Y145_SLICE_X9Y145_DLUT (
.I0(CLBLM_R_X5Y145_SLICE_X6Y145_AQ),
.I1(CLBLM_L_X10Y146_SLICE_X12Y146_BO6),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X7Y149_SLICE_X9Y149_CO6),
.I4(CLBLM_R_X7Y147_SLICE_X9Y147_DO6),
.I5(CLBLM_L_X8Y145_SLICE_X10Y145_BO6),
.O5(CLBLM_R_X7Y145_SLICE_X9Y145_DO5),
.O6(CLBLM_R_X7Y145_SLICE_X9Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0eef0fff044f000)
  ) CLBLM_R_X7Y145_SLICE_X9Y145_CLUT (
.I0(CLBLM_L_X8Y150_SLICE_X11Y150_B5Q),
.I1(CLBLM_R_X7Y145_SLICE_X9Y145_CQ),
.I2(CLBLM_R_X3Y146_SLICE_X3Y146_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X5Y149_SLICE_X6Y149_D5Q),
.I5(CLBLM_L_X8Y145_SLICE_X10Y145_AQ),
.O5(CLBLM_R_X7Y145_SLICE_X9Y145_CO5),
.O6(CLBLM_R_X7Y145_SLICE_X9Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0eeee00ee)
  ) CLBLM_R_X7Y145_SLICE_X9Y145_BLUT (
.I0(CLBLM_R_X7Y153_SLICE_X8Y153_AQ),
.I1(CLBLM_R_X7Y145_SLICE_X9Y145_BQ),
.I2(CLBLM_R_X7Y145_SLICE_X9Y145_AQ),
.I3(CLBLM_R_X5Y149_SLICE_X7Y149_DQ),
.I4(CLBLM_L_X8Y142_SLICE_X11Y142_CQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X7Y145_SLICE_X9Y145_BO5),
.O6(CLBLM_R_X7Y145_SLICE_X9Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00fafa5050)
  ) CLBLM_R_X7Y145_SLICE_X9Y145_ALUT (
.I0(CLBLM_L_X10Y143_SLICE_X12Y143_BO5),
.I1(1'b1),
.I2(CLBLM_R_X7Y145_SLICE_X9Y145_AQ),
.I3(CLBLM_R_X7Y145_SLICE_X9Y145_CQ),
.I4(CLBLM_R_X7Y145_SLICE_X8Y145_AQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X7Y145_SLICE_X9Y145_AO5),
.O6(CLBLM_R_X7Y145_SLICE_X9Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y146_SLICE_X8Y146_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_R_X3Y144_SLICE_X3Y144_CQ),
.Q(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y146_SLICE_X8Y146_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_L_X8Y144_SLICE_X10Y144_A5Q),
.Q(CLBLM_R_X7Y146_SLICE_X8Y146_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff75ff30ff75ff30)
  ) CLBLM_R_X7Y146_SLICE_X8Y146_DLUT (
.I0(CLBLM_L_X8Y145_SLICE_X10Y145_CO5),
.I1(CLBLM_L_X8Y142_SLICE_X10Y142_BO5),
.I2(CLBLM_R_X7Y149_SLICE_X8Y149_DQ),
.I3(CLBLM_R_X7Y146_SLICE_X8Y146_AO5),
.I4(CLBLM_R_X5Y147_SLICE_X7Y147_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X7Y146_SLICE_X8Y146_DO5),
.O6(CLBLM_R_X7Y146_SLICE_X8Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff0faf00aa)
  ) CLBLM_R_X7Y146_SLICE_X8Y146_CLUT (
.I0(CLBLM_R_X7Y147_SLICE_X8Y147_AQ),
.I1(1'b1),
.I2(CLBLM_L_X10Y143_SLICE_X12Y143_BO5),
.I3(CLBLM_L_X10Y143_SLICE_X12Y143_AO6),
.I4(CLBLM_R_X7Y147_SLICE_X8Y147_CQ),
.I5(CLBLM_L_X12Y149_SLICE_X16Y149_CO6),
.O5(CLBLM_R_X7Y146_SLICE_X8Y146_CO5),
.O6(CLBLM_R_X7Y146_SLICE_X8Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffffae)
  ) CLBLM_R_X7Y146_SLICE_X8Y146_BLUT (
.I0(CLBLM_R_X7Y146_SLICE_X8Y146_DO6),
.I1(CLBLM_R_X5Y147_SLICE_X7Y147_C5Q),
.I2(CLBLM_R_X5Y145_SLICE_X7Y145_BO6),
.I3(CLBLM_R_X7Y148_SLICE_X8Y148_BO6),
.I4(CLBLM_R_X7Y146_SLICE_X8Y146_CO6),
.I5(CLBLL_L_X4Y142_SLICE_X5Y142_DO6),
.O5(CLBLM_R_X7Y146_SLICE_X8Y146_BO5),
.O6(CLBLM_R_X7Y146_SLICE_X8Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55ffff00e40000)
  ) CLBLM_R_X7Y146_SLICE_X8Y146_ALUT (
.I0(CLBLM_R_X11Y149_SLICE_X14Y149_AQ),
.I1(CLBLM_R_X5Y147_SLICE_X7Y147_A5Q),
.I2(CLBLM_R_X5Y147_SLICE_X7Y147_BQ),
.I3(CLBLM_L_X8Y150_SLICE_X10Y150_A5Q),
.I4(CLBLM_L_X10Y143_SLICE_X13Y143_AO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y146_SLICE_X8Y146_AO5),
.O6(CLBLM_R_X7Y146_SLICE_X8Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y146_SLICE_X9Y146_B5_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y146_SLICE_X9Y146_BO5),
.Q(CLBLM_R_X7Y146_SLICE_X9Y146_B5Q),
.S(CLBLM_R_X11Y148_SLICE_X14Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y146_SLICE_X9Y146_B_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y146_SLICE_X9Y146_BO6),
.Q(CLBLM_R_X7Y146_SLICE_X9Y146_BQ),
.S(CLBLM_R_X11Y148_SLICE_X14Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7d7d7d7dbebebebe)
  ) CLBLM_R_X7Y146_SLICE_X9Y146_DLUT (
.I0(CLBLM_R_X5Y150_SLICE_X6Y150_DQ),
.I1(CLBLM_R_X5Y146_SLICE_X6Y146_AQ),
.I2(CLBLM_R_X3Y150_SLICE_X2Y150_DQ),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X8Y146_SLICE_X11Y146_AQ),
.O5(CLBLM_R_X7Y146_SLICE_X9Y146_DO5),
.O6(CLBLM_R_X7Y146_SLICE_X9Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00ccf0fc)
  ) CLBLM_R_X7Y146_SLICE_X9Y146_CLUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y146_SLICE_X4Y146_DQ),
.I2(CLBLL_L_X2Y143_SLICE_X1Y143_DQ),
.I3(CLBLM_L_X10Y143_SLICE_X12Y143_DO5),
.I4(CLBLM_L_X8Y142_SLICE_X10Y142_BO5),
.I5(CLBLM_L_X8Y147_SLICE_X10Y147_DO6),
.O5(CLBLM_R_X7Y146_SLICE_X9Y146_CO5),
.O6(CLBLM_R_X7Y146_SLICE_X9Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00000aaaa0000)
  ) CLBLM_R_X7Y146_SLICE_X9Y146_BLUT (
.I0(CLBLM_R_X7Y144_SLICE_X9Y144_DQ),
.I1(1'b1),
.I2(CLBLL_L_X2Y149_SLICE_X0Y149_AQ),
.I3(1'b1),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y146_SLICE_X9Y146_BO5),
.O6(CLBLM_R_X7Y146_SLICE_X9Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa003cffff3c)
  ) CLBLM_R_X7Y146_SLICE_X9Y146_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X3Y150_SLICE_X2Y150_DQ),
.I2(CLBLL_L_X4Y144_SLICE_X5Y144_DQ),
.I3(CLBLM_R_X5Y150_SLICE_X6Y150_DQ),
.I4(CLBLM_L_X8Y144_SLICE_X10Y144_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X7Y146_SLICE_X9Y146_AO5),
.O6(CLBLM_R_X7Y146_SLICE_X9Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y147_SLICE_X8Y147_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y147_SLICE_X8Y147_DO5),
.Q(CLBLM_R_X7Y147_SLICE_X8Y147_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y147_SLICE_X8Y147_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y147_SLICE_X8Y147_AO6),
.Q(CLBLM_R_X7Y147_SLICE_X8Y147_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y147_SLICE_X8Y147_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y147_SLICE_X8Y147_BO6),
.Q(CLBLM_R_X7Y147_SLICE_X8Y147_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y147_SLICE_X8Y147_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y147_SLICE_X8Y147_CO6),
.Q(CLBLM_R_X7Y147_SLICE_X8Y147_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y147_SLICE_X8Y147_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y147_SLICE_X8Y147_DO6),
.Q(CLBLM_R_X7Y147_SLICE_X8Y147_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8dd88dd8f5f5a0a0)
  ) CLBLM_R_X7Y147_SLICE_X8Y147_DLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X11Y151_SLICE_X15Y151_A5Q),
.I2(CLBLM_R_X5Y147_SLICE_X7Y147_B5Q),
.I3(CLBLM_R_X5Y144_SLICE_X7Y144_CQ),
.I4(CLBLM_L_X8Y148_SLICE_X11Y148_DQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y147_SLICE_X8Y147_DO5),
.O6(CLBLM_R_X7Y147_SLICE_X8Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ee44f0f0ff00)
  ) CLBLM_R_X7Y147_SLICE_X8Y147_CLUT (
.I0(CLBLM_R_X5Y144_SLICE_X6Y144_CQ),
.I1(CLBLM_R_X7Y147_SLICE_X8Y147_CQ),
.I2(CLBLM_R_X7Y141_SLICE_X8Y141_AQ),
.I3(CLBLL_L_X2Y148_SLICE_X1Y148_AQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X3Y147_SLICE_X3Y147_BQ),
.O5(CLBLM_R_X7Y147_SLICE_X8Y147_CO5),
.O6(CLBLM_R_X7Y147_SLICE_X8Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfaeefaee50445044)
  ) CLBLM_R_X7Y147_SLICE_X8Y147_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X7Y147_SLICE_X8Y147_BQ),
.I2(CLBLM_R_X5Y147_SLICE_X6Y147_DQ),
.I3(CLBLM_R_X11Y145_SLICE_X15Y145_BO5),
.I4(1'b1),
.I5(CLBLM_R_X3Y153_SLICE_X3Y153_A5Q),
.O5(CLBLM_R_X7Y147_SLICE_X8Y147_BO5),
.O6(CLBLM_R_X7Y147_SLICE_X8Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffd00fdff200020)
  ) CLBLM_R_X7Y147_SLICE_X8Y147_ALUT (
.I0(CLBLM_R_X5Y149_SLICE_X6Y149_D5Q),
.I1(CLBLM_L_X8Y150_SLICE_X11Y150_B5Q),
.I2(CLBLM_R_X7Y147_SLICE_X8Y147_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X7Y147_SLICE_X9Y147_AQ),
.I5(CLBLL_L_X2Y148_SLICE_X1Y148_A5Q),
.O5(CLBLM_R_X7Y147_SLICE_X8Y147_AO5),
.O6(CLBLM_R_X7Y147_SLICE_X8Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y147_SLICE_X9Y147_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y147_SLICE_X9Y147_CO5),
.Q(CLBLM_R_X7Y147_SLICE_X9Y147_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y147_SLICE_X9Y147_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y147_SLICE_X9Y147_AO6),
.Q(CLBLM_R_X7Y147_SLICE_X9Y147_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y147_SLICE_X9Y147_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y147_SLICE_X9Y147_BO6),
.Q(CLBLM_R_X7Y147_SLICE_X9Y147_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y147_SLICE_X9Y147_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y147_SLICE_X9Y147_CO6),
.Q(CLBLM_R_X7Y147_SLICE_X9Y147_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5ff5affa88888888)
  ) CLBLM_R_X7Y147_SLICE_X9Y147_DLUT (
.I0(CLBLM_R_X5Y148_SLICE_X6Y148_AQ),
.I1(CLBLM_L_X10Y142_SLICE_X12Y142_CO6),
.I2(CLBLL_L_X4Y147_SLICE_X5Y147_AQ),
.I3(CLBLM_R_X11Y147_SLICE_X14Y147_AQ),
.I4(CLBLM_R_X3Y146_SLICE_X3Y146_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y147_SLICE_X9Y147_DO5),
.O6(CLBLM_R_X7Y147_SLICE_X9Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff00f00cacacaca)
  ) CLBLM_R_X7Y147_SLICE_X9Y147_CLUT (
.I0(CLBLL_L_X4Y143_SLICE_X5Y143_DQ),
.I1(CLBLM_R_X7Y147_SLICE_X9Y147_CQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X5Y147_SLICE_X7Y147_CQ),
.I4(CLBLL_L_X4Y147_SLICE_X5Y147_CQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y147_SLICE_X9Y147_CO5),
.O6(CLBLM_R_X7Y147_SLICE_X9Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcffc0330cffc0330)
  ) CLBLM_R_X7Y147_SLICE_X9Y147_BLUT (
.I0(1'b1),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X7Y144_SLICE_X8Y144_BQ),
.I3(CLBLL_L_X4Y151_SLICE_X5Y151_AQ),
.I4(CLBLM_L_X10Y149_SLICE_X12Y149_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X7Y147_SLICE_X9Y147_BO5),
.O6(CLBLM_R_X7Y147_SLICE_X9Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff008d8dd8d8)
  ) CLBLM_R_X7Y147_SLICE_X9Y147_ALUT (
.I0(CLBLM_L_X8Y149_SLICE_X11Y149_BQ),
.I1(CLBLM_L_X10Y147_SLICE_X12Y147_BQ),
.I2(CLBLM_R_X7Y147_SLICE_X9Y147_AQ),
.I3(CLBLM_R_X7Y145_SLICE_X9Y145_BQ),
.I4(CLBLL_L_X4Y146_SLICE_X5Y146_DO6),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X7Y147_SLICE_X9Y147_AO5),
.O6(CLBLM_R_X7Y147_SLICE_X9Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y148_SLICE_X8Y148_A_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y148_SLICE_X8Y148_AO6),
.Q(CLBLM_R_X7Y148_SLICE_X8Y148_AQ),
.S(CLBLM_R_X11Y148_SLICE_X15Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000000a0000)
  ) CLBLM_R_X7Y148_SLICE_X8Y148_DLUT (
.I0(CLBLM_R_X3Y148_SLICE_X3Y148_CO5),
.I1(1'b1),
.I2(CLBLL_L_X4Y148_SLICE_X4Y148_BO5),
.I3(CLBLM_L_X10Y151_SLICE_X12Y151_BO6),
.I4(CLBLM_R_X7Y152_SLICE_X8Y152_DO6),
.I5(CLBLM_L_X10Y143_SLICE_X12Y143_AO5),
.O5(CLBLM_R_X7Y148_SLICE_X8Y148_DO5),
.O6(CLBLM_R_X7Y148_SLICE_X8Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7530550055005500)
  ) CLBLM_R_X7Y148_SLICE_X8Y148_CLUT (
.I0(CLBLM_R_X5Y145_SLICE_X7Y145_BO6),
.I1(CLBLM_L_X8Y150_SLICE_X10Y150_A5Q),
.I2(CLBLM_R_X11Y149_SLICE_X14Y149_AQ),
.I3(CLBLM_L_X8Y146_SLICE_X11Y146_A5Q),
.I4(CLBLM_L_X10Y144_SLICE_X13Y144_CO6),
.I5(CLBLM_R_X5Y149_SLICE_X7Y149_C5Q),
.O5(CLBLM_R_X7Y148_SLICE_X8Y148_CO5),
.O6(CLBLM_R_X7Y148_SLICE_X8Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00d00080afffafff)
  ) CLBLM_R_X7Y148_SLICE_X8Y148_BLUT (
.I0(CLBLM_R_X11Y149_SLICE_X14Y149_AQ),
.I1(CLBLM_R_X3Y147_SLICE_X2Y147_C5Q),
.I2(CLBLM_L_X10Y144_SLICE_X13Y144_CO6),
.I3(CLBLM_L_X8Y150_SLICE_X10Y150_A5Q),
.I4(CLBLM_R_X7Y148_SLICE_X9Y148_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y148_SLICE_X8Y148_BO5),
.O6(CLBLM_R_X7Y148_SLICE_X8Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0000000000)
  ) CLBLM_R_X7Y148_SLICE_X8Y148_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(1'b1),
.I5(CLBLL_L_X4Y148_SLICE_X5Y148_DQ),
.O5(CLBLM_R_X7Y148_SLICE_X8Y148_AO5),
.O6(CLBLM_R_X7Y148_SLICE_X8Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y148_SLICE_X9Y148_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y148_SLICE_X9Y148_BO5),
.Q(CLBLM_R_X7Y148_SLICE_X9Y148_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y148_SLICE_X9Y148_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y148_SLICE_X9Y148_CO5),
.Q(CLBLM_R_X7Y148_SLICE_X9Y148_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y148_SLICE_X9Y148_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y148_SLICE_X9Y148_AO6),
.Q(CLBLM_R_X7Y148_SLICE_X9Y148_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y148_SLICE_X9Y148_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y148_SLICE_X9Y148_BO6),
.Q(CLBLM_R_X7Y148_SLICE_X9Y148_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y148_SLICE_X9Y148_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y148_SLICE_X9Y148_CO6),
.Q(CLBLM_R_X7Y148_SLICE_X9Y148_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333333300000000)
  ) CLBLM_R_X7Y148_SLICE_X9Y148_DLUT (
.I0(1'b1),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLL_L_X4Y151_SLICE_X5Y151_AQ),
.O5(CLBLM_R_X7Y148_SLICE_X9Y148_DO5),
.O6(CLBLM_R_X7Y148_SLICE_X9Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaa00f0ccf0cc)
  ) CLBLM_R_X7Y148_SLICE_X9Y148_CLUT (
.I0(CLBLM_R_X7Y149_SLICE_X9Y149_BQ),
.I1(CLBLM_R_X3Y149_SLICE_X3Y149_DQ),
.I2(CLBLL_L_X2Y146_SLICE_X1Y146_A5Q),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X5Y150_SLICE_X7Y150_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y148_SLICE_X9Y148_CO5),
.O6(CLBLM_R_X7Y148_SLICE_X9Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f055aaccccf0f0)
  ) CLBLM_R_X7Y148_SLICE_X9Y148_BLUT (
.I0(CLBLM_L_X8Y147_SLICE_X11Y147_AQ),
.I1(CLBLM_R_X3Y148_SLICE_X2Y148_C5Q),
.I2(CLBLL_L_X4Y147_SLICE_X5Y147_AQ),
.I3(CLBLL_L_X4Y151_SLICE_X5Y151_AQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y148_SLICE_X9Y148_BO5),
.O6(CLBLM_R_X7Y148_SLICE_X9Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0050500000cccc)
  ) CLBLM_R_X7Y148_SLICE_X9Y148_ALUT (
.I0(CLBLM_L_X8Y146_SLICE_X10Y146_CQ),
.I1(CLBLM_L_X10Y147_SLICE_X13Y147_A5Q),
.I2(CLBLM_R_X7Y148_SLICE_X9Y148_AQ),
.I3(CLBLM_R_X5Y146_SLICE_X7Y146_BQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y148_SLICE_X9Y148_AO5),
.O6(CLBLM_R_X7Y148_SLICE_X9Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y149_SLICE_X8Y149_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y149_SLICE_X8Y149_AO6),
.Q(CLBLM_R_X7Y149_SLICE_X8Y149_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y149_SLICE_X8Y149_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y149_SLICE_X8Y149_BO6),
.Q(CLBLM_R_X7Y149_SLICE_X8Y149_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y149_SLICE_X8Y149_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y149_SLICE_X8Y149_CO6),
.Q(CLBLM_R_X7Y149_SLICE_X8Y149_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y149_SLICE_X8Y149_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y149_SLICE_X8Y149_DO6),
.Q(CLBLM_R_X7Y149_SLICE_X8Y149_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccaaf0aaf0)
  ) CLBLM_R_X7Y149_SLICE_X8Y149_DLUT (
.I0(CLBLM_R_X7Y143_SLICE_X8Y143_AQ),
.I1(CLBLM_R_X7Y149_SLICE_X8Y149_CQ),
.I2(CLBLM_R_X7Y149_SLICE_X8Y149_DQ),
.I3(CLBLM_L_X10Y143_SLICE_X12Y143_BO5),
.I4(1'b1),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X7Y149_SLICE_X8Y149_DO5),
.O6(CLBLM_R_X7Y149_SLICE_X8Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0066666666)
  ) CLBLM_R_X7Y149_SLICE_X8Y149_CLUT (
.I0(CLBLM_R_X5Y142_SLICE_X7Y142_BQ),
.I1(CLBLM_R_X3Y151_SLICE_X3Y151_BQ),
.I2(1'b1),
.I3(CLBLM_L_X12Y149_SLICE_X16Y149_BQ),
.I4(1'b1),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X7Y149_SLICE_X8Y149_CO5),
.O6(CLBLM_R_X7Y149_SLICE_X8Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0ffa0af505f000)
  ) CLBLM_R_X7Y149_SLICE_X8Y149_BLUT (
.I0(CLBLM_L_X10Y143_SLICE_X12Y143_AO6),
.I1(1'b1),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLL_L_X4Y151_SLICE_X5Y151_AQ),
.I4(CLBLM_R_X7Y149_SLICE_X8Y149_BQ),
.I5(CLBLM_R_X7Y150_SLICE_X9Y150_AQ),
.O5(CLBLM_R_X7Y149_SLICE_X8Y149_BO5),
.O6(CLBLM_R_X7Y149_SLICE_X8Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa00003cf0)
  ) CLBLM_R_X7Y149_SLICE_X8Y149_ALUT (
.I0(CLBLM_R_X7Y150_SLICE_X8Y150_DQ),
.I1(CLBLM_R_X7Y150_SLICE_X8Y150_CQ),
.I2(CLBLM_R_X7Y149_SLICE_X8Y149_AQ),
.I3(CLBLM_R_X7Y150_SLICE_X8Y150_AQ),
.I4(CLBLM_R_X3Y146_SLICE_X3Y146_CQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X7Y149_SLICE_X8Y149_AO5),
.O6(CLBLM_R_X7Y149_SLICE_X8Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y149_SLICE_X9Y149_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_L_X8Y149_SLICE_X10Y149_A5Q),
.Q(CLBLM_R_X7Y149_SLICE_X9Y149_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y149_SLICE_X9Y149_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_R_X5Y148_SLICE_X6Y148_AQ),
.Q(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y149_SLICE_X9Y149_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_R_X3Y152_SLICE_X2Y152_BQ),
.Q(CLBLM_R_X7Y149_SLICE_X9Y149_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y149_SLICE_X9Y149_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_R_X7Y149_SLICE_X9Y149_CO5),
.Q(CLBLM_R_X7Y149_SLICE_X9Y149_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y149_SLICE_X9Y149_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLL_L_X4Y149_SLICE_X4Y149_CQ),
.Q(CLBLM_R_X7Y149_SLICE_X9Y149_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfef0fafccee00aa)
  ) CLBLM_R_X7Y149_SLICE_X9Y149_DLUT (
.I0(CLBLM_R_X7Y152_SLICE_X8Y152_AQ),
.I1(CLBLM_L_X10Y142_SLICE_X12Y142_CO6),
.I2(CLBLM_R_X7Y148_SLICE_X8Y148_BO5),
.I3(CLBLM_L_X10Y143_SLICE_X12Y143_DO6),
.I4(CLBLM_L_X8Y149_SLICE_X10Y149_A5Q),
.I5(CLBLM_R_X7Y147_SLICE_X8Y147_D5Q),
.O5(CLBLM_R_X7Y149_SLICE_X9Y149_DO5),
.O6(CLBLM_R_X7Y149_SLICE_X9Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7bde7bdeffff0000)
  ) CLBLM_R_X7Y149_SLICE_X9Y149_CLUT (
.I0(CLBLM_R_X7Y149_SLICE_X8Y149_AQ),
.I1(CLBLM_R_X3Y147_SLICE_X3Y147_AQ),
.I2(CLBLM_L_X8Y149_SLICE_X10Y149_A5Q),
.I3(CLBLM_R_X7Y150_SLICE_X8Y150_DQ),
.I4(CLBLM_R_X7Y143_SLICE_X9Y143_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y149_SLICE_X9Y149_CO5),
.O6(CLBLM_R_X7Y149_SLICE_X9Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7733550030303030)
  ) CLBLM_R_X7Y149_SLICE_X9Y149_BLUT (
.I0(CLBLM_R_X7Y148_SLICE_X8Y148_BO5),
.I1(CLBLM_L_X10Y143_SLICE_X12Y143_DO6),
.I2(CLBLL_L_X4Y146_SLICE_X4Y146_AQ),
.I3(CLBLL_L_X2Y149_SLICE_X1Y149_A5Q),
.I4(CLBLM_R_X5Y152_SLICE_X7Y152_CQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y149_SLICE_X9Y149_BO5),
.O6(CLBLM_R_X7Y149_SLICE_X9Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00000000010001)
  ) CLBLM_R_X7Y149_SLICE_X9Y149_ALUT (
.I0(CLBLM_R_X7Y151_SLICE_X9Y151_CQ),
.I1(CLBLM_R_X7Y152_SLICE_X8Y152_BQ),
.I2(CLBLM_R_X7Y145_SLICE_X8Y145_AQ),
.I3(CLBLL_L_X2Y151_SLICE_X1Y151_BQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y149_SLICE_X9Y149_AO5),
.O6(CLBLM_R_X7Y149_SLICE_X9Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y150_SLICE_X8Y150_C5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y150_SLICE_X8Y150_CO5),
.Q(CLBLM_R_X7Y150_SLICE_X8Y150_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y150_SLICE_X8Y150_D5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y150_SLICE_X8Y150_DO5),
.Q(CLBLM_R_X7Y150_SLICE_X8Y150_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y150_SLICE_X8Y150_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y150_SLICE_X8Y150_AO6),
.Q(CLBLM_R_X7Y150_SLICE_X8Y150_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y150_SLICE_X8Y150_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y150_SLICE_X8Y150_BO6),
.Q(CLBLM_R_X7Y150_SLICE_X8Y150_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y150_SLICE_X8Y150_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y150_SLICE_X8Y150_CO6),
.Q(CLBLM_R_X7Y150_SLICE_X8Y150_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y150_SLICE_X8Y150_D_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y150_SLICE_X8Y150_DO6),
.Q(CLBLM_R_X7Y150_SLICE_X8Y150_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccf0f0ff00f0f0)
  ) CLBLM_R_X7Y150_SLICE_X8Y150_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y154_SLICE_X8Y154_BQ),
.I2(CLBLM_R_X3Y148_SLICE_X2Y148_C5Q),
.I3(CLBLM_R_X7Y150_SLICE_X8Y150_BQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y150_SLICE_X8Y150_DO5),
.O6(CLBLM_R_X7Y150_SLICE_X8Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff003333ccccf0f0)
  ) CLBLM_R_X7Y150_SLICE_X8Y150_CLUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y152_SLICE_X4Y152_C5Q),
.I2(CLBLM_L_X8Y145_SLICE_X11Y145_CO6),
.I3(CLBLL_L_X2Y149_SLICE_X1Y149_A5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y150_SLICE_X8Y150_CO5),
.O6(CLBLM_R_X7Y150_SLICE_X8Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0ff0cccc0ff0)
  ) CLBLM_R_X7Y150_SLICE_X8Y150_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y152_SLICE_X13Y152_AQ),
.I2(CLBLM_R_X3Y144_SLICE_X3Y144_CQ),
.I3(CLBLM_R_X5Y142_SLICE_X7Y142_B5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y150_SLICE_X8Y150_BO5),
.O6(CLBLM_R_X7Y150_SLICE_X8Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h888888888dd88dd8)
  ) CLBLM_R_X7Y150_SLICE_X8Y150_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X8Y147_SLICE_X11Y147_A5Q),
.I2(CLBLM_R_X7Y150_SLICE_X8Y150_AQ),
.I3(CLBLM_R_X7Y150_SLICE_X8Y150_CQ),
.I4(1'b1),
.I5(CLBLM_R_X3Y146_SLICE_X3Y146_CQ),
.O5(CLBLM_R_X7Y150_SLICE_X8Y150_AO5),
.O6(CLBLM_R_X7Y150_SLICE_X8Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y150_SLICE_X9Y150_B5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y150_SLICE_X9Y150_BO5),
.Q(CLBLM_R_X7Y150_SLICE_X9Y150_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y150_SLICE_X9Y150_C5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y150_SLICE_X9Y150_CO5),
.Q(CLBLM_R_X7Y150_SLICE_X9Y150_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y150_SLICE_X9Y150_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y150_SLICE_X9Y150_AO6),
.Q(CLBLM_R_X7Y150_SLICE_X9Y150_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y150_SLICE_X9Y150_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y150_SLICE_X9Y150_BO6),
.Q(CLBLM_R_X7Y150_SLICE_X9Y150_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y150_SLICE_X9Y150_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y150_SLICE_X9Y150_CO6),
.Q(CLBLM_R_X7Y150_SLICE_X9Y150_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y150_SLICE_X9Y150_D_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y150_SLICE_X9Y150_DO6),
.Q(CLBLM_R_X7Y150_SLICE_X9Y150_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ff00f0f0aaaa)
  ) CLBLM_R_X7Y150_SLICE_X9Y150_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y106_I),
.I1(1'b1),
.I2(CLBLM_R_X7Y149_SLICE_X8Y149_AQ),
.I3(CLBLM_R_X3Y152_SLICE_X3Y152_A5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X7Y149_SLICE_X9Y149_C5Q),
.O5(CLBLM_R_X7Y150_SLICE_X9Y150_DO5),
.O6(CLBLM_R_X7Y150_SLICE_X9Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'he4e4e4e4fafa5050)
  ) CLBLM_R_X7Y150_SLICE_X9Y150_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X8Y146_SLICE_X10Y146_AQ),
.I2(CLBLM_R_X7Y144_SLICE_X9Y144_B5Q),
.I3(1'b1),
.I4(CLBLM_L_X10Y147_SLICE_X12Y147_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y150_SLICE_X9Y150_CO5),
.O6(CLBLM_R_X7Y150_SLICE_X9Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc5050ff00cccc)
  ) CLBLM_R_X7Y150_SLICE_X9Y150_BLUT (
.I0(CLBLL_L_X4Y150_SLICE_X4Y150_AQ),
.I1(CLBLM_R_X7Y150_SLICE_X9Y150_DQ),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(CLBLL_L_X4Y151_SLICE_X5Y151_BQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y150_SLICE_X9Y150_BO5),
.O6(CLBLM_R_X7Y150_SLICE_X9Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccaaffcccca0f0)
  ) CLBLM_R_X7Y150_SLICE_X9Y150_ALUT (
.I0(CLBLM_L_X8Y150_SLICE_X11Y150_B5Q),
.I1(CLBLM_L_X8Y143_SLICE_X11Y143_CQ),
.I2(CLBLM_R_X7Y150_SLICE_X9Y150_AQ),
.I3(CLBLM_R_X5Y149_SLICE_X6Y149_D5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X5Y151_SLICE_X7Y151_AQ),
.O5(CLBLM_R_X7Y150_SLICE_X9Y150_AO5),
.O6(CLBLM_R_X7Y150_SLICE_X9Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y151_SLICE_X8Y151_C5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y151_SLICE_X8Y151_CO5),
.Q(CLBLM_R_X7Y151_SLICE_X8Y151_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y151_SLICE_X8Y151_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y151_SLICE_X8Y151_AO6),
.Q(CLBLM_R_X7Y151_SLICE_X8Y151_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y151_SLICE_X8Y151_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y151_SLICE_X8Y151_BO6),
.Q(CLBLM_R_X7Y151_SLICE_X8Y151_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y151_SLICE_X8Y151_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y151_SLICE_X8Y151_CO6),
.Q(CLBLM_R_X7Y151_SLICE_X8Y151_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff00f0000000101)
  ) CLBLM_R_X7Y151_SLICE_X8Y151_DLUT (
.I0(CLBLM_R_X7Y151_SLICE_X8Y151_C5Q),
.I1(CLBLM_R_X7Y151_SLICE_X8Y151_AQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X5Y152_SLICE_X6Y152_DQ),
.I4(CLBLM_R_X5Y152_SLICE_X7Y152_D5Q),
.I5(1'b1),
.O5(CLBLM_R_X7Y151_SLICE_X8Y151_DO5),
.O6(CLBLM_R_X7Y151_SLICE_X8Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfc303088bbbb88)
  ) CLBLM_R_X7Y151_SLICE_X8Y151_CLUT (
.I0(CLBLM_R_X5Y152_SLICE_X7Y152_BQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_L_X10Y150_SLICE_X13Y150_A5Q),
.I3(CLBLM_R_X3Y151_SLICE_X3Y151_AQ),
.I4(CLBLM_R_X5Y147_SLICE_X7Y147_BQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y151_SLICE_X8Y151_CO5),
.O6(CLBLM_R_X7Y151_SLICE_X8Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaafcfcaaaa00fc)
  ) CLBLM_R_X7Y151_SLICE_X8Y151_BLUT (
.I0(CLBLM_R_X5Y153_SLICE_X6Y153_AQ),
.I1(CLBLM_R_X7Y151_SLICE_X8Y151_BQ),
.I2(CLBLM_R_X5Y153_SLICE_X7Y153_AQ),
.I3(CLBLM_R_X3Y148_SLICE_X2Y148_D5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X5Y144_SLICE_X6Y144_DQ),
.O5(CLBLM_R_X7Y151_SLICE_X8Y151_BO5),
.O6(CLBLM_R_X7Y151_SLICE_X8Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa00ffaaaaff00)
  ) CLBLM_R_X7Y151_SLICE_X8Y151_ALUT (
.I0(CLBLM_R_X5Y143_SLICE_X6Y143_CQ),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_L_X8Y146_SLICE_X11Y146_A5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X7Y144_SLICE_X9Y144_AQ),
.O5(CLBLM_R_X7Y151_SLICE_X8Y151_AO5),
.O6(CLBLM_R_X7Y151_SLICE_X8Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y151_SLICE_X9Y151_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y151_SLICE_X9Y151_AO6),
.Q(CLBLM_R_X7Y151_SLICE_X9Y151_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y151_SLICE_X9Y151_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y151_SLICE_X9Y151_BO6),
.Q(CLBLM_R_X7Y151_SLICE_X9Y151_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y151_SLICE_X9Y151_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y151_SLICE_X9Y151_CO6),
.Q(CLBLM_R_X7Y151_SLICE_X9Y151_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y151_SLICE_X9Y151_D_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y151_SLICE_X9Y151_DO6),
.Q(CLBLM_R_X7Y151_SLICE_X9Y151_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff82a0000082a0)
  ) CLBLM_R_X7Y151_SLICE_X9Y151_DLUT (
.I0(CLBLM_R_X3Y152_SLICE_X2Y152_BQ),
.I1(CLBLM_L_X8Y152_SLICE_X11Y152_CO6),
.I2(CLBLM_R_X7Y151_SLICE_X9Y151_DQ),
.I3(CLBLM_L_X8Y151_SLICE_X10Y151_DQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X7Y147_SLICE_X8Y147_AQ),
.O5(CLBLM_R_X7Y151_SLICE_X9Y151_DO5),
.O6(CLBLM_R_X7Y151_SLICE_X9Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hddddd8d8ddddd8d8)
  ) CLBLM_R_X7Y151_SLICE_X9Y151_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X5Y142_SLICE_X7Y142_BQ),
.I2(CLBLM_L_X8Y151_SLICE_X10Y151_CO5),
.I3(1'b1),
.I4(CLBLM_R_X5Y151_SLICE_X7Y151_BO5),
.I5(1'b1),
.O5(CLBLM_R_X7Y151_SLICE_X9Y151_CO5),
.O6(CLBLM_R_X7Y151_SLICE_X9Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00000f0f40004)
  ) CLBLM_R_X7Y151_SLICE_X9Y151_BLUT (
.I0(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I1(CLBLM_R_X5Y149_SLICE_X7Y149_D5Q),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(RIOB33_X105Y101_IOB_X1Y102_I),
.I4(CLBLM_L_X8Y146_SLICE_X10Y146_AQ),
.I5(CLBLM_R_X5Y153_SLICE_X7Y153_CO6),
.O5(CLBLM_R_X7Y151_SLICE_X9Y151_BO5),
.O6(CLBLM_R_X7Y151_SLICE_X9Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a3a0a3a0a0a0a0)
  ) CLBLM_R_X7Y151_SLICE_X9Y151_ALUT (
.I0(CLBLM_R_X3Y148_SLICE_X2Y148_DQ),
.I1(CLBLM_R_X7Y146_SLICE_X8Y146_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X7Y153_SLICE_X8Y153_DO6),
.I4(1'b1),
.I5(CLBLM_L_X10Y150_SLICE_X12Y150_CQ),
.O5(CLBLM_R_X7Y151_SLICE_X9Y151_AO5),
.O6(CLBLM_R_X7Y151_SLICE_X9Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y152_SLICE_X8Y152_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y152_SLICE_X8Y152_AO6),
.Q(CLBLM_R_X7Y152_SLICE_X8Y152_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y152_SLICE_X8Y152_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y152_SLICE_X8Y152_BO6),
.Q(CLBLM_R_X7Y152_SLICE_X8Y152_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y152_SLICE_X8Y152_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y152_SLICE_X8Y152_CO6),
.Q(CLBLM_R_X7Y152_SLICE_X8Y152_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000800)
  ) CLBLM_R_X7Y152_SLICE_X8Y152_DLUT (
.I0(CLBLM_R_X7Y149_SLICE_X8Y149_BQ),
.I1(CLBLM_L_X8Y152_SLICE_X11Y152_AQ),
.I2(CLBLM_L_X8Y153_SLICE_X10Y153_CQ),
.I3(CLBLM_R_X7Y149_SLICE_X9Y149_AO5),
.I4(CLBLM_R_X7Y153_SLICE_X9Y153_BQ),
.I5(CLBLM_R_X7Y153_SLICE_X9Y153_AQ),
.O5(CLBLM_R_X7Y152_SLICE_X8Y152_DO5),
.O6(CLBLM_R_X7Y152_SLICE_X8Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'heb41aa00eb41aa00)
  ) CLBLM_R_X7Y152_SLICE_X8Y152_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X7Y152_SLICE_X8Y152_CQ),
.I2(CLBLM_R_X7Y154_SLICE_X8Y154_DO6),
.I3(CLBLM_R_X5Y152_SLICE_X6Y152_AQ),
.I4(CLBLM_R_X3Y152_SLICE_X2Y152_BQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y152_SLICE_X8Y152_CO5),
.O6(CLBLM_R_X7Y152_SLICE_X8Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ff33f0f0ff33)
  ) CLBLM_R_X7Y152_SLICE_X8Y152_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y152_SLICE_X8Y152_BQ),
.I2(CLBLM_R_X7Y151_SLICE_X8Y151_CQ),
.I3(CLBLL_L_X2Y148_SLICE_X0Y148_B5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y152_SLICE_X8Y152_BO5),
.O6(CLBLM_R_X7Y152_SLICE_X8Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff33fc30cc00fc30)
  ) CLBLM_R_X7Y152_SLICE_X8Y152_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X7Y152_SLICE_X8Y152_AQ),
.I3(CLBLM_L_X8Y152_SLICE_X10Y152_CQ),
.I4(CLBLM_L_X10Y143_SLICE_X12Y143_BO6),
.I5(CLBLM_L_X8Y146_SLICE_X10Y146_BQ),
.O5(CLBLM_R_X7Y152_SLICE_X8Y152_AO5),
.O6(CLBLM_R_X7Y152_SLICE_X8Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y152_SLICE_X9Y152_C5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y152_SLICE_X9Y152_CO5),
.Q(CLBLM_R_X7Y152_SLICE_X9Y152_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y152_SLICE_X9Y152_D5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y152_SLICE_X9Y152_DO5),
.Q(CLBLM_R_X7Y152_SLICE_X9Y152_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y152_SLICE_X9Y152_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y152_SLICE_X9Y152_AO6),
.Q(CLBLM_R_X7Y152_SLICE_X9Y152_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y152_SLICE_X9Y152_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y152_SLICE_X9Y152_BO6),
.Q(CLBLM_R_X7Y152_SLICE_X9Y152_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y152_SLICE_X9Y152_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y152_SLICE_X9Y152_CO6),
.Q(CLBLM_R_X7Y152_SLICE_X9Y152_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y152_SLICE_X9Y152_D_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y152_SLICE_X9Y152_DO6),
.Q(CLBLM_R_X7Y152_SLICE_X9Y152_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55aa008d8d8d8d)
  ) CLBLM_R_X7Y152_SLICE_X9Y152_DLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X8Y144_SLICE_X10Y144_B5Q),
.I2(CLBLM_R_X7Y145_SLICE_X8Y145_B5Q),
.I3(CLBLM_R_X5Y151_SLICE_X6Y151_CQ),
.I4(CLBLM_R_X7Y149_SLICE_X9Y149_CQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y152_SLICE_X9Y152_DO5),
.O6(CLBLM_R_X7Y152_SLICE_X9Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd88dd88e4e4e4e4)
  ) CLBLM_R_X7Y152_SLICE_X9Y152_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X7Y150_SLICE_X9Y150_BQ),
.I2(CLBLM_R_X5Y152_SLICE_X7Y152_AQ),
.I3(CLBLM_R_X5Y152_SLICE_X6Y152_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y152_SLICE_X9Y152_CO5),
.O6(CLBLM_R_X7Y152_SLICE_X9Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaf3fcfcfc)
  ) CLBLM_R_X7Y152_SLICE_X9Y152_BLUT (
.I0(CLBLM_L_X8Y142_SLICE_X10Y142_AQ),
.I1(CLBLM_R_X7Y152_SLICE_X9Y152_BQ),
.I2(CLBLM_R_X5Y152_SLICE_X6Y152_C5Q),
.I3(CLBLM_R_X7Y154_SLICE_X8Y154_BQ),
.I4(CLBLM_R_X7Y155_SLICE_X8Y155_AQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X7Y152_SLICE_X9Y152_BO5),
.O6(CLBLM_R_X7Y152_SLICE_X9Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hef23fe32ef23fe32)
  ) CLBLM_R_X7Y152_SLICE_X9Y152_ALUT (
.I0(CLBLM_R_X3Y148_SLICE_X2Y148_B5Q),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X7Y152_SLICE_X9Y152_AQ),
.I3(CLBLM_R_X3Y152_SLICE_X3Y152_AQ),
.I4(CLBLM_L_X10Y151_SLICE_X12Y151_AO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y152_SLICE_X9Y152_AO5),
.O6(CLBLM_R_X7Y152_SLICE_X9Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y153_SLICE_X8Y153_A_FDSE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y153_SLICE_X8Y153_AO6),
.Q(CLBLM_R_X7Y153_SLICE_X8Y153_AQ),
.S(CLBLM_R_X5Y153_SLICE_X7Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0ffffffbbbbffff)
  ) CLBLM_R_X7Y153_SLICE_X8Y153_DLUT (
.I0(CLBLM_R_X3Y150_SLICE_X2Y150_CO5),
.I1(CLBLM_R_X7Y153_SLICE_X9Y153_A5Q),
.I2(CLBLM_R_X7Y152_SLICE_X9Y152_DQ),
.I3(CLBLM_R_X7Y154_SLICE_X8Y154_AQ),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y153_SLICE_X8Y153_DO5),
.O6(CLBLM_R_X7Y153_SLICE_X8Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00aa00aaf300ff00)
  ) CLBLM_R_X7Y153_SLICE_X8Y153_CLUT (
.I0(CLBLM_R_X7Y149_SLICE_X9Y149_DQ),
.I1(CLBLM_R_X3Y151_SLICE_X3Y151_C5Q),
.I2(CLBLL_L_X4Y154_SLICE_X4Y154_AQ),
.I3(CLBLM_L_X10Y150_SLICE_X12Y150_CQ),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y153_SLICE_X8Y153_CO5),
.O6(CLBLM_R_X7Y153_SLICE_X8Y153_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0a000000c0cfc0cf)
  ) CLBLM_R_X7Y153_SLICE_X8Y153_BLUT (
.I0(CLBLM_R_X7Y152_SLICE_X9Y152_DQ),
.I1(CLBLM_R_X11Y149_SLICE_X15Y149_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_L_X10Y150_SLICE_X12Y150_CQ),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y153_SLICE_X8Y153_BO5),
.O6(CLBLM_R_X7Y153_SLICE_X8Y153_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0c0c0c0c0)
  ) CLBLM_R_X7Y153_SLICE_X8Y153_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y153_SLICE_X10Y153_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y153_SLICE_X8Y153_AO5),
.O6(CLBLM_R_X7Y153_SLICE_X8Y153_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y153_SLICE_X9Y153_A5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y153_SLICE_X11Y153_AO6),
.Q(CLBLM_R_X7Y153_SLICE_X9Y153_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y153_SLICE_X9Y153_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y153_SLICE_X9Y153_AO6),
.Q(CLBLM_R_X7Y153_SLICE_X9Y153_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y153_SLICE_X9Y153_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y153_SLICE_X9Y153_BO6),
.Q(CLBLM_R_X7Y153_SLICE_X9Y153_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y153_SLICE_X9Y153_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y153_SLICE_X9Y153_CO6),
.Q(CLBLM_R_X7Y153_SLICE_X9Y153_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'heeeeeeeeff0fff4f)
  ) CLBLM_R_X7Y153_SLICE_X9Y153_DLUT (
.I0(CLBLM_R_X7Y153_SLICE_X9Y153_BQ),
.I1(CLBLM_L_X8Y153_SLICE_X10Y153_CQ),
.I2(CLBLM_R_X7Y153_SLICE_X8Y153_DO6),
.I3(CLBLM_L_X10Y151_SLICE_X12Y151_CO6),
.I4(CLBLM_R_X7Y153_SLICE_X9Y153_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y153_SLICE_X9Y153_DO5),
.O6(CLBLM_R_X7Y153_SLICE_X9Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcfcacacacfcfca)
  ) CLBLM_R_X7Y153_SLICE_X9Y153_CLUT (
.I0(CLBLM_R_X5Y152_SLICE_X6Y152_C5Q),
.I1(CLBLM_L_X8Y149_SLICE_X10Y149_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X7Y155_SLICE_X9Y155_AO5),
.I4(CLBLM_R_X7Y153_SLICE_X9Y153_CQ),
.I5(CLBLM_R_X7Y152_SLICE_X9Y152_BQ),
.O5(CLBLM_R_X7Y153_SLICE_X9Y153_CO5),
.O6(CLBLM_R_X7Y153_SLICE_X9Y153_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf4f0f0f404000004)
  ) CLBLM_R_X7Y153_SLICE_X9Y153_BLUT (
.I0(CLBLM_R_X7Y152_SLICE_X9Y152_DQ),
.I1(CLBLM_R_X7Y154_SLICE_X9Y154_BO6),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_L_X8Y153_SLICE_X10Y153_CQ),
.I4(CLBLM_R_X7Y153_SLICE_X9Y153_BQ),
.I5(CLBLM_R_X5Y149_SLICE_X7Y149_DQ),
.O5(CLBLM_R_X7Y153_SLICE_X9Y153_BO5),
.O6(CLBLM_R_X7Y153_SLICE_X9Y153_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffeccccccceccc)
  ) CLBLM_R_X7Y153_SLICE_X9Y153_ALUT (
.I0(CLBLM_R_X7Y153_SLICE_X9Y153_DO6),
.I1(CLBLM_R_X7Y153_SLICE_X8Y153_BO6),
.I2(CLBLM_R_X7Y153_SLICE_X9Y153_AQ),
.I3(CLBLM_R_X7Y154_SLICE_X9Y154_BO6),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X3Y151_SLICE_X3Y151_DQ),
.O5(CLBLM_R_X7Y153_SLICE_X9Y153_AO5),
.O6(CLBLM_R_X7Y153_SLICE_X9Y153_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y154_SLICE_X8Y154_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y154_SLICE_X8Y154_AO6),
.Q(CLBLM_R_X7Y154_SLICE_X8Y154_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y154_SLICE_X8Y154_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y154_SLICE_X8Y154_BO6),
.Q(CLBLM_R_X7Y154_SLICE_X8Y154_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y154_SLICE_X8Y154_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y154_SLICE_X8Y154_CO6),
.Q(CLBLM_R_X7Y154_SLICE_X8Y154_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fffffff55ffffff)
  ) CLBLM_R_X7Y154_SLICE_X8Y154_DLUT (
.I0(CLBLM_L_X8Y153_SLICE_X11Y153_BQ),
.I1(CLBLM_R_X7Y154_SLICE_X8Y154_CQ),
.I2(CLBLM_L_X8Y154_SLICE_X10Y154_AQ),
.I3(CLBLM_R_X3Y154_SLICE_X3Y154_AQ),
.I4(CLBLM_R_X5Y154_SLICE_X7Y154_DQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y154_SLICE_X8Y154_DO5),
.O6(CLBLM_R_X7Y154_SLICE_X8Y154_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0099990000)
  ) CLBLM_R_X7Y154_SLICE_X8Y154_CLUT (
.I0(CLBLM_R_X7Y154_SLICE_X8Y154_DO5),
.I1(CLBLM_R_X7Y154_SLICE_X8Y154_CQ),
.I2(1'b1),
.I3(CLBLM_R_X7Y151_SLICE_X8Y151_AQ),
.I4(CLBLM_R_X3Y152_SLICE_X2Y152_BQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X7Y154_SLICE_X8Y154_CO5),
.O6(CLBLM_R_X7Y154_SLICE_X8Y154_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc0500050a)
  ) CLBLM_R_X7Y154_SLICE_X8Y154_BLUT (
.I0(CLBLM_R_X7Y154_SLICE_X8Y154_BQ),
.I1(CLBLL_L_X4Y149_SLICE_X4Y149_D5Q),
.I2(CLBLM_R_X5Y152_SLICE_X6Y152_C5Q),
.I3(CLBLM_R_X7Y155_SLICE_X8Y155_BQ),
.I4(CLBLM_R_X7Y155_SLICE_X8Y155_AQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X7Y154_SLICE_X8Y154_BO5),
.O6(CLBLM_R_X7Y154_SLICE_X8Y154_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffc400c4ffcc00cc)
  ) CLBLM_R_X7Y154_SLICE_X8Y154_ALUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(CLBLM_R_X7Y153_SLICE_X9Y153_DO5),
.I2(CLBLM_R_X3Y150_SLICE_X2Y150_CO5),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X3Y151_SLICE_X3Y151_BQ),
.I5(CLBLM_R_X3Y153_SLICE_X3Y153_A5Q),
.O5(CLBLM_R_X7Y154_SLICE_X8Y154_AO5),
.O6(CLBLM_R_X7Y154_SLICE_X8Y154_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y154_SLICE_X9Y154_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y154_SLICE_X9Y154_DO5),
.O6(CLBLM_R_X7Y154_SLICE_X9Y154_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff0020ffffffff)
  ) CLBLM_R_X7Y154_SLICE_X9Y154_CLUT (
.I0(CLBLM_R_X7Y154_SLICE_X8Y154_AQ),
.I1(CLBLM_R_X7Y152_SLICE_X9Y152_DQ),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(CLBLM_R_X7Y154_SLICE_X9Y154_AO5),
.I4(RIOB33_X105Y101_IOB_X1Y101_I),
.I5(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.O5(CLBLM_R_X7Y154_SLICE_X9Y154_CO5),
.O6(CLBLM_R_X7Y154_SLICE_X9Y154_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff550000fc540000)
  ) CLBLM_R_X7Y154_SLICE_X9Y154_BLUT (
.I0(CLBLM_R_X7Y153_SLICE_X8Y153_DO6),
.I1(CLBLM_L_X8Y153_SLICE_X10Y153_CQ),
.I2(CLBLM_R_X7Y153_SLICE_X9Y153_BQ),
.I3(CLBLM_L_X10Y150_SLICE_X12Y150_CQ),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(CLBLM_R_X7Y153_SLICE_X9Y153_AQ),
.O5(CLBLM_R_X7Y154_SLICE_X9Y154_BO5),
.O6(CLBLM_R_X7Y154_SLICE_X9Y154_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0c0c0000ff5dff55)
  ) CLBLM_R_X7Y154_SLICE_X9Y154_ALUT (
.I0(CLBLM_R_X7Y153_SLICE_X8Y153_DO5),
.I1(CLBLM_R_X3Y151_SLICE_X3Y151_C5Q),
.I2(CLBLL_L_X4Y154_SLICE_X4Y154_AQ),
.I3(CLBLM_R_X7Y151_SLICE_X9Y151_AQ),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y154_SLICE_X9Y154_AO5),
.O6(CLBLM_R_X7Y154_SLICE_X9Y154_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y155_SLICE_X8Y155_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y155_SLICE_X8Y155_AO6),
.Q(CLBLM_R_X7Y155_SLICE_X8Y155_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y155_SLICE_X8Y155_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y155_SLICE_X8Y155_BO6),
.Q(CLBLM_R_X7Y155_SLICE_X8Y155_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y155_SLICE_X8Y155_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y155_SLICE_X8Y155_DO5),
.O6(CLBLM_R_X7Y155_SLICE_X8Y155_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y155_SLICE_X8Y155_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y155_SLICE_X8Y155_CO5),
.O6(CLBLM_R_X7Y155_SLICE_X8Y155_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaaffaaf3aa33)
  ) CLBLM_R_X7Y155_SLICE_X8Y155_BLUT (
.I0(CLBLM_L_X8Y146_SLICE_X11Y146_A5Q),
.I1(CLBLM_R_X7Y155_SLICE_X8Y155_BQ),
.I2(CLBLM_R_X7Y155_SLICE_X8Y155_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X7Y154_SLICE_X8Y154_BQ),
.I5(CLBLM_R_X5Y152_SLICE_X6Y152_C5Q),
.O5(CLBLM_R_X7Y155_SLICE_X8Y155_BO5),
.O6(CLBLM_R_X7Y155_SLICE_X8Y155_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00ae04fa50)
  ) CLBLM_R_X7Y155_SLICE_X8Y155_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X7Y155_SLICE_X8Y155_BQ),
.I2(CLBLM_R_X7Y155_SLICE_X8Y155_AQ),
.I3(CLBLM_R_X5Y150_SLICE_X6Y150_AQ),
.I4(CLBLM_R_X7Y154_SLICE_X8Y154_BQ),
.I5(CLBLM_R_X5Y152_SLICE_X6Y152_C5Q),
.O5(CLBLM_R_X7Y155_SLICE_X8Y155_AO5),
.O6(CLBLM_R_X7Y155_SLICE_X8Y155_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y155_SLICE_X9Y155_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y155_SLICE_X9Y155_DO5),
.O6(CLBLM_R_X7Y155_SLICE_X9Y155_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y155_SLICE_X9Y155_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y155_SLICE_X9Y155_CO5),
.O6(CLBLM_R_X7Y155_SLICE_X9Y155_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y155_SLICE_X9Y155_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y155_SLICE_X9Y155_BO5),
.O6(CLBLM_R_X7Y155_SLICE_X9Y155_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000fffff0f00000)
  ) CLBLM_R_X7Y155_SLICE_X9Y155_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X7Y154_SLICE_X8Y154_BQ),
.I3(1'b1),
.I4(CLBLM_R_X7Y155_SLICE_X8Y155_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y155_SLICE_X9Y155_AO5),
.O6(CLBLM_R_X7Y155_SLICE_X9Y155_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y142_SLICE_X14Y142_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y142_SLICE_X14Y142_AO6),
.Q(CLBLM_R_X11Y142_SLICE_X14Y142_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000200000000000)
  ) CLBLM_R_X11Y142_SLICE_X14Y142_DLUT (
.I0(CLBLM_R_X5Y142_SLICE_X7Y142_C5Q),
.I1(CLBLM_R_X11Y146_SLICE_X14Y146_AQ),
.I2(CLBLM_L_X8Y144_SLICE_X11Y144_A5Q),
.I3(CLBLM_L_X8Y144_SLICE_X10Y144_B5Q),
.I4(CLBLM_R_X7Y146_SLICE_X9Y146_B5Q),
.I5(CLBLM_R_X7Y144_SLICE_X8Y144_AQ),
.O5(CLBLM_R_X11Y142_SLICE_X14Y142_DO5),
.O6(CLBLM_R_X11Y142_SLICE_X14Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0080008000800000)
  ) CLBLM_R_X11Y142_SLICE_X14Y142_CLUT (
.I0(CLBLM_R_X11Y149_SLICE_X14Y149_AQ),
.I1(CLBLM_L_X8Y144_SLICE_X11Y144_A5Q),
.I2(CLBLM_R_X7Y146_SLICE_X9Y146_B5Q),
.I3(CLBLM_L_X8Y150_SLICE_X10Y150_A5Q),
.I4(CLBLM_R_X11Y142_SLICE_X14Y142_BO5),
.I5(1'b1),
.O5(CLBLM_R_X11Y142_SLICE_X14Y142_CO5),
.O6(CLBLM_R_X11Y142_SLICE_X14Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000100000c00000)
  ) CLBLM_R_X11Y142_SLICE_X14Y142_BLUT (
.I0(CLBLM_L_X8Y144_SLICE_X11Y144_A5Q),
.I1(CLBLM_R_X7Y144_SLICE_X8Y144_AQ),
.I2(CLBLM_R_X5Y142_SLICE_X7Y142_C5Q),
.I3(CLBLM_R_X11Y146_SLICE_X14Y146_AQ),
.I4(CLBLM_L_X8Y144_SLICE_X10Y144_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X11Y142_SLICE_X14Y142_BO5),
.O6(CLBLM_R_X11Y142_SLICE_X14Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffd800d8ffd800d8)
  ) CLBLM_R_X11Y142_SLICE_X14Y142_ALUT (
.I0(CLBLM_R_X11Y145_SLICE_X15Y145_BO5),
.I1(CLBLM_L_X10Y147_SLICE_X13Y147_CQ),
.I2(CLBLM_R_X11Y142_SLICE_X14Y142_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X11Y146_SLICE_X15Y146_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y142_SLICE_X14Y142_AO5),
.O6(CLBLM_R_X11Y142_SLICE_X14Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y142_SLICE_X15Y142_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y142_SLICE_X15Y142_DO5),
.O6(CLBLM_R_X11Y142_SLICE_X15Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y142_SLICE_X15Y142_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y142_SLICE_X15Y142_CO5),
.O6(CLBLM_R_X11Y142_SLICE_X15Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y142_SLICE_X15Y142_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y142_SLICE_X15Y142_BO5),
.O6(CLBLM_R_X11Y142_SLICE_X15Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y142_SLICE_X15Y142_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y142_SLICE_X15Y142_AO5),
.O6(CLBLM_R_X11Y142_SLICE_X15Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y143_SLICE_X14Y143_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y143_SLICE_X14Y143_AO6),
.Q(CLBLM_R_X11Y143_SLICE_X14Y143_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf888f888f888f888)
  ) CLBLM_R_X11Y143_SLICE_X14Y143_DLUT (
.I0(CLBLM_R_X11Y148_SLICE_X14Y148_AQ),
.I1(RIOB33_X105Y139_IOB_X1Y140_I),
.I2(CLBLM_R_X11Y145_SLICE_X14Y145_AQ),
.I3(RIOB33_X105Y141_IOB_X1Y141_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y143_SLICE_X14Y143_DO5),
.O6(CLBLM_R_X11Y143_SLICE_X14Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0800000000000011)
  ) CLBLM_R_X11Y143_SLICE_X14Y143_CLUT (
.I0(CLBLM_R_X5Y142_SLICE_X7Y142_C5Q),
.I1(CLBLM_L_X8Y144_SLICE_X10Y144_B5Q),
.I2(CLBLM_R_X7Y146_SLICE_X9Y146_B5Q),
.I3(CLBLM_R_X7Y144_SLICE_X8Y144_AQ),
.I4(CLBLM_L_X8Y144_SLICE_X11Y144_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X11Y143_SLICE_X14Y143_CO5),
.O6(CLBLM_R_X11Y143_SLICE_X14Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h08000000f7fff7ff)
  ) CLBLM_R_X11Y143_SLICE_X14Y143_BLUT (
.I0(CLBLM_L_X8Y150_SLICE_X10Y150_A5Q),
.I1(CLBLM_R_X11Y143_SLICE_X14Y143_CO6),
.I2(CLBLM_R_X11Y149_SLICE_X14Y149_AQ),
.I3(CLBLM_R_X11Y146_SLICE_X14Y146_AQ),
.I4(CLBLM_R_X11Y149_SLICE_X15Y149_CQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y143_SLICE_X14Y143_BO5),
.O6(CLBLM_R_X11Y143_SLICE_X14Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffccfaccfaccfa)
  ) CLBLM_R_X11Y143_SLICE_X14Y143_ALUT (
.I0(CLBLM_R_X11Y143_SLICE_X14Y143_DO6),
.I1(CLBLM_R_X7Y144_SLICE_X9Y144_CQ),
.I2(CLBLM_L_X12Y144_SLICE_X16Y144_BO6),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(RIOB33_X105Y139_IOB_X1Y139_I),
.I5(CLBLM_L_X10Y143_SLICE_X12Y143_AQ),
.O5(CLBLM_R_X11Y143_SLICE_X14Y143_AO5),
.O6(CLBLM_R_X11Y143_SLICE_X14Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff88ff88ff888888)
  ) CLBLM_R_X11Y143_SLICE_X15Y143_DLUT (
.I0(CLBLM_R_X11Y142_SLICE_X14Y142_CO6),
.I1(CLBLM_R_X11Y142_SLICE_X14Y142_BO5),
.I2(1'b1),
.I3(CLBLM_L_X10Y148_SLICE_X13Y148_BO6),
.I4(CLBLM_R_X11Y143_SLICE_X14Y143_CO6),
.I5(CLBLM_R_X11Y142_SLICE_X14Y142_BO6),
.O5(CLBLM_R_X11Y143_SLICE_X15Y143_DO5),
.O6(CLBLM_R_X11Y143_SLICE_X15Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf888f00088880000)
  ) CLBLM_R_X11Y143_SLICE_X15Y143_CLUT (
.I0(CLBLM_R_X11Y142_SLICE_X14Y142_CO6),
.I1(CLBLM_R_X11Y142_SLICE_X14Y142_BO5),
.I2(CLBLM_R_X11Y142_SLICE_X14Y142_DO6),
.I3(CLBLM_L_X10Y148_SLICE_X13Y148_BO6),
.I4(LIOB33_SING_X0Y50_IOB_X0Y50_I),
.I5(RIOB33_X105Y135_IOB_X1Y136_I),
.O5(CLBLM_R_X11Y143_SLICE_X15Y143_CO5),
.O6(CLBLM_R_X11Y143_SLICE_X15Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'heaaac000c000c000)
  ) CLBLM_R_X11Y143_SLICE_X15Y143_BLUT (
.I0(CLBLM_R_X11Y142_SLICE_X14Y142_DO6),
.I1(CLBLM_R_X11Y142_SLICE_X14Y142_BO5),
.I2(RIOB33_X105Y133_IOB_X1Y134_I),
.I3(CLBLM_R_X11Y142_SLICE_X14Y142_CO6),
.I4(CLBLM_R_X11Y148_SLICE_X14Y148_AQ),
.I5(CLBLM_L_X8Y144_SLICE_X10Y144_CO6),
.O5(CLBLM_R_X11Y143_SLICE_X15Y143_BO5),
.O6(CLBLM_R_X11Y143_SLICE_X15Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffefffeeffcfffcc)
  ) CLBLM_R_X11Y143_SLICE_X15Y143_ALUT (
.I0(CLBLM_L_X10Y142_SLICE_X13Y142_AQ),
.I1(CLBLM_R_X11Y143_SLICE_X14Y143_BO6),
.I2(CLBLM_L_X12Y145_SLICE_X16Y145_AO6),
.I3(CLBLM_R_X11Y143_SLICE_X15Y143_BO6),
.I4(RIOB33_X105Y139_IOB_X1Y140_I),
.I5(CLBLM_R_X11Y145_SLICE_X15Y145_BO5),
.O5(CLBLM_R_X11Y143_SLICE_X15Y143_AO5),
.O6(CLBLM_R_X11Y143_SLICE_X15Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y144_SLICE_X14Y144_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_R_X11Y142_SLICE_X14Y142_AQ),
.Q(CLBLM_R_X11Y144_SLICE_X14Y144_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haa000c0000000000)
  ) CLBLM_R_X11Y144_SLICE_X14Y144_DLUT (
.I0(CLBLM_R_X3Y145_SLICE_X2Y145_BQ),
.I1(CLBLM_R_X7Y150_SLICE_X8Y150_C5Q),
.I2(CLBLM_R_X7Y146_SLICE_X9Y146_B5Q),
.I3(CLBLM_L_X8Y150_SLICE_X10Y150_A5Q),
.I4(CLBLM_R_X11Y149_SLICE_X14Y149_AQ),
.I5(CLBLM_R_X11Y142_SLICE_X14Y142_BO6),
.O5(CLBLM_R_X11Y144_SLICE_X14Y144_DO5),
.O6(CLBLM_R_X11Y144_SLICE_X14Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0100000000000000)
  ) CLBLM_R_X11Y144_SLICE_X14Y144_CLUT (
.I0(CLBLM_R_X11Y142_SLICE_X14Y142_CO5),
.I1(CLBLM_R_X11Y144_SLICE_X15Y144_AO5),
.I2(CLBLM_R_X11Y145_SLICE_X15Y145_BO5),
.I3(CLBLM_R_X11Y143_SLICE_X14Y143_BO5),
.I4(CLBLM_L_X12Y145_SLICE_X16Y145_AO6),
.I5(CLBLM_R_X11Y144_SLICE_X15Y144_CO6),
.O5(CLBLM_R_X11Y144_SLICE_X14Y144_CO5),
.O6(CLBLM_R_X11Y144_SLICE_X14Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0c0f0c0f0f0f0e)
  ) CLBLM_R_X11Y144_SLICE_X14Y144_BLUT (
.I0(CLBLM_L_X12Y144_SLICE_X16Y144_DO6),
.I1(CLBLM_L_X10Y145_SLICE_X13Y145_BO6),
.I2(CLBLM_R_X11Y143_SLICE_X14Y143_CO5),
.I3(CLBLM_R_X11Y145_SLICE_X14Y145_BO6),
.I4(CLBLM_R_X11Y144_SLICE_X14Y144_AO6),
.I5(CLBLM_L_X10Y142_SLICE_X13Y142_BO6),
.O5(CLBLM_R_X11Y144_SLICE_X14Y144_BO5),
.O6(CLBLM_R_X11Y144_SLICE_X14Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffdfcfdfcfdfc)
  ) CLBLM_R_X11Y144_SLICE_X14Y144_ALUT (
.I0(CLBLM_L_X12Y145_SLICE_X16Y145_AO6),
.I1(CLBLM_L_X10Y143_SLICE_X13Y143_BO6),
.I2(CLBLM_R_X11Y144_SLICE_X15Y144_AO6),
.I3(RIOB33_X105Y139_IOB_X1Y139_I),
.I4(CLBLM_L_X10Y147_SLICE_X13Y147_DQ),
.I5(CLBLM_R_X11Y145_SLICE_X15Y145_BO5),
.O5(CLBLM_R_X11Y144_SLICE_X14Y144_AO5),
.O6(CLBLM_R_X11Y144_SLICE_X14Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hdddddddfcccccccf)
  ) CLBLM_R_X11Y144_SLICE_X15Y144_DLUT (
.I0(CLBLM_R_X11Y144_SLICE_X15Y144_CO6),
.I1(CLBLM_R_X11Y143_SLICE_X15Y143_CO6),
.I2(CLBLM_R_X11Y143_SLICE_X15Y143_DO6),
.I3(CLBLM_R_X11Y144_SLICE_X15Y144_AO5),
.I4(CLBLM_R_X11Y145_SLICE_X15Y145_BO5),
.I5(CLBLM_R_X11Y142_SLICE_X14Y142_AQ),
.O5(CLBLM_R_X11Y144_SLICE_X15Y144_DO5),
.O6(CLBLM_R_X11Y144_SLICE_X15Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffdffffffffffff)
  ) CLBLM_R_X11Y144_SLICE_X15Y144_CLUT (
.I0(CLBLM_R_X11Y146_SLICE_X14Y146_AQ),
.I1(CLBLM_R_X7Y144_SLICE_X8Y144_AQ),
.I2(CLBLM_L_X8Y144_SLICE_X11Y144_A5Q),
.I3(CLBLM_L_X8Y144_SLICE_X10Y144_B5Q),
.I4(CLBLM_R_X5Y142_SLICE_X7Y142_C5Q),
.I5(CLBLM_L_X10Y148_SLICE_X13Y148_BO6),
.O5(CLBLM_R_X11Y144_SLICE_X15Y144_CO5),
.O6(CLBLM_R_X11Y144_SLICE_X15Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ffff0000afae)
  ) CLBLM_R_X11Y144_SLICE_X15Y144_BLUT (
.I0(CLBLM_L_X10Y144_SLICE_X12Y144_BO6),
.I1(CLBLM_R_X11Y143_SLICE_X15Y143_AO6),
.I2(CLBLM_L_X10Y142_SLICE_X13Y142_BO6),
.I3(CLBLM_L_X12Y144_SLICE_X16Y144_CO6),
.I4(CLBLM_R_X11Y143_SLICE_X14Y143_CO5),
.I5(CLBLM_R_X11Y145_SLICE_X15Y145_CO6),
.O5(CLBLM_R_X11Y144_SLICE_X15Y144_BO5),
.O6(CLBLM_R_X11Y144_SLICE_X15Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h2000000010d010d0)
  ) CLBLM_R_X11Y144_SLICE_X15Y144_ALUT (
.I0(CLBLM_L_X8Y150_SLICE_X10Y150_A5Q),
.I1(CLBLM_R_X11Y149_SLICE_X14Y149_AQ),
.I2(CLBLM_R_X11Y143_SLICE_X14Y143_CO6),
.I3(CLBLM_R_X11Y146_SLICE_X14Y146_AQ),
.I4(CLBLM_R_X11Y149_SLICE_X15Y149_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y144_SLICE_X15Y144_AO5),
.O6(CLBLM_R_X11Y144_SLICE_X15Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y145_SLICE_X14Y145_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_R_X3Y145_SLICE_X2Y145_AQ),
.Q(CLBLM_R_X11Y145_SLICE_X14Y145_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y145_SLICE_X14Y145_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_R_X7Y147_SLICE_X9Y147_BQ),
.Q(CLBLM_R_X11Y145_SLICE_X14Y145_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y145_SLICE_X14Y145_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_R_X11Y147_SLICE_X14Y147_A5Q),
.Q(CLBLM_R_X11Y145_SLICE_X14Y145_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y145_SLICE_X14Y145_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_R_X11Y145_SLICE_X14Y145_CQ),
.Q(CLBLM_R_X11Y145_SLICE_X14Y145_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbaabbaa33003300)
  ) CLBLM_R_X11Y145_SLICE_X14Y145_DLUT (
.I0(CLBLM_R_X11Y142_SLICE_X14Y142_CO5),
.I1(CLBLM_L_X12Y145_SLICE_X16Y145_AO6),
.I2(1'b1),
.I3(RIOB33_X105Y141_IOB_X1Y141_I),
.I4(1'b1),
.I5(RIOB33_X105Y147_IOB_X1Y147_I),
.O5(CLBLM_R_X11Y145_SLICE_X14Y145_DO5),
.O6(CLBLM_R_X11Y145_SLICE_X14Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5544f5f45544f5f4)
  ) CLBLM_R_X11Y145_SLICE_X14Y145_CLUT (
.I0(CLBLM_L_X10Y142_SLICE_X13Y142_BO6),
.I1(CLBLM_R_X11Y145_SLICE_X15Y145_AO5),
.I2(CLBLM_R_X11Y147_SLICE_X14Y147_AQ),
.I3(CLBLM_L_X12Y145_SLICE_X16Y145_DO6),
.I4(CLBLM_R_X11Y145_SLICE_X14Y145_BO5),
.I5(1'b1),
.O5(CLBLM_R_X11Y145_SLICE_X14Y145_CO5),
.O6(CLBLM_R_X11Y145_SLICE_X14Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h20200000eeeeffff)
  ) CLBLM_R_X11Y145_SLICE_X14Y145_BLUT (
.I0(CLBLM_R_X11Y149_SLICE_X14Y149_AQ),
.I1(CLBLM_L_X12Y143_SLICE_X16Y143_AO6),
.I2(CLBLM_R_X7Y149_SLICE_X9Y149_C5Q),
.I3(1'b1),
.I4(CLBLM_L_X8Y150_SLICE_X10Y150_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X11Y145_SLICE_X14Y145_BO5),
.O6(CLBLM_R_X11Y145_SLICE_X14Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000ababaaaa)
  ) CLBLM_R_X11Y145_SLICE_X14Y145_ALUT (
.I0(CLBLM_R_X11Y144_SLICE_X14Y144_DO6),
.I1(CLBLM_L_X10Y142_SLICE_X13Y142_BO6),
.I2(CLBLM_R_X11Y146_SLICE_X15Y146_CO5),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X11Y145_SLICE_X15Y145_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y145_SLICE_X14Y145_AO5),
.O6(CLBLM_R_X11Y145_SLICE_X14Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y145_SLICE_X15Y145_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_L_X10Y146_SLICE_X13Y146_AQ),
.Q(CLBLM_R_X11Y145_SLICE_X15Y145_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00ff44ff44)
  ) CLBLM_R_X11Y145_SLICE_X15Y145_DLUT (
.I0(CLBLM_R_X11Y146_SLICE_X15Y146_CO5),
.I1(CLBLM_R_X11Y144_SLICE_X14Y144_AQ),
.I2(1'b1),
.I3(CLBLM_L_X12Y145_SLICE_X16Y145_CO6),
.I4(1'b1),
.I5(CLBLM_L_X10Y142_SLICE_X13Y142_BO6),
.O5(CLBLM_R_X11Y145_SLICE_X15Y145_DO5),
.O6(CLBLM_R_X11Y145_SLICE_X15Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h400040004000ffff)
  ) CLBLM_R_X11Y145_SLICE_X15Y145_CLUT (
.I0(CLBLM_L_X12Y143_SLICE_X16Y143_AO6),
.I1(CLBLL_L_X4Y145_SLICE_X5Y145_BQ),
.I2(CLBLM_R_X11Y149_SLICE_X14Y149_AQ),
.I3(CLBLM_L_X8Y150_SLICE_X10Y150_A5Q),
.I4(CLBLM_L_X8Y152_SLICE_X11Y152_A5Q),
.I5(CLBLM_R_X11Y145_SLICE_X15Y145_BO6),
.O5(CLBLM_R_X11Y145_SLICE_X15Y145_CO5),
.O6(CLBLM_R_X11Y145_SLICE_X15Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffafff01000000)
  ) CLBLM_R_X11Y145_SLICE_X15Y145_BLUT (
.I0(CLBLM_R_X11Y149_SLICE_X14Y149_AQ),
.I1(CLBLM_L_X12Y149_SLICE_X16Y149_CO6),
.I2(CLBLM_L_X8Y150_SLICE_X10Y150_A5Q),
.I3(CLBLM_R_X11Y142_SLICE_X14Y142_BO6),
.I4(CLBLM_R_X7Y146_SLICE_X9Y146_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X11Y145_SLICE_X15Y145_BO5),
.O6(CLBLM_R_X11Y145_SLICE_X15Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00aeae0c0c)
  ) CLBLM_R_X11Y145_SLICE_X15Y145_ALUT (
.I0(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.I1(CLBLM_L_X10Y145_SLICE_X12Y145_AQ),
.I2(CLBLM_R_X11Y146_SLICE_X15Y146_CO5),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X11Y142_SLICE_X14Y142_CO5),
.I5(1'b1),
.O5(CLBLM_R_X11Y145_SLICE_X15Y145_AO5),
.O6(CLBLM_R_X11Y145_SLICE_X15Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y146_SLICE_X14Y146_A_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y145_SLICE_X14Y145_AO6),
.Q(CLBLM_R_X11Y146_SLICE_X14Y146_AQ),
.S(CLBLM_R_X11Y148_SLICE_X15Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h33223322f3f2f3f2)
  ) CLBLM_R_X11Y146_SLICE_X14Y146_DLUT (
.I0(CLBLM_L_X12Y145_SLICE_X17Y145_CO6),
.I1(CLBLM_L_X10Y142_SLICE_X13Y142_BO6),
.I2(CLBLM_R_X7Y150_SLICE_X8Y150_DQ),
.I3(CLBLM_L_X12Y146_SLICE_X16Y146_BO6),
.I4(1'b1),
.I5(CLBLM_R_X11Y145_SLICE_X14Y145_BO5),
.O5(CLBLM_R_X11Y146_SLICE_X14Y146_DO5),
.O6(CLBLM_R_X11Y146_SLICE_X14Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdfdfdfdfdfdfdfc)
  ) CLBLM_R_X11Y146_SLICE_X14Y146_CLUT (
.I0(CLBLM_L_X10Y142_SLICE_X13Y142_BO6),
.I1(CLBLM_L_X8Y148_SLICE_X10Y148_BO5),
.I2(CLBLM_R_X11Y147_SLICE_X15Y147_BO6),
.I3(CLBLM_L_X12Y145_SLICE_X16Y145_AO5),
.I4(CLBLM_L_X10Y146_SLICE_X12Y146_CO5),
.I5(CLBLM_R_X11Y144_SLICE_X14Y144_CO6),
.O5(CLBLM_R_X11Y146_SLICE_X14Y146_CO5),
.O6(CLBLM_R_X11Y146_SLICE_X14Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffeeffffffeefe)
  ) CLBLM_R_X11Y146_SLICE_X14Y146_BLUT (
.I0(CLBLM_R_X11Y147_SLICE_X14Y147_DO6),
.I1(CLBLM_R_X5Y145_SLICE_X7Y145_CO6),
.I2(CLBLM_R_X11Y146_SLICE_X14Y146_DO6),
.I3(CLBLM_R_X11Y143_SLICE_X14Y143_CO5),
.I4(CLBLM_L_X8Y145_SLICE_X10Y145_DO6),
.I5(CLBLM_R_X11Y146_SLICE_X14Y146_CO6),
.O5(CLBLM_R_X11Y146_SLICE_X14Y146_BO5),
.O6(CLBLM_R_X11Y146_SLICE_X14Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ff000000cccc)
  ) CLBLM_R_X11Y146_SLICE_X14Y146_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y144_SLICE_X10Y144_A5Q),
.I2(1'b1),
.I3(CLBLM_L_X8Y147_SLICE_X11Y147_A5Q),
.I4(CLBLM_L_X10Y145_SLICE_X12Y145_AO6),
.I5(1'b1),
.O5(CLBLM_R_X11Y146_SLICE_X14Y146_AO5),
.O6(CLBLM_R_X11Y146_SLICE_X14Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y146_SLICE_X15Y146_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y146_SLICE_X15Y146_AO6),
.Q(CLBLM_R_X11Y146_SLICE_X15Y146_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0fffff0f0fbfa)
  ) CLBLM_R_X11Y146_SLICE_X15Y146_DLUT (
.I0(CLBLM_R_X11Y146_SLICE_X14Y146_AO6),
.I1(CLBLM_L_X10Y142_SLICE_X13Y142_BO6),
.I2(CLBLM_L_X10Y146_SLICE_X12Y146_BO5),
.I3(CLBLM_R_X11Y144_SLICE_X15Y144_DO6),
.I4(CLBLM_R_X11Y143_SLICE_X14Y143_CO5),
.I5(CLBLM_R_X11Y145_SLICE_X15Y145_DO6),
.O5(CLBLM_R_X11Y146_SLICE_X15Y146_DO5),
.O6(CLBLM_R_X11Y146_SLICE_X15Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00e2000033ffffff)
  ) CLBLM_R_X11Y146_SLICE_X15Y146_CLUT (
.I0(RIOB33_X105Y145_IOB_X1Y145_I),
.I1(CLBLM_R_X11Y149_SLICE_X14Y149_AQ),
.I2(CLBLM_R_X11Y148_SLICE_X14Y148_CQ),
.I3(CLBLM_L_X8Y150_SLICE_X10Y150_A5Q),
.I4(CLBLM_R_X11Y142_SLICE_X14Y142_DO6),
.I5(1'b1),
.O5(CLBLM_R_X11Y146_SLICE_X15Y146_CO5),
.O6(CLBLM_R_X11Y146_SLICE_X15Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0eeccaa00)
  ) CLBLM_R_X11Y146_SLICE_X15Y146_BLUT (
.I0(CLBLM_R_X11Y148_SLICE_X14Y148_CQ),
.I1(CLBLM_R_X11Y145_SLICE_X14Y145_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(RIOB33_X105Y145_IOB_X1Y145_I),
.I4(CLBLM_R_X5Y151_SLICE_X6Y151_BQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y146_SLICE_X15Y146_BO5),
.O6(CLBLM_R_X11Y146_SLICE_X15Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff8d008dffd800d8)
  ) CLBLM_R_X11Y146_SLICE_X15Y146_ALUT (
.I0(CLBLM_L_X8Y149_SLICE_X11Y149_BQ),
.I1(CLBLM_L_X8Y151_SLICE_X10Y151_BQ),
.I2(CLBLM_R_X11Y146_SLICE_X15Y146_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X12Y149_SLICE_X16Y149_AQ),
.I5(CLBLM_R_X5Y146_SLICE_X7Y146_AQ),
.O5(CLBLM_R_X11Y146_SLICE_X15Y146_AO5),
.O6(CLBLM_R_X11Y146_SLICE_X15Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y147_SLICE_X14Y147_A5_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y147_SLICE_X14Y147_AO5),
.Q(CLBLM_R_X11Y147_SLICE_X14Y147_A5Q),
.S(CLBLM_R_X11Y148_SLICE_X15Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y147_SLICE_X14Y147_A_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y147_SLICE_X14Y147_AO6),
.Q(CLBLM_R_X11Y147_SLICE_X14Y147_AQ),
.S(CLBLM_R_X11Y148_SLICE_X15Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00aa00aa00aa00aa)
  ) CLBLM_R_X11Y147_SLICE_X14Y147_DLUT (
.I0(CLBLM_R_X5Y145_SLICE_X7Y145_AQ),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_L_X10Y144_SLICE_X12Y144_AO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y147_SLICE_X14Y147_DO5),
.O6(CLBLM_R_X11Y147_SLICE_X14Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffff00fffe)
  ) CLBLM_R_X11Y147_SLICE_X14Y147_CLUT (
.I0(CLBLM_L_X10Y147_SLICE_X12Y147_DO5),
.I1(CLBLM_R_X11Y144_SLICE_X14Y144_CO6),
.I2(CLBLM_R_X11Y145_SLICE_X14Y145_DO6),
.I3(CLBLM_R_X11Y146_SLICE_X14Y146_AO5),
.I4(CLBLM_L_X10Y142_SLICE_X13Y142_BO6),
.I5(CLBLM_L_X10Y145_SLICE_X13Y145_AO5),
.O5(CLBLM_R_X11Y147_SLICE_X14Y147_CO5),
.O6(CLBLM_R_X11Y147_SLICE_X14Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffeeffffffeefe)
  ) CLBLM_R_X11Y147_SLICE_X14Y147_BLUT (
.I0(CLBLM_L_X8Y144_SLICE_X11Y144_DO6),
.I1(CLBLM_R_X7Y146_SLICE_X9Y146_CO6),
.I2(CLBLM_R_X11Y147_SLICE_X15Y147_CO6),
.I3(CLBLM_R_X11Y143_SLICE_X14Y143_CO5),
.I4(CLBLM_R_X7Y149_SLICE_X9Y149_BO5),
.I5(CLBLM_R_X11Y147_SLICE_X14Y147_CO6),
.O5(CLBLM_R_X11Y147_SLICE_X14Y147_BO5),
.O6(CLBLM_R_X11Y147_SLICE_X14Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000cccc0000)
  ) CLBLM_R_X11Y147_SLICE_X14Y147_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y142_SLICE_X9Y142_CQ),
.I2(1'b1),
.I3(CLBLM_L_X10Y149_SLICE_X12Y149_CQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y147_SLICE_X14Y147_AO5),
.O6(CLBLM_R_X11Y147_SLICE_X14Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y147_SLICE_X15Y147_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y147_SLICE_X15Y147_AO6),
.Q(CLBLM_R_X11Y147_SLICE_X15Y147_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0c0c0c0c0c0c0c0c)
  ) CLBLM_R_X11Y147_SLICE_X15Y147_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y147_SLICE_X14Y147_A5Q),
.I2(CLBLM_L_X10Y145_SLICE_X12Y145_AO6),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y147_SLICE_X15Y147_DO5),
.O6(CLBLM_R_X11Y147_SLICE_X15Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0537050500330000)
  ) CLBLM_R_X11Y147_SLICE_X15Y147_CLUT (
.I0(CLBLM_R_X11Y146_SLICE_X15Y146_CO5),
.I1(CLBLM_R_X7Y146_SLICE_X9Y146_B5Q),
.I2(CLBLM_L_X10Y142_SLICE_X13Y142_BO6),
.I3(CLBLM_R_X11Y144_SLICE_X15Y144_CO6),
.I4(CLBLM_L_X10Y147_SLICE_X13Y147_A5Q),
.I5(CLBLM_R_X11Y145_SLICE_X14Y145_AQ),
.O5(CLBLM_R_X11Y147_SLICE_X15Y147_CO5),
.O6(CLBLM_R_X11Y147_SLICE_X15Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha000a00030000000)
  ) CLBLM_R_X11Y147_SLICE_X15Y147_BLUT (
.I0(CLBLL_L_X4Y147_SLICE_X5Y147_BQ),
.I1(CLBLM_R_X7Y146_SLICE_X9Y146_B5Q),
.I2(CLBLM_R_X11Y142_SLICE_X14Y142_BO6),
.I3(CLBLM_L_X8Y150_SLICE_X10Y150_A5Q),
.I4(CLBLM_R_X3Y148_SLICE_X2Y148_C5Q),
.I5(CLBLM_R_X11Y149_SLICE_X14Y149_AQ),
.O5(CLBLM_R_X11Y147_SLICE_X15Y147_BO5),
.O6(CLBLM_R_X11Y147_SLICE_X15Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa3faa30aa3faa30)
  ) CLBLM_R_X11Y147_SLICE_X15Y147_ALUT (
.I0(CLBLM_L_X10Y148_SLICE_X13Y148_AQ),
.I1(CLBLL_L_X4Y152_SLICE_X5Y152_B5Q),
.I2(CLBLM_R_X11Y147_SLICE_X15Y147_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y147_SLICE_X15Y147_AO5),
.O6(CLBLM_R_X11Y147_SLICE_X15Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y148_SLICE_X14Y148_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.Q(CLBLM_R_X11Y148_SLICE_X14Y148_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y148_SLICE_X14Y148_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLL_L_X4Y152_SLICE_X4Y152_BQ),
.Q(CLBLM_R_X11Y148_SLICE_X14Y148_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y148_SLICE_X14Y148_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_R_X11Y148_SLICE_X14Y148_BQ),
.Q(CLBLM_R_X11Y148_SLICE_X14Y148_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y148_SLICE_X14Y148_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_R_X7Y151_SLICE_X8Y151_C5Q),
.Q(CLBLM_R_X11Y148_SLICE_X14Y148_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0505050505050505)
  ) CLBLM_R_X11Y148_SLICE_X14Y148_DLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(1'b1),
.I2(CLBLM_L_X10Y150_SLICE_X13Y150_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y148_SLICE_X14Y148_DO5),
.O6(CLBLM_R_X11Y148_SLICE_X14Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000055555555)
  ) CLBLM_R_X11Y148_SLICE_X14Y148_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X10Y150_SLICE_X13Y150_A5Q),
.O5(CLBLM_R_X11Y148_SLICE_X14Y148_CO5),
.O6(CLBLM_R_X11Y148_SLICE_X14Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6699669999669966)
  ) CLBLM_R_X11Y148_SLICE_X14Y148_BLUT (
.I0(CLBLM_L_X8Y152_SLICE_X11Y152_A5Q),
.I1(CLBLM_R_X3Y148_SLICE_X2Y148_C5Q),
.I2(1'b1),
.I3(CLBLM_L_X10Y150_SLICE_X13Y150_A5Q),
.I4(1'b1),
.I5(CLBLM_L_X10Y150_SLICE_X13Y150_AQ),
.O5(CLBLM_R_X11Y148_SLICE_X14Y148_BO5),
.O6(CLBLM_R_X11Y148_SLICE_X14Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc33c3cc33cc3c33c)
  ) CLBLM_R_X11Y148_SLICE_X14Y148_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y150_SLICE_X8Y150_C5Q),
.I2(CLBLM_L_X10Y147_SLICE_X13Y147_AQ),
.I3(CLBLM_R_X11Y148_SLICE_X14Y148_BO6),
.I4(CLBLM_L_X10Y147_SLICE_X13Y147_A5Q),
.I5(CLBLM_L_X8Y152_SLICE_X11Y152_AQ),
.O5(CLBLM_R_X11Y148_SLICE_X14Y148_AO5),
.O6(CLBLM_R_X11Y148_SLICE_X14Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y148_SLICE_X15Y148_A_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y146_SLICE_X15Y146_BO6),
.Q(CLBLM_R_X11Y148_SLICE_X15Y148_AQ),
.S(CLBLM_R_X11Y150_SLICE_X14Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y148_SLICE_X15Y148_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y148_SLICE_X15Y148_DO5),
.O6(CLBLM_R_X11Y148_SLICE_X15Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0505050505050505)
  ) CLBLM_R_X11Y148_SLICE_X15Y148_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(1'b1),
.I2(CLBLM_L_X8Y152_SLICE_X11Y152_A5Q),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y148_SLICE_X15Y148_CO5),
.O6(CLBLM_R_X11Y148_SLICE_X15Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000333300003333)
  ) CLBLM_R_X11Y148_SLICE_X15Y148_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y152_SLICE_X11Y152_AQ),
.I2(1'b1),
.I3(1'b1),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y148_SLICE_X15Y148_BO5),
.O6(CLBLM_R_X11Y148_SLICE_X15Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00f000f000f000f0)
  ) CLBLM_R_X11Y148_SLICE_X15Y148_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_L_X10Y147_SLICE_X13Y147_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y148_SLICE_X15Y148_AO5),
.O6(CLBLM_R_X11Y148_SLICE_X15Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y149_SLICE_X14Y149_A_FDSE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y149_SLICE_X13Y149_BO6),
.Q(CLBLM_R_X11Y149_SLICE_X14Y149_AQ),
.S(CLBLM_R_X11Y148_SLICE_X14Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y149_SLICE_X14Y149_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y149_SLICE_X14Y149_DO5),
.O6(CLBLM_R_X11Y149_SLICE_X14Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3bfbfb3b37f7f737)
  ) CLBLM_R_X11Y149_SLICE_X14Y149_CLUT (
.I0(CLBLM_R_X11Y148_SLICE_X14Y148_AO6),
.I1(CLBLM_R_X3Y151_SLICE_X3Y151_D5Q),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(CLBLM_R_X11Y149_SLICE_X14Y149_AO5),
.I4(CLBLM_R_X11Y149_SLICE_X14Y149_BO5),
.I5(CLBLM_R_X11Y149_SLICE_X15Y149_BQ),
.O5(CLBLM_R_X11Y149_SLICE_X14Y149_CO5),
.O6(CLBLM_R_X11Y149_SLICE_X14Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0f0f99666699)
  ) CLBLM_R_X11Y149_SLICE_X14Y149_BLUT (
.I0(CLBLM_L_X10Y145_SLICE_X13Y145_CO6),
.I1(CLBLM_R_X11Y147_SLICE_X14Y147_BO6),
.I2(CLBLM_R_X3Y151_SLICE_X3Y151_D5Q),
.I3(CLBLM_L_X8Y145_SLICE_X11Y145_CO6),
.I4(CLBLM_L_X8Y147_SLICE_X11Y147_BO6),
.I5(1'b1),
.O5(CLBLM_R_X11Y149_SLICE_X14Y149_BO5),
.O6(CLBLM_R_X11Y149_SLICE_X14Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hafafafaf66999966)
  ) CLBLM_R_X11Y149_SLICE_X14Y149_ALUT (
.I0(CLBLM_L_X10Y149_SLICE_X13Y149_CO6),
.I1(CLBLM_R_X11Y146_SLICE_X14Y146_BO6),
.I2(CLBLM_R_X3Y151_SLICE_X3Y151_D5Q),
.I3(CLBLM_L_X10Y148_SLICE_X13Y148_CO6),
.I4(CLBLM_L_X10Y145_SLICE_X12Y145_BO6),
.I5(1'b1),
.O5(CLBLM_R_X11Y149_SLICE_X14Y149_AO5),
.O6(CLBLM_R_X11Y149_SLICE_X14Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y149_SLICE_X15Y149_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y149_SLICE_X15Y149_AO6),
.Q(CLBLM_R_X11Y149_SLICE_X15Y149_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y149_SLICE_X15Y149_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y149_SLICE_X15Y149_BO6),
.Q(CLBLM_R_X11Y149_SLICE_X15Y149_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y149_SLICE_X15Y149_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y149_SLICE_X15Y149_CO6),
.Q(CLBLM_R_X11Y149_SLICE_X15Y149_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000ff00000001)
  ) CLBLM_R_X11Y149_SLICE_X15Y149_DLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(RIOB33_X105Y131_IOB_X1Y132_I),
.I2(RIOB33_X105Y133_IOB_X1Y133_I),
.I3(RIOB33_X105Y129_IOB_X1Y129_I),
.I4(RIOB33_X105Y129_IOB_X1Y130_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y149_SLICE_X15Y149_DO5),
.O6(CLBLM_R_X11Y149_SLICE_X15Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hef45ee44ee44ee44)
  ) CLBLM_R_X11Y149_SLICE_X15Y149_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X11Y149_SLICE_X15Y149_CQ),
.I2(RIOB33_X105Y133_IOB_X1Y133_I),
.I3(CLBLM_R_X11Y145_SLICE_X14Y145_AQ),
.I4(CLBLM_R_X11Y149_SLICE_X15Y149_DO6),
.I5(CLBLM_L_X12Y149_SLICE_X16Y149_AQ),
.O5(CLBLM_R_X11Y149_SLICE_X15Y149_CO5),
.O6(CLBLM_R_X11Y149_SLICE_X15Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffcc5accffcc00)
  ) CLBLM_R_X11Y149_SLICE_X15Y149_BLUT (
.I0(CLBLM_R_X11Y149_SLICE_X14Y149_AO5),
.I1(CLBLM_R_X3Y146_SLICE_X2Y146_BQ),
.I2(CLBLM_R_X11Y149_SLICE_X14Y149_BO5),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X12Y149_SLICE_X16Y149_DO6),
.I5(RIOB33_X105Y131_IOB_X1Y132_I),
.O5(CLBLM_R_X11Y149_SLICE_X15Y149_BO5),
.O6(CLBLM_R_X11Y149_SLICE_X15Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffccdeccffcccccc)
  ) CLBLM_R_X11Y149_SLICE_X15Y149_ALUT (
.I0(CLBLM_R_X11Y149_SLICE_X14Y149_AO5),
.I1(CLBLM_L_X10Y149_SLICE_X13Y149_BO5),
.I2(CLBLM_R_X11Y149_SLICE_X14Y149_BO5),
.I3(CLBLM_R_X11Y149_SLICE_X15Y149_DO5),
.I4(CLBLM_L_X12Y149_SLICE_X16Y149_DO6),
.I5(RIOB33_X105Y131_IOB_X1Y132_I),
.O5(CLBLM_R_X11Y149_SLICE_X15Y149_AO5),
.O6(CLBLM_R_X11Y149_SLICE_X15Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y150_SLICE_X14Y150_A_FDSE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y150_SLICE_X14Y150_AO6),
.Q(CLBLM_R_X11Y150_SLICE_X14Y150_AQ),
.S(CLBLM_R_X11Y150_SLICE_X14Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000ff00ff00)
  ) CLBLM_R_X11Y150_SLICE_X14Y150_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X5Y153_SLICE_X6Y153_AQ),
.I4(1'b1),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X11Y150_SLICE_X14Y150_DO5),
.O6(CLBLM_R_X11Y150_SLICE_X14Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hdffddffdeffeeffe)
  ) CLBLM_R_X11Y150_SLICE_X14Y150_CLUT (
.I0(CLBLM_R_X7Y152_SLICE_X8Y152_CQ),
.I1(CLBLM_L_X10Y150_SLICE_X13Y150_DO5),
.I2(CLBLM_L_X8Y147_SLICE_X11Y147_A5Q),
.I3(CLBLM_R_X7Y151_SLICE_X9Y151_DQ),
.I4(1'b1),
.I5(CLBLM_R_X11Y147_SLICE_X14Y147_A5Q),
.O5(CLBLM_R_X11Y150_SLICE_X14Y150_CO5),
.O6(CLBLM_R_X11Y150_SLICE_X14Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fff0ffccffccff)
  ) CLBLM_R_X11Y150_SLICE_X14Y150_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y147_SLICE_X14Y147_BO6),
.I2(CLBLM_L_X8Y145_SLICE_X11Y145_CO6),
.I3(CLBLM_R_X3Y151_SLICE_X3Y151_D5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y150_SLICE_X14Y150_BO5),
.O6(CLBLM_R_X11Y150_SLICE_X14Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa00000000)
  ) CLBLM_R_X11Y150_SLICE_X14Y150_ALUT (
.I0(CLBLM_R_X11Y145_SLICE_X14Y145_DQ),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X11Y150_SLICE_X14Y150_AO5),
.O6(CLBLM_R_X11Y150_SLICE_X14Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y150_SLICE_X15Y150_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y150_SLICE_X15Y150_AO6),
.Q(CLBLM_R_X11Y150_SLICE_X15Y150_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y150_SLICE_X15Y150_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y150_SLICE_X15Y150_DO5),
.O6(CLBLM_R_X11Y150_SLICE_X15Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y150_SLICE_X15Y150_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y150_SLICE_X15Y150_CO5),
.O6(CLBLM_R_X11Y150_SLICE_X15Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y150_SLICE_X15Y150_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y150_SLICE_X15Y150_BO5),
.O6(CLBLM_R_X11Y150_SLICE_X15Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000ff5a005a)
  ) CLBLM_R_X11Y150_SLICE_X15Y150_ALUT (
.I0(CLBLM_L_X8Y146_SLICE_X10Y146_A5Q),
.I1(1'b1),
.I2(CLBLM_R_X11Y150_SLICE_X15Y150_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X11Y148_SLICE_X14Y148_AQ),
.I5(CLBLM_R_X3Y148_SLICE_X2Y148_B5Q),
.O5(CLBLM_R_X11Y150_SLICE_X15Y150_AO5),
.O6(CLBLM_R_X11Y150_SLICE_X15Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y151_SLICE_X14Y151_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y151_SLICE_X14Y151_AO6),
.Q(CLBLM_R_X11Y151_SLICE_X14Y151_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y151_SLICE_X14Y151_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y151_SLICE_X14Y151_BO6),
.Q(CLBLM_R_X11Y151_SLICE_X14Y151_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0ffffffffffffff)
  ) CLBLM_R_X11Y151_SLICE_X14Y151_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_L_X10Y153_SLICE_X12Y153_DO6),
.I3(CLBLM_R_X11Y151_SLICE_X14Y151_AQ),
.I4(CLBLM_R_X11Y152_SLICE_X14Y152_A5Q),
.I5(CLBLM_L_X10Y152_SLICE_X12Y152_AQ),
.O5(CLBLM_R_X11Y151_SLICE_X14Y151_DO5),
.O6(CLBLM_R_X11Y151_SLICE_X14Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffefffefe)
  ) CLBLM_R_X11Y151_SLICE_X14Y151_CLUT (
.I0(CLBLM_L_X10Y149_SLICE_X12Y149_AQ),
.I1(CLBLM_R_X11Y151_SLICE_X15Y151_A5Q),
.I2(CLBLM_L_X10Y150_SLICE_X13Y150_C5Q),
.I3(CLBLM_L_X10Y151_SLICE_X13Y151_CO6),
.I4(CLBLM_R_X11Y151_SLICE_X15Y151_BQ),
.I5(CLBLM_L_X10Y149_SLICE_X12Y149_BQ),
.O5(CLBLM_R_X11Y151_SLICE_X14Y151_CO5),
.O6(CLBLM_R_X11Y151_SLICE_X14Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffeebb0000eebb)
  ) CLBLM_R_X11Y151_SLICE_X14Y151_BLUT (
.I0(CLBLM_R_X3Y148_SLICE_X2Y148_B5Q),
.I1(CLBLM_R_X11Y151_SLICE_X14Y151_BQ),
.I2(1'b1),
.I3(CLBLM_L_X10Y151_SLICE_X13Y151_BO5),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_L_X10Y147_SLICE_X13Y147_B5Q),
.O5(CLBLM_R_X11Y151_SLICE_X14Y151_BO5),
.O6(CLBLM_R_X11Y151_SLICE_X14Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccca5f00000)
  ) CLBLM_R_X11Y151_SLICE_X14Y151_ALUT (
.I0(CLBLM_L_X10Y153_SLICE_X12Y153_DO6),
.I1(CLBLM_L_X8Y149_SLICE_X11Y149_B5Q),
.I2(CLBLM_R_X11Y151_SLICE_X14Y151_AQ),
.I3(CLBLM_L_X10Y151_SLICE_X12Y151_DO6),
.I4(CLBLM_L_X10Y152_SLICE_X13Y152_CO5),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X11Y151_SLICE_X14Y151_AO5),
.O6(CLBLM_R_X11Y151_SLICE_X14Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y151_SLICE_X15Y151_A5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y151_SLICE_X15Y151_CO5),
.Q(CLBLM_R_X11Y151_SLICE_X15Y151_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y151_SLICE_X15Y151_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y151_SLICE_X15Y151_AO6),
.Q(CLBLM_R_X11Y151_SLICE_X15Y151_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y151_SLICE_X15Y151_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y151_SLICE_X15Y151_BO6),
.Q(CLBLM_R_X11Y151_SLICE_X15Y151_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y151_SLICE_X15Y151_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y151_SLICE_X15Y151_DO5),
.O6(CLBLM_R_X11Y151_SLICE_X15Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccffffaa30aa30)
  ) CLBLM_R_X11Y151_SLICE_X15Y151_CLUT (
.I0(CLBLM_L_X12Y151_SLICE_X16Y151_AQ),
.I1(CLBLM_L_X10Y151_SLICE_X13Y151_CO6),
.I2(CLBLM_R_X11Y151_SLICE_X15Y151_BQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X8Y146_SLICE_X10Y146_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X11Y151_SLICE_X15Y151_CO5),
.O6(CLBLM_R_X11Y151_SLICE_X15Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff441400004414)
  ) CLBLM_R_X11Y151_SLICE_X15Y151_BLUT (
.I0(CLBLM_R_X3Y148_SLICE_X2Y148_B5Q),
.I1(CLBLM_R_X11Y151_SLICE_X15Y151_BQ),
.I2(CLBLM_L_X8Y146_SLICE_X10Y146_A5Q),
.I3(CLBLM_L_X10Y151_SLICE_X13Y151_CO6),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X11Y148_SLICE_X14Y148_CQ),
.O5(CLBLM_R_X11Y151_SLICE_X15Y151_BO5),
.O6(CLBLM_R_X11Y151_SLICE_X15Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff33fe32ff33ee22)
  ) CLBLM_R_X11Y151_SLICE_X15Y151_ALUT (
.I0(CLBLM_R_X3Y148_SLICE_X2Y148_B5Q),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X11Y151_SLICE_X15Y151_AQ),
.I3(CLBLM_R_X5Y151_SLICE_X6Y151_BQ),
.I4(CLBLM_L_X10Y151_SLICE_X13Y151_DO6),
.I5(CLBLM_R_X11Y151_SLICE_X15Y151_CO6),
.O5(CLBLM_R_X11Y151_SLICE_X15Y151_AO5),
.O6(CLBLM_R_X11Y151_SLICE_X15Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y152_SLICE_X14Y152_A5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y152_SLICE_X14Y152_AO5),
.Q(CLBLM_R_X11Y152_SLICE_X14Y152_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y152_SLICE_X14Y152_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y152_SLICE_X14Y152_AO6),
.Q(CLBLM_R_X11Y152_SLICE_X14Y152_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff7fffffffffff)
  ) CLBLM_R_X11Y152_SLICE_X14Y152_DLUT (
.I0(CLBLM_L_X12Y151_SLICE_X16Y151_AQ),
.I1(CLBLM_L_X10Y152_SLICE_X12Y152_BQ),
.I2(CLBLM_R_X11Y152_SLICE_X14Y152_AQ),
.I3(CLBLM_L_X10Y152_SLICE_X13Y152_AQ),
.I4(CLBLM_R_X11Y151_SLICE_X14Y151_DO6),
.I5(CLBLM_L_X12Y151_SLICE_X16Y151_BQ),
.O5(CLBLM_R_X11Y152_SLICE_X14Y152_DO5),
.O6(CLBLM_R_X11Y152_SLICE_X14Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf7ffffffffffffff)
  ) CLBLM_R_X11Y152_SLICE_X14Y152_CLUT (
.I0(CLBLM_L_X12Y151_SLICE_X16Y151_AQ),
.I1(CLBLM_R_X11Y152_SLICE_X14Y152_AQ),
.I2(CLBLM_L_X10Y153_SLICE_X12Y153_DO6),
.I3(CLBLM_R_X11Y152_SLICE_X14Y152_A5Q),
.I4(CLBLM_R_X11Y151_SLICE_X14Y151_AQ),
.I5(CLBLM_L_X10Y152_SLICE_X12Y152_AQ),
.O5(CLBLM_R_X11Y152_SLICE_X14Y152_CO5),
.O6(CLBLM_R_X11Y152_SLICE_X14Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3323ffff00100000)
  ) CLBLM_R_X11Y152_SLICE_X14Y152_BLUT (
.I0(CLBLM_L_X10Y153_SLICE_X12Y153_DO6),
.I1(CLBLM_L_X8Y153_SLICE_X10Y153_AQ),
.I2(CLBLM_R_X11Y151_SLICE_X14Y151_AQ),
.I3(CLBLM_R_X3Y150_SLICE_X3Y150_BQ),
.I4(CLBLM_R_X7Y145_SLICE_X8Y145_B5Q),
.I5(CLBLM_R_X11Y152_SLICE_X14Y152_A5Q),
.O5(CLBLM_R_X11Y152_SLICE_X14Y152_BO5),
.O6(CLBLM_R_X11Y152_SLICE_X14Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hb8b8b8b8ffcc3300)
  ) CLBLM_R_X11Y152_SLICE_X14Y152_ALUT (
.I0(CLBLM_R_X5Y150_SLICE_X7Y150_AQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X11Y152_SLICE_X15Y152_AO6),
.I3(CLBLM_R_X11Y152_SLICE_X14Y152_BO6),
.I4(CLBLM_R_X11Y150_SLICE_X14Y150_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y152_SLICE_X14Y152_AO5),
.O6(CLBLM_R_X11Y152_SLICE_X14Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y152_SLICE_X15Y152_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y152_SLICE_X15Y152_DO5),
.O6(CLBLM_R_X11Y152_SLICE_X15Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y152_SLICE_X15Y152_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y152_SLICE_X15Y152_CO5),
.O6(CLBLM_R_X11Y152_SLICE_X15Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3233ffff3333ffff)
  ) CLBLM_R_X11Y152_SLICE_X15Y152_BLUT (
.I0(CLBLM_L_X12Y151_SLICE_X16Y151_DO6),
.I1(CLBLM_L_X8Y153_SLICE_X10Y153_AQ),
.I2(CLBLM_R_X3Y150_SLICE_X3Y150_BQ),
.I3(CLBLM_L_X12Y151_SLICE_X16Y151_BQ),
.I4(CLBLM_R_X7Y145_SLICE_X8Y145_B5Q),
.I5(CLBLM_L_X10Y152_SLICE_X13Y152_AQ),
.O5(CLBLM_R_X11Y152_SLICE_X15Y152_BO5),
.O6(CLBLM_R_X11Y152_SLICE_X15Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00efffff00100000)
  ) CLBLM_R_X11Y152_SLICE_X15Y152_ALUT (
.I0(CLBLM_R_X11Y151_SLICE_X14Y151_DO6),
.I1(CLBLM_R_X3Y150_SLICE_X3Y150_BQ),
.I2(CLBLM_L_X12Y151_SLICE_X16Y151_AQ),
.I3(CLBLM_L_X8Y153_SLICE_X10Y153_AQ),
.I4(CLBLM_R_X7Y145_SLICE_X8Y145_B5Q),
.I5(CLBLM_R_X11Y152_SLICE_X14Y152_AQ),
.O5(CLBLM_R_X11Y152_SLICE_X15Y152_AO5),
.O6(CLBLM_R_X11Y152_SLICE_X15Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y153_SLICE_X14Y153_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y153_SLICE_X14Y153_DO5),
.O6(CLBLM_R_X11Y153_SLICE_X14Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y153_SLICE_X14Y153_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y153_SLICE_X14Y153_CO5),
.O6(CLBLM_R_X11Y153_SLICE_X14Y153_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y153_SLICE_X14Y153_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y153_SLICE_X14Y153_BO5),
.O6(CLBLM_R_X11Y153_SLICE_X14Y153_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff33ff33bbbbbbbb)
  ) CLBLM_R_X11Y153_SLICE_X14Y153_ALUT (
.I0(CLBLM_L_X10Y145_SLICE_X13Y145_CO6),
.I1(CLBLM_R_X3Y151_SLICE_X3Y151_D5Q),
.I2(1'b1),
.I3(CLBLM_L_X10Y148_SLICE_X13Y148_CO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y153_SLICE_X14Y153_AO5),
.O6(CLBLM_R_X11Y153_SLICE_X14Y153_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y153_SLICE_X15Y153_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y153_SLICE_X15Y153_DO5),
.O6(CLBLM_R_X11Y153_SLICE_X15Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y153_SLICE_X15Y153_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y153_SLICE_X15Y153_CO5),
.O6(CLBLM_R_X11Y153_SLICE_X15Y153_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y153_SLICE_X15Y153_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y153_SLICE_X15Y153_BO5),
.O6(CLBLM_R_X11Y153_SLICE_X15Y153_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y153_SLICE_X15Y153_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y153_SLICE_X15Y153_AO5),
.O6(CLBLM_R_X11Y153_SLICE_X15Y153_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y145_SLICE_X18Y145_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y145_SLICE_X18Y145_DO5),
.O6(CLBLM_R_X13Y145_SLICE_X18Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y145_SLICE_X18Y145_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y145_SLICE_X18Y145_CO5),
.O6(CLBLM_R_X13Y145_SLICE_X18Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y145_SLICE_X18Y145_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y145_SLICE_X18Y145_BO5),
.O6(CLBLM_R_X13Y145_SLICE_X18Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfaf0aa00faf0aa00)
  ) CLBLM_R_X13Y145_SLICE_X18Y145_ALUT (
.I0(CLBLM_R_X11Y148_SLICE_X14Y148_DQ),
.I1(1'b1),
.I2(CLBLM_R_X11Y148_SLICE_X14Y148_BQ),
.I3(RIOB33_X105Y143_IOB_X1Y144_I),
.I4(RIOB33_X105Y143_IOB_X1Y143_I),
.I5(1'b1),
.O5(CLBLM_R_X13Y145_SLICE_X18Y145_AO5),
.O6(CLBLM_R_X13Y145_SLICE_X18Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y145_SLICE_X19Y145_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y145_SLICE_X19Y145_DO5),
.O6(CLBLM_R_X13Y145_SLICE_X19Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y145_SLICE_X19Y145_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y145_SLICE_X19Y145_CO5),
.O6(CLBLM_R_X13Y145_SLICE_X19Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y145_SLICE_X19Y145_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y145_SLICE_X19Y145_BO5),
.O6(CLBLM_R_X13Y145_SLICE_X19Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y145_SLICE_X19Y145_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y145_SLICE_X19Y145_AO5),
.O6(CLBLM_R_X13Y145_SLICE_X19Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y178_SLICE_X162Y178_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y178_SLICE_X162Y178_DO5),
.O6(CLBLM_R_X103Y178_SLICE_X162Y178_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y178_SLICE_X162Y178_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y178_SLICE_X162Y178_CO5),
.O6(CLBLM_R_X103Y178_SLICE_X162Y178_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y178_SLICE_X162Y178_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y178_SLICE_X162Y178_BO5),
.O6(CLBLM_R_X103Y178_SLICE_X162Y178_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y178_SLICE_X162Y178_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y178_SLICE_X162Y178_AO5),
.O6(CLBLM_R_X103Y178_SLICE_X162Y178_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y178_SLICE_X163Y178_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y178_SLICE_X163Y178_DO5),
.O6(CLBLM_R_X103Y178_SLICE_X163Y178_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y178_SLICE_X163Y178_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y178_SLICE_X163Y178_CO5),
.O6(CLBLM_R_X103Y178_SLICE_X163Y178_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y178_SLICE_X163Y178_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y178_SLICE_X163Y178_BO5),
.O6(CLBLM_R_X103Y178_SLICE_X163Y178_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd88dd88dd88dd88)
  ) CLBLM_R_X103Y178_SLICE_X163Y178_ALUT (
.I0(RIOB33_X105Y127_IOB_X1Y127_I),
.I1(RIOB33_X105Y125_IOB_X1Y125_I),
.I2(1'b1),
.I3(RIOB33_X105Y125_IOB_X1Y126_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y178_SLICE_X163Y178_AO5),
.O6(CLBLM_R_X103Y178_SLICE_X163Y178_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFGCTRL" *)
  BUFGCTRL #(
    .INIT_OUT(0),
    .IS_CE0_INVERTED(0),
    .IS_CE1_INVERTED(1),
    .IS_IGNORE0_INVERTED(1),
    .IS_IGNORE1_INVERTED(0),
    .IS_S0_INVERTED(0),
    .IS_S1_INVERTED(1),
    .PRESELECT_I0("TRUE"),
    .PRESELECT_I1("FALSE")
  ) CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_BUFGCTRL (
.CE0(1'b1),
.CE1(1'b1),
.I0(LIOB33_X0Y77_IOB_X0Y78_I),
.I1(1'b1),
.IGNORE0(1'b1),
.IGNORE1(1'b1),
.O(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.S0(1'b1),
.S1(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFHCE" *)
  BUFHCE #(
    .CE_TYPE("SYNC"),
    .INIT_OUT(0),
    .IS_CE_INVERTED(0)
  ) CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_BUFHCE (
.CE(1'b1),
.I(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.O(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFHCE" *)
  BUFHCE #(
    .CE_TYPE("SYNC"),
    .INIT_OUT(0),
    .IS_CE_INVERTED(0)
  ) CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_BUFHCE (
.CE(1'b1),
.I(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.O(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y51_IOB_X0Y51_IBUF (
.I(LIOB33_X0Y51_IOB_X0Y51_IPAD),
.O(LIOB33_X0Y51_IOB_X0Y51_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y51_IOB_X0Y52_IBUF (
.I(LIOB33_X0Y51_IOB_X0Y52_IPAD),
.O(LIOB33_X0Y51_IOB_X0Y52_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y53_IOB_X0Y53_IBUF (
.I(LIOB33_X0Y53_IOB_X0Y53_IPAD),
.O(LIOB33_X0Y53_IOB_X0Y53_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y53_IOB_X0Y54_IBUF (
.I(LIOB33_X0Y53_IOB_X0Y54_IPAD),
.O(LIOB33_X0Y53_IOB_X0Y54_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y55_IOB_X0Y55_IBUF (
.I(LIOB33_X0Y55_IOB_X0Y55_IPAD),
.O(LIOB33_X0Y55_IOB_X0Y55_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y55_IOB_X0Y56_IBUF (
.I(LIOB33_X0Y55_IOB_X0Y56_IPAD),
.O(LIOB33_X0Y55_IOB_X0Y56_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y57_IOB_X0Y57_IBUF (
.I(LIOB33_X0Y57_IOB_X0Y57_IPAD),
.O(LIOB33_X0Y57_IOB_X0Y57_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y57_IOB_X0Y58_IBUF (
.I(LIOB33_X0Y57_IOB_X0Y58_IPAD),
.O(LIOB33_X0Y57_IOB_X0Y58_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y59_IOB_X0Y59_IBUF (
.I(LIOB33_X0Y59_IOB_X0Y59_IPAD),
.O(LIOB33_X0Y59_IOB_X0Y59_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y59_IOB_X0Y60_IBUF (
.I(LIOB33_X0Y59_IOB_X0Y60_IPAD),
.O(LIOB33_X0Y59_IOB_X0Y60_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y61_IOB_X0Y61_IBUF (
.I(LIOB33_X0Y61_IOB_X0Y61_IPAD),
.O(LIOB33_X0Y61_IOB_X0Y61_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y61_IOB_X0Y62_IBUF (
.I(LIOB33_X0Y61_IOB_X0Y62_IPAD),
.O(LIOB33_X0Y61_IOB_X0Y62_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y63_IOB_X0Y63_IBUF (
.I(LIOB33_X0Y63_IOB_X0Y63_IPAD),
.O(LIOB33_X0Y63_IOB_X0Y63_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y63_IOB_X0Y64_OBUF (
.I(CLBLL_L_X4Y140_SLICE_X5Y140_BO6),
.O(LIOB33_X0Y63_IOB_X0Y64_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y65_IOB_X0Y65_OBUF (
.I(CLBLL_L_X4Y140_SLICE_X5Y140_CO6),
.O(LIOB33_X0Y65_IOB_X0Y65_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y65_IOB_X0Y66_OBUF (
.I(CLBLM_R_X7Y152_SLICE_X9Y152_DQ),
.O(LIOB33_X0Y65_IOB_X0Y66_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y77_IOB_X0Y78_IBUF (
.I(LIOB33_X0Y77_IOB_X0Y78_IPAD),
.O(LIOB33_X0Y77_IOB_X0Y78_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y101_IOB_X0Y101_OBUF (
.I(CLBLM_R_X3Y142_SLICE_X2Y142_B5Q),
.O(LIOB33_X0Y101_IOB_X0Y101_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y101_IOB_X0Y102_OBUF (
.I(CLBLM_R_X5Y140_SLICE_X7Y140_BQ),
.O(LIOB33_X0Y101_IOB_X0Y102_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y103_IOB_X0Y103_OBUF (
.I(CLBLL_L_X4Y150_SLICE_X5Y150_DQ),
.O(LIOB33_X0Y103_IOB_X0Y103_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y103_IOB_X0Y104_OBUF (
.I(CLBLM_R_X7Y144_SLICE_X9Y144_C5Q),
.O(LIOB33_X0Y103_IOB_X0Y104_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y105_IOB_X0Y105_OBUF (
.I(CLBLM_R_X5Y144_SLICE_X6Y144_B5Q),
.O(LIOB33_X0Y105_IOB_X0Y105_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y105_IOB_X0Y106_OBUF (
.I(CLBLL_L_X4Y147_SLICE_X5Y147_DQ),
.O(LIOB33_X0Y105_IOB_X0Y106_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y107_IOB_X0Y107_OBUF (
.I(CLBLM_R_X3Y145_SLICE_X2Y145_C5Q),
.O(LIOB33_X0Y107_IOB_X0Y107_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y107_IOB_X0Y108_OBUF (
.I(CLBLL_L_X4Y143_SLICE_X5Y143_C5Q),
.O(LIOB33_X0Y107_IOB_X0Y108_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y109_IOB_X0Y109_OBUF (
.I(CLBLL_L_X2Y153_SLICE_X1Y153_AQ),
.O(LIOB33_X0Y109_IOB_X0Y109_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y109_IOB_X0Y110_OBUF (
.I(CLBLM_R_X5Y143_SLICE_X6Y143_DQ),
.O(LIOB33_X0Y109_IOB_X0Y110_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y111_IOB_X0Y111_OBUF (
.I(CLBLM_R_X3Y145_SLICE_X2Y145_CQ),
.O(LIOB33_X0Y111_IOB_X0Y111_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y111_IOB_X0Y112_OBUF (
.I(CLBLM_R_X3Y145_SLICE_X2Y145_B5Q),
.O(LIOB33_X0Y111_IOB_X0Y112_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y113_IOB_X0Y113_OBUF (
.I(CLBLM_R_X3Y146_SLICE_X2Y146_CQ),
.O(LIOB33_X0Y113_IOB_X0Y113_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y113_IOB_X0Y114_OBUF (
.I(CLBLL_L_X4Y153_SLICE_X4Y153_A5Q),
.O(LIOB33_X0Y113_IOB_X0Y114_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y115_IOB_X0Y115_OBUF (
.I(CLBLM_R_X3Y151_SLICE_X3Y151_CQ),
.O(LIOB33_X0Y115_IOB_X0Y115_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y115_IOB_X0Y116_OBUF (
.I(CLBLM_R_X5Y152_SLICE_X6Y152_CQ),
.O(LIOB33_X0Y115_IOB_X0Y116_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y117_IOB_X0Y117_OBUF (
.I(CLBLM_R_X7Y144_SLICE_X9Y144_B5Q),
.O(LIOB33_X0Y117_IOB_X0Y117_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y117_IOB_X0Y118_OBUF (
.I(CLBLM_R_X11Y147_SLICE_X15Y147_AQ),
.O(LIOB33_X0Y117_IOB_X0Y118_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y119_IOB_X0Y119_OBUF (
.I(CLBLM_R_X3Y149_SLICE_X2Y149_CQ),
.O(LIOB33_X0Y119_IOB_X0Y119_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y119_IOB_X0Y120_OBUF (
.I(CLBLM_R_X3Y150_SLICE_X3Y150_AQ),
.O(LIOB33_X0Y119_IOB_X0Y120_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y121_IOB_X0Y121_OBUF (
.I(CLBLM_L_X8Y146_SLICE_X10Y146_AQ),
.O(LIOB33_X0Y121_IOB_X0Y121_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y121_IOB_X0Y122_OBUF (
.I(CLBLL_L_X4Y149_SLICE_X4Y149_D5Q),
.O(LIOB33_X0Y121_IOB_X0Y122_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y123_IOB_X0Y123_OBUF (
.I(CLBLM_R_X3Y149_SLICE_X2Y149_CQ),
.O(LIOB33_X0Y123_IOB_X0Y123_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y123_IOB_X0Y124_OBUF (
.I(CLBLM_R_X7Y152_SLICE_X9Y152_DQ),
.O(LIOB33_X0Y123_IOB_X0Y124_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y125_IOB_X0Y125_OBUF (
.I(CLBLM_R_X5Y144_SLICE_X6Y144_DQ),
.O(LIOB33_X0Y125_IOB_X0Y125_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y125_IOB_X0Y126_OBUF (
.I(CLBLM_R_X5Y144_SLICE_X6Y144_CQ),
.O(LIOB33_X0Y125_IOB_X0Y126_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y127_IOB_X0Y127_OBUF (
.I(CLBLM_L_X8Y150_SLICE_X11Y150_B5Q),
.O(LIOB33_X0Y127_IOB_X0Y127_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y127_IOB_X0Y128_OBUF (
.I(CLBLM_L_X8Y142_SLICE_X11Y142_CQ),
.O(LIOB33_X0Y127_IOB_X0Y128_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y129_IOB_X0Y129_OBUF (
.I(CLBLM_R_X3Y149_SLICE_X2Y149_CQ),
.O(LIOB33_X0Y129_IOB_X0Y129_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y129_IOB_X0Y130_OBUF (
.I(CLBLM_R_X3Y149_SLICE_X2Y149_BQ),
.O(LIOB33_X0Y129_IOB_X0Y130_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y131_IOB_X0Y131_OBUF (
.I(CLBLL_L_X2Y75_SLICE_X0Y75_AO6),
.O(LIOB33_X0Y131_IOB_X0Y131_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y131_IOB_X0Y132_OBUF (
.I(CLBLL_L_X4Y142_SLICE_X4Y142_BO5),
.O(LIOB33_X0Y131_IOB_X0Y132_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y133_IOB_X0Y133_OBUF (
.I(CLBLM_R_X3Y142_SLICE_X2Y142_CO5),
.O(LIOB33_X0Y133_IOB_X0Y133_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y133_IOB_X0Y134_OBUF (
.I(CLBLM_R_X3Y149_SLICE_X2Y149_BQ),
.O(LIOB33_X0Y133_IOB_X0Y134_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y135_IOB_X0Y135_OBUF (
.I(CLBLM_R_X3Y149_SLICE_X2Y149_BQ),
.O(LIOB33_X0Y135_IOB_X0Y135_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y135_IOB_X0Y136_OBUF (
.I(CLBLM_L_X8Y153_SLICE_X10Y153_AQ),
.O(LIOB33_X0Y135_IOB_X0Y136_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y137_IOB_X0Y137_OBUF (
.I(CLBLM_R_X7Y150_SLICE_X9Y150_B5Q),
.O(LIOB33_X0Y137_IOB_X0Y137_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y137_IOB_X0Y138_OBUF (
.I(CLBLM_R_X3Y144_SLICE_X3Y144_A5Q),
.O(LIOB33_X0Y137_IOB_X0Y138_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y139_IOB_X0Y139_OBUF (
.I(CLBLL_L_X2Y148_SLICE_X0Y148_AQ),
.O(LIOB33_X0Y139_IOB_X0Y139_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y139_IOB_X0Y140_OBUF (
.I(CLBLL_L_X2Y147_SLICE_X0Y147_BQ),
.O(LIOB33_X0Y139_IOB_X0Y140_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y141_IOB_X0Y141_OBUF (
.I(CLBLL_L_X2Y150_SLICE_X1Y150_C5Q),
.O(LIOB33_X0Y141_IOB_X0Y141_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y141_IOB_X0Y142_OBUF (
.I(CLBLM_R_X3Y149_SLICE_X2Y149_CQ),
.O(LIOB33_X0Y141_IOB_X0Y142_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y143_IOB_X0Y143_OBUF (
.I(CLBLL_L_X2Y150_SLICE_X1Y150_DO5),
.O(LIOB33_X0Y143_IOB_X0Y143_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y145_IOB_X0Y145_OBUF (
.I(CLBLL_L_X2Y146_SLICE_X1Y146_CO6),
.O(LIOB33_X0Y145_IOB_X0Y145_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y145_IOB_X0Y146_OBUF (
.I(CLBLL_L_X2Y148_SLICE_X1Y148_BO6),
.O(LIOB33_X0Y145_IOB_X0Y146_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y147_IOB_X0Y147_OBUF (
.I(CLBLM_R_X5Y147_SLICE_X7Y147_DO6),
.O(LIOB33_X0Y147_IOB_X0Y147_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y147_IOB_X0Y148_OBUF (
.I(CLBLM_R_X3Y149_SLICE_X2Y149_DO6),
.O(LIOB33_X0Y147_IOB_X0Y148_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y151_IOB_X0Y151_OBUF (
.I(CLBLM_R_X3Y149_SLICE_X2Y149_CQ),
.O(LIOB33_X0Y151_IOB_X0Y151_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y151_IOB_X0Y152_OBUF (
.I(CLBLM_R_X3Y150_SLICE_X2Y150_B5Q),
.O(LIOB33_X0Y151_IOB_X0Y152_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y153_IOB_X0Y153_OBUF (
.I(CLBLM_L_X10Y153_SLICE_X13Y153_AQ),
.O(LIOB33_X0Y153_IOB_X0Y153_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y153_IOB_X0Y154_OBUF (
.I(CLBLM_L_X8Y152_SLICE_X10Y152_DQ),
.O(LIOB33_X0Y153_IOB_X0Y154_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y155_IOB_X0Y155_OBUF (
.I(CLBLM_L_X8Y150_SLICE_X11Y150_CQ),
.O(LIOB33_X0Y155_IOB_X0Y155_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y155_IOB_X0Y156_OBUF (
.I(CLBLM_R_X7Y152_SLICE_X9Y152_BQ),
.O(LIOB33_X0Y155_IOB_X0Y156_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y157_IOB_X0Y157_OBUF (
.I(CLBLM_R_X7Y153_SLICE_X9Y153_CQ),
.O(LIOB33_X0Y157_IOB_X0Y157_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y157_IOB_X0Y158_OBUF (
.I(RIOB33_X105Y133_IOB_X1Y134_I),
.O(LIOB33_X0Y157_IOB_X0Y158_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y159_IOB_X0Y159_OBUF (
.I(CLBLM_R_X3Y149_SLICE_X2Y149_CQ),
.O(LIOB33_X0Y159_IOB_X0Y159_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y159_IOB_X0Y160_OBUF (
.I(CLBLL_L_X4Y145_SLICE_X5Y145_AQ),
.O(LIOB33_X0Y159_IOB_X0Y160_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y161_IOB_X0Y161_OBUF (
.I(CLBLM_R_X5Y151_SLICE_X6Y151_CQ),
.O(LIOB33_X0Y161_IOB_X0Y161_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y161_IOB_X0Y162_OBUF (
.I(CLBLM_R_X3Y153_SLICE_X3Y153_CO6),
.O(LIOB33_X0Y161_IOB_X0Y162_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y163_IOB_X0Y163_OBUF (
.I(CLBLM_R_X5Y159_SLICE_X6Y159_AO6),
.O(LIOB33_X0Y163_IOB_X0Y163_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y163_IOB_X0Y164_OBUF (
.I(RIOB33_X105Y101_IOB_X1Y102_I),
.O(LIOB33_X0Y163_IOB_X0Y164_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y165_IOB_X0Y165_OBUF (
.I(LIOB33_X0Y57_IOB_X0Y57_I),
.O(LIOB33_X0Y165_IOB_X0Y165_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y165_IOB_X0Y166_OBUF (
.I(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.O(LIOB33_X0Y165_IOB_X0Y166_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y167_IOB_X0Y167_OBUF (
.I(RIOB33_X105Y105_IOB_X1Y106_I),
.O(LIOB33_X0Y167_IOB_X0Y167_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y167_IOB_X0Y168_OBUF (
.I(RIOB33_X105Y101_IOB_X1Y101_I),
.O(LIOB33_X0Y167_IOB_X0Y168_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y169_IOB_X0Y169_OBUF (
.I(RIOB33_X105Y117_IOB_X1Y117_I),
.O(LIOB33_X0Y169_IOB_X0Y169_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y169_IOB_X0Y170_OBUF (
.I(RIOB33_X105Y117_IOB_X1Y118_I),
.O(LIOB33_X0Y169_IOB_X0Y170_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y171_IOB_X0Y171_OBUF (
.I(RIOB33_X105Y119_IOB_X1Y119_I),
.O(LIOB33_X0Y171_IOB_X0Y171_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y171_IOB_X0Y172_OBUF (
.I(RIOB33_X105Y119_IOB_X1Y120_I),
.O(LIOB33_X0Y171_IOB_X0Y172_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y173_IOB_X0Y173_OBUF (
.I(RIOB33_X105Y121_IOB_X1Y121_I),
.O(LIOB33_X0Y173_IOB_X0Y173_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y173_IOB_X0Y174_OBUF (
.I(RIOB33_X105Y121_IOB_X1Y122_I),
.O(LIOB33_X0Y173_IOB_X0Y174_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y175_IOB_X0Y175_OBUF (
.I(RIOB33_X105Y123_IOB_X1Y123_I),
.O(LIOB33_X0Y175_IOB_X0Y175_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y175_IOB_X0Y176_OBUF (
.I(RIOB33_X105Y115_IOB_X1Y116_I),
.O(LIOB33_X0Y175_IOB_X0Y176_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y177_IOB_X0Y177_OBUF (
.I(RIOB33_X105Y123_IOB_X1Y124_I),
.O(LIOB33_X0Y177_IOB_X0Y177_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y177_IOB_X0Y178_OBUF (
.I(RIOB33_X105Y125_IOB_X1Y125_I),
.O(LIOB33_X0Y177_IOB_X0Y178_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y179_IOB_X0Y179_OBUF (
.I(RIOB33_X105Y125_IOB_X1Y126_I),
.O(LIOB33_X0Y179_IOB_X0Y179_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y179_IOB_X0Y180_OBUF (
.I(RIOB33_X105Y127_IOB_X1Y127_I),
.O(LIOB33_X0Y179_IOB_X0Y180_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y181_IOB_X0Y181_OBUF (
.I(RIOB33_X105Y127_IOB_X1Y128_I),
.O(LIOB33_X0Y181_IOB_X0Y181_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y181_IOB_X0Y182_OBUF (
.I(RIOB33_X105Y129_IOB_X1Y129_I),
.O(LIOB33_X0Y181_IOB_X0Y182_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y183_IOB_X0Y183_OBUF (
.I(RIOB33_X105Y129_IOB_X1Y130_I),
.O(LIOB33_X0Y183_IOB_X0Y183_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y183_IOB_X0Y184_OBUF (
.I(RIOB33_X105Y131_IOB_X1Y132_I),
.O(LIOB33_X0Y183_IOB_X0Y184_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y185_IOB_X0Y185_OBUF (
.I(RIOB33_X105Y133_IOB_X1Y133_I),
.O(LIOB33_X0Y185_IOB_X0Y185_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y185_IOB_X0Y186_OBUF (
.I(RIOB33_X105Y119_IOB_X1Y120_I),
.O(LIOB33_X0Y185_IOB_X0Y186_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y187_IOB_X0Y187_OBUF (
.I(CLBLM_L_X10Y150_SLICE_X12Y150_CQ),
.O(LIOB33_X0Y187_IOB_X0Y187_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y187_IOB_X0Y188_OBUF (
.I(CLBLM_R_X3Y150_SLICE_X3Y150_BQ),
.O(LIOB33_X0Y187_IOB_X0Y188_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y189_IOB_X0Y189_OBUF (
.I(CLBLM_R_X3Y149_SLICE_X3Y149_DQ),
.O(LIOB33_X0Y189_IOB_X0Y189_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y189_IOB_X0Y190_OBUF (
.I(CLBLM_R_X7Y155_SLICE_X9Y155_AO6),
.O(LIOB33_X0Y189_IOB_X0Y190_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y191_IOB_X0Y191_OBUF (
.I(CLBLL_L_X4Y145_SLICE_X4Y145_BO6),
.O(LIOB33_X0Y191_IOB_X0Y191_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y191_IOB_X0Y192_OBUF (
.I(CLBLL_L_X4Y154_SLICE_X4Y154_AO5),
.O(LIOB33_X0Y191_IOB_X0Y192_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y193_IOB_X0Y193_OBUF (
.I(CLBLL_L_X2Y166_SLICE_X0Y166_AO6),
.O(LIOB33_X0Y193_IOB_X0Y193_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y193_IOB_X0Y194_OBUF (
.I(RIOB33_X105Y103_IOB_X1Y103_I),
.O(LIOB33_X0Y193_IOB_X0Y194_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y195_IOB_X0Y195_OBUF (
.I(CLBLL_L_X2Y152_SLICE_X1Y152_AO6),
.O(LIOB33_X0Y195_IOB_X0Y195_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y195_IOB_X0Y196_OBUF (
.I(CLBLL_L_X4Y154_SLICE_X5Y154_AO6),
.O(LIOB33_X0Y195_IOB_X0Y196_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y197_IOB_X0Y197_OBUF (
.I(CLBLM_R_X3Y153_SLICE_X3Y153_BO5),
.O(LIOB33_X0Y197_IOB_X0Y197_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y197_IOB_X0Y198_OBUF (
.I(1'b1),
.O(LIOB33_X0Y197_IOB_X0Y198_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_SING_X0Y50_IOB_X0Y50_IBUF (
.I(LIOB33_SING_X0Y50_IOB_X0Y50_IPAD),
.O(LIOB33_SING_X0Y50_IOB_X0Y50_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y100_IOB_X0Y100_OBUF (
.I(CLBLM_R_X3Y149_SLICE_X2Y149_AQ),
.O(LIOB33_SING_X0Y100_IOB_X0Y100_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y149_IOB_X0Y149_OBUF (
.I(RIOB33_X105Y115_IOB_X1Y115_I),
.O(LIOB33_SING_X0Y149_IOB_X0Y149_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y150_IOB_X0Y150_OBUF (
.I(CLBLL_L_X4Y142_SLICE_X4Y142_DO5),
.O(LIOB33_SING_X0Y150_IOB_X0Y150_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y199_IOB_X0Y199_OBUF (
.I(1'b1),
.O(LIOB33_SING_X0Y199_IOB_X0Y199_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y101_IOB_X1Y101_IBUF (
.I(RIOB33_X105Y101_IOB_X1Y101_IPAD),
.O(RIOB33_X105Y101_IOB_X1Y101_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y101_IOB_X1Y102_IBUF (
.I(RIOB33_X105Y101_IOB_X1Y102_IPAD),
.O(RIOB33_X105Y101_IOB_X1Y102_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y103_IOB_X1Y103_IBUF (
.I(RIOB33_X105Y103_IOB_X1Y103_IPAD),
.O(RIOB33_X105Y103_IOB_X1Y103_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y103_IOB_X1Y104_IBUF (
.I(RIOB33_X105Y103_IOB_X1Y104_IPAD),
.O(RIOB33_X105Y103_IOB_X1Y104_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y105_IOB_X1Y105_IBUF (
.I(RIOB33_X105Y105_IOB_X1Y105_IPAD),
.O(RIOB33_X105Y105_IOB_X1Y105_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y105_IOB_X1Y106_IBUF (
.I(RIOB33_X105Y105_IOB_X1Y106_IPAD),
.O(RIOB33_X105Y105_IOB_X1Y106_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y107_IOB_X1Y107_IBUF (
.I(RIOB33_X105Y107_IOB_X1Y107_IPAD),
.O(RIOB33_X105Y107_IOB_X1Y107_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y107_IOB_X1Y108_IBUF (
.I(RIOB33_X105Y107_IOB_X1Y108_IPAD),
.O(RIOB33_X105Y107_IOB_X1Y108_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y109_IOB_X1Y109_IBUF (
.I(RIOB33_X105Y109_IOB_X1Y109_IPAD),
.O(RIOB33_X105Y109_IOB_X1Y109_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y109_IOB_X1Y110_IBUF (
.I(RIOB33_X105Y109_IOB_X1Y110_IPAD),
.O(RIOB33_X105Y109_IOB_X1Y110_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y111_IOB_X1Y111_IBUF (
.I(RIOB33_X105Y111_IOB_X1Y111_IPAD),
.O(RIOB33_X105Y111_IOB_X1Y111_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y111_IOB_X1Y112_IBUF (
.I(RIOB33_X105Y111_IOB_X1Y112_IPAD),
.O(RIOB33_X105Y111_IOB_X1Y112_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y113_IOB_X1Y113_IBUF (
.I(RIOB33_X105Y113_IOB_X1Y113_IPAD),
.O(RIOB33_X105Y113_IOB_X1Y113_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y113_IOB_X1Y114_IBUF (
.I(RIOB33_X105Y113_IOB_X1Y114_IPAD),
.O(RIOB33_X105Y113_IOB_X1Y114_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y115_IOB_X1Y115_IBUF (
.I(RIOB33_X105Y115_IOB_X1Y115_IPAD),
.O(RIOB33_X105Y115_IOB_X1Y115_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y115_IOB_X1Y116_IBUF (
.I(RIOB33_X105Y115_IOB_X1Y116_IPAD),
.O(RIOB33_X105Y115_IOB_X1Y116_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y117_IOB_X1Y117_IBUF (
.I(RIOB33_X105Y117_IOB_X1Y117_IPAD),
.O(RIOB33_X105Y117_IOB_X1Y117_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y117_IOB_X1Y118_IBUF (
.I(RIOB33_X105Y117_IOB_X1Y118_IPAD),
.O(RIOB33_X105Y117_IOB_X1Y118_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y119_IOB_X1Y119_IBUF (
.I(RIOB33_X105Y119_IOB_X1Y119_IPAD),
.O(RIOB33_X105Y119_IOB_X1Y119_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y119_IOB_X1Y120_IBUF (
.I(RIOB33_X105Y119_IOB_X1Y120_IPAD),
.O(RIOB33_X105Y119_IOB_X1Y120_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y121_IOB_X1Y121_IBUF (
.I(RIOB33_X105Y121_IOB_X1Y121_IPAD),
.O(RIOB33_X105Y121_IOB_X1Y121_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y121_IOB_X1Y122_IBUF (
.I(RIOB33_X105Y121_IOB_X1Y122_IPAD),
.O(RIOB33_X105Y121_IOB_X1Y122_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y123_IOB_X1Y123_IBUF (
.I(RIOB33_X105Y123_IOB_X1Y123_IPAD),
.O(RIOB33_X105Y123_IOB_X1Y123_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y123_IOB_X1Y124_IBUF (
.I(RIOB33_X105Y123_IOB_X1Y124_IPAD),
.O(RIOB33_X105Y123_IOB_X1Y124_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y125_IOB_X1Y125_IBUF (
.I(RIOB33_X105Y125_IOB_X1Y125_IPAD),
.O(RIOB33_X105Y125_IOB_X1Y125_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y125_IOB_X1Y126_IBUF (
.I(RIOB33_X105Y125_IOB_X1Y126_IPAD),
.O(RIOB33_X105Y125_IOB_X1Y126_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y127_IOB_X1Y127_IBUF (
.I(RIOB33_X105Y127_IOB_X1Y127_IPAD),
.O(RIOB33_X105Y127_IOB_X1Y127_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y127_IOB_X1Y128_IBUF (
.I(RIOB33_X105Y127_IOB_X1Y128_IPAD),
.O(RIOB33_X105Y127_IOB_X1Y128_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y129_IOB_X1Y129_IBUF (
.I(RIOB33_X105Y129_IOB_X1Y129_IPAD),
.O(RIOB33_X105Y129_IOB_X1Y129_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y129_IOB_X1Y130_IBUF (
.I(RIOB33_X105Y129_IOB_X1Y130_IPAD),
.O(RIOB33_X105Y129_IOB_X1Y130_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y131_IOB_X1Y131_IBUF (
.I(RIOB33_X105Y131_IOB_X1Y131_IPAD),
.O(RIOB33_X105Y131_IOB_X1Y131_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y131_IOB_X1Y132_IBUF (
.I(RIOB33_X105Y131_IOB_X1Y132_IPAD),
.O(RIOB33_X105Y131_IOB_X1Y132_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y133_IOB_X1Y133_IBUF (
.I(RIOB33_X105Y133_IOB_X1Y133_IPAD),
.O(RIOB33_X105Y133_IOB_X1Y133_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y133_IOB_X1Y134_IBUF (
.I(RIOB33_X105Y133_IOB_X1Y134_IPAD),
.O(RIOB33_X105Y133_IOB_X1Y134_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y135_IOB_X1Y135_IBUF (
.I(RIOB33_X105Y135_IOB_X1Y135_IPAD),
.O(RIOB33_X105Y135_IOB_X1Y135_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y135_IOB_X1Y136_IBUF (
.I(RIOB33_X105Y135_IOB_X1Y136_IPAD),
.O(RIOB33_X105Y135_IOB_X1Y136_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y137_IOB_X1Y137_IBUF (
.I(RIOB33_X105Y137_IOB_X1Y137_IPAD),
.O(RIOB33_X105Y137_IOB_X1Y137_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y137_IOB_X1Y138_IBUF (
.I(RIOB33_X105Y137_IOB_X1Y138_IPAD),
.O(RIOB33_X105Y137_IOB_X1Y138_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y139_IOB_X1Y139_IBUF (
.I(RIOB33_X105Y139_IOB_X1Y139_IPAD),
.O(RIOB33_X105Y139_IOB_X1Y139_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y139_IOB_X1Y140_IBUF (
.I(RIOB33_X105Y139_IOB_X1Y140_IPAD),
.O(RIOB33_X105Y139_IOB_X1Y140_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y141_IOB_X1Y141_IBUF (
.I(RIOB33_X105Y141_IOB_X1Y141_IPAD),
.O(RIOB33_X105Y141_IOB_X1Y141_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y141_IOB_X1Y142_IBUF (
.I(RIOB33_X105Y141_IOB_X1Y142_IPAD),
.O(RIOB33_X105Y141_IOB_X1Y142_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y143_IOB_X1Y143_IBUF (
.I(RIOB33_X105Y143_IOB_X1Y143_IPAD),
.O(RIOB33_X105Y143_IOB_X1Y143_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y143_IOB_X1Y144_IBUF (
.I(RIOB33_X105Y143_IOB_X1Y144_IPAD),
.O(RIOB33_X105Y143_IOB_X1Y144_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y145_IOB_X1Y145_IBUF (
.I(RIOB33_X105Y145_IOB_X1Y145_IPAD),
.O(RIOB33_X105Y145_IOB_X1Y145_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y145_IOB_X1Y146_IBUF (
.I(RIOB33_X105Y145_IOB_X1Y146_IPAD),
.O(RIOB33_X105Y145_IOB_X1Y146_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y147_IOB_X1Y147_IBUF (
.I(RIOB33_X105Y147_IOB_X1Y147_IPAD),
.O(RIOB33_X105Y147_IOB_X1Y147_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y147_IOB_X1Y148_IBUF (
.I(RIOB33_X105Y147_IOB_X1Y148_IPAD),
.O(RIOB33_X105Y147_IOB_X1Y148_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y151_IOB_X1Y151_OBUF (
.I(1'b1),
.O(RIOB33_X105Y151_IOB_X1Y151_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y151_IOB_X1Y152_OBUF (
.I(1'b1),
.O(RIOB33_X105Y151_IOB_X1Y152_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y153_IOB_X1Y153_OBUF (
.I(1'b1),
.O(RIOB33_X105Y153_IOB_X1Y153_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y153_IOB_X1Y154_OBUF (
.I(1'b1),
.O(RIOB33_X105Y153_IOB_X1Y154_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y155_IOB_X1Y155_OBUF (
.I(1'b1),
.O(RIOB33_X105Y155_IOB_X1Y155_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y155_IOB_X1Y156_OBUF (
.I(1'b1),
.O(RIOB33_X105Y155_IOB_X1Y156_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y157_IOB_X1Y157_OBUF (
.I(1'b1),
.O(RIOB33_X105Y157_IOB_X1Y157_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y157_IOB_X1Y158_OBUF (
.I(1'b1),
.O(RIOB33_X105Y157_IOB_X1Y158_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y159_IOB_X1Y159_OBUF (
.I(1'b1),
.O(RIOB33_X105Y159_IOB_X1Y159_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y159_IOB_X1Y160_OBUF (
.I(1'b1),
.O(RIOB33_X105Y159_IOB_X1Y160_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y161_IOB_X1Y161_OBUF (
.I(CLBLM_L_X8Y153_SLICE_X11Y153_AO5),
.O(RIOB33_X105Y161_IOB_X1Y161_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y161_IOB_X1Y162_OBUF (
.I(CLBLM_L_X10Y150_SLICE_X13Y150_C5Q),
.O(RIOB33_X105Y161_IOB_X1Y162_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y163_IOB_X1Y163_OBUF (
.I(CLBLM_L_X10Y149_SLICE_X12Y149_BQ),
.O(RIOB33_X105Y163_IOB_X1Y163_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y163_IOB_X1Y164_OBUF (
.I(CLBLM_R_X11Y151_SLICE_X15Y151_A5Q),
.O(RIOB33_X105Y163_IOB_X1Y164_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y165_IOB_X1Y165_OBUF (
.I(CLBLM_R_X3Y153_SLICE_X2Y153_AO5),
.O(RIOB33_X105Y165_IOB_X1Y165_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y165_IOB_X1Y166_OBUF (
.I(CLBLM_L_X10Y153_SLICE_X13Y153_AQ),
.O(RIOB33_X105Y165_IOB_X1Y166_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y167_IOB_X1Y167_OBUF (
.I(CLBLM_L_X8Y152_SLICE_X10Y152_DQ),
.O(RIOB33_X105Y167_IOB_X1Y167_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y167_IOB_X1Y168_OBUF (
.I(CLBLM_L_X8Y150_SLICE_X11Y150_CQ),
.O(RIOB33_X105Y167_IOB_X1Y168_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y169_IOB_X1Y169_OBUF (
.I(CLBLM_R_X7Y152_SLICE_X9Y152_BQ),
.O(RIOB33_X105Y169_IOB_X1Y169_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y169_IOB_X1Y170_OBUF (
.I(CLBLM_R_X7Y153_SLICE_X9Y153_CQ),
.O(RIOB33_X105Y169_IOB_X1Y170_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y171_IOB_X1Y171_OBUF (
.I(CLBLM_R_X7Y153_SLICE_X8Y153_CO5),
.O(RIOB33_X105Y171_IOB_X1Y171_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y171_IOB_X1Y172_OBUF (
.I(CLBLL_L_X4Y145_SLICE_X5Y145_AQ),
.O(RIOB33_X105Y171_IOB_X1Y172_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y173_IOB_X1Y173_OBUF (
.I(CLBLM_R_X5Y151_SLICE_X6Y151_CQ),
.O(RIOB33_X105Y173_IOB_X1Y173_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y173_IOB_X1Y174_OBUF (
.I(CLBLM_R_X5Y159_SLICE_X6Y159_AO6),
.O(RIOB33_X105Y173_IOB_X1Y174_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y175_IOB_X1Y175_OBUF (
.I(CLBLM_R_X3Y153_SLICE_X3Y153_CO6),
.O(RIOB33_X105Y175_IOB_X1Y175_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y175_IOB_X1Y176_OBUF (
.I(CLBLL_L_X2Y151_SLICE_X1Y151_CO6),
.O(RIOB33_X105Y175_IOB_X1Y176_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y177_IOB_X1Y177_OBUF (
.I(CLBLM_L_X10Y142_SLICE_X12Y142_AQ),
.O(RIOB33_X105Y177_IOB_X1Y177_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y177_IOB_X1Y178_OBUF (
.I(CLBLM_R_X3Y150_SLICE_X3Y150_BQ),
.O(RIOB33_X105Y177_IOB_X1Y178_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y179_IOB_X1Y179_OBUF (
.I(CLBLM_R_X3Y149_SLICE_X3Y149_DQ),
.O(RIOB33_X105Y179_IOB_X1Y179_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y179_IOB_X1Y180_OBUF (
.I(CLBLM_L_X10Y150_SLICE_X12Y150_CQ),
.O(RIOB33_X105Y179_IOB_X1Y180_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y181_IOB_X1Y181_OBUF (
.I(CLBLM_R_X7Y155_SLICE_X9Y155_AO6),
.O(RIOB33_X105Y181_IOB_X1Y181_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y181_IOB_X1Y182_OBUF (
.I(CLBLM_R_X7Y153_SLICE_X8Y153_DO6),
.O(RIOB33_X105Y181_IOB_X1Y182_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y183_IOB_X1Y183_OBUF (
.I(1'b0),
.O(RIOB33_X105Y183_IOB_X1Y183_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y183_IOB_X1Y184_OBUF (
.I(CLBLL_L_X4Y154_SLICE_X5Y154_AO6),
.O(RIOB33_X105Y183_IOB_X1Y184_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y185_IOB_X1Y185_OBUF (
.I(CLBLM_L_X8Y154_SLICE_X10Y154_BO6),
.O(RIOB33_X105Y185_IOB_X1Y185_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y185_IOB_X1Y186_OBUF (
.I(CLBLM_R_X7Y154_SLICE_X9Y154_CO6),
.O(RIOB33_X105Y185_IOB_X1Y186_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y187_IOB_X1Y187_OBUF (
.I(CLBLM_R_X103Y178_SLICE_X163Y178_AO6),
.O(RIOB33_X105Y187_IOB_X1Y187_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y187_IOB_X1Y188_OBUF (
.I(CLBLM_R_X7Y153_SLICE_X8Y153_DO6),
.O(RIOB33_X105Y187_IOB_X1Y188_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y189_IOB_X1Y189_OBUF (
.I(CLBLM_R_X103Y178_SLICE_X163Y178_AO6),
.O(RIOB33_X105Y189_IOB_X1Y189_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y189_IOB_X1Y190_OBUF (
.I(CLBLM_R_X11Y153_SLICE_X14Y153_AO6),
.O(RIOB33_X105Y189_IOB_X1Y190_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y191_IOB_X1Y191_OBUF (
.I(CLBLM_R_X11Y149_SLICE_X14Y149_AO6),
.O(RIOB33_X105Y191_IOB_X1Y191_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y191_IOB_X1Y192_OBUF (
.I(CLBLM_L_X12Y151_SLICE_X16Y151_CO6),
.O(RIOB33_X105Y191_IOB_X1Y192_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y193_IOB_X1Y193_OBUF (
.I(CLBLM_R_X11Y153_SLICE_X14Y153_AO5),
.O(RIOB33_X105Y193_IOB_X1Y193_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y193_IOB_X1Y194_OBUF (
.I(CLBLM_L_X12Y151_SLICE_X16Y151_CO5),
.O(RIOB33_X105Y193_IOB_X1Y194_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y195_IOB_X1Y195_OBUF (
.I(CLBLM_R_X11Y149_SLICE_X14Y149_BO6),
.O(RIOB33_X105Y195_IOB_X1Y195_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y195_IOB_X1Y196_OBUF (
.I(CLBLM_R_X11Y150_SLICE_X14Y150_BO6),
.O(RIOB33_X105Y195_IOB_X1Y196_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y197_IOB_X1Y197_OBUF (
.I(CLBLM_R_X11Y150_SLICE_X14Y150_BO5),
.O(RIOB33_X105Y197_IOB_X1Y197_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y197_IOB_X1Y198_OBUF (
.I(CLBLM_R_X11Y149_SLICE_X14Y149_CO6),
.O(RIOB33_X105Y197_IOB_X1Y198_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_SING_X105Y100_IOB_X1Y100_IBUF (
.I(RIOB33_SING_X105Y100_IOB_X1Y100_IPAD),
.O(RIOB33_SING_X105Y100_IOB_X1Y100_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_SING_X105Y149_IOB_X1Y149_IBUF (
.I(RIOB33_SING_X105Y149_IOB_X1Y149_IPAD),
.O(RIOB33_SING_X105Y149_IOB_X1Y149_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_SING_X105Y150_IOB_X1Y150_OBUF (
.I(1'b1),
.O(RIOB33_SING_X105Y150_IOB_X1Y150_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_SING_X105Y199_IOB_X1Y199_OBUF (
.I(CLBLM_R_X11Y149_SLICE_X14Y149_AQ),
.O(RIOB33_SING_X105Y199_IOB_X1Y199_OPAD)
  );
  assign CLBLL_L_X2Y75_SLICE_X0Y75_A = CLBLL_L_X2Y75_SLICE_X0Y75_AO6;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_B = CLBLL_L_X2Y75_SLICE_X0Y75_BO6;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_C = CLBLL_L_X2Y75_SLICE_X0Y75_CO6;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_D = CLBLL_L_X2Y75_SLICE_X0Y75_DO6;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_A = CLBLL_L_X2Y75_SLICE_X1Y75_AO6;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_B = CLBLL_L_X2Y75_SLICE_X1Y75_BO6;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_C = CLBLL_L_X2Y75_SLICE_X1Y75_CO6;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_D = CLBLL_L_X2Y75_SLICE_X1Y75_DO6;
  assign CLBLL_L_X2Y143_SLICE_X0Y143_A = CLBLL_L_X2Y143_SLICE_X0Y143_AO6;
  assign CLBLL_L_X2Y143_SLICE_X0Y143_B = CLBLL_L_X2Y143_SLICE_X0Y143_BO6;
  assign CLBLL_L_X2Y143_SLICE_X0Y143_C = CLBLL_L_X2Y143_SLICE_X0Y143_CO6;
  assign CLBLL_L_X2Y143_SLICE_X0Y143_D = CLBLL_L_X2Y143_SLICE_X0Y143_DO6;
  assign CLBLL_L_X2Y143_SLICE_X1Y143_A = CLBLL_L_X2Y143_SLICE_X1Y143_AO6;
  assign CLBLL_L_X2Y143_SLICE_X1Y143_B = CLBLL_L_X2Y143_SLICE_X1Y143_BO6;
  assign CLBLL_L_X2Y143_SLICE_X1Y143_C = CLBLL_L_X2Y143_SLICE_X1Y143_CO6;
  assign CLBLL_L_X2Y143_SLICE_X1Y143_D = CLBLL_L_X2Y143_SLICE_X1Y143_DO6;
  assign CLBLL_L_X2Y144_SLICE_X0Y144_A = CLBLL_L_X2Y144_SLICE_X0Y144_AO6;
  assign CLBLL_L_X2Y144_SLICE_X0Y144_B = CLBLL_L_X2Y144_SLICE_X0Y144_BO6;
  assign CLBLL_L_X2Y144_SLICE_X0Y144_C = CLBLL_L_X2Y144_SLICE_X0Y144_CO6;
  assign CLBLL_L_X2Y144_SLICE_X0Y144_D = CLBLL_L_X2Y144_SLICE_X0Y144_DO6;
  assign CLBLL_L_X2Y144_SLICE_X1Y144_A = CLBLL_L_X2Y144_SLICE_X1Y144_AO6;
  assign CLBLL_L_X2Y144_SLICE_X1Y144_B = CLBLL_L_X2Y144_SLICE_X1Y144_BO6;
  assign CLBLL_L_X2Y144_SLICE_X1Y144_C = CLBLL_L_X2Y144_SLICE_X1Y144_CO6;
  assign CLBLL_L_X2Y144_SLICE_X1Y144_D = CLBLL_L_X2Y144_SLICE_X1Y144_DO6;
  assign CLBLL_L_X2Y144_SLICE_X1Y144_AMUX = CLBLL_L_X2Y144_SLICE_X1Y144_A5Q;
  assign CLBLL_L_X2Y144_SLICE_X1Y144_BMUX = CLBLL_L_X2Y144_SLICE_X1Y144_B5Q;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_A = CLBLL_L_X2Y145_SLICE_X0Y145_AO6;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_B = CLBLL_L_X2Y145_SLICE_X0Y145_BO6;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_C = CLBLL_L_X2Y145_SLICE_X0Y145_CO6;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_D = CLBLL_L_X2Y145_SLICE_X0Y145_DO6;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_A = CLBLL_L_X2Y145_SLICE_X1Y145_AO6;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_B = CLBLL_L_X2Y145_SLICE_X1Y145_BO6;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_C = CLBLL_L_X2Y145_SLICE_X1Y145_CO6;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_D = CLBLL_L_X2Y145_SLICE_X1Y145_DO6;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_AMUX = CLBLL_L_X2Y145_SLICE_X1Y145_A5Q;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_A = CLBLL_L_X2Y146_SLICE_X0Y146_AO6;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_B = CLBLL_L_X2Y146_SLICE_X0Y146_BO6;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_C = CLBLL_L_X2Y146_SLICE_X0Y146_CO6;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_D = CLBLL_L_X2Y146_SLICE_X0Y146_DO6;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_A = CLBLL_L_X2Y146_SLICE_X1Y146_AO6;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_B = CLBLL_L_X2Y146_SLICE_X1Y146_BO6;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_C = CLBLL_L_X2Y146_SLICE_X1Y146_CO6;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_D = CLBLL_L_X2Y146_SLICE_X1Y146_DO6;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_AMUX = CLBLL_L_X2Y146_SLICE_X1Y146_A5Q;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_A = CLBLL_L_X2Y147_SLICE_X0Y147_AO6;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_B = CLBLL_L_X2Y147_SLICE_X0Y147_BO6;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_C = CLBLL_L_X2Y147_SLICE_X0Y147_CO6;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_D = CLBLL_L_X2Y147_SLICE_X0Y147_DO6;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_BMUX = CLBLL_L_X2Y147_SLICE_X0Y147_B5Q;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_A = CLBLL_L_X2Y147_SLICE_X1Y147_AO6;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_B = CLBLL_L_X2Y147_SLICE_X1Y147_BO6;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_C = CLBLL_L_X2Y147_SLICE_X1Y147_CO6;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_D = CLBLL_L_X2Y147_SLICE_X1Y147_DO6;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_AMUX = CLBLL_L_X2Y147_SLICE_X1Y147_A5Q;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_A = CLBLL_L_X2Y148_SLICE_X0Y148_AO6;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_B = CLBLL_L_X2Y148_SLICE_X0Y148_BO6;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_C = CLBLL_L_X2Y148_SLICE_X0Y148_CO6;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_D = CLBLL_L_X2Y148_SLICE_X0Y148_DO6;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_AMUX = CLBLL_L_X2Y148_SLICE_X0Y148_A5Q;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_BMUX = CLBLL_L_X2Y148_SLICE_X0Y148_B5Q;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_A = CLBLL_L_X2Y148_SLICE_X1Y148_AO6;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_B = CLBLL_L_X2Y148_SLICE_X1Y148_BO6;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_C = CLBLL_L_X2Y148_SLICE_X1Y148_CO6;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_D = CLBLL_L_X2Y148_SLICE_X1Y148_DO6;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_AMUX = CLBLL_L_X2Y148_SLICE_X1Y148_A5Q;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_BMUX = CLBLL_L_X2Y148_SLICE_X1Y148_BO5;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_A = CLBLL_L_X2Y149_SLICE_X0Y149_AO6;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_B = CLBLL_L_X2Y149_SLICE_X0Y149_BO6;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_C = CLBLL_L_X2Y149_SLICE_X0Y149_CO6;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_D = CLBLL_L_X2Y149_SLICE_X0Y149_DO6;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_A = CLBLL_L_X2Y149_SLICE_X1Y149_AO6;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_B = CLBLL_L_X2Y149_SLICE_X1Y149_BO6;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_C = CLBLL_L_X2Y149_SLICE_X1Y149_CO6;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_D = CLBLL_L_X2Y149_SLICE_X1Y149_DO6;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_AMUX = CLBLL_L_X2Y149_SLICE_X1Y149_A5Q;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_A = CLBLL_L_X2Y150_SLICE_X0Y150_AO6;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_B = CLBLL_L_X2Y150_SLICE_X0Y150_BO6;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_C = CLBLL_L_X2Y150_SLICE_X0Y150_CO6;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_D = CLBLL_L_X2Y150_SLICE_X0Y150_DO6;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_A = CLBLL_L_X2Y150_SLICE_X1Y150_AO6;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_B = CLBLL_L_X2Y150_SLICE_X1Y150_BO6;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_C = CLBLL_L_X2Y150_SLICE_X1Y150_CO6;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_D = CLBLL_L_X2Y150_SLICE_X1Y150_DO6;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_AMUX = CLBLL_L_X2Y150_SLICE_X1Y150_A5Q;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_BMUX = CLBLL_L_X2Y150_SLICE_X1Y150_BO5;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_CMUX = CLBLL_L_X2Y150_SLICE_X1Y150_C5Q;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_DMUX = CLBLL_L_X2Y150_SLICE_X1Y150_DO5;
  assign CLBLL_L_X2Y151_SLICE_X0Y151_A = CLBLL_L_X2Y151_SLICE_X0Y151_AO6;
  assign CLBLL_L_X2Y151_SLICE_X0Y151_B = CLBLL_L_X2Y151_SLICE_X0Y151_BO6;
  assign CLBLL_L_X2Y151_SLICE_X0Y151_C = CLBLL_L_X2Y151_SLICE_X0Y151_CO6;
  assign CLBLL_L_X2Y151_SLICE_X0Y151_D = CLBLL_L_X2Y151_SLICE_X0Y151_DO6;
  assign CLBLL_L_X2Y151_SLICE_X1Y151_A = CLBLL_L_X2Y151_SLICE_X1Y151_AO6;
  assign CLBLL_L_X2Y151_SLICE_X1Y151_B = CLBLL_L_X2Y151_SLICE_X1Y151_BO6;
  assign CLBLL_L_X2Y151_SLICE_X1Y151_C = CLBLL_L_X2Y151_SLICE_X1Y151_CO6;
  assign CLBLL_L_X2Y151_SLICE_X1Y151_D = CLBLL_L_X2Y151_SLICE_X1Y151_DO6;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_A = CLBLL_L_X2Y152_SLICE_X0Y152_AO6;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_B = CLBLL_L_X2Y152_SLICE_X0Y152_BO6;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_C = CLBLL_L_X2Y152_SLICE_X0Y152_CO6;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_D = CLBLL_L_X2Y152_SLICE_X0Y152_DO6;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_A = CLBLL_L_X2Y152_SLICE_X1Y152_AO6;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_B = CLBLL_L_X2Y152_SLICE_X1Y152_BO6;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_C = CLBLL_L_X2Y152_SLICE_X1Y152_CO6;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_D = CLBLL_L_X2Y152_SLICE_X1Y152_DO6;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_A = CLBLL_L_X2Y153_SLICE_X0Y153_AO6;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_B = CLBLL_L_X2Y153_SLICE_X0Y153_BO6;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_C = CLBLL_L_X2Y153_SLICE_X0Y153_CO6;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_D = CLBLL_L_X2Y153_SLICE_X0Y153_DO6;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_A = CLBLL_L_X2Y153_SLICE_X1Y153_AO6;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_B = CLBLL_L_X2Y153_SLICE_X1Y153_BO6;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_C = CLBLL_L_X2Y153_SLICE_X1Y153_CO6;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_D = CLBLL_L_X2Y153_SLICE_X1Y153_DO6;
  assign CLBLL_L_X2Y166_SLICE_X0Y166_A = CLBLL_L_X2Y166_SLICE_X0Y166_AO6;
  assign CLBLL_L_X2Y166_SLICE_X0Y166_B = CLBLL_L_X2Y166_SLICE_X0Y166_BO6;
  assign CLBLL_L_X2Y166_SLICE_X0Y166_C = CLBLL_L_X2Y166_SLICE_X0Y166_CO6;
  assign CLBLL_L_X2Y166_SLICE_X0Y166_D = CLBLL_L_X2Y166_SLICE_X0Y166_DO6;
  assign CLBLL_L_X2Y166_SLICE_X1Y166_A = CLBLL_L_X2Y166_SLICE_X1Y166_AO6;
  assign CLBLL_L_X2Y166_SLICE_X1Y166_B = CLBLL_L_X2Y166_SLICE_X1Y166_BO6;
  assign CLBLL_L_X2Y166_SLICE_X1Y166_C = CLBLL_L_X2Y166_SLICE_X1Y166_CO6;
  assign CLBLL_L_X2Y166_SLICE_X1Y166_D = CLBLL_L_X2Y166_SLICE_X1Y166_DO6;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_A = CLBLL_L_X4Y140_SLICE_X4Y140_AO6;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_B = CLBLL_L_X4Y140_SLICE_X4Y140_BO6;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_C = CLBLL_L_X4Y140_SLICE_X4Y140_CO6;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_D = CLBLL_L_X4Y140_SLICE_X4Y140_DO6;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_A = CLBLL_L_X4Y140_SLICE_X5Y140_AO6;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_B = CLBLL_L_X4Y140_SLICE_X5Y140_BO6;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_C = CLBLL_L_X4Y140_SLICE_X5Y140_CO6;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_D = CLBLL_L_X4Y140_SLICE_X5Y140_DO6;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_A = CLBLL_L_X4Y141_SLICE_X4Y141_AO6;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_B = CLBLL_L_X4Y141_SLICE_X4Y141_BO6;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_C = CLBLL_L_X4Y141_SLICE_X4Y141_CO6;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_D = CLBLL_L_X4Y141_SLICE_X4Y141_DO6;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_A = CLBLL_L_X4Y141_SLICE_X5Y141_AO6;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_B = CLBLL_L_X4Y141_SLICE_X5Y141_BO6;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_C = CLBLL_L_X4Y141_SLICE_X5Y141_CO6;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_D = CLBLL_L_X4Y141_SLICE_X5Y141_DO6;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_AMUX = CLBLL_L_X4Y141_SLICE_X5Y141_A5Q;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_BMUX = CLBLL_L_X4Y141_SLICE_X5Y141_BO5;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_A = CLBLL_L_X4Y142_SLICE_X4Y142_AO6;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_B = CLBLL_L_X4Y142_SLICE_X4Y142_BO6;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_C = CLBLL_L_X4Y142_SLICE_X4Y142_CO6;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_D = CLBLL_L_X4Y142_SLICE_X4Y142_DO6;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_AMUX = CLBLL_L_X4Y142_SLICE_X4Y142_A5Q;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_BMUX = CLBLL_L_X4Y142_SLICE_X4Y142_BO5;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_CMUX = CLBLL_L_X4Y142_SLICE_X4Y142_CO5;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_DMUX = CLBLL_L_X4Y142_SLICE_X4Y142_DO5;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_A = CLBLL_L_X4Y142_SLICE_X5Y142_AO6;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_B = CLBLL_L_X4Y142_SLICE_X5Y142_BO6;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_C = CLBLL_L_X4Y142_SLICE_X5Y142_CO6;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_D = CLBLL_L_X4Y142_SLICE_X5Y142_DO6;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_AMUX = CLBLL_L_X4Y142_SLICE_X5Y142_A5Q;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_A = CLBLL_L_X4Y143_SLICE_X4Y143_AO6;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_B = CLBLL_L_X4Y143_SLICE_X4Y143_BO6;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_C = CLBLL_L_X4Y143_SLICE_X4Y143_CO6;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_D = CLBLL_L_X4Y143_SLICE_X4Y143_DO6;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_A = CLBLL_L_X4Y143_SLICE_X5Y143_AO6;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_B = CLBLL_L_X4Y143_SLICE_X5Y143_BO6;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_C = CLBLL_L_X4Y143_SLICE_X5Y143_CO6;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_D = CLBLL_L_X4Y143_SLICE_X5Y143_DO6;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_CMUX = CLBLL_L_X4Y143_SLICE_X5Y143_C5Q;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_A = CLBLL_L_X4Y144_SLICE_X4Y144_AO6;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_B = CLBLL_L_X4Y144_SLICE_X4Y144_BO6;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_C = CLBLL_L_X4Y144_SLICE_X4Y144_CO6;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_D = CLBLL_L_X4Y144_SLICE_X4Y144_DO6;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_BMUX = CLBLL_L_X4Y144_SLICE_X4Y144_BO6;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_A = CLBLL_L_X4Y144_SLICE_X5Y144_AO6;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_B = CLBLL_L_X4Y144_SLICE_X5Y144_BO6;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_C = CLBLL_L_X4Y144_SLICE_X5Y144_CO6;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_D = CLBLL_L_X4Y144_SLICE_X5Y144_DO6;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_BMUX = CLBLL_L_X4Y144_SLICE_X5Y144_B5Q;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_CMUX = CLBLL_L_X4Y144_SLICE_X5Y144_C5Q;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_DMUX = CLBLL_L_X4Y144_SLICE_X5Y144_D5Q;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_A = CLBLL_L_X4Y145_SLICE_X4Y145_AO6;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_B = CLBLL_L_X4Y145_SLICE_X4Y145_BO6;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_C = CLBLL_L_X4Y145_SLICE_X4Y145_CO6;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_D = CLBLL_L_X4Y145_SLICE_X4Y145_DO6;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_AMUX = CLBLL_L_X4Y145_SLICE_X4Y145_A5Q;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_A = CLBLL_L_X4Y145_SLICE_X5Y145_AO6;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_B = CLBLL_L_X4Y145_SLICE_X5Y145_BO6;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_C = CLBLL_L_X4Y145_SLICE_X5Y145_CO6;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_D = CLBLL_L_X4Y145_SLICE_X5Y145_DO6;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_A = CLBLL_L_X4Y146_SLICE_X4Y146_AO6;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_B = CLBLL_L_X4Y146_SLICE_X4Y146_BO6;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_C = CLBLL_L_X4Y146_SLICE_X4Y146_CO6;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_D = CLBLL_L_X4Y146_SLICE_X4Y146_DO6;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_A = CLBLL_L_X4Y146_SLICE_X5Y146_AO6;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_B = CLBLL_L_X4Y146_SLICE_X5Y146_BO6;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_C = CLBLL_L_X4Y146_SLICE_X5Y146_CO6;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_D = CLBLL_L_X4Y146_SLICE_X5Y146_DO6;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_AMUX = CLBLL_L_X4Y146_SLICE_X5Y146_A5Q;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_BMUX = CLBLL_L_X4Y146_SLICE_X5Y146_B5Q;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_CMUX = CLBLL_L_X4Y146_SLICE_X5Y146_CO6;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_A = CLBLL_L_X4Y147_SLICE_X4Y147_AO6;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_B = CLBLL_L_X4Y147_SLICE_X4Y147_BO6;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_C = CLBLL_L_X4Y147_SLICE_X4Y147_CO6;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_D = CLBLL_L_X4Y147_SLICE_X4Y147_DO6;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_CMUX = CLBLL_L_X4Y147_SLICE_X4Y147_C5Q;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_DMUX = CLBLL_L_X4Y147_SLICE_X4Y147_D5Q;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_A = CLBLL_L_X4Y147_SLICE_X5Y147_AO6;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_B = CLBLL_L_X4Y147_SLICE_X5Y147_BO6;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_C = CLBLL_L_X4Y147_SLICE_X5Y147_CO6;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_D = CLBLL_L_X4Y147_SLICE_X5Y147_DO6;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_BMUX = CLBLL_L_X4Y147_SLICE_X5Y147_B5Q;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_CMUX = CLBLL_L_X4Y147_SLICE_X5Y147_C5Q;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_A = CLBLL_L_X4Y148_SLICE_X4Y148_AO6;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_B = CLBLL_L_X4Y148_SLICE_X4Y148_BO6;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_C = CLBLL_L_X4Y148_SLICE_X4Y148_CO6;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_D = CLBLL_L_X4Y148_SLICE_X4Y148_DO6;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_AMUX = CLBLL_L_X4Y148_SLICE_X4Y148_A5Q;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_BMUX = CLBLL_L_X4Y148_SLICE_X4Y148_BO5;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_CMUX = CLBLL_L_X4Y148_SLICE_X4Y148_CO5;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_A = CLBLL_L_X4Y148_SLICE_X5Y148_AO6;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_B = CLBLL_L_X4Y148_SLICE_X5Y148_BO6;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_C = CLBLL_L_X4Y148_SLICE_X5Y148_CO6;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_D = CLBLL_L_X4Y148_SLICE_X5Y148_DO6;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_BMUX = CLBLL_L_X4Y148_SLICE_X5Y148_B5Q;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_A = CLBLL_L_X4Y149_SLICE_X4Y149_AO6;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_B = CLBLL_L_X4Y149_SLICE_X4Y149_BO6;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_C = CLBLL_L_X4Y149_SLICE_X4Y149_CO6;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_D = CLBLL_L_X4Y149_SLICE_X4Y149_DO6;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_BMUX = CLBLL_L_X4Y149_SLICE_X4Y149_B5Q;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_CMUX = CLBLL_L_X4Y149_SLICE_X4Y149_C5Q;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_DMUX = CLBLL_L_X4Y149_SLICE_X4Y149_D5Q;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_A = CLBLL_L_X4Y149_SLICE_X5Y149_AO6;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_B = CLBLL_L_X4Y149_SLICE_X5Y149_BO6;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_C = CLBLL_L_X4Y149_SLICE_X5Y149_CO6;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_D = CLBLL_L_X4Y149_SLICE_X5Y149_DO6;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_A = CLBLL_L_X4Y150_SLICE_X4Y150_AO6;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_B = CLBLL_L_X4Y150_SLICE_X4Y150_BO6;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_C = CLBLL_L_X4Y150_SLICE_X4Y150_CO6;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_D = CLBLL_L_X4Y150_SLICE_X4Y150_DO6;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_AMUX = CLBLL_L_X4Y150_SLICE_X4Y150_AO5;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_BMUX = CLBLL_L_X4Y150_SLICE_X4Y150_BO6;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_A = CLBLL_L_X4Y150_SLICE_X5Y150_AO6;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_B = CLBLL_L_X4Y150_SLICE_X5Y150_BO6;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_C = CLBLL_L_X4Y150_SLICE_X5Y150_CO6;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_D = CLBLL_L_X4Y150_SLICE_X5Y150_DO6;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_CMUX = CLBLL_L_X4Y150_SLICE_X5Y150_C5Q;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_DMUX = CLBLL_L_X4Y150_SLICE_X5Y150_D5Q;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_A = CLBLL_L_X4Y151_SLICE_X4Y151_AO6;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_B = CLBLL_L_X4Y151_SLICE_X4Y151_BO6;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_C = CLBLL_L_X4Y151_SLICE_X4Y151_CO6;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_D = CLBLL_L_X4Y151_SLICE_X4Y151_DO6;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_AMUX = CLBLL_L_X4Y151_SLICE_X4Y151_AO5;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_BMUX = CLBLL_L_X4Y151_SLICE_X4Y151_BO5;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_A = CLBLL_L_X4Y151_SLICE_X5Y151_AO6;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_B = CLBLL_L_X4Y151_SLICE_X5Y151_BO6;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_C = CLBLL_L_X4Y151_SLICE_X5Y151_CO6;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_D = CLBLL_L_X4Y151_SLICE_X5Y151_DO6;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_AMUX = CLBLL_L_X4Y151_SLICE_X5Y151_A5Q;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_A = CLBLL_L_X4Y152_SLICE_X4Y152_AO6;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_B = CLBLL_L_X4Y152_SLICE_X4Y152_BO6;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_C = CLBLL_L_X4Y152_SLICE_X4Y152_CO6;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_D = CLBLL_L_X4Y152_SLICE_X4Y152_DO6;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_CMUX = CLBLL_L_X4Y152_SLICE_X4Y152_C5Q;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_A = CLBLL_L_X4Y152_SLICE_X5Y152_AO6;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_B = CLBLL_L_X4Y152_SLICE_X5Y152_BO6;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_C = CLBLL_L_X4Y152_SLICE_X5Y152_CO6;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_D = CLBLL_L_X4Y152_SLICE_X5Y152_DO6;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_BMUX = CLBLL_L_X4Y152_SLICE_X5Y152_B5Q;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_CMUX = CLBLL_L_X4Y152_SLICE_X5Y152_C5Q;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_A = CLBLL_L_X4Y153_SLICE_X4Y153_AO6;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_B = CLBLL_L_X4Y153_SLICE_X4Y153_BO6;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_C = CLBLL_L_X4Y153_SLICE_X4Y153_CO6;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_D = CLBLL_L_X4Y153_SLICE_X4Y153_DO6;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_AMUX = CLBLL_L_X4Y153_SLICE_X4Y153_A5Q;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_DMUX = CLBLL_L_X4Y153_SLICE_X4Y153_DO5;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_A = CLBLL_L_X4Y153_SLICE_X5Y153_AO6;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_B = CLBLL_L_X4Y153_SLICE_X5Y153_BO6;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_C = CLBLL_L_X4Y153_SLICE_X5Y153_CO6;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_D = CLBLL_L_X4Y153_SLICE_X5Y153_DO6;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_DMUX = CLBLL_L_X4Y153_SLICE_X5Y153_DO6;
  assign CLBLL_L_X4Y154_SLICE_X4Y154_A = CLBLL_L_X4Y154_SLICE_X4Y154_AO6;
  assign CLBLL_L_X4Y154_SLICE_X4Y154_B = CLBLL_L_X4Y154_SLICE_X4Y154_BO6;
  assign CLBLL_L_X4Y154_SLICE_X4Y154_C = CLBLL_L_X4Y154_SLICE_X4Y154_CO6;
  assign CLBLL_L_X4Y154_SLICE_X4Y154_D = CLBLL_L_X4Y154_SLICE_X4Y154_DO6;
  assign CLBLL_L_X4Y154_SLICE_X4Y154_AMUX = CLBLL_L_X4Y154_SLICE_X4Y154_AO5;
  assign CLBLL_L_X4Y154_SLICE_X4Y154_BMUX = CLBLL_L_X4Y154_SLICE_X4Y154_BO5;
  assign CLBLL_L_X4Y154_SLICE_X5Y154_A = CLBLL_L_X4Y154_SLICE_X5Y154_AO6;
  assign CLBLL_L_X4Y154_SLICE_X5Y154_B = CLBLL_L_X4Y154_SLICE_X5Y154_BO6;
  assign CLBLL_L_X4Y154_SLICE_X5Y154_C = CLBLL_L_X4Y154_SLICE_X5Y154_CO6;
  assign CLBLL_L_X4Y154_SLICE_X5Y154_D = CLBLL_L_X4Y154_SLICE_X5Y154_DO6;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_A = CLBLM_L_X8Y140_SLICE_X10Y140_AO6;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_B = CLBLM_L_X8Y140_SLICE_X10Y140_BO6;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_C = CLBLM_L_X8Y140_SLICE_X10Y140_CO6;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_D = CLBLM_L_X8Y140_SLICE_X10Y140_DO6;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_AMUX = CLBLM_L_X8Y140_SLICE_X10Y140_A5Q;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_A = CLBLM_L_X8Y140_SLICE_X11Y140_AO6;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_B = CLBLM_L_X8Y140_SLICE_X11Y140_BO6;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_C = CLBLM_L_X8Y140_SLICE_X11Y140_CO6;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_D = CLBLM_L_X8Y140_SLICE_X11Y140_DO6;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_A = CLBLM_L_X8Y141_SLICE_X10Y141_AO6;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_B = CLBLM_L_X8Y141_SLICE_X10Y141_BO6;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_C = CLBLM_L_X8Y141_SLICE_X10Y141_CO6;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_D = CLBLM_L_X8Y141_SLICE_X10Y141_DO6;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_A = CLBLM_L_X8Y141_SLICE_X11Y141_AO6;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_B = CLBLM_L_X8Y141_SLICE_X11Y141_BO6;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_C = CLBLM_L_X8Y141_SLICE_X11Y141_CO6;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_D = CLBLM_L_X8Y141_SLICE_X11Y141_DO6;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_A = CLBLM_L_X8Y142_SLICE_X10Y142_AO6;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_B = CLBLM_L_X8Y142_SLICE_X10Y142_BO6;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_C = CLBLM_L_X8Y142_SLICE_X10Y142_CO6;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_D = CLBLM_L_X8Y142_SLICE_X10Y142_DO6;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_AMUX = CLBLM_L_X8Y142_SLICE_X10Y142_A5Q;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_BMUX = CLBLM_L_X8Y142_SLICE_X10Y142_BO5;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_CMUX = CLBLM_L_X8Y142_SLICE_X10Y142_C5Q;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_DMUX = CLBLM_L_X8Y142_SLICE_X10Y142_DO5;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_A = CLBLM_L_X8Y142_SLICE_X11Y142_AO6;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_B = CLBLM_L_X8Y142_SLICE_X11Y142_BO6;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_C = CLBLM_L_X8Y142_SLICE_X11Y142_CO6;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_D = CLBLM_L_X8Y142_SLICE_X11Y142_DO6;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_CMUX = CLBLM_L_X8Y142_SLICE_X11Y142_C5Q;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_A = CLBLM_L_X8Y143_SLICE_X10Y143_AO6;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_B = CLBLM_L_X8Y143_SLICE_X10Y143_BO6;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_C = CLBLM_L_X8Y143_SLICE_X10Y143_CO6;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_D = CLBLM_L_X8Y143_SLICE_X10Y143_DO6;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_A = CLBLM_L_X8Y143_SLICE_X11Y143_AO6;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_B = CLBLM_L_X8Y143_SLICE_X11Y143_BO6;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_C = CLBLM_L_X8Y143_SLICE_X11Y143_CO6;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_D = CLBLM_L_X8Y143_SLICE_X11Y143_DO6;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_AMUX = CLBLM_L_X8Y143_SLICE_X11Y143_A5Q;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_A = CLBLM_L_X8Y144_SLICE_X10Y144_AO6;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_B = CLBLM_L_X8Y144_SLICE_X10Y144_BO6;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_C = CLBLM_L_X8Y144_SLICE_X10Y144_CO6;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_D = CLBLM_L_X8Y144_SLICE_X10Y144_DO6;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_AMUX = CLBLM_L_X8Y144_SLICE_X10Y144_A5Q;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_BMUX = CLBLM_L_X8Y144_SLICE_X10Y144_B5Q;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_CMUX = CLBLM_L_X8Y144_SLICE_X10Y144_CO5;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_A = CLBLM_L_X8Y144_SLICE_X11Y144_AO6;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_B = CLBLM_L_X8Y144_SLICE_X11Y144_BO6;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_C = CLBLM_L_X8Y144_SLICE_X11Y144_CO6;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_D = CLBLM_L_X8Y144_SLICE_X11Y144_DO6;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_AMUX = CLBLM_L_X8Y144_SLICE_X11Y144_A5Q;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_A = CLBLM_L_X8Y145_SLICE_X10Y145_AO6;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_B = CLBLM_L_X8Y145_SLICE_X10Y145_BO6;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_C = CLBLM_L_X8Y145_SLICE_X10Y145_CO6;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_D = CLBLM_L_X8Y145_SLICE_X10Y145_DO6;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_AMUX = CLBLM_L_X8Y145_SLICE_X10Y145_AO5;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_BMUX = CLBLM_L_X8Y145_SLICE_X10Y145_BO5;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_CMUX = CLBLM_L_X8Y145_SLICE_X10Y145_CO5;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_A = CLBLM_L_X8Y145_SLICE_X11Y145_AO6;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_B = CLBLM_L_X8Y145_SLICE_X11Y145_BO6;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_C = CLBLM_L_X8Y145_SLICE_X11Y145_CO6;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_D = CLBLM_L_X8Y145_SLICE_X11Y145_DO6;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_AMUX = CLBLM_L_X8Y145_SLICE_X11Y145_AO5;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_BMUX = CLBLM_L_X8Y145_SLICE_X11Y145_BO6;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_A = CLBLM_L_X8Y146_SLICE_X10Y146_AO6;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_B = CLBLM_L_X8Y146_SLICE_X10Y146_BO6;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_C = CLBLM_L_X8Y146_SLICE_X10Y146_CO6;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_D = CLBLM_L_X8Y146_SLICE_X10Y146_DO6;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_AMUX = CLBLM_L_X8Y146_SLICE_X10Y146_A5Q;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_CMUX = CLBLM_L_X8Y146_SLICE_X10Y146_C5Q;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_A = CLBLM_L_X8Y146_SLICE_X11Y146_AO6;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_B = CLBLM_L_X8Y146_SLICE_X11Y146_BO6;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_C = CLBLM_L_X8Y146_SLICE_X11Y146_CO6;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_D = CLBLM_L_X8Y146_SLICE_X11Y146_DO6;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_AMUX = CLBLM_L_X8Y146_SLICE_X11Y146_A5Q;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_CMUX = CLBLM_L_X8Y146_SLICE_X11Y146_CO6;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_A = CLBLM_L_X8Y147_SLICE_X10Y147_AO6;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_B = CLBLM_L_X8Y147_SLICE_X10Y147_BO6;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_C = CLBLM_L_X8Y147_SLICE_X10Y147_CO6;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_D = CLBLM_L_X8Y147_SLICE_X10Y147_DO6;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_AMUX = CLBLM_L_X8Y147_SLICE_X10Y147_A5Q;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_BMUX = CLBLM_L_X8Y147_SLICE_X10Y147_B5Q;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_A = CLBLM_L_X8Y147_SLICE_X11Y147_AO6;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_B = CLBLM_L_X8Y147_SLICE_X11Y147_BO6;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_C = CLBLM_L_X8Y147_SLICE_X11Y147_CO6;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_D = CLBLM_L_X8Y147_SLICE_X11Y147_DO6;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_AMUX = CLBLM_L_X8Y147_SLICE_X11Y147_A5Q;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_A = CLBLM_L_X8Y148_SLICE_X10Y148_AO6;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_B = CLBLM_L_X8Y148_SLICE_X10Y148_BO6;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_C = CLBLM_L_X8Y148_SLICE_X10Y148_CO6;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_D = CLBLM_L_X8Y148_SLICE_X10Y148_DO6;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_AMUX = CLBLM_L_X8Y148_SLICE_X10Y148_A5Q;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_BMUX = CLBLM_L_X8Y148_SLICE_X10Y148_BO5;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_CMUX = CLBLM_L_X8Y148_SLICE_X10Y148_CO5;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_A = CLBLM_L_X8Y148_SLICE_X11Y148_AO6;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_B = CLBLM_L_X8Y148_SLICE_X11Y148_BO6;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_C = CLBLM_L_X8Y148_SLICE_X11Y148_CO6;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_D = CLBLM_L_X8Y148_SLICE_X11Y148_DO6;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_BMUX = CLBLM_L_X8Y148_SLICE_X11Y148_B5Q;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_CMUX = CLBLM_L_X8Y148_SLICE_X11Y148_C5Q;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_A = CLBLM_L_X8Y149_SLICE_X10Y149_AO6;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_B = CLBLM_L_X8Y149_SLICE_X10Y149_BO6;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_C = CLBLM_L_X8Y149_SLICE_X10Y149_CO6;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_D = CLBLM_L_X8Y149_SLICE_X10Y149_DO6;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_AMUX = CLBLM_L_X8Y149_SLICE_X10Y149_A5Q;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_BMUX = CLBLM_L_X8Y149_SLICE_X10Y149_B5Q;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_A = CLBLM_L_X8Y149_SLICE_X11Y149_AO6;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_B = CLBLM_L_X8Y149_SLICE_X11Y149_BO6;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_C = CLBLM_L_X8Y149_SLICE_X11Y149_CO6;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_D = CLBLM_L_X8Y149_SLICE_X11Y149_DO6;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_BMUX = CLBLM_L_X8Y149_SLICE_X11Y149_B5Q;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_A = CLBLM_L_X8Y150_SLICE_X10Y150_AO6;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_B = CLBLM_L_X8Y150_SLICE_X10Y150_BO6;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_C = CLBLM_L_X8Y150_SLICE_X10Y150_CO6;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_D = CLBLM_L_X8Y150_SLICE_X10Y150_DO6;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_AMUX = CLBLM_L_X8Y150_SLICE_X10Y150_A5Q;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_A = CLBLM_L_X8Y150_SLICE_X11Y150_AO6;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_B = CLBLM_L_X8Y150_SLICE_X11Y150_BO6;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_C = CLBLM_L_X8Y150_SLICE_X11Y150_CO6;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_D = CLBLM_L_X8Y150_SLICE_X11Y150_DO6;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_BMUX = CLBLM_L_X8Y150_SLICE_X11Y150_B5Q;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_A = CLBLM_L_X8Y151_SLICE_X10Y151_AO6;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_B = CLBLM_L_X8Y151_SLICE_X10Y151_BO6;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_C = CLBLM_L_X8Y151_SLICE_X10Y151_CO6;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_D = CLBLM_L_X8Y151_SLICE_X10Y151_DO6;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_BMUX = CLBLM_L_X8Y151_SLICE_X10Y151_B5Q;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_CMUX = CLBLM_L_X8Y151_SLICE_X10Y151_CO5;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_A = CLBLM_L_X8Y151_SLICE_X11Y151_AO6;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_B = CLBLM_L_X8Y151_SLICE_X11Y151_BO6;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_C = CLBLM_L_X8Y151_SLICE_X11Y151_CO6;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_D = CLBLM_L_X8Y151_SLICE_X11Y151_DO6;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_AMUX = CLBLM_L_X8Y151_SLICE_X11Y151_A5Q;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_BMUX = CLBLM_L_X8Y151_SLICE_X11Y151_BO5;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_A = CLBLM_L_X8Y152_SLICE_X10Y152_AO6;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_B = CLBLM_L_X8Y152_SLICE_X10Y152_BO6;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_C = CLBLM_L_X8Y152_SLICE_X10Y152_CO6;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_D = CLBLM_L_X8Y152_SLICE_X10Y152_DO6;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_DMUX = CLBLM_L_X8Y152_SLICE_X10Y152_D5Q;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_A = CLBLM_L_X8Y152_SLICE_X11Y152_AO6;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_B = CLBLM_L_X8Y152_SLICE_X11Y152_BO6;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_C = CLBLM_L_X8Y152_SLICE_X11Y152_CO6;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_D = CLBLM_L_X8Y152_SLICE_X11Y152_DO6;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_AMUX = CLBLM_L_X8Y152_SLICE_X11Y152_A5Q;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_BMUX = CLBLM_L_X8Y152_SLICE_X11Y152_B5Q;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_A = CLBLM_L_X8Y153_SLICE_X10Y153_AO6;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_B = CLBLM_L_X8Y153_SLICE_X10Y153_BO6;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_C = CLBLM_L_X8Y153_SLICE_X10Y153_CO6;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_D = CLBLM_L_X8Y153_SLICE_X10Y153_DO6;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_DMUX = CLBLM_L_X8Y153_SLICE_X10Y153_DO5;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_A = CLBLM_L_X8Y153_SLICE_X11Y153_AO6;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_B = CLBLM_L_X8Y153_SLICE_X11Y153_BO6;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_C = CLBLM_L_X8Y153_SLICE_X11Y153_CO6;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_D = CLBLM_L_X8Y153_SLICE_X11Y153_DO6;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_AMUX = CLBLM_L_X8Y153_SLICE_X11Y153_AO5;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_A = CLBLM_L_X8Y154_SLICE_X10Y154_AO6;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_B = CLBLM_L_X8Y154_SLICE_X10Y154_BO6;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_C = CLBLM_L_X8Y154_SLICE_X10Y154_CO6;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_D = CLBLM_L_X8Y154_SLICE_X10Y154_DO6;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_A = CLBLM_L_X8Y154_SLICE_X11Y154_AO6;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_B = CLBLM_L_X8Y154_SLICE_X11Y154_BO6;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_C = CLBLM_L_X8Y154_SLICE_X11Y154_CO6;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_D = CLBLM_L_X8Y154_SLICE_X11Y154_DO6;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_A = CLBLM_L_X10Y141_SLICE_X12Y141_AO6;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_B = CLBLM_L_X10Y141_SLICE_X12Y141_BO6;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_C = CLBLM_L_X10Y141_SLICE_X12Y141_CO6;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_D = CLBLM_L_X10Y141_SLICE_X12Y141_DO6;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_A = CLBLM_L_X10Y141_SLICE_X13Y141_AO6;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_B = CLBLM_L_X10Y141_SLICE_X13Y141_BO6;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_C = CLBLM_L_X10Y141_SLICE_X13Y141_CO6;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_D = CLBLM_L_X10Y141_SLICE_X13Y141_DO6;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_A = CLBLM_L_X10Y142_SLICE_X12Y142_AO6;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_B = CLBLM_L_X10Y142_SLICE_X12Y142_BO6;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_C = CLBLM_L_X10Y142_SLICE_X12Y142_CO6;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_D = CLBLM_L_X10Y142_SLICE_X12Y142_DO6;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_AMUX = CLBLM_L_X10Y142_SLICE_X12Y142_AO5;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_BMUX = CLBLM_L_X10Y142_SLICE_X12Y142_BO6;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_A = CLBLM_L_X10Y142_SLICE_X13Y142_AO6;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_B = CLBLM_L_X10Y142_SLICE_X13Y142_BO6;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_C = CLBLM_L_X10Y142_SLICE_X13Y142_CO6;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_D = CLBLM_L_X10Y142_SLICE_X13Y142_DO6;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_A = CLBLM_L_X10Y143_SLICE_X12Y143_AO6;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_B = CLBLM_L_X10Y143_SLICE_X12Y143_BO6;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_C = CLBLM_L_X10Y143_SLICE_X12Y143_CO6;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_D = CLBLM_L_X10Y143_SLICE_X12Y143_DO6;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_AMUX = CLBLM_L_X10Y143_SLICE_X12Y143_AO5;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_BMUX = CLBLM_L_X10Y143_SLICE_X12Y143_BO5;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_CMUX = CLBLM_L_X10Y143_SLICE_X12Y143_CO5;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_DMUX = CLBLM_L_X10Y143_SLICE_X12Y143_DO5;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_A = CLBLM_L_X10Y143_SLICE_X13Y143_AO6;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_B = CLBLM_L_X10Y143_SLICE_X13Y143_BO6;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_C = CLBLM_L_X10Y143_SLICE_X13Y143_CO6;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_D = CLBLM_L_X10Y143_SLICE_X13Y143_DO6;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_A = CLBLM_L_X10Y144_SLICE_X12Y144_AO6;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_B = CLBLM_L_X10Y144_SLICE_X12Y144_BO6;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_C = CLBLM_L_X10Y144_SLICE_X12Y144_CO6;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_D = CLBLM_L_X10Y144_SLICE_X12Y144_DO6;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_AMUX = CLBLM_L_X10Y144_SLICE_X12Y144_AO5;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_A = CLBLM_L_X10Y144_SLICE_X13Y144_AO6;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_B = CLBLM_L_X10Y144_SLICE_X13Y144_BO6;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_C = CLBLM_L_X10Y144_SLICE_X13Y144_CO6;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_D = CLBLM_L_X10Y144_SLICE_X13Y144_DO6;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_BMUX = CLBLM_L_X10Y144_SLICE_X13Y144_BO6;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_DMUX = CLBLM_L_X10Y144_SLICE_X13Y144_DO6;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_A = CLBLM_L_X10Y145_SLICE_X12Y145_AO6;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_B = CLBLM_L_X10Y145_SLICE_X12Y145_BO6;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_C = CLBLM_L_X10Y145_SLICE_X12Y145_CO6;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_D = CLBLM_L_X10Y145_SLICE_X12Y145_DO6;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_AMUX = CLBLM_L_X10Y145_SLICE_X12Y145_AO5;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_CMUX = CLBLM_L_X10Y145_SLICE_X12Y145_CO6;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_A = CLBLM_L_X10Y145_SLICE_X13Y145_AO6;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_B = CLBLM_L_X10Y145_SLICE_X13Y145_BO6;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_C = CLBLM_L_X10Y145_SLICE_X13Y145_CO6;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_D = CLBLM_L_X10Y145_SLICE_X13Y145_DO6;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_AMUX = CLBLM_L_X10Y145_SLICE_X13Y145_AO5;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_BMUX = CLBLM_L_X10Y145_SLICE_X13Y145_BO5;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_A = CLBLM_L_X10Y146_SLICE_X12Y146_AO6;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_B = CLBLM_L_X10Y146_SLICE_X12Y146_BO6;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_C = CLBLM_L_X10Y146_SLICE_X12Y146_CO6;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_D = CLBLM_L_X10Y146_SLICE_X12Y146_DO6;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_AMUX = CLBLM_L_X10Y146_SLICE_X12Y146_AO5;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_BMUX = CLBLM_L_X10Y146_SLICE_X12Y146_BO5;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_CMUX = CLBLM_L_X10Y146_SLICE_X12Y146_CO5;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_A = CLBLM_L_X10Y146_SLICE_X13Y146_AO6;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_B = CLBLM_L_X10Y146_SLICE_X13Y146_BO6;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_C = CLBLM_L_X10Y146_SLICE_X13Y146_CO6;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_D = CLBLM_L_X10Y146_SLICE_X13Y146_DO6;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_BMUX = CLBLM_L_X10Y146_SLICE_X13Y146_BO5;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_DMUX = CLBLM_L_X10Y146_SLICE_X13Y146_DO6;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_A = CLBLM_L_X10Y147_SLICE_X12Y147_AO6;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_B = CLBLM_L_X10Y147_SLICE_X12Y147_BO6;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_C = CLBLM_L_X10Y147_SLICE_X12Y147_CO6;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_D = CLBLM_L_X10Y147_SLICE_X12Y147_DO6;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_BMUX = CLBLM_L_X10Y147_SLICE_X12Y147_B5Q;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_CMUX = CLBLM_L_X10Y147_SLICE_X12Y147_C5Q;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_DMUX = CLBLM_L_X10Y147_SLICE_X12Y147_DO5;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_A = CLBLM_L_X10Y147_SLICE_X13Y147_AO6;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_B = CLBLM_L_X10Y147_SLICE_X13Y147_BO6;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_C = CLBLM_L_X10Y147_SLICE_X13Y147_CO6;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_D = CLBLM_L_X10Y147_SLICE_X13Y147_DO6;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_AMUX = CLBLM_L_X10Y147_SLICE_X13Y147_A5Q;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_BMUX = CLBLM_L_X10Y147_SLICE_X13Y147_B5Q;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_A = CLBLM_L_X10Y148_SLICE_X12Y148_AO6;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_B = CLBLM_L_X10Y148_SLICE_X12Y148_BO6;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_C = CLBLM_L_X10Y148_SLICE_X12Y148_CO6;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_D = CLBLM_L_X10Y148_SLICE_X12Y148_DO6;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_AMUX = CLBLM_L_X10Y148_SLICE_X12Y148_A5Q;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_BMUX = CLBLM_L_X10Y148_SLICE_X12Y148_BO5;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_A = CLBLM_L_X10Y148_SLICE_X13Y148_AO6;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_B = CLBLM_L_X10Y148_SLICE_X13Y148_BO6;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_C = CLBLM_L_X10Y148_SLICE_X13Y148_CO6;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_D = CLBLM_L_X10Y148_SLICE_X13Y148_DO6;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_AMUX = CLBLM_L_X10Y148_SLICE_X13Y148_AO5;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_BMUX = CLBLM_L_X10Y148_SLICE_X13Y148_BO5;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_A = CLBLM_L_X10Y149_SLICE_X12Y149_AO6;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_B = CLBLM_L_X10Y149_SLICE_X12Y149_BO6;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_C = CLBLM_L_X10Y149_SLICE_X12Y149_CO6;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_D = CLBLM_L_X10Y149_SLICE_X12Y149_DO6;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_AMUX = CLBLM_L_X10Y149_SLICE_X12Y149_A5Q;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_BMUX = CLBLM_L_X10Y149_SLICE_X12Y149_B5Q;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_A = CLBLM_L_X10Y149_SLICE_X13Y149_AO6;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_B = CLBLM_L_X10Y149_SLICE_X13Y149_BO6;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_C = CLBLM_L_X10Y149_SLICE_X13Y149_CO6;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_D = CLBLM_L_X10Y149_SLICE_X13Y149_DO6;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_AMUX = CLBLM_L_X10Y149_SLICE_X13Y149_A5Q;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_BMUX = CLBLM_L_X10Y149_SLICE_X13Y149_BO5;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_A = CLBLM_L_X10Y150_SLICE_X12Y150_AO6;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_B = CLBLM_L_X10Y150_SLICE_X12Y150_BO6;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_C = CLBLM_L_X10Y150_SLICE_X12Y150_CO6;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_D = CLBLM_L_X10Y150_SLICE_X12Y150_DO6;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_AMUX = CLBLM_L_X10Y150_SLICE_X12Y150_A5Q;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_DMUX = CLBLM_L_X10Y150_SLICE_X12Y150_DO5;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_A = CLBLM_L_X10Y150_SLICE_X13Y150_AO6;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_B = CLBLM_L_X10Y150_SLICE_X13Y150_BO6;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_C = CLBLM_L_X10Y150_SLICE_X13Y150_CO6;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_D = CLBLM_L_X10Y150_SLICE_X13Y150_DO6;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_AMUX = CLBLM_L_X10Y150_SLICE_X13Y150_A5Q;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_BMUX = CLBLM_L_X10Y150_SLICE_X13Y150_B5Q;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_CMUX = CLBLM_L_X10Y150_SLICE_X13Y150_C5Q;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_DMUX = CLBLM_L_X10Y150_SLICE_X13Y150_DO5;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_A = CLBLM_L_X10Y151_SLICE_X12Y151_AO6;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_B = CLBLM_L_X10Y151_SLICE_X12Y151_BO6;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_C = CLBLM_L_X10Y151_SLICE_X12Y151_CO6;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_D = CLBLM_L_X10Y151_SLICE_X12Y151_DO6;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_AMUX = CLBLM_L_X10Y151_SLICE_X12Y151_AO5;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_A = CLBLM_L_X10Y151_SLICE_X13Y151_AO6;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_B = CLBLM_L_X10Y151_SLICE_X13Y151_BO6;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_C = CLBLM_L_X10Y151_SLICE_X13Y151_CO6;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_D = CLBLM_L_X10Y151_SLICE_X13Y151_DO6;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_BMUX = CLBLM_L_X10Y151_SLICE_X13Y151_BO5;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_DMUX = CLBLM_L_X10Y151_SLICE_X13Y151_DO6;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_A = CLBLM_L_X10Y152_SLICE_X12Y152_AO6;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_B = CLBLM_L_X10Y152_SLICE_X12Y152_BO6;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_C = CLBLM_L_X10Y152_SLICE_X12Y152_CO6;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_D = CLBLM_L_X10Y152_SLICE_X12Y152_DO6;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_A = CLBLM_L_X10Y152_SLICE_X13Y152_AO6;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_B = CLBLM_L_X10Y152_SLICE_X13Y152_BO6;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_C = CLBLM_L_X10Y152_SLICE_X13Y152_CO6;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_D = CLBLM_L_X10Y152_SLICE_X13Y152_DO6;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_CMUX = CLBLM_L_X10Y152_SLICE_X13Y152_CO5;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_A = CLBLM_L_X10Y153_SLICE_X12Y153_AO6;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_B = CLBLM_L_X10Y153_SLICE_X12Y153_BO6;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_C = CLBLM_L_X10Y153_SLICE_X12Y153_CO6;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_D = CLBLM_L_X10Y153_SLICE_X12Y153_DO6;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_DMUX = CLBLM_L_X10Y153_SLICE_X12Y153_DO5;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_A = CLBLM_L_X10Y153_SLICE_X13Y153_AO6;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_B = CLBLM_L_X10Y153_SLICE_X13Y153_BO6;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_C = CLBLM_L_X10Y153_SLICE_X13Y153_CO6;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_D = CLBLM_L_X10Y153_SLICE_X13Y153_DO6;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_A = CLBLM_L_X12Y143_SLICE_X16Y143_AO6;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_B = CLBLM_L_X12Y143_SLICE_X16Y143_BO6;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_C = CLBLM_L_X12Y143_SLICE_X16Y143_CO6;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_D = CLBLM_L_X12Y143_SLICE_X16Y143_DO6;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_A = CLBLM_L_X12Y143_SLICE_X17Y143_AO6;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_B = CLBLM_L_X12Y143_SLICE_X17Y143_BO6;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_C = CLBLM_L_X12Y143_SLICE_X17Y143_CO6;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_D = CLBLM_L_X12Y143_SLICE_X17Y143_DO6;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_A = CLBLM_L_X12Y144_SLICE_X16Y144_AO6;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_B = CLBLM_L_X12Y144_SLICE_X16Y144_BO6;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_C = CLBLM_L_X12Y144_SLICE_X16Y144_CO6;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_D = CLBLM_L_X12Y144_SLICE_X16Y144_DO6;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_AMUX = CLBLM_L_X12Y144_SLICE_X16Y144_AO5;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_A = CLBLM_L_X12Y144_SLICE_X17Y144_AO6;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_B = CLBLM_L_X12Y144_SLICE_X17Y144_BO6;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_C = CLBLM_L_X12Y144_SLICE_X17Y144_CO6;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_D = CLBLM_L_X12Y144_SLICE_X17Y144_DO6;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_A = CLBLM_L_X12Y145_SLICE_X16Y145_AO6;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_B = CLBLM_L_X12Y145_SLICE_X16Y145_BO6;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_C = CLBLM_L_X12Y145_SLICE_X16Y145_CO6;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_D = CLBLM_L_X12Y145_SLICE_X16Y145_DO6;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_AMUX = CLBLM_L_X12Y145_SLICE_X16Y145_AO5;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_DMUX = CLBLM_L_X12Y145_SLICE_X16Y145_DO6;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_A = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_B = CLBLM_L_X12Y145_SLICE_X17Y145_BO6;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_C = CLBLM_L_X12Y145_SLICE_X17Y145_CO6;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_D = CLBLM_L_X12Y145_SLICE_X17Y145_DO6;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_CMUX = CLBLM_L_X12Y145_SLICE_X17Y145_CO6;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_A = CLBLM_L_X12Y146_SLICE_X16Y146_AO6;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_B = CLBLM_L_X12Y146_SLICE_X16Y146_BO6;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_C = CLBLM_L_X12Y146_SLICE_X16Y146_CO6;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_D = CLBLM_L_X12Y146_SLICE_X16Y146_DO6;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_A = CLBLM_L_X12Y146_SLICE_X17Y146_AO6;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_B = CLBLM_L_X12Y146_SLICE_X17Y146_BO6;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_C = CLBLM_L_X12Y146_SLICE_X17Y146_CO6;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_D = CLBLM_L_X12Y146_SLICE_X17Y146_DO6;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_A = CLBLM_L_X12Y149_SLICE_X16Y149_AO6;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_B = CLBLM_L_X12Y149_SLICE_X16Y149_BO6;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_C = CLBLM_L_X12Y149_SLICE_X16Y149_CO6;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_D = CLBLM_L_X12Y149_SLICE_X16Y149_DO6;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_DMUX = CLBLM_L_X12Y149_SLICE_X16Y149_DO6;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_A = CLBLM_L_X12Y149_SLICE_X17Y149_AO6;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_B = CLBLM_L_X12Y149_SLICE_X17Y149_BO6;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_C = CLBLM_L_X12Y149_SLICE_X17Y149_CO6;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_D = CLBLM_L_X12Y149_SLICE_X17Y149_DO6;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_A = CLBLM_L_X12Y151_SLICE_X16Y151_AO6;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_B = CLBLM_L_X12Y151_SLICE_X16Y151_BO6;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_C = CLBLM_L_X12Y151_SLICE_X16Y151_CO6;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_D = CLBLM_L_X12Y151_SLICE_X16Y151_DO6;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_CMUX = CLBLM_L_X12Y151_SLICE_X16Y151_CO5;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_A = CLBLM_L_X12Y151_SLICE_X17Y151_AO6;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_B = CLBLM_L_X12Y151_SLICE_X17Y151_BO6;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_C = CLBLM_L_X12Y151_SLICE_X17Y151_CO6;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_D = CLBLM_L_X12Y151_SLICE_X17Y151_DO6;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_A = CLBLM_R_X3Y141_SLICE_X2Y141_AO6;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_B = CLBLM_R_X3Y141_SLICE_X2Y141_BO6;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_C = CLBLM_R_X3Y141_SLICE_X2Y141_CO6;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_D = CLBLM_R_X3Y141_SLICE_X2Y141_DO6;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_AMUX = CLBLM_R_X3Y141_SLICE_X2Y141_AO5;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_A = CLBLM_R_X3Y141_SLICE_X3Y141_AO6;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_B = CLBLM_R_X3Y141_SLICE_X3Y141_BO6;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_C = CLBLM_R_X3Y141_SLICE_X3Y141_CO6;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_D = CLBLM_R_X3Y141_SLICE_X3Y141_DO6;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_A = CLBLM_R_X3Y142_SLICE_X2Y142_AO6;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_B = CLBLM_R_X3Y142_SLICE_X2Y142_BO6;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_C = CLBLM_R_X3Y142_SLICE_X2Y142_CO6;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_D = CLBLM_R_X3Y142_SLICE_X2Y142_DO6;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_AMUX = CLBLM_R_X3Y142_SLICE_X2Y142_A5Q;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_BMUX = CLBLM_R_X3Y142_SLICE_X2Y142_B5Q;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_CMUX = CLBLM_R_X3Y142_SLICE_X2Y142_CO5;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_A = CLBLM_R_X3Y142_SLICE_X3Y142_AO6;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_B = CLBLM_R_X3Y142_SLICE_X3Y142_BO6;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_C = CLBLM_R_X3Y142_SLICE_X3Y142_CO6;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_D = CLBLM_R_X3Y142_SLICE_X3Y142_DO6;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_DMUX = CLBLM_R_X3Y142_SLICE_X3Y142_DO6;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_A = CLBLM_R_X3Y143_SLICE_X2Y143_AO6;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_B = CLBLM_R_X3Y143_SLICE_X2Y143_BO6;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_C = CLBLM_R_X3Y143_SLICE_X2Y143_CO6;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_D = CLBLM_R_X3Y143_SLICE_X2Y143_DO6;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_A = CLBLM_R_X3Y143_SLICE_X3Y143_AO6;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_B = CLBLM_R_X3Y143_SLICE_X3Y143_BO6;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_C = CLBLM_R_X3Y143_SLICE_X3Y143_CO6;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_D = CLBLM_R_X3Y143_SLICE_X3Y143_DO6;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_BMUX = CLBLM_R_X3Y143_SLICE_X3Y143_BO5;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_CMUX = CLBLM_R_X3Y143_SLICE_X3Y143_CO5;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_DMUX = CLBLM_R_X3Y143_SLICE_X3Y143_DO6;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_A = CLBLM_R_X3Y144_SLICE_X2Y144_AO6;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_B = CLBLM_R_X3Y144_SLICE_X2Y144_BO6;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_C = CLBLM_R_X3Y144_SLICE_X2Y144_CO6;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_D = CLBLM_R_X3Y144_SLICE_X2Y144_DO6;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_AMUX = CLBLM_R_X3Y144_SLICE_X2Y144_A5Q;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_BMUX = CLBLM_R_X3Y144_SLICE_X2Y144_BO5;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_A = CLBLM_R_X3Y144_SLICE_X3Y144_AO6;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_B = CLBLM_R_X3Y144_SLICE_X3Y144_BO6;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_C = CLBLM_R_X3Y144_SLICE_X3Y144_CO6;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_D = CLBLM_R_X3Y144_SLICE_X3Y144_DO6;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_AMUX = CLBLM_R_X3Y144_SLICE_X3Y144_A5Q;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_DMUX = CLBLM_R_X3Y144_SLICE_X3Y144_D5Q;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_A = CLBLM_R_X3Y145_SLICE_X2Y145_AO6;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_B = CLBLM_R_X3Y145_SLICE_X2Y145_BO6;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_C = CLBLM_R_X3Y145_SLICE_X2Y145_CO6;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_D = CLBLM_R_X3Y145_SLICE_X2Y145_DO6;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_BMUX = CLBLM_R_X3Y145_SLICE_X2Y145_B5Q;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_CMUX = CLBLM_R_X3Y145_SLICE_X2Y145_C5Q;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_A = CLBLM_R_X3Y145_SLICE_X3Y145_AO6;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_B = CLBLM_R_X3Y145_SLICE_X3Y145_BO6;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_C = CLBLM_R_X3Y145_SLICE_X3Y145_CO6;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_D = CLBLM_R_X3Y145_SLICE_X3Y145_DO6;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_AMUX = CLBLM_R_X3Y145_SLICE_X3Y145_A5Q;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_A = CLBLM_R_X3Y146_SLICE_X2Y146_AO6;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_B = CLBLM_R_X3Y146_SLICE_X2Y146_BO6;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_C = CLBLM_R_X3Y146_SLICE_X2Y146_CO6;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_D = CLBLM_R_X3Y146_SLICE_X2Y146_DO6;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_BMUX = CLBLM_R_X3Y146_SLICE_X2Y146_B5Q;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_CMUX = CLBLM_R_X3Y146_SLICE_X2Y146_C5Q;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_A = CLBLM_R_X3Y146_SLICE_X3Y146_AO6;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_B = CLBLM_R_X3Y146_SLICE_X3Y146_BO6;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_C = CLBLM_R_X3Y146_SLICE_X3Y146_CO6;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_D = CLBLM_R_X3Y146_SLICE_X3Y146_DO6;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_CMUX = CLBLM_R_X3Y146_SLICE_X3Y146_C5Q;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_A = CLBLM_R_X3Y147_SLICE_X2Y147_AO6;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_B = CLBLM_R_X3Y147_SLICE_X2Y147_BO6;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_C = CLBLM_R_X3Y147_SLICE_X2Y147_CO6;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_D = CLBLM_R_X3Y147_SLICE_X2Y147_DO6;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_CMUX = CLBLM_R_X3Y147_SLICE_X2Y147_C5Q;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_DMUX = CLBLM_R_X3Y147_SLICE_X2Y147_DO5;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_A = CLBLM_R_X3Y147_SLICE_X3Y147_AO6;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_B = CLBLM_R_X3Y147_SLICE_X3Y147_BO6;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_C = CLBLM_R_X3Y147_SLICE_X3Y147_CO6;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_D = CLBLM_R_X3Y147_SLICE_X3Y147_DO6;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_AMUX = CLBLM_R_X3Y147_SLICE_X3Y147_A5Q;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_BMUX = CLBLM_R_X3Y147_SLICE_X3Y147_B5Q;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_CMUX = CLBLM_R_X3Y147_SLICE_X3Y147_CO5;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_A = CLBLM_R_X3Y148_SLICE_X2Y148_AO6;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_B = CLBLM_R_X3Y148_SLICE_X2Y148_BO6;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_C = CLBLM_R_X3Y148_SLICE_X2Y148_CO6;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_D = CLBLM_R_X3Y148_SLICE_X2Y148_DO6;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_BMUX = CLBLM_R_X3Y148_SLICE_X2Y148_B5Q;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_CMUX = CLBLM_R_X3Y148_SLICE_X2Y148_C5Q;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_DMUX = CLBLM_R_X3Y148_SLICE_X2Y148_D5Q;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_A = CLBLM_R_X3Y148_SLICE_X3Y148_AO6;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_B = CLBLM_R_X3Y148_SLICE_X3Y148_BO6;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_C = CLBLM_R_X3Y148_SLICE_X3Y148_CO6;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_D = CLBLM_R_X3Y148_SLICE_X3Y148_DO6;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_AMUX = CLBLM_R_X3Y148_SLICE_X3Y148_A5Q;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_BMUX = CLBLM_R_X3Y148_SLICE_X3Y148_BO5;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_CMUX = CLBLM_R_X3Y148_SLICE_X3Y148_CO5;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_DMUX = CLBLM_R_X3Y148_SLICE_X3Y148_DO6;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_A = CLBLM_R_X3Y149_SLICE_X2Y149_AO6;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_B = CLBLM_R_X3Y149_SLICE_X2Y149_BO6;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_C = CLBLM_R_X3Y149_SLICE_X2Y149_CO6;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_D = CLBLM_R_X3Y149_SLICE_X2Y149_DO6;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_AMUX = CLBLM_R_X3Y149_SLICE_X2Y149_A5Q;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_A = CLBLM_R_X3Y149_SLICE_X3Y149_AO6;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_B = CLBLM_R_X3Y149_SLICE_X3Y149_BO6;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_C = CLBLM_R_X3Y149_SLICE_X3Y149_CO6;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_D = CLBLM_R_X3Y149_SLICE_X3Y149_DO6;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_A = CLBLM_R_X3Y150_SLICE_X2Y150_AO6;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_B = CLBLM_R_X3Y150_SLICE_X2Y150_BO6;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_C = CLBLM_R_X3Y150_SLICE_X2Y150_CO6;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_D = CLBLM_R_X3Y150_SLICE_X2Y150_DO6;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_BMUX = CLBLM_R_X3Y150_SLICE_X2Y150_B5Q;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_CMUX = CLBLM_R_X3Y150_SLICE_X2Y150_CO5;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_A = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_B = CLBLM_R_X3Y150_SLICE_X3Y150_BO6;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_C = CLBLM_R_X3Y150_SLICE_X3Y150_CO6;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_D = CLBLM_R_X3Y150_SLICE_X3Y150_DO6;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_A = CLBLM_R_X3Y151_SLICE_X2Y151_AO6;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_B = CLBLM_R_X3Y151_SLICE_X2Y151_BO6;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_C = CLBLM_R_X3Y151_SLICE_X2Y151_CO6;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_D = CLBLM_R_X3Y151_SLICE_X2Y151_DO6;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_AMUX = CLBLM_R_X3Y151_SLICE_X2Y151_A5Q;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_CMUX = CLBLM_R_X3Y151_SLICE_X2Y151_CO5;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_A = CLBLM_R_X3Y151_SLICE_X3Y151_AO6;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_B = CLBLM_R_X3Y151_SLICE_X3Y151_BO6;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_C = CLBLM_R_X3Y151_SLICE_X3Y151_CO6;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_D = CLBLM_R_X3Y151_SLICE_X3Y151_DO6;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_CMUX = CLBLM_R_X3Y151_SLICE_X3Y151_C5Q;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_DMUX = CLBLM_R_X3Y151_SLICE_X3Y151_D5Q;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_A = CLBLM_R_X3Y152_SLICE_X2Y152_AO6;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_B = CLBLM_R_X3Y152_SLICE_X2Y152_BO6;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_C = CLBLM_R_X3Y152_SLICE_X2Y152_CO6;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_D = CLBLM_R_X3Y152_SLICE_X2Y152_DO6;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_A = CLBLM_R_X3Y152_SLICE_X3Y152_AO6;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_B = CLBLM_R_X3Y152_SLICE_X3Y152_BO6;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_C = CLBLM_R_X3Y152_SLICE_X3Y152_CO6;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_D = CLBLM_R_X3Y152_SLICE_X3Y152_DO6;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_AMUX = CLBLM_R_X3Y152_SLICE_X3Y152_A5Q;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_CMUX = CLBLM_R_X3Y152_SLICE_X3Y152_CO6;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_A = CLBLM_R_X3Y153_SLICE_X2Y153_AO6;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_B = CLBLM_R_X3Y153_SLICE_X2Y153_BO6;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_C = CLBLM_R_X3Y153_SLICE_X2Y153_CO6;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_D = CLBLM_R_X3Y153_SLICE_X2Y153_DO6;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_AMUX = CLBLM_R_X3Y153_SLICE_X2Y153_AO5;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_A = CLBLM_R_X3Y153_SLICE_X3Y153_AO6;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_B = CLBLM_R_X3Y153_SLICE_X3Y153_BO6;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_C = CLBLM_R_X3Y153_SLICE_X3Y153_CO6;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_D = CLBLM_R_X3Y153_SLICE_X3Y153_DO6;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_AMUX = CLBLM_R_X3Y153_SLICE_X3Y153_A5Q;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_BMUX = CLBLM_R_X3Y153_SLICE_X3Y153_BO5;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_CMUX = CLBLM_R_X3Y153_SLICE_X3Y153_CO5;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_A = CLBLM_R_X3Y154_SLICE_X2Y154_AO6;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_B = CLBLM_R_X3Y154_SLICE_X2Y154_BO6;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_C = CLBLM_R_X3Y154_SLICE_X2Y154_CO6;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_D = CLBLM_R_X3Y154_SLICE_X2Y154_DO6;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_A = CLBLM_R_X3Y154_SLICE_X3Y154_AO6;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_B = CLBLM_R_X3Y154_SLICE_X3Y154_BO6;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_C = CLBLM_R_X3Y154_SLICE_X3Y154_CO6;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_D = CLBLM_R_X3Y154_SLICE_X3Y154_DO6;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_A = CLBLM_R_X5Y140_SLICE_X6Y140_AO6;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_B = CLBLM_R_X5Y140_SLICE_X6Y140_BO6;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_C = CLBLM_R_X5Y140_SLICE_X6Y140_CO6;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_D = CLBLM_R_X5Y140_SLICE_X6Y140_DO6;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_A = CLBLM_R_X5Y140_SLICE_X7Y140_AO6;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_B = CLBLM_R_X5Y140_SLICE_X7Y140_BO6;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_C = CLBLM_R_X5Y140_SLICE_X7Y140_CO6;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_D = CLBLM_R_X5Y140_SLICE_X7Y140_DO6;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_BMUX = CLBLM_R_X5Y140_SLICE_X7Y140_B5Q;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_A = CLBLM_R_X5Y141_SLICE_X6Y141_AO6;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_B = CLBLM_R_X5Y141_SLICE_X6Y141_BO6;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_C = CLBLM_R_X5Y141_SLICE_X6Y141_CO6;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_D = CLBLM_R_X5Y141_SLICE_X6Y141_DO6;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_A = CLBLM_R_X5Y141_SLICE_X7Y141_AO6;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_B = CLBLM_R_X5Y141_SLICE_X7Y141_BO6;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_C = CLBLM_R_X5Y141_SLICE_X7Y141_CO6;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_D = CLBLM_R_X5Y141_SLICE_X7Y141_DO6;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_AMUX = CLBLM_R_X5Y141_SLICE_X7Y141_A5Q;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_A = CLBLM_R_X5Y142_SLICE_X6Y142_AO6;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_B = CLBLM_R_X5Y142_SLICE_X6Y142_BO6;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_C = CLBLM_R_X5Y142_SLICE_X6Y142_CO6;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_D = CLBLM_R_X5Y142_SLICE_X6Y142_DO6;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_CMUX = CLBLM_R_X5Y142_SLICE_X6Y142_C5Q;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_A = CLBLM_R_X5Y142_SLICE_X7Y142_AO6;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_B = CLBLM_R_X5Y142_SLICE_X7Y142_BO6;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_C = CLBLM_R_X5Y142_SLICE_X7Y142_CO6;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_D = CLBLM_R_X5Y142_SLICE_X7Y142_DO6;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_AMUX = CLBLM_R_X5Y142_SLICE_X7Y142_AO5;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_BMUX = CLBLM_R_X5Y142_SLICE_X7Y142_B5Q;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_CMUX = CLBLM_R_X5Y142_SLICE_X7Y142_C5Q;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_A = CLBLM_R_X5Y143_SLICE_X6Y143_AO6;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_B = CLBLM_R_X5Y143_SLICE_X6Y143_BO6;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_C = CLBLM_R_X5Y143_SLICE_X6Y143_CO6;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_D = CLBLM_R_X5Y143_SLICE_X6Y143_DO6;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_DMUX = CLBLM_R_X5Y143_SLICE_X6Y143_D5Q;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_A = CLBLM_R_X5Y143_SLICE_X7Y143_AO6;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_B = CLBLM_R_X5Y143_SLICE_X7Y143_BO6;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_C = CLBLM_R_X5Y143_SLICE_X7Y143_CO6;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_D = CLBLM_R_X5Y143_SLICE_X7Y143_DO6;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_A = CLBLM_R_X5Y144_SLICE_X6Y144_AO6;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_B = CLBLM_R_X5Y144_SLICE_X6Y144_BO6;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_C = CLBLM_R_X5Y144_SLICE_X6Y144_CO6;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_D = CLBLM_R_X5Y144_SLICE_X6Y144_DO6;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_BMUX = CLBLM_R_X5Y144_SLICE_X6Y144_B5Q;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_CMUX = CLBLM_R_X5Y144_SLICE_X6Y144_C5Q;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_DMUX = CLBLM_R_X5Y144_SLICE_X6Y144_D5Q;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_A = CLBLM_R_X5Y144_SLICE_X7Y144_AO6;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_B = CLBLM_R_X5Y144_SLICE_X7Y144_BO6;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_C = CLBLM_R_X5Y144_SLICE_X7Y144_CO6;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_D = CLBLM_R_X5Y144_SLICE_X7Y144_DO6;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_A = CLBLM_R_X5Y145_SLICE_X6Y145_AO6;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_B = CLBLM_R_X5Y145_SLICE_X6Y145_BO6;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_C = CLBLM_R_X5Y145_SLICE_X6Y145_CO6;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_D = CLBLM_R_X5Y145_SLICE_X6Y145_DO6;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_BMUX = CLBLM_R_X5Y145_SLICE_X6Y145_B5Q;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_A = CLBLM_R_X5Y145_SLICE_X7Y145_AO6;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_B = CLBLM_R_X5Y145_SLICE_X7Y145_BO6;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_C = CLBLM_R_X5Y145_SLICE_X7Y145_CO6;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_D = CLBLM_R_X5Y145_SLICE_X7Y145_DO6;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_AMUX = CLBLM_R_X5Y145_SLICE_X7Y145_A5Q;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_BMUX = CLBLM_R_X5Y145_SLICE_X7Y145_BO5;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_A = CLBLM_R_X5Y146_SLICE_X6Y146_AO6;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_B = CLBLM_R_X5Y146_SLICE_X6Y146_BO6;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_C = CLBLM_R_X5Y146_SLICE_X6Y146_CO6;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_D = CLBLM_R_X5Y146_SLICE_X6Y146_DO6;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_BMUX = CLBLM_R_X5Y146_SLICE_X6Y146_B5Q;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_CMUX = CLBLM_R_X5Y146_SLICE_X6Y146_CO6;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_A = CLBLM_R_X5Y146_SLICE_X7Y146_AO6;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_B = CLBLM_R_X5Y146_SLICE_X7Y146_BO6;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_C = CLBLM_R_X5Y146_SLICE_X7Y146_CO6;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_D = CLBLM_R_X5Y146_SLICE_X7Y146_DO6;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_BMUX = CLBLM_R_X5Y146_SLICE_X7Y146_B5Q;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_A = CLBLM_R_X5Y147_SLICE_X6Y147_AO6;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_B = CLBLM_R_X5Y147_SLICE_X6Y147_BO6;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_C = CLBLM_R_X5Y147_SLICE_X6Y147_CO6;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_D = CLBLM_R_X5Y147_SLICE_X6Y147_DO6;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_BMUX = CLBLM_R_X5Y147_SLICE_X6Y147_B5Q;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_A = CLBLM_R_X5Y147_SLICE_X7Y147_AO6;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_B = CLBLM_R_X5Y147_SLICE_X7Y147_BO6;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_C = CLBLM_R_X5Y147_SLICE_X7Y147_CO6;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_D = CLBLM_R_X5Y147_SLICE_X7Y147_DO6;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_AMUX = CLBLM_R_X5Y147_SLICE_X7Y147_A5Q;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_BMUX = CLBLM_R_X5Y147_SLICE_X7Y147_B5Q;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_CMUX = CLBLM_R_X5Y147_SLICE_X7Y147_C5Q;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_A = CLBLM_R_X5Y148_SLICE_X6Y148_AO6;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_B = CLBLM_R_X5Y148_SLICE_X6Y148_BO6;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_C = CLBLM_R_X5Y148_SLICE_X6Y148_CO6;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_D = CLBLM_R_X5Y148_SLICE_X6Y148_DO6;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_AMUX = CLBLM_R_X5Y148_SLICE_X6Y148_AO5;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_BMUX = CLBLM_R_X5Y148_SLICE_X6Y148_B5Q;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_CMUX = CLBLM_R_X5Y148_SLICE_X6Y148_CO5;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_A = CLBLM_R_X5Y148_SLICE_X7Y148_AO6;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_B = CLBLM_R_X5Y148_SLICE_X7Y148_BO6;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_C = CLBLM_R_X5Y148_SLICE_X7Y148_CO6;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_D = CLBLM_R_X5Y148_SLICE_X7Y148_DO6;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_A = CLBLM_R_X5Y149_SLICE_X6Y149_AO6;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_B = CLBLM_R_X5Y149_SLICE_X6Y149_BO6;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_C = CLBLM_R_X5Y149_SLICE_X6Y149_CO6;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_D = CLBLM_R_X5Y149_SLICE_X6Y149_DO6;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_AMUX = CLBLM_R_X5Y149_SLICE_X6Y149_A5Q;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_DMUX = CLBLM_R_X5Y149_SLICE_X6Y149_D5Q;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_A = CLBLM_R_X5Y149_SLICE_X7Y149_AO6;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_B = CLBLM_R_X5Y149_SLICE_X7Y149_BO6;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_C = CLBLM_R_X5Y149_SLICE_X7Y149_CO6;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_D = CLBLM_R_X5Y149_SLICE_X7Y149_DO6;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_BMUX = CLBLM_R_X5Y149_SLICE_X7Y149_B5Q;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_CMUX = CLBLM_R_X5Y149_SLICE_X7Y149_C5Q;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_DMUX = CLBLM_R_X5Y149_SLICE_X7Y149_D5Q;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_A = CLBLM_R_X5Y150_SLICE_X6Y150_AO6;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_B = CLBLM_R_X5Y150_SLICE_X6Y150_BO6;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_C = CLBLM_R_X5Y150_SLICE_X6Y150_CO6;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_D = CLBLM_R_X5Y150_SLICE_X6Y150_DO6;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_AMUX = CLBLM_R_X5Y150_SLICE_X6Y150_A5Q;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_CMUX = CLBLM_R_X5Y150_SLICE_X6Y150_C5Q;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_A = CLBLM_R_X5Y150_SLICE_X7Y150_AO6;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_B = CLBLM_R_X5Y150_SLICE_X7Y150_BO6;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_C = CLBLM_R_X5Y150_SLICE_X7Y150_CO6;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_D = CLBLM_R_X5Y150_SLICE_X7Y150_DO6;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_AMUX = CLBLM_R_X5Y150_SLICE_X7Y150_A5Q;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_BMUX = CLBLM_R_X5Y150_SLICE_X7Y150_BO5;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_A = CLBLM_R_X5Y151_SLICE_X6Y151_AO6;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_B = CLBLM_R_X5Y151_SLICE_X6Y151_BO6;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_C = CLBLM_R_X5Y151_SLICE_X6Y151_CO6;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_D = CLBLM_R_X5Y151_SLICE_X6Y151_DO6;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_AMUX = CLBLM_R_X5Y151_SLICE_X6Y151_A5Q;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_BMUX = CLBLM_R_X5Y151_SLICE_X6Y151_B5Q;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_DMUX = CLBLM_R_X5Y151_SLICE_X6Y151_D5Q;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_A = CLBLM_R_X5Y151_SLICE_X7Y151_AO6;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_B = CLBLM_R_X5Y151_SLICE_X7Y151_BO6;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_C = CLBLM_R_X5Y151_SLICE_X7Y151_CO6;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_D = CLBLM_R_X5Y151_SLICE_X7Y151_DO6;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_AMUX = CLBLM_R_X5Y151_SLICE_X7Y151_A5Q;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_BMUX = CLBLM_R_X5Y151_SLICE_X7Y151_BO5;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_A = CLBLM_R_X5Y152_SLICE_X6Y152_AO6;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_B = CLBLM_R_X5Y152_SLICE_X6Y152_BO6;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_C = CLBLM_R_X5Y152_SLICE_X6Y152_CO6;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_D = CLBLM_R_X5Y152_SLICE_X6Y152_DO6;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_AMUX = CLBLM_R_X5Y152_SLICE_X6Y152_A5Q;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_BMUX = CLBLM_R_X5Y152_SLICE_X6Y152_B5Q;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_CMUX = CLBLM_R_X5Y152_SLICE_X6Y152_C5Q;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_A = CLBLM_R_X5Y152_SLICE_X7Y152_AO6;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_B = CLBLM_R_X5Y152_SLICE_X7Y152_BO6;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_C = CLBLM_R_X5Y152_SLICE_X7Y152_CO6;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_D = CLBLM_R_X5Y152_SLICE_X7Y152_DO6;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_DMUX = CLBLM_R_X5Y152_SLICE_X7Y152_D5Q;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_A = CLBLM_R_X5Y153_SLICE_X6Y153_AO6;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_B = CLBLM_R_X5Y153_SLICE_X6Y153_BO6;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_C = CLBLM_R_X5Y153_SLICE_X6Y153_CO6;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_D = CLBLM_R_X5Y153_SLICE_X6Y153_DO6;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_A = CLBLM_R_X5Y153_SLICE_X7Y153_AO6;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_B = CLBLM_R_X5Y153_SLICE_X7Y153_BO6;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_C = CLBLM_R_X5Y153_SLICE_X7Y153_CO6;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_D = CLBLM_R_X5Y153_SLICE_X7Y153_DO6;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_AMUX = CLBLM_R_X5Y153_SLICE_X7Y153_A5Q;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_A = CLBLM_R_X5Y154_SLICE_X6Y154_AO6;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_B = CLBLM_R_X5Y154_SLICE_X6Y154_BO6;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_C = CLBLM_R_X5Y154_SLICE_X6Y154_CO6;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_D = CLBLM_R_X5Y154_SLICE_X6Y154_DO6;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_A = CLBLM_R_X5Y154_SLICE_X7Y154_AO6;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_B = CLBLM_R_X5Y154_SLICE_X7Y154_BO6;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_C = CLBLM_R_X5Y154_SLICE_X7Y154_CO6;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_D = CLBLM_R_X5Y154_SLICE_X7Y154_DO6;
  assign CLBLM_R_X5Y159_SLICE_X6Y159_A = CLBLM_R_X5Y159_SLICE_X6Y159_AO6;
  assign CLBLM_R_X5Y159_SLICE_X6Y159_B = CLBLM_R_X5Y159_SLICE_X6Y159_BO6;
  assign CLBLM_R_X5Y159_SLICE_X6Y159_C = CLBLM_R_X5Y159_SLICE_X6Y159_CO6;
  assign CLBLM_R_X5Y159_SLICE_X6Y159_D = CLBLM_R_X5Y159_SLICE_X6Y159_DO6;
  assign CLBLM_R_X5Y159_SLICE_X7Y159_A = CLBLM_R_X5Y159_SLICE_X7Y159_AO6;
  assign CLBLM_R_X5Y159_SLICE_X7Y159_B = CLBLM_R_X5Y159_SLICE_X7Y159_BO6;
  assign CLBLM_R_X5Y159_SLICE_X7Y159_C = CLBLM_R_X5Y159_SLICE_X7Y159_CO6;
  assign CLBLM_R_X5Y159_SLICE_X7Y159_D = CLBLM_R_X5Y159_SLICE_X7Y159_DO6;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_A = CLBLM_R_X7Y141_SLICE_X8Y141_AO6;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_B = CLBLM_R_X7Y141_SLICE_X8Y141_BO6;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_C = CLBLM_R_X7Y141_SLICE_X8Y141_CO6;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_D = CLBLM_R_X7Y141_SLICE_X8Y141_DO6;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_A = CLBLM_R_X7Y141_SLICE_X9Y141_AO6;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_B = CLBLM_R_X7Y141_SLICE_X9Y141_BO6;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_C = CLBLM_R_X7Y141_SLICE_X9Y141_CO6;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_D = CLBLM_R_X7Y141_SLICE_X9Y141_DO6;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_A = CLBLM_R_X7Y142_SLICE_X8Y142_AO6;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_B = CLBLM_R_X7Y142_SLICE_X8Y142_BO6;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_C = CLBLM_R_X7Y142_SLICE_X8Y142_CO6;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_D = CLBLM_R_X7Y142_SLICE_X8Y142_DO6;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_AMUX = CLBLM_R_X7Y142_SLICE_X8Y142_A5Q;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_BMUX = CLBLM_R_X7Y142_SLICE_X8Y142_B5Q;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_A = CLBLM_R_X7Y142_SLICE_X9Y142_AO6;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_B = CLBLM_R_X7Y142_SLICE_X9Y142_BO6;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_C = CLBLM_R_X7Y142_SLICE_X9Y142_CO6;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_D = CLBLM_R_X7Y142_SLICE_X9Y142_DO6;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_AMUX = CLBLM_R_X7Y142_SLICE_X9Y142_A5Q;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_DMUX = CLBLM_R_X7Y142_SLICE_X9Y142_D5Q;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_A = CLBLM_R_X7Y143_SLICE_X8Y143_AO6;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_B = CLBLM_R_X7Y143_SLICE_X8Y143_BO6;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_C = CLBLM_R_X7Y143_SLICE_X8Y143_CO6;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_D = CLBLM_R_X7Y143_SLICE_X8Y143_DO6;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_A = CLBLM_R_X7Y143_SLICE_X9Y143_AO6;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_B = CLBLM_R_X7Y143_SLICE_X9Y143_BO6;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_C = CLBLM_R_X7Y143_SLICE_X9Y143_CO6;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_D = CLBLM_R_X7Y143_SLICE_X9Y143_DO6;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_A = CLBLM_R_X7Y144_SLICE_X8Y144_AO6;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_B = CLBLM_R_X7Y144_SLICE_X8Y144_BO6;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_C = CLBLM_R_X7Y144_SLICE_X8Y144_CO6;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_D = CLBLM_R_X7Y144_SLICE_X8Y144_DO6;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_AMUX = CLBLM_R_X7Y144_SLICE_X8Y144_A5Q;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_A = CLBLM_R_X7Y144_SLICE_X9Y144_AO6;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_B = CLBLM_R_X7Y144_SLICE_X9Y144_BO6;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_C = CLBLM_R_X7Y144_SLICE_X9Y144_CO6;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_D = CLBLM_R_X7Y144_SLICE_X9Y144_DO6;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_AMUX = CLBLM_R_X7Y144_SLICE_X9Y144_A5Q;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_BMUX = CLBLM_R_X7Y144_SLICE_X9Y144_B5Q;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_CMUX = CLBLM_R_X7Y144_SLICE_X9Y144_C5Q;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_DMUX = CLBLM_R_X7Y144_SLICE_X9Y144_D5Q;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_A = CLBLM_R_X7Y145_SLICE_X8Y145_AO6;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_B = CLBLM_R_X7Y145_SLICE_X8Y145_BO6;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_C = CLBLM_R_X7Y145_SLICE_X8Y145_CO6;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_D = CLBLM_R_X7Y145_SLICE_X8Y145_DO6;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_BMUX = CLBLM_R_X7Y145_SLICE_X8Y145_B5Q;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_CMUX = CLBLM_R_X7Y145_SLICE_X8Y145_C5Q;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_A = CLBLM_R_X7Y145_SLICE_X9Y145_AO6;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_B = CLBLM_R_X7Y145_SLICE_X9Y145_BO6;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_C = CLBLM_R_X7Y145_SLICE_X9Y145_CO6;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_D = CLBLM_R_X7Y145_SLICE_X9Y145_DO6;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_A = CLBLM_R_X7Y146_SLICE_X8Y146_AO6;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_B = CLBLM_R_X7Y146_SLICE_X8Y146_BO6;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_C = CLBLM_R_X7Y146_SLICE_X8Y146_CO6;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_D = CLBLM_R_X7Y146_SLICE_X8Y146_DO6;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_AMUX = CLBLM_R_X7Y146_SLICE_X8Y146_AO5;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_CMUX = CLBLM_R_X7Y146_SLICE_X8Y146_CO6;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_A = CLBLM_R_X7Y146_SLICE_X9Y146_AO6;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_B = CLBLM_R_X7Y146_SLICE_X9Y146_BO6;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_C = CLBLM_R_X7Y146_SLICE_X9Y146_CO6;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_D = CLBLM_R_X7Y146_SLICE_X9Y146_DO6;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_AMUX = CLBLM_R_X7Y146_SLICE_X9Y146_AO5;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_BMUX = CLBLM_R_X7Y146_SLICE_X9Y146_B5Q;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_A = CLBLM_R_X7Y147_SLICE_X8Y147_AO6;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_B = CLBLM_R_X7Y147_SLICE_X8Y147_BO6;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_C = CLBLM_R_X7Y147_SLICE_X8Y147_CO6;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_D = CLBLM_R_X7Y147_SLICE_X8Y147_DO6;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_DMUX = CLBLM_R_X7Y147_SLICE_X8Y147_D5Q;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_A = CLBLM_R_X7Y147_SLICE_X9Y147_AO6;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_B = CLBLM_R_X7Y147_SLICE_X9Y147_BO6;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_C = CLBLM_R_X7Y147_SLICE_X9Y147_CO6;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_D = CLBLM_R_X7Y147_SLICE_X9Y147_DO6;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_CMUX = CLBLM_R_X7Y147_SLICE_X9Y147_C5Q;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_DMUX = CLBLM_R_X7Y147_SLICE_X9Y147_DO5;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_A = CLBLM_R_X7Y148_SLICE_X8Y148_AO6;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_B = CLBLM_R_X7Y148_SLICE_X8Y148_BO6;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_C = CLBLM_R_X7Y148_SLICE_X8Y148_CO6;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_D = CLBLM_R_X7Y148_SLICE_X8Y148_DO6;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_BMUX = CLBLM_R_X7Y148_SLICE_X8Y148_BO5;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_A = CLBLM_R_X7Y148_SLICE_X9Y148_AO6;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_B = CLBLM_R_X7Y148_SLICE_X9Y148_BO6;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_C = CLBLM_R_X7Y148_SLICE_X9Y148_CO6;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_D = CLBLM_R_X7Y148_SLICE_X9Y148_DO6;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_AMUX = CLBLM_R_X7Y148_SLICE_X9Y148_AO5;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_BMUX = CLBLM_R_X7Y148_SLICE_X9Y148_B5Q;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_CMUX = CLBLM_R_X7Y148_SLICE_X9Y148_C5Q;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_A = CLBLM_R_X7Y149_SLICE_X8Y149_AO6;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_B = CLBLM_R_X7Y149_SLICE_X8Y149_BO6;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_C = CLBLM_R_X7Y149_SLICE_X8Y149_CO6;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_D = CLBLM_R_X7Y149_SLICE_X8Y149_DO6;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_A = CLBLM_R_X7Y149_SLICE_X9Y149_AO6;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_B = CLBLM_R_X7Y149_SLICE_X9Y149_BO6;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_C = CLBLM_R_X7Y149_SLICE_X9Y149_CO6;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_D = CLBLM_R_X7Y149_SLICE_X9Y149_DO6;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_AMUX = CLBLM_R_X7Y149_SLICE_X9Y149_AO5;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_BMUX = CLBLM_R_X7Y149_SLICE_X9Y149_BO5;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_CMUX = CLBLM_R_X7Y149_SLICE_X9Y149_C5Q;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_A = CLBLM_R_X7Y150_SLICE_X8Y150_AO6;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_B = CLBLM_R_X7Y150_SLICE_X8Y150_BO6;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_C = CLBLM_R_X7Y150_SLICE_X8Y150_CO6;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_D = CLBLM_R_X7Y150_SLICE_X8Y150_DO6;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_CMUX = CLBLM_R_X7Y150_SLICE_X8Y150_C5Q;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_DMUX = CLBLM_R_X7Y150_SLICE_X8Y150_D5Q;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_A = CLBLM_R_X7Y150_SLICE_X9Y150_AO6;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_B = CLBLM_R_X7Y150_SLICE_X9Y150_BO6;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_C = CLBLM_R_X7Y150_SLICE_X9Y150_CO6;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_D = CLBLM_R_X7Y150_SLICE_X9Y150_DO6;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_BMUX = CLBLM_R_X7Y150_SLICE_X9Y150_B5Q;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_CMUX = CLBLM_R_X7Y150_SLICE_X9Y150_C5Q;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_A = CLBLM_R_X7Y151_SLICE_X8Y151_AO6;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_B = CLBLM_R_X7Y151_SLICE_X8Y151_BO6;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_C = CLBLM_R_X7Y151_SLICE_X8Y151_CO6;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_D = CLBLM_R_X7Y151_SLICE_X8Y151_DO6;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_CMUX = CLBLM_R_X7Y151_SLICE_X8Y151_C5Q;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_DMUX = CLBLM_R_X7Y151_SLICE_X8Y151_DO5;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_A = CLBLM_R_X7Y151_SLICE_X9Y151_AO6;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_B = CLBLM_R_X7Y151_SLICE_X9Y151_BO6;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_C = CLBLM_R_X7Y151_SLICE_X9Y151_CO6;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_D = CLBLM_R_X7Y151_SLICE_X9Y151_DO6;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_A = CLBLM_R_X7Y152_SLICE_X8Y152_AO6;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_B = CLBLM_R_X7Y152_SLICE_X8Y152_BO6;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_C = CLBLM_R_X7Y152_SLICE_X8Y152_CO6;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_D = CLBLM_R_X7Y152_SLICE_X8Y152_DO6;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_A = CLBLM_R_X7Y152_SLICE_X9Y152_AO6;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_B = CLBLM_R_X7Y152_SLICE_X9Y152_BO6;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_C = CLBLM_R_X7Y152_SLICE_X9Y152_CO6;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_D = CLBLM_R_X7Y152_SLICE_X9Y152_DO6;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_CMUX = CLBLM_R_X7Y152_SLICE_X9Y152_C5Q;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_DMUX = CLBLM_R_X7Y152_SLICE_X9Y152_D5Q;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_A = CLBLM_R_X7Y153_SLICE_X8Y153_AO6;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_B = CLBLM_R_X7Y153_SLICE_X8Y153_BO6;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_C = CLBLM_R_X7Y153_SLICE_X8Y153_CO6;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_D = CLBLM_R_X7Y153_SLICE_X8Y153_DO6;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_BMUX = CLBLM_R_X7Y153_SLICE_X8Y153_BO5;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_CMUX = CLBLM_R_X7Y153_SLICE_X8Y153_CO5;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_DMUX = CLBLM_R_X7Y153_SLICE_X8Y153_DO5;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_A = CLBLM_R_X7Y153_SLICE_X9Y153_AO6;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_B = CLBLM_R_X7Y153_SLICE_X9Y153_BO6;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_C = CLBLM_R_X7Y153_SLICE_X9Y153_CO6;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_D = CLBLM_R_X7Y153_SLICE_X9Y153_DO6;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_AMUX = CLBLM_R_X7Y153_SLICE_X9Y153_A5Q;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_DMUX = CLBLM_R_X7Y153_SLICE_X9Y153_DO5;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_A = CLBLM_R_X7Y154_SLICE_X8Y154_AO6;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_B = CLBLM_R_X7Y154_SLICE_X8Y154_BO6;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_C = CLBLM_R_X7Y154_SLICE_X8Y154_CO6;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_D = CLBLM_R_X7Y154_SLICE_X8Y154_DO6;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_DMUX = CLBLM_R_X7Y154_SLICE_X8Y154_DO5;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_A = CLBLM_R_X7Y154_SLICE_X9Y154_AO6;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_B = CLBLM_R_X7Y154_SLICE_X9Y154_BO6;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_C = CLBLM_R_X7Y154_SLICE_X9Y154_CO6;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_D = CLBLM_R_X7Y154_SLICE_X9Y154_DO6;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_AMUX = CLBLM_R_X7Y154_SLICE_X9Y154_AO5;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_A = CLBLM_R_X7Y155_SLICE_X8Y155_AO6;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_B = CLBLM_R_X7Y155_SLICE_X8Y155_BO6;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_C = CLBLM_R_X7Y155_SLICE_X8Y155_CO6;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_D = CLBLM_R_X7Y155_SLICE_X8Y155_DO6;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_A = CLBLM_R_X7Y155_SLICE_X9Y155_AO6;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_B = CLBLM_R_X7Y155_SLICE_X9Y155_BO6;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_C = CLBLM_R_X7Y155_SLICE_X9Y155_CO6;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_D = CLBLM_R_X7Y155_SLICE_X9Y155_DO6;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_AMUX = CLBLM_R_X7Y155_SLICE_X9Y155_AO5;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_A = CLBLM_R_X11Y142_SLICE_X14Y142_AO6;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_B = CLBLM_R_X11Y142_SLICE_X14Y142_BO6;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_C = CLBLM_R_X11Y142_SLICE_X14Y142_CO6;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_D = CLBLM_R_X11Y142_SLICE_X14Y142_DO6;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_BMUX = CLBLM_R_X11Y142_SLICE_X14Y142_BO5;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_CMUX = CLBLM_R_X11Y142_SLICE_X14Y142_CO5;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_A = CLBLM_R_X11Y142_SLICE_X15Y142_AO6;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_B = CLBLM_R_X11Y142_SLICE_X15Y142_BO6;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_C = CLBLM_R_X11Y142_SLICE_X15Y142_CO6;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_D = CLBLM_R_X11Y142_SLICE_X15Y142_DO6;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_A = CLBLM_R_X11Y143_SLICE_X14Y143_AO6;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_B = CLBLM_R_X11Y143_SLICE_X14Y143_BO6;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_C = CLBLM_R_X11Y143_SLICE_X14Y143_CO6;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_D = CLBLM_R_X11Y143_SLICE_X14Y143_DO6;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_BMUX = CLBLM_R_X11Y143_SLICE_X14Y143_BO5;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_CMUX = CLBLM_R_X11Y143_SLICE_X14Y143_CO5;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_A = CLBLM_R_X11Y143_SLICE_X15Y143_AO6;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_B = CLBLM_R_X11Y143_SLICE_X15Y143_BO6;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_C = CLBLM_R_X11Y143_SLICE_X15Y143_CO6;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_D = CLBLM_R_X11Y143_SLICE_X15Y143_DO6;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_A = CLBLM_R_X11Y144_SLICE_X14Y144_AO6;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_B = CLBLM_R_X11Y144_SLICE_X14Y144_BO6;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_C = CLBLM_R_X11Y144_SLICE_X14Y144_CO6;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_D = CLBLM_R_X11Y144_SLICE_X14Y144_DO6;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_A = CLBLM_R_X11Y144_SLICE_X15Y144_AO6;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_B = CLBLM_R_X11Y144_SLICE_X15Y144_BO6;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_C = CLBLM_R_X11Y144_SLICE_X15Y144_CO6;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_D = CLBLM_R_X11Y144_SLICE_X15Y144_DO6;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_AMUX = CLBLM_R_X11Y144_SLICE_X15Y144_AO5;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_CMUX = CLBLM_R_X11Y144_SLICE_X15Y144_CO6;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_A = CLBLM_R_X11Y145_SLICE_X14Y145_AO6;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_B = CLBLM_R_X11Y145_SLICE_X14Y145_BO6;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_C = CLBLM_R_X11Y145_SLICE_X14Y145_CO6;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_D = CLBLM_R_X11Y145_SLICE_X14Y145_DO6;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_AMUX = CLBLM_R_X11Y145_SLICE_X14Y145_AO5;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_BMUX = CLBLM_R_X11Y145_SLICE_X14Y145_BO5;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_A = CLBLM_R_X11Y145_SLICE_X15Y145_AO6;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_B = CLBLM_R_X11Y145_SLICE_X15Y145_BO6;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_C = CLBLM_R_X11Y145_SLICE_X15Y145_CO6;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_D = CLBLM_R_X11Y145_SLICE_X15Y145_DO6;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_AMUX = CLBLM_R_X11Y145_SLICE_X15Y145_AO5;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_BMUX = CLBLM_R_X11Y145_SLICE_X15Y145_BO5;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_A = CLBLM_R_X11Y146_SLICE_X14Y146_AO6;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_B = CLBLM_R_X11Y146_SLICE_X14Y146_BO6;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_C = CLBLM_R_X11Y146_SLICE_X14Y146_CO6;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_D = CLBLM_R_X11Y146_SLICE_X14Y146_DO6;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_AMUX = CLBLM_R_X11Y146_SLICE_X14Y146_AO5;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_A = CLBLM_R_X11Y146_SLICE_X15Y146_AO6;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_B = CLBLM_R_X11Y146_SLICE_X15Y146_BO6;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_C = CLBLM_R_X11Y146_SLICE_X15Y146_CO6;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_D = CLBLM_R_X11Y146_SLICE_X15Y146_DO6;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_BMUX = CLBLM_R_X11Y146_SLICE_X15Y146_BO5;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_CMUX = CLBLM_R_X11Y146_SLICE_X15Y146_CO5;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_A = CLBLM_R_X11Y147_SLICE_X14Y147_AO6;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_B = CLBLM_R_X11Y147_SLICE_X14Y147_BO6;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_C = CLBLM_R_X11Y147_SLICE_X14Y147_CO6;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_D = CLBLM_R_X11Y147_SLICE_X14Y147_DO6;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_AMUX = CLBLM_R_X11Y147_SLICE_X14Y147_A5Q;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_A = CLBLM_R_X11Y147_SLICE_X15Y147_AO6;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_B = CLBLM_R_X11Y147_SLICE_X15Y147_BO6;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_C = CLBLM_R_X11Y147_SLICE_X15Y147_CO6;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_D = CLBLM_R_X11Y147_SLICE_X15Y147_DO6;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_CMUX = CLBLM_R_X11Y147_SLICE_X15Y147_CO6;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_A = CLBLM_R_X11Y148_SLICE_X14Y148_AO6;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_B = CLBLM_R_X11Y148_SLICE_X14Y148_BO6;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_C = CLBLM_R_X11Y148_SLICE_X14Y148_CO6;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_D = CLBLM_R_X11Y148_SLICE_X14Y148_DO6;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_A = CLBLM_R_X11Y148_SLICE_X15Y148_AO6;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_B = CLBLM_R_X11Y148_SLICE_X15Y148_BO6;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_C = CLBLM_R_X11Y148_SLICE_X15Y148_CO6;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_D = CLBLM_R_X11Y148_SLICE_X15Y148_DO6;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_AMUX = CLBLM_R_X11Y148_SLICE_X15Y148_AO6;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_A = CLBLM_R_X11Y149_SLICE_X14Y149_AO6;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_B = CLBLM_R_X11Y149_SLICE_X14Y149_BO6;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_C = CLBLM_R_X11Y149_SLICE_X14Y149_CO6;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_D = CLBLM_R_X11Y149_SLICE_X14Y149_DO6;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_AMUX = CLBLM_R_X11Y149_SLICE_X14Y149_AO5;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_BMUX = CLBLM_R_X11Y149_SLICE_X14Y149_BO5;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_A = CLBLM_R_X11Y149_SLICE_X15Y149_AO6;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_B = CLBLM_R_X11Y149_SLICE_X15Y149_BO6;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_C = CLBLM_R_X11Y149_SLICE_X15Y149_CO6;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_D = CLBLM_R_X11Y149_SLICE_X15Y149_DO6;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_DMUX = CLBLM_R_X11Y149_SLICE_X15Y149_DO5;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_A = CLBLM_R_X11Y150_SLICE_X14Y150_AO6;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_B = CLBLM_R_X11Y150_SLICE_X14Y150_BO6;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_C = CLBLM_R_X11Y150_SLICE_X14Y150_CO6;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_D = CLBLM_R_X11Y150_SLICE_X14Y150_DO6;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_BMUX = CLBLM_R_X11Y150_SLICE_X14Y150_BO5;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_A = CLBLM_R_X11Y150_SLICE_X15Y150_AO6;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_B = CLBLM_R_X11Y150_SLICE_X15Y150_BO6;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_C = CLBLM_R_X11Y150_SLICE_X15Y150_CO6;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_D = CLBLM_R_X11Y150_SLICE_X15Y150_DO6;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_A = CLBLM_R_X11Y151_SLICE_X14Y151_AO6;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_B = CLBLM_R_X11Y151_SLICE_X14Y151_BO6;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_C = CLBLM_R_X11Y151_SLICE_X14Y151_CO6;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_D = CLBLM_R_X11Y151_SLICE_X14Y151_DO6;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_CMUX = CLBLM_R_X11Y151_SLICE_X14Y151_CO6;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_A = CLBLM_R_X11Y151_SLICE_X15Y151_AO6;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_B = CLBLM_R_X11Y151_SLICE_X15Y151_BO6;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_C = CLBLM_R_X11Y151_SLICE_X15Y151_CO6;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_D = CLBLM_R_X11Y151_SLICE_X15Y151_DO6;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_AMUX = CLBLM_R_X11Y151_SLICE_X15Y151_A5Q;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_CMUX = CLBLM_R_X11Y151_SLICE_X15Y151_CO5;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_A = CLBLM_R_X11Y152_SLICE_X14Y152_AO6;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_B = CLBLM_R_X11Y152_SLICE_X14Y152_BO6;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_C = CLBLM_R_X11Y152_SLICE_X14Y152_CO6;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_D = CLBLM_R_X11Y152_SLICE_X14Y152_DO6;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_AMUX = CLBLM_R_X11Y152_SLICE_X14Y152_A5Q;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_A = CLBLM_R_X11Y152_SLICE_X15Y152_AO6;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_B = CLBLM_R_X11Y152_SLICE_X15Y152_BO6;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_C = CLBLM_R_X11Y152_SLICE_X15Y152_CO6;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_D = CLBLM_R_X11Y152_SLICE_X15Y152_DO6;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_A = CLBLM_R_X11Y153_SLICE_X14Y153_AO6;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_B = CLBLM_R_X11Y153_SLICE_X14Y153_BO6;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_C = CLBLM_R_X11Y153_SLICE_X14Y153_CO6;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_D = CLBLM_R_X11Y153_SLICE_X14Y153_DO6;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_AMUX = CLBLM_R_X11Y153_SLICE_X14Y153_AO5;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_A = CLBLM_R_X11Y153_SLICE_X15Y153_AO6;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_B = CLBLM_R_X11Y153_SLICE_X15Y153_BO6;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_C = CLBLM_R_X11Y153_SLICE_X15Y153_CO6;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_D = CLBLM_R_X11Y153_SLICE_X15Y153_DO6;
  assign CLBLM_R_X13Y145_SLICE_X18Y145_A = CLBLM_R_X13Y145_SLICE_X18Y145_AO6;
  assign CLBLM_R_X13Y145_SLICE_X18Y145_B = CLBLM_R_X13Y145_SLICE_X18Y145_BO6;
  assign CLBLM_R_X13Y145_SLICE_X18Y145_C = CLBLM_R_X13Y145_SLICE_X18Y145_CO6;
  assign CLBLM_R_X13Y145_SLICE_X18Y145_D = CLBLM_R_X13Y145_SLICE_X18Y145_DO6;
  assign CLBLM_R_X13Y145_SLICE_X19Y145_A = CLBLM_R_X13Y145_SLICE_X19Y145_AO6;
  assign CLBLM_R_X13Y145_SLICE_X19Y145_B = CLBLM_R_X13Y145_SLICE_X19Y145_BO6;
  assign CLBLM_R_X13Y145_SLICE_X19Y145_C = CLBLM_R_X13Y145_SLICE_X19Y145_CO6;
  assign CLBLM_R_X13Y145_SLICE_X19Y145_D = CLBLM_R_X13Y145_SLICE_X19Y145_DO6;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_A = CLBLM_R_X103Y178_SLICE_X162Y178_AO6;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_B = CLBLM_R_X103Y178_SLICE_X162Y178_BO6;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_C = CLBLM_R_X103Y178_SLICE_X162Y178_CO6;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_D = CLBLM_R_X103Y178_SLICE_X162Y178_DO6;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_A = CLBLM_R_X103Y178_SLICE_X163Y178_AO6;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_B = CLBLM_R_X103Y178_SLICE_X163Y178_BO6;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_C = CLBLM_R_X103Y178_SLICE_X163Y178_CO6;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_D = CLBLM_R_X103Y178_SLICE_X163Y178_DO6;
  assign LIOI3_X0Y51_ILOGIC_X0Y52_O = LIOB33_X0Y51_IOB_X0Y52_I;
  assign LIOI3_X0Y51_ILOGIC_X0Y51_O = LIOB33_X0Y51_IOB_X0Y51_I;
  assign LIOI3_X0Y53_ILOGIC_X0Y54_O = LIOB33_X0Y53_IOB_X0Y54_I;
  assign LIOI3_X0Y53_ILOGIC_X0Y53_O = LIOB33_X0Y53_IOB_X0Y53_I;
  assign LIOI3_X0Y55_ILOGIC_X0Y56_O = LIOB33_X0Y55_IOB_X0Y56_I;
  assign LIOI3_X0Y55_ILOGIC_X0Y55_O = LIOB33_X0Y55_IOB_X0Y55_I;
  assign LIOI3_X0Y59_ILOGIC_X0Y60_O = LIOB33_X0Y59_IOB_X0Y60_I;
  assign LIOI3_X0Y59_ILOGIC_X0Y59_O = LIOB33_X0Y59_IOB_X0Y59_I;
  assign LIOI3_X0Y61_ILOGIC_X0Y62_O = LIOB33_X0Y61_IOB_X0Y62_I;
  assign LIOI3_X0Y61_ILOGIC_X0Y61_O = LIOB33_X0Y61_IOB_X0Y61_I;
  assign LIOI3_X0Y65_OLOGIC_X0Y66_OQ = CLBLM_R_X7Y152_SLICE_X9Y152_DQ;
  assign LIOI3_X0Y65_OLOGIC_X0Y66_TQ = 1'b1;
  assign LIOI3_X0Y65_OLOGIC_X0Y65_OQ = CLBLL_L_X4Y140_SLICE_X5Y140_CO6;
  assign LIOI3_X0Y65_OLOGIC_X0Y65_TQ = 1'b1;
  assign LIOI3_X0Y77_ILOGIC_X0Y78_O = LIOB33_X0Y77_IOB_X0Y78_I;
  assign LIOI3_X0Y101_OLOGIC_X0Y102_OQ = CLBLM_R_X5Y140_SLICE_X7Y140_BQ;
  assign LIOI3_X0Y101_OLOGIC_X0Y102_TQ = 1'b1;
  assign LIOI3_X0Y101_OLOGIC_X0Y101_OQ = CLBLM_R_X3Y142_SLICE_X2Y142_B5Q;
  assign LIOI3_X0Y101_OLOGIC_X0Y101_TQ = 1'b1;
  assign LIOI3_X0Y103_OLOGIC_X0Y104_OQ = CLBLM_R_X7Y144_SLICE_X9Y144_C5Q;
  assign LIOI3_X0Y103_OLOGIC_X0Y104_TQ = 1'b1;
  assign LIOI3_X0Y103_OLOGIC_X0Y103_OQ = CLBLL_L_X4Y150_SLICE_X5Y150_DQ;
  assign LIOI3_X0Y103_OLOGIC_X0Y103_TQ = 1'b1;
  assign LIOI3_X0Y105_OLOGIC_X0Y106_OQ = CLBLL_L_X4Y147_SLICE_X5Y147_DQ;
  assign LIOI3_X0Y105_OLOGIC_X0Y106_TQ = 1'b1;
  assign LIOI3_X0Y105_OLOGIC_X0Y105_OQ = CLBLM_R_X5Y144_SLICE_X6Y144_B5Q;
  assign LIOI3_X0Y105_OLOGIC_X0Y105_TQ = 1'b1;
  assign LIOI3_X0Y109_OLOGIC_X0Y110_OQ = CLBLM_R_X5Y143_SLICE_X6Y143_DQ;
  assign LIOI3_X0Y109_OLOGIC_X0Y110_TQ = 1'b1;
  assign LIOI3_X0Y109_OLOGIC_X0Y109_OQ = CLBLL_L_X2Y153_SLICE_X1Y153_AQ;
  assign LIOI3_X0Y109_OLOGIC_X0Y109_TQ = 1'b1;
  assign LIOI3_X0Y111_OLOGIC_X0Y112_OQ = CLBLM_R_X3Y145_SLICE_X2Y145_B5Q;
  assign LIOI3_X0Y111_OLOGIC_X0Y112_TQ = 1'b1;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_OQ = CLBLM_R_X3Y145_SLICE_X2Y145_CQ;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_TQ = 1'b1;
  assign LIOI3_X0Y115_OLOGIC_X0Y116_OQ = CLBLM_R_X5Y152_SLICE_X6Y152_CQ;
  assign LIOI3_X0Y115_OLOGIC_X0Y116_TQ = 1'b1;
  assign LIOI3_X0Y115_OLOGIC_X0Y115_OQ = CLBLM_R_X3Y151_SLICE_X3Y151_CQ;
  assign LIOI3_X0Y115_OLOGIC_X0Y115_TQ = 1'b1;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_OQ = CLBLM_R_X11Y147_SLICE_X15Y147_AQ;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_TQ = 1'b1;
  assign LIOI3_X0Y117_OLOGIC_X0Y117_OQ = CLBLM_R_X7Y144_SLICE_X9Y144_B5Q;
  assign LIOI3_X0Y117_OLOGIC_X0Y117_TQ = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_OQ = CLBLL_L_X4Y149_SLICE_X4Y149_D5Q;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_TQ = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_OQ = CLBLM_L_X8Y146_SLICE_X10Y146_AQ;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_TQ = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_OQ = CLBLM_R_X7Y152_SLICE_X9Y152_DQ;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_TQ = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_OQ = CLBLM_R_X3Y149_SLICE_X2Y149_CQ;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_TQ = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_OQ = CLBLM_R_X5Y144_SLICE_X6Y144_CQ;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_TQ = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_OQ = CLBLM_R_X5Y144_SLICE_X6Y144_DQ;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_TQ = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_OQ = CLBLM_L_X8Y142_SLICE_X11Y142_CQ;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_TQ = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_OQ = CLBLM_L_X8Y150_SLICE_X11Y150_B5Q;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_TQ = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_OQ = CLBLM_R_X3Y149_SLICE_X2Y149_BQ;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_TQ = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_OQ = CLBLM_R_X3Y149_SLICE_X2Y149_CQ;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_TQ = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_OQ = CLBLM_R_X3Y149_SLICE_X2Y149_BQ;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_TQ = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_OQ = CLBLM_R_X3Y142_SLICE_X2Y142_CO5;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_TQ = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_OQ = CLBLM_L_X8Y153_SLICE_X10Y153_AQ;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_TQ = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_OQ = CLBLM_R_X3Y149_SLICE_X2Y149_BQ;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_TQ = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_OQ = CLBLL_L_X2Y147_SLICE_X0Y147_BQ;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_TQ = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_OQ = CLBLL_L_X2Y148_SLICE_X0Y148_AQ;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_TQ = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_OQ = CLBLM_R_X3Y149_SLICE_X2Y149_CQ;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_TQ = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_OQ = CLBLL_L_X2Y150_SLICE_X1Y150_C5Q;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_TQ = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_OQ = CLBLL_L_X2Y148_SLICE_X1Y148_BO6;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_TQ = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_OQ = CLBLL_L_X2Y146_SLICE_X1Y146_CO6;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_TQ = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_OQ = CLBLM_R_X3Y149_SLICE_X2Y149_DO6;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_TQ = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_OQ = CLBLM_R_X5Y147_SLICE_X7Y147_DO6;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_TQ = 1'b1;
  assign LIOI3_X0Y151_OLOGIC_X0Y152_OQ = CLBLM_R_X3Y150_SLICE_X2Y150_B5Q;
  assign LIOI3_X0Y151_OLOGIC_X0Y152_TQ = 1'b1;
  assign LIOI3_X0Y151_OLOGIC_X0Y151_OQ = CLBLM_R_X3Y149_SLICE_X2Y149_CQ;
  assign LIOI3_X0Y151_OLOGIC_X0Y151_TQ = 1'b1;
  assign LIOI3_X0Y153_OLOGIC_X0Y154_OQ = CLBLM_L_X8Y152_SLICE_X10Y152_DQ;
  assign LIOI3_X0Y153_OLOGIC_X0Y154_TQ = 1'b1;
  assign LIOI3_X0Y153_OLOGIC_X0Y153_OQ = CLBLM_L_X10Y153_SLICE_X13Y153_AQ;
  assign LIOI3_X0Y153_OLOGIC_X0Y153_TQ = 1'b1;
  assign LIOI3_X0Y155_OLOGIC_X0Y156_OQ = CLBLM_R_X7Y152_SLICE_X9Y152_BQ;
  assign LIOI3_X0Y155_OLOGIC_X0Y156_TQ = 1'b1;
  assign LIOI3_X0Y155_OLOGIC_X0Y155_OQ = CLBLM_L_X8Y150_SLICE_X11Y150_CQ;
  assign LIOI3_X0Y155_OLOGIC_X0Y155_TQ = 1'b1;
  assign LIOI3_X0Y159_OLOGIC_X0Y160_OQ = CLBLL_L_X4Y145_SLICE_X5Y145_AQ;
  assign LIOI3_X0Y159_OLOGIC_X0Y160_TQ = 1'b1;
  assign LIOI3_X0Y159_OLOGIC_X0Y159_OQ = CLBLM_R_X3Y149_SLICE_X2Y149_CQ;
  assign LIOI3_X0Y159_OLOGIC_X0Y159_TQ = 1'b1;
  assign LIOI3_X0Y161_OLOGIC_X0Y162_OQ = CLBLM_R_X3Y153_SLICE_X3Y153_CO6;
  assign LIOI3_X0Y161_OLOGIC_X0Y162_TQ = 1'b1;
  assign LIOI3_X0Y161_OLOGIC_X0Y161_OQ = CLBLM_R_X5Y151_SLICE_X6Y151_CQ;
  assign LIOI3_X0Y161_OLOGIC_X0Y161_TQ = 1'b1;
  assign LIOI3_X0Y165_OLOGIC_X0Y166_OQ = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign LIOI3_X0Y165_OLOGIC_X0Y166_TQ = 1'b1;
  assign LIOI3_X0Y165_OLOGIC_X0Y165_OQ = LIOB33_X0Y57_IOB_X0Y57_I;
  assign LIOI3_X0Y165_OLOGIC_X0Y165_TQ = 1'b1;
  assign LIOI3_X0Y167_OLOGIC_X0Y168_OQ = RIOB33_X105Y101_IOB_X1Y101_I;
  assign LIOI3_X0Y167_OLOGIC_X0Y168_TQ = 1'b1;
  assign LIOI3_X0Y167_OLOGIC_X0Y167_OQ = RIOB33_X105Y105_IOB_X1Y106_I;
  assign LIOI3_X0Y167_OLOGIC_X0Y167_TQ = 1'b1;
  assign LIOI3_X0Y171_OLOGIC_X0Y172_OQ = RIOB33_X105Y119_IOB_X1Y120_I;
  assign LIOI3_X0Y171_OLOGIC_X0Y172_TQ = 1'b1;
  assign LIOI3_X0Y171_OLOGIC_X0Y171_OQ = RIOB33_X105Y119_IOB_X1Y119_I;
  assign LIOI3_X0Y171_OLOGIC_X0Y171_TQ = 1'b1;
  assign LIOI3_X0Y173_OLOGIC_X0Y174_OQ = RIOB33_X105Y121_IOB_X1Y122_I;
  assign LIOI3_X0Y173_OLOGIC_X0Y174_TQ = 1'b1;
  assign LIOI3_X0Y173_OLOGIC_X0Y173_OQ = RIOB33_X105Y121_IOB_X1Y121_I;
  assign LIOI3_X0Y173_OLOGIC_X0Y173_TQ = 1'b1;
  assign LIOI3_X0Y175_OLOGIC_X0Y176_OQ = RIOB33_X105Y115_IOB_X1Y116_I;
  assign LIOI3_X0Y175_OLOGIC_X0Y176_TQ = 1'b1;
  assign LIOI3_X0Y175_OLOGIC_X0Y175_OQ = RIOB33_X105Y123_IOB_X1Y123_I;
  assign LIOI3_X0Y175_OLOGIC_X0Y175_TQ = 1'b1;
  assign LIOI3_X0Y177_OLOGIC_X0Y178_OQ = RIOB33_X105Y125_IOB_X1Y125_I;
  assign LIOI3_X0Y177_OLOGIC_X0Y178_TQ = 1'b1;
  assign LIOI3_X0Y177_OLOGIC_X0Y177_OQ = RIOB33_X105Y123_IOB_X1Y124_I;
  assign LIOI3_X0Y177_OLOGIC_X0Y177_TQ = 1'b1;
  assign LIOI3_X0Y179_OLOGIC_X0Y180_OQ = RIOB33_X105Y127_IOB_X1Y127_I;
  assign LIOI3_X0Y179_OLOGIC_X0Y180_TQ = 1'b1;
  assign LIOI3_X0Y179_OLOGIC_X0Y179_OQ = RIOB33_X105Y125_IOB_X1Y126_I;
  assign LIOI3_X0Y179_OLOGIC_X0Y179_TQ = 1'b1;
  assign LIOI3_X0Y183_OLOGIC_X0Y184_OQ = RIOB33_X105Y131_IOB_X1Y132_I;
  assign LIOI3_X0Y183_OLOGIC_X0Y184_TQ = 1'b1;
  assign LIOI3_X0Y183_OLOGIC_X0Y183_OQ = RIOB33_X105Y129_IOB_X1Y130_I;
  assign LIOI3_X0Y183_OLOGIC_X0Y183_TQ = 1'b1;
  assign LIOI3_X0Y185_OLOGIC_X0Y186_OQ = RIOB33_X105Y119_IOB_X1Y120_I;
  assign LIOI3_X0Y185_OLOGIC_X0Y186_TQ = 1'b1;
  assign LIOI3_X0Y185_OLOGIC_X0Y185_OQ = RIOB33_X105Y133_IOB_X1Y133_I;
  assign LIOI3_X0Y185_OLOGIC_X0Y185_TQ = 1'b1;
  assign LIOI3_X0Y189_OLOGIC_X0Y190_OQ = CLBLM_R_X7Y155_SLICE_X9Y155_AO6;
  assign LIOI3_X0Y189_OLOGIC_X0Y190_TQ = 1'b1;
  assign LIOI3_X0Y189_OLOGIC_X0Y189_OQ = CLBLM_R_X3Y149_SLICE_X3Y149_DQ;
  assign LIOI3_X0Y189_OLOGIC_X0Y189_TQ = 1'b1;
  assign LIOI3_X0Y191_OLOGIC_X0Y192_OQ = CLBLL_L_X4Y154_SLICE_X4Y154_AO5;
  assign LIOI3_X0Y191_OLOGIC_X0Y192_TQ = 1'b1;
  assign LIOI3_X0Y191_OLOGIC_X0Y191_OQ = CLBLL_L_X4Y145_SLICE_X4Y145_BO6;
  assign LIOI3_X0Y191_OLOGIC_X0Y191_TQ = 1'b1;
  assign LIOI3_X0Y195_OLOGIC_X0Y196_OQ = CLBLL_L_X4Y154_SLICE_X5Y154_AO6;
  assign LIOI3_X0Y195_OLOGIC_X0Y196_TQ = 1'b1;
  assign LIOI3_X0Y195_OLOGIC_X0Y195_OQ = CLBLL_L_X2Y152_SLICE_X1Y152_AO6;
  assign LIOI3_X0Y195_OLOGIC_X0Y195_TQ = 1'b1;
  assign LIOI3_X0Y197_OLOGIC_X0Y198_OQ = 1'b1;
  assign LIOI3_X0Y197_OLOGIC_X0Y198_TQ = 1'b1;
  assign LIOI3_X0Y197_OLOGIC_X0Y197_OQ = CLBLM_R_X3Y153_SLICE_X3Y153_BO5;
  assign LIOI3_X0Y197_OLOGIC_X0Y197_TQ = 1'b1;
  assign LIOI3_SING_X0Y50_ILOGIC_X0Y50_O = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign LIOI3_SING_X0Y100_OLOGIC_X0Y100_OQ = CLBLM_R_X3Y149_SLICE_X2Y149_AQ;
  assign LIOI3_SING_X0Y100_OLOGIC_X0Y100_TQ = 1'b1;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_OQ = RIOB33_X105Y115_IOB_X1Y115_I;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_TQ = 1'b1;
  assign LIOI3_SING_X0Y150_OLOGIC_X0Y150_OQ = CLBLL_L_X4Y142_SLICE_X4Y142_DO5;
  assign LIOI3_SING_X0Y150_OLOGIC_X0Y150_TQ = 1'b1;
  assign LIOI3_SING_X0Y199_OLOGIC_X0Y199_OQ = 1'b1;
  assign LIOI3_SING_X0Y199_OLOGIC_X0Y199_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y58_O = LIOB33_X0Y57_IOB_X0Y58_I;
  assign LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y57_O = LIOB33_X0Y57_IOB_X0Y57_I;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_OQ = CLBLL_L_X4Y143_SLICE_X5Y143_C5Q;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_OQ = CLBLM_R_X3Y145_SLICE_X2Y145_C5Q;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_OQ = CLBLM_R_X3Y150_SLICE_X3Y150_AQ;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_OQ = CLBLM_R_X3Y149_SLICE_X2Y149_CQ;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_OQ = CLBLL_L_X4Y142_SLICE_X4Y142_BO5;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_OQ = CLBLL_L_X2Y75_SLICE_X0Y75_AO6;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_OQ = CLBLM_R_X3Y144_SLICE_X2Y144_CO6;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_OQ = CLBLL_L_X2Y150_SLICE_X1Y150_DO5;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_OQ = RIOB33_X105Y133_IOB_X1Y134_I;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_OQ = CLBLM_R_X7Y153_SLICE_X9Y153_CQ;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_OQ = RIOB33_X105Y117_IOB_X1Y118_I;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_OQ = RIOB33_X105Y117_IOB_X1Y117_I;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_OQ = RIOB33_X105Y129_IOB_X1Y129_I;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_OQ = RIOB33_X105Y127_IOB_X1Y128_I;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_OQ = RIOB33_X105Y103_IOB_X1Y103_I;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_OQ = CLBLL_L_X2Y166_SLICE_X0Y166_AO6;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y63_O = LIOB33_X0Y63_IOB_X0Y63_I;
  assign LIOI3_TBYTETERM_X0Y63_OLOGIC_X0Y64_OQ = CLBLL_L_X4Y140_SLICE_X5Y140_BO6;
  assign LIOI3_TBYTETERM_X0Y63_OLOGIC_X0Y64_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_OQ = CLBLL_L_X4Y153_SLICE_X4Y153_A5Q;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_OQ = CLBLM_R_X3Y146_SLICE_X2Y146_CQ;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_OQ = CLBLM_R_X3Y144_SLICE_X3Y144_A5Q;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_OQ = CLBLM_R_X7Y150_SLICE_X9Y150_B5Q;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_OQ = RIOB33_X105Y101_IOB_X1Y102_I;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_OQ = CLBLM_R_X5Y159_SLICE_X6Y159_AO6;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_OQ = CLBLM_R_X3Y150_SLICE_X3Y150_BQ;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_OQ = CLBLM_L_X10Y150_SLICE_X12Y150_CQ;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_TQ = 1'b1;
  assign RIOI3_X105Y101_ILOGIC_X1Y102_O = RIOB33_X105Y101_IOB_X1Y102_I;
  assign RIOI3_X105Y101_ILOGIC_X1Y101_O = RIOB33_X105Y101_IOB_X1Y101_I;
  assign RIOI3_X105Y103_ILOGIC_X1Y104_O = RIOB33_X105Y103_IOB_X1Y104_I;
  assign RIOI3_X105Y103_ILOGIC_X1Y103_O = RIOB33_X105Y103_IOB_X1Y103_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y106_O = RIOB33_X105Y105_IOB_X1Y106_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y105_O = RIOB33_X105Y105_IOB_X1Y105_I;
  assign RIOI3_X105Y109_ILOGIC_X1Y110_O = RIOB33_X105Y109_IOB_X1Y110_I;
  assign RIOI3_X105Y109_ILOGIC_X1Y109_O = RIOB33_X105Y109_IOB_X1Y109_I;
  assign RIOI3_X105Y111_ILOGIC_X1Y112_O = RIOB33_X105Y111_IOB_X1Y112_I;
  assign RIOI3_X105Y111_ILOGIC_X1Y111_O = RIOB33_X105Y111_IOB_X1Y111_I;
  assign RIOI3_X105Y115_ILOGIC_X1Y116_O = RIOB33_X105Y115_IOB_X1Y116_I;
  assign RIOI3_X105Y115_ILOGIC_X1Y115_O = RIOB33_X105Y115_IOB_X1Y115_I;
  assign RIOI3_X105Y117_ILOGIC_X1Y118_O = RIOB33_X105Y117_IOB_X1Y118_I;
  assign RIOI3_X105Y117_ILOGIC_X1Y117_O = RIOB33_X105Y117_IOB_X1Y117_I;
  assign RIOI3_X105Y121_ILOGIC_X1Y122_O = RIOB33_X105Y121_IOB_X1Y122_I;
  assign RIOI3_X105Y121_ILOGIC_X1Y121_O = RIOB33_X105Y121_IOB_X1Y121_I;
  assign RIOI3_X105Y123_ILOGIC_X1Y124_O = RIOB33_X105Y123_IOB_X1Y124_I;
  assign RIOI3_X105Y123_ILOGIC_X1Y123_O = RIOB33_X105Y123_IOB_X1Y123_I;
  assign RIOI3_X105Y125_ILOGIC_X1Y126_O = RIOB33_X105Y125_IOB_X1Y126_I;
  assign RIOI3_X105Y125_ILOGIC_X1Y125_O = RIOB33_X105Y125_IOB_X1Y125_I;
  assign RIOI3_X105Y127_ILOGIC_X1Y128_O = RIOB33_X105Y127_IOB_X1Y128_I;
  assign RIOI3_X105Y127_ILOGIC_X1Y127_O = RIOB33_X105Y127_IOB_X1Y127_I;
  assign RIOI3_X105Y129_ILOGIC_X1Y130_O = RIOB33_X105Y129_IOB_X1Y130_I;
  assign RIOI3_X105Y129_ILOGIC_X1Y129_O = RIOB33_X105Y129_IOB_X1Y129_I;
  assign RIOI3_X105Y133_ILOGIC_X1Y134_O = RIOB33_X105Y133_IOB_X1Y134_I;
  assign RIOI3_X105Y133_ILOGIC_X1Y133_O = RIOB33_X105Y133_IOB_X1Y133_I;
  assign RIOI3_X105Y135_ILOGIC_X1Y136_O = RIOB33_X105Y135_IOB_X1Y136_I;
  assign RIOI3_X105Y135_ILOGIC_X1Y135_O = RIOB33_X105Y135_IOB_X1Y135_I;
  assign RIOI3_X105Y139_ILOGIC_X1Y140_O = RIOB33_X105Y139_IOB_X1Y140_I;
  assign RIOI3_X105Y139_ILOGIC_X1Y139_O = RIOB33_X105Y139_IOB_X1Y139_I;
  assign RIOI3_X105Y141_ILOGIC_X1Y142_O = RIOB33_X105Y141_IOB_X1Y142_I;
  assign RIOI3_X105Y141_ILOGIC_X1Y141_O = RIOB33_X105Y141_IOB_X1Y141_I;
  assign RIOI3_X105Y145_ILOGIC_X1Y146_O = RIOB33_X105Y145_IOB_X1Y146_I;
  assign RIOI3_X105Y145_ILOGIC_X1Y145_O = RIOB33_X105Y145_IOB_X1Y145_I;
  assign RIOI3_X105Y147_ILOGIC_X1Y148_O = RIOB33_X105Y147_IOB_X1Y148_I;
  assign RIOI3_X105Y147_ILOGIC_X1Y147_O = RIOB33_X105Y147_IOB_X1Y147_I;
  assign RIOI3_X105Y151_OLOGIC_X1Y152_OQ = 1'b1;
  assign RIOI3_X105Y151_OLOGIC_X1Y152_TQ = 1'b1;
  assign RIOI3_X105Y151_OLOGIC_X1Y151_OQ = 1'b1;
  assign RIOI3_X105Y151_OLOGIC_X1Y151_TQ = 1'b1;
  assign RIOI3_X105Y153_OLOGIC_X1Y154_OQ = 1'b1;
  assign RIOI3_X105Y153_OLOGIC_X1Y154_TQ = 1'b1;
  assign RIOI3_X105Y153_OLOGIC_X1Y153_OQ = 1'b1;
  assign RIOI3_X105Y153_OLOGIC_X1Y153_TQ = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y156_OQ = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y156_TQ = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y155_OQ = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y155_TQ = 1'b1;
  assign RIOI3_X105Y159_OLOGIC_X1Y160_OQ = 1'b1;
  assign RIOI3_X105Y159_OLOGIC_X1Y160_TQ = 1'b1;
  assign RIOI3_X105Y159_OLOGIC_X1Y159_OQ = 1'b1;
  assign RIOI3_X105Y159_OLOGIC_X1Y159_TQ = 1'b1;
  assign RIOI3_X105Y161_OLOGIC_X1Y162_OQ = CLBLM_L_X10Y150_SLICE_X13Y150_C5Q;
  assign RIOI3_X105Y161_OLOGIC_X1Y162_TQ = 1'b1;
  assign RIOI3_X105Y161_OLOGIC_X1Y161_OQ = CLBLM_L_X8Y153_SLICE_X11Y153_AO5;
  assign RIOI3_X105Y161_OLOGIC_X1Y161_TQ = 1'b1;
  assign RIOI3_X105Y165_OLOGIC_X1Y166_OQ = CLBLM_L_X10Y153_SLICE_X13Y153_AQ;
  assign RIOI3_X105Y165_OLOGIC_X1Y166_TQ = 1'b1;
  assign RIOI3_X105Y165_OLOGIC_X1Y165_OQ = CLBLM_R_X3Y153_SLICE_X2Y153_AO5;
  assign RIOI3_X105Y165_OLOGIC_X1Y165_TQ = 1'b1;
  assign RIOI3_X105Y167_OLOGIC_X1Y168_OQ = CLBLM_L_X8Y150_SLICE_X11Y150_CQ;
  assign RIOI3_X105Y167_OLOGIC_X1Y168_TQ = 1'b1;
  assign RIOI3_X105Y167_OLOGIC_X1Y167_OQ = CLBLM_L_X8Y152_SLICE_X10Y152_DQ;
  assign RIOI3_X105Y167_OLOGIC_X1Y167_TQ = 1'b1;
  assign RIOI3_X105Y171_OLOGIC_X1Y172_OQ = CLBLL_L_X4Y145_SLICE_X5Y145_AQ;
  assign RIOI3_X105Y171_OLOGIC_X1Y172_TQ = 1'b1;
  assign RIOI3_X105Y171_OLOGIC_X1Y171_OQ = CLBLM_R_X7Y153_SLICE_X8Y153_CO5;
  assign RIOI3_X105Y171_OLOGIC_X1Y171_TQ = 1'b1;
  assign RIOI3_X105Y173_OLOGIC_X1Y174_OQ = CLBLM_R_X5Y159_SLICE_X6Y159_AO6;
  assign RIOI3_X105Y173_OLOGIC_X1Y174_TQ = 1'b1;
  assign RIOI3_X105Y173_OLOGIC_X1Y173_OQ = CLBLM_R_X5Y151_SLICE_X6Y151_CQ;
  assign RIOI3_X105Y173_OLOGIC_X1Y173_TQ = 1'b1;
  assign RIOI3_X105Y175_OLOGIC_X1Y176_OQ = CLBLL_L_X2Y151_SLICE_X1Y151_CO6;
  assign RIOI3_X105Y175_OLOGIC_X1Y176_TQ = 1'b1;
  assign RIOI3_X105Y175_OLOGIC_X1Y175_OQ = CLBLM_R_X3Y153_SLICE_X3Y153_CO6;
  assign RIOI3_X105Y175_OLOGIC_X1Y175_TQ = 1'b1;
  assign RIOI3_X105Y177_OLOGIC_X1Y178_OQ = CLBLM_R_X3Y150_SLICE_X3Y150_BQ;
  assign RIOI3_X105Y177_OLOGIC_X1Y178_TQ = 1'b1;
  assign RIOI3_X105Y177_OLOGIC_X1Y177_OQ = CLBLM_L_X10Y142_SLICE_X12Y142_AQ;
  assign RIOI3_X105Y177_OLOGIC_X1Y177_TQ = 1'b1;
  assign RIOI3_X105Y179_OLOGIC_X1Y180_OQ = CLBLM_L_X10Y150_SLICE_X12Y150_CQ;
  assign RIOI3_X105Y179_OLOGIC_X1Y180_TQ = 1'b1;
  assign RIOI3_X105Y179_OLOGIC_X1Y179_OQ = CLBLM_R_X3Y149_SLICE_X3Y149_DQ;
  assign RIOI3_X105Y179_OLOGIC_X1Y179_TQ = 1'b1;
  assign RIOI3_X105Y183_OLOGIC_X1Y184_OQ = CLBLL_L_X4Y154_SLICE_X5Y154_AO6;
  assign RIOI3_X105Y183_OLOGIC_X1Y184_TQ = 1'b1;
  assign RIOI3_X105Y183_OLOGIC_X1Y183_OQ = 1'b0;
  assign RIOI3_X105Y183_OLOGIC_X1Y183_TQ = 1'b1;
  assign RIOI3_X105Y185_OLOGIC_X1Y186_OQ = CLBLM_R_X7Y154_SLICE_X9Y154_CO6;
  assign RIOI3_X105Y185_OLOGIC_X1Y186_TQ = 1'b1;
  assign RIOI3_X105Y185_OLOGIC_X1Y185_OQ = CLBLM_L_X8Y154_SLICE_X10Y154_BO6;
  assign RIOI3_X105Y185_OLOGIC_X1Y185_TQ = 1'b1;
  assign RIOI3_X105Y189_OLOGIC_X1Y190_OQ = CLBLM_R_X11Y153_SLICE_X14Y153_AO6;
  assign RIOI3_X105Y189_OLOGIC_X1Y190_TQ = 1'b1;
  assign RIOI3_X105Y189_OLOGIC_X1Y189_OQ = CLBLM_R_X103Y178_SLICE_X163Y178_AO6;
  assign RIOI3_X105Y189_OLOGIC_X1Y189_TQ = 1'b1;
  assign RIOI3_X105Y191_OLOGIC_X1Y192_OQ = CLBLM_L_X12Y151_SLICE_X16Y151_CO6;
  assign RIOI3_X105Y191_OLOGIC_X1Y192_TQ = 1'b1;
  assign RIOI3_X105Y191_OLOGIC_X1Y191_OQ = CLBLM_R_X11Y149_SLICE_X14Y149_AO6;
  assign RIOI3_X105Y191_OLOGIC_X1Y191_TQ = 1'b1;
  assign RIOI3_X105Y195_OLOGIC_X1Y196_OQ = CLBLM_R_X11Y150_SLICE_X14Y150_BO6;
  assign RIOI3_X105Y195_OLOGIC_X1Y196_TQ = 1'b1;
  assign RIOI3_X105Y195_OLOGIC_X1Y195_OQ = CLBLM_R_X11Y149_SLICE_X14Y149_BO6;
  assign RIOI3_X105Y195_OLOGIC_X1Y195_TQ = 1'b1;
  assign RIOI3_X105Y197_OLOGIC_X1Y198_OQ = CLBLM_R_X11Y149_SLICE_X14Y149_CO6;
  assign RIOI3_X105Y197_OLOGIC_X1Y198_TQ = 1'b1;
  assign RIOI3_X105Y197_OLOGIC_X1Y197_OQ = CLBLM_R_X11Y150_SLICE_X14Y150_BO5;
  assign RIOI3_X105Y197_OLOGIC_X1Y197_TQ = 1'b1;
  assign RIOI3_SING_X105Y100_ILOGIC_X1Y100_O = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign RIOI3_SING_X105Y149_ILOGIC_X1Y149_O = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign RIOI3_SING_X105Y150_OLOGIC_X1Y150_OQ = 1'b1;
  assign RIOI3_SING_X105Y150_OLOGIC_X1Y150_TQ = 1'b1;
  assign RIOI3_SING_X105Y199_OLOGIC_X1Y199_OQ = CLBLM_R_X11Y149_SLICE_X14Y149_AQ;
  assign RIOI3_SING_X105Y199_OLOGIC_X1Y199_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_O = RIOB33_X105Y107_IOB_X1Y108_I;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_O = RIOB33_X105Y107_IOB_X1Y107_I;
  assign RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y120_O = RIOB33_X105Y119_IOB_X1Y120_I;
  assign RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_O = RIOB33_X105Y119_IOB_X1Y119_I;
  assign RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y132_O = RIOB33_X105Y131_IOB_X1Y132_I;
  assign RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y131_O = RIOB33_X105Y131_IOB_X1Y131_I;
  assign RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y144_O = RIOB33_X105Y143_IOB_X1Y144_I;
  assign RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y143_O = RIOB33_X105Y143_IOB_X1Y143_I;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_OQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_OQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_OQ = CLBLM_R_X7Y153_SLICE_X9Y153_CQ;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_OQ = CLBLM_R_X7Y152_SLICE_X9Y152_BQ;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_OQ = CLBLM_R_X7Y153_SLICE_X8Y153_DO6;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_OQ = CLBLM_R_X7Y155_SLICE_X9Y155_AO6;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_OQ = CLBLM_L_X12Y151_SLICE_X16Y151_CO5;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_OQ = CLBLM_R_X11Y153_SLICE_X14Y153_AO5;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_O = RIOB33_X105Y113_IOB_X1Y113_I;
  assign RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y138_O = RIOB33_X105Y137_IOB_X1Y138_I;
  assign RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y137_O = RIOB33_X105Y137_IOB_X1Y137_I;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_OQ = CLBLM_R_X11Y151_SLICE_X15Y151_A5Q;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_OQ = CLBLM_L_X10Y149_SLICE_X12Y149_BQ;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_OQ = CLBLM_R_X7Y153_SLICE_X8Y153_DO6;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_OQ = CLBLM_R_X103Y178_SLICE_X163Y178_AO6;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_TQ = 1'b1;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_B1 = CLBLM_R_X7Y150_SLICE_X8Y150_AQ;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_B2 = CLBLM_L_X10Y142_SLICE_X12Y142_CO6;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_B3 = CLBLM_R_X3Y148_SLICE_X2Y148_AQ;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_B4 = CLBLM_L_X8Y140_SLICE_X10Y140_AQ;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_B5 = CLBLM_L_X8Y144_SLICE_X10Y144_BQ;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_B6 = 1'b1;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_BX = CLBLM_L_X8Y145_SLICE_X10Y145_AO6;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_C1 = CLBLM_L_X10Y143_SLICE_X13Y143_AO6;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_C2 = CLBLM_L_X8Y150_SLICE_X10Y150_A5Q;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_C3 = CLBLM_R_X5Y146_SLICE_X6Y146_B5Q;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_C4 = CLBLM_R_X11Y149_SLICE_X14Y149_AQ;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_C5 = CLBLM_R_X7Y146_SLICE_X9Y146_BQ;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_C6 = 1'b1;
  assign LIOB33_X0Y147_IOB_X0Y147_O = CLBLM_R_X5Y147_SLICE_X7Y147_DO6;
  assign LIOB33_X0Y147_IOB_X0Y148_O = CLBLM_R_X3Y149_SLICE_X2Y149_DO6;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_D1 = CLBLM_L_X8Y144_SLICE_X10Y144_CO5;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_D2 = 1'b1;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_D3 = CLBLM_L_X10Y143_SLICE_X12Y143_DO6;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_D4 = CLBLM_L_X10Y143_SLICE_X12Y143_DO5;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_D5 = CLBLM_R_X5Y145_SLICE_X6Y145_CQ;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_D6 = CLBLM_R_X7Y145_SLICE_X8Y145_DQ;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_SR = CLBLL_L_X4Y145_SLICE_X4Y145_DO6;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_A1 = CLBLM_R_X11Y149_SLICE_X14Y149_AO5;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_A2 = CLBLM_L_X10Y149_SLICE_X13Y149_BO5;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_A3 = CLBLM_R_X11Y149_SLICE_X14Y149_BO5;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_A4 = CLBLM_R_X11Y149_SLICE_X15Y149_DO5;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_A5 = CLBLM_L_X12Y149_SLICE_X16Y149_DO6;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_A6 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_B1 = CLBLM_R_X11Y149_SLICE_X14Y149_AO5;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_B2 = CLBLM_R_X3Y146_SLICE_X2Y146_BQ;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_B3 = CLBLM_R_X11Y149_SLICE_X14Y149_BO5;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_B5 = CLBLM_L_X12Y149_SLICE_X16Y149_DO6;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_B6 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign LIOI3_X0Y155_OLOGIC_X0Y156_D1 = CLBLM_R_X7Y152_SLICE_X9Y152_BQ;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_C2 = CLBLM_R_X11Y149_SLICE_X15Y149_CQ;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_C3 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_C4 = CLBLM_R_X11Y145_SLICE_X14Y145_AQ;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_C5 = CLBLM_R_X11Y149_SLICE_X15Y149_DO6;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_A1 = CLBLL_L_X4Y153_SLICE_X4Y153_DO6;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_A2 = 1'b1;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_A3 = CLBLL_L_X4Y152_SLICE_X4Y152_AQ;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_A5 = CLBLL_L_X4Y145_SLICE_X4Y145_AQ;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_A6 = CLBLM_R_X5Y153_SLICE_X7Y153_BO6;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_C6 = CLBLM_L_X12Y149_SLICE_X16Y149_AQ;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_B2 = CLBLM_R_X7Y144_SLICE_X9Y144_AQ;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_B3 = 1'b1;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_B4 = CLBLM_R_X7Y152_SLICE_X8Y152_BQ;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_B5 = CLBLM_R_X5Y151_SLICE_X7Y151_A5Q;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_B6 = CLBLL_L_X4Y150_SLICE_X4Y150_AO5;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_D1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_D2 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_D3 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_C1 = CLBLM_R_X5Y151_SLICE_X6Y151_D5Q;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_C2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_C3 = CLBLL_L_X4Y152_SLICE_X4Y152_BQ;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_C4 = CLBLL_L_X4Y150_SLICE_X4Y150_CO6;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_C5 = CLBLM_R_X3Y153_SLICE_X3Y153_BQ;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_C6 = 1'b1;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_A1 = CLBLM_L_X10Y149_SLICE_X13Y149_CO6;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_A2 = CLBLM_R_X11Y146_SLICE_X14Y146_BO6;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_A3 = CLBLM_R_X3Y151_SLICE_X3Y151_D5Q;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_A4 = CLBLM_L_X10Y148_SLICE_X13Y148_CO6;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_A5 = CLBLM_L_X10Y145_SLICE_X12Y145_BO6;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_A6 = 1'b1;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_AX = CLBLM_L_X10Y149_SLICE_X13Y149_BO6;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_D1 = CLBLM_R_X3Y145_SLICE_X2Y145_DQ;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_D2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_D3 = CLBLM_R_X3Y143_SLICE_X2Y143_AQ;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_D4 = CLBLM_R_X3Y151_SLICE_X2Y151_BQ;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_D5 = CLBLM_L_X8Y152_SLICE_X11Y152_AQ;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_D6 = CLBLM_R_X5Y154_SLICE_X7Y154_BQ;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_B3 = CLBLM_R_X3Y151_SLICE_X3Y151_D5Q;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_B4 = CLBLM_L_X8Y145_SLICE_X11Y145_CO6;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_B5 = CLBLM_L_X8Y147_SLICE_X11Y147_BO6;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_B6 = 1'b1;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_C1 = CLBLM_R_X11Y148_SLICE_X14Y148_AO6;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_C2 = CLBLM_R_X3Y151_SLICE_X3Y151_D5Q;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_C3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_C4 = CLBLM_R_X11Y149_SLICE_X14Y149_AO5;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_C5 = CLBLM_R_X11Y149_SLICE_X14Y149_BO5;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_C6 = CLBLM_R_X11Y149_SLICE_X15Y149_BQ;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_D1 = 1'b1;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_D2 = 1'b1;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_D3 = 1'b1;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_D4 = 1'b1;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_D5 = 1'b1;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_D6 = 1'b1;
  assign RIOB33_SING_X105Y150_IOB_X1Y150_O = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_A3 = CLBLM_R_X5Y143_SLICE_X7Y143_CQ;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_D1 = CLBLM_R_X7Y153_SLICE_X8Y153_DO6;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_A2 = CLBLL_L_X4Y152_SLICE_X5Y152_BQ;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_A3 = CLBLL_L_X4Y152_SLICE_X5Y152_AQ;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_A4 = CLBLL_L_X4Y146_SLICE_X5Y146_BQ;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_A5 = CLBLM_R_X5Y144_SLICE_X6Y144_CQ;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_A6 = CLBLM_R_X3Y147_SLICE_X3Y147_BQ;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_A4 = CLBLM_R_X7Y147_SLICE_X8Y147_DQ;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_B2 = CLBLL_L_X4Y150_SLICE_X4Y150_DO6;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_B3 = CLBLM_R_X5Y152_SLICE_X6Y152_B5Q;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_B4 = CLBLL_L_X4Y152_SLICE_X4Y152_C5Q;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_B5 = CLBLL_L_X4Y152_SLICE_X5Y152_DQ;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_B6 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_A6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_T1 = 1'b1;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_C1 = 1'b1;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_C2 = CLBLL_L_X4Y152_SLICE_X4Y152_C5Q;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_C3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_C4 = CLBLM_R_X5Y141_SLICE_X6Y141_AQ;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_C5 = CLBLM_L_X8Y150_SLICE_X11Y150_CQ;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_C6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_D1 = CLBLM_R_X7Y155_SLICE_X9Y155_AO6;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_D1 = CLBLM_R_X3Y145_SLICE_X2Y145_DQ;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_D2 = CLBLM_L_X10Y150_SLICE_X13Y150_A5Q;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_D3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_D4 = CLBLM_R_X3Y143_SLICE_X2Y143_AQ;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_D5 = CLBLL_L_X4Y152_SLICE_X4Y152_DQ;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_D6 = CLBLL_L_X4Y152_SLICE_X5Y152_AQ;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_B1 = CLBLM_R_X5Y142_SLICE_X7Y142_CQ;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_T1 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_B2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_A2 = 1'b1;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_A3 = CLBLL_L_X4Y150_SLICE_X5Y150_C5Q;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_A4 = CLBLL_L_X4Y146_SLICE_X4Y146_CQ;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_A5 = 1'b1;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_A6 = 1'b1;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_B1 = CLBLM_L_X8Y150_SLICE_X10Y150_A5Q;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_B2 = CLBLM_L_X8Y140_SLICE_X10Y140_A5Q;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_B3 = CLBLM_L_X10Y142_SLICE_X12Y142_DO6;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_B4 = CLBLM_R_X11Y149_SLICE_X14Y149_AQ;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_B5 = CLBLM_L_X10Y143_SLICE_X12Y143_DO5;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_B6 = CLBLL_L_X4Y146_SLICE_X4Y146_CQ;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_C1 = CLBLM_L_X10Y143_SLICE_X12Y143_DO5;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_C2 = CLBLM_L_X10Y142_SLICE_X12Y142_DO6;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_C3 = CLBLM_L_X8Y146_SLICE_X11Y146_AQ;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_C4 = CLBLM_L_X8Y150_SLICE_X10Y150_A5Q;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_C5 = CLBLM_L_X8Y146_SLICE_X10Y146_DQ;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_C6 = CLBLM_R_X11Y149_SLICE_X14Y149_AQ;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_D1 = 1'b1;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_D2 = 1'b1;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_D3 = 1'b1;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_D4 = 1'b1;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_D5 = 1'b1;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_D6 = 1'b1;
  assign LIOB33_X0Y151_IOB_X0Y151_O = CLBLM_R_X3Y149_SLICE_X2Y149_CQ;
  assign LIOB33_X0Y151_IOB_X0Y152_O = CLBLM_R_X3Y150_SLICE_X2Y150_B5Q;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_SR = CLBLM_R_X11Y148_SLICE_X14Y148_DO6;
  assign LIOI3_SING_X0Y199_OLOGIC_X0Y199_D1 = 1'b1;
  assign RIOB33_SING_X105Y199_IOB_X1Y199_O = CLBLM_R_X11Y149_SLICE_X14Y149_AQ;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_A2 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_A3 = CLBLM_L_X8Y143_SLICE_X10Y143_CQ;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_A4 = CLBLL_L_X4Y149_SLICE_X4Y149_C5Q;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_A5 = CLBLM_R_X7Y149_SLICE_X8Y149_DQ;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_A6 = 1'b1;
  assign LIOI3_SING_X0Y199_OLOGIC_X0Y199_T1 = 1'b1;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_B1 = CLBLL_L_X4Y146_SLICE_X5Y146_B5Q;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_B2 = CLBLM_L_X8Y146_SLICE_X10Y146_BQ;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_B3 = CLBLM_R_X5Y144_SLICE_X6Y144_DQ;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_B4 = CLBLM_R_X3Y148_SLICE_X2Y148_D5Q;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_B5 = CLBLM_L_X8Y141_SLICE_X10Y141_BQ;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_B6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign RIOI3_X105Y139_ILOGIC_X1Y140_D = RIOB33_X105Y139_IOB_X1Y140_I;
  assign RIOI3_X105Y139_ILOGIC_X1Y139_D = RIOB33_X105Y139_IOB_X1Y139_I;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_C1 = CLBLL_L_X4Y144_SLICE_X5Y144_B5Q;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_C2 = CLBLL_L_X4Y141_SLICE_X5Y141_A5Q;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_C3 = CLBLM_L_X10Y150_SLICE_X13Y150_AQ;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_C5 = 1'b1;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_C6 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_D1 = 1'b1;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_D3 = 1'b1;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_D1 = CLBLL_L_X4Y145_SLICE_X5Y145_AQ;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_D2 = CLBLM_L_X8Y143_SLICE_X10Y143_CQ;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_D3 = CLBLM_L_X8Y146_SLICE_X10Y146_DQ;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_D4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_D5 = CLBLM_L_X10Y143_SLICE_X12Y143_AO6;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_D6 = 1'b1;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_A1 = CLBLM_L_X8Y146_SLICE_X10Y146_A5Q;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_A2 = 1'b1;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_A3 = CLBLM_R_X11Y150_SLICE_X15Y150_AQ;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_A5 = CLBLM_R_X11Y148_SLICE_X14Y148_AQ;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_A6 = CLBLM_R_X3Y148_SLICE_X2Y148_B5Q;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_B1 = 1'b1;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_B2 = 1'b1;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_B3 = 1'b1;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_B4 = 1'b1;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_B5 = 1'b1;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_B6 = 1'b1;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_A1 = CLBLL_L_X4Y153_SLICE_X4Y153_CQ;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_A2 = CLBLM_R_X5Y154_SLICE_X6Y154_AQ;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_A3 = CLBLL_L_X4Y153_SLICE_X4Y153_AQ;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_A5 = CLBLM_R_X5Y153_SLICE_X7Y153_BO6;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_A6 = CLBLM_R_X3Y153_SLICE_X3Y153_DO6;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_C1 = 1'b1;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_C2 = 1'b1;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_AX = CLBLL_L_X4Y154_SLICE_X4Y154_BO5;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_C3 = 1'b1;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_B1 = CLBLL_L_X4Y149_SLICE_X5Y149_DQ;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_B2 = CLBLL_L_X4Y153_SLICE_X4Y153_BQ;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_B4 = CLBLL_L_X4Y153_SLICE_X4Y153_DO5;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_B5 = 1'b1;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_B6 = CLBLM_R_X5Y153_SLICE_X7Y153_BO6;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_D1 = 1'b1;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_C1 = CLBLM_R_X11Y149_SLICE_X15Y149_CQ;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_C2 = CLBLL_L_X4Y153_SLICE_X4Y153_CQ;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_C3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_C4 = CLBLM_R_X5Y153_SLICE_X7Y153_BO6;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_C5 = 1'b1;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_C6 = CLBLM_R_X3Y153_SLICE_X3Y153_DO6;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_D3 = 1'b1;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_D4 = 1'b1;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_A1 = CLBLM_R_X11Y145_SLICE_X14Y145_DQ;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_A2 = 1'b1;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_A3 = 1'b1;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_A4 = 1'b1;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_A5 = 1'b1;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_D1 = CLBLL_L_X4Y153_SLICE_X4Y153_BQ;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_D2 = CLBLL_L_X4Y153_SLICE_X4Y153_CQ;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_D3 = CLBLL_L_X4Y153_SLICE_X4Y153_AQ;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_D4 = CLBLM_R_X3Y153_SLICE_X3Y153_DO6;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_D5 = 1'b1;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_D6 = 1'b1;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_B1 = 1'b1;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_B2 = CLBLM_R_X11Y147_SLICE_X14Y147_BO6;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_B3 = CLBLM_L_X8Y145_SLICE_X11Y145_CO6;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_B4 = CLBLM_R_X3Y151_SLICE_X3Y151_D5Q;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_B5 = 1'b1;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_B6 = 1'b1;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_C1 = CLBLM_R_X7Y152_SLICE_X8Y152_CQ;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_C2 = CLBLM_L_X10Y150_SLICE_X13Y150_DO5;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_C1 = 1'b1;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_C3 = CLBLM_L_X8Y147_SLICE_X11Y147_A5Q;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_C4 = CLBLM_R_X7Y151_SLICE_X9Y151_DQ;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_C5 = 1'b1;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_C6 = CLBLM_R_X11Y147_SLICE_X14Y147_A5Q;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_C2 = 1'b1;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_D1 = 1'b1;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_D2 = 1'b1;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_D3 = 1'b1;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_D4 = CLBLM_R_X5Y153_SLICE_X6Y153_AQ;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_A1 = CLBLM_R_X5Y149_SLICE_X6Y149_CQ;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_A2 = CLBLM_R_X7Y153_SLICE_X8Y153_CO6;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_A3 = CLBLM_R_X7Y144_SLICE_X9Y144_B5Q;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_A5 = CLBLL_L_X4Y153_SLICE_X5Y153_AQ;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_A6 = CLBLL_L_X4Y153_SLICE_X5Y153_CO6;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_D5 = 1'b1;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_D6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_B1 = CLBLL_L_X2Y148_SLICE_X0Y148_B5Q;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_B2 = CLBLL_L_X4Y153_SLICE_X5Y153_BQ;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_B3 = CLBLM_R_X5Y153_SLICE_X6Y153_AQ;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_B5 = CLBLM_R_X3Y152_SLICE_X2Y152_DO6;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_B6 = CLBLM_L_X10Y152_SLICE_X13Y152_BQ;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_C1 = CLBLL_L_X4Y153_SLICE_X4Y153_AQ;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_C2 = CLBLM_R_X3Y153_SLICE_X3Y153_BQ;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_C3 = CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_C4 = CLBLL_L_X4Y153_SLICE_X4Y153_CQ;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_C5 = CLBLL_L_X4Y150_SLICE_X5Y150_D5Q;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_C6 = CLBLL_L_X4Y153_SLICE_X5Y153_DO6;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_D1 = CLBLL_L_X4Y152_SLICE_X4Y152_AQ;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_D2 = CLBLM_R_X7Y153_SLICE_X8Y153_CO6;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_D3 = CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_D4 = CLBLM_R_X3Y148_SLICE_X3Y148_BO6;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_D5 = CLBLM_R_X3Y149_SLICE_X3Y149_AQ;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_D6 = CLBLL_L_X4Y153_SLICE_X4Y153_BQ;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_C2 = CLBLM_R_X7Y150_SLICE_X9Y150_B5Q;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_D3 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_D4 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_A2 = CLBLM_R_X5Y145_SLICE_X6Y145_CQ;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_A3 = 1'b1;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_A4 = CLBLM_R_X7Y151_SLICE_X9Y151_BQ;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_A5 = 1'b1;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_A6 = 1'b1;
  assign LIOB33_X0Y153_IOB_X0Y154_O = CLBLM_L_X8Y152_SLICE_X10Y152_DQ;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_B1 = CLBLM_L_X8Y147_SLICE_X11Y147_DO6;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_B2 = CLBLM_R_X7Y144_SLICE_X8Y144_CO6;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_B3 = CLBLM_R_X11Y146_SLICE_X15Y146_DO6;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_B4 = CLBLM_R_X7Y144_SLICE_X8Y144_A5Q;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_B5 = CLBLM_L_X10Y148_SLICE_X12Y148_BO5;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_B6 = CLBLM_L_X8Y147_SLICE_X11Y147_CO6;
  assign LIOB33_X0Y153_IOB_X0Y153_O = CLBLM_L_X10Y153_SLICE_X13Y153_AQ;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_C1 = CLBLM_L_X10Y144_SLICE_X12Y144_AO6;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_C2 = CLBLM_R_X7Y148_SLICE_X8Y148_BO5;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_C3 = CLBLM_R_X5Y154_SLICE_X6Y154_AQ;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_C4 = CLBLM_L_X10Y143_SLICE_X12Y143_DO5;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_C5 = CLBLM_L_X8Y149_SLICE_X11Y149_B5Q;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_C6 = CLBLM_L_X10Y146_SLICE_X13Y146_AQ;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_D3 = CLBLM_R_X7Y144_SLICE_X9Y144_C5Q;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_D1 = CLBLM_L_X10Y143_SLICE_X12Y143_AO5;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_D2 = 1'b1;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_D3 = CLBLM_R_X7Y149_SLICE_X9Y149_DQ;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_D4 = CLBLM_L_X8Y148_SLICE_X10Y148_CO6;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_D5 = CLBLM_L_X10Y149_SLICE_X12Y149_CQ;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_D6 = CLBLM_L_X8Y147_SLICE_X10Y147_CO6;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_SR = CLBLM_R_X11Y148_SLICE_X15Y148_AO6;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_A2 = 1'b1;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_A3 = CLBLM_R_X7Y150_SLICE_X9Y150_AQ;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_A4 = CLBLM_R_X5Y154_SLICE_X7Y154_AQ;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_A5 = 1'b1;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_A6 = 1'b1;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_B2 = CLBLM_L_X8Y145_SLICE_X10Y145_BQ;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_B3 = 1'b1;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_B4 = 1'b1;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_B5 = CLBLM_R_X7Y147_SLICE_X8Y147_BQ;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_B6 = 1'b1;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_C1 = 1'b1;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_C1 = CLBLL_L_X4Y144_SLICE_X5Y144_AQ;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_C2 = CLBLM_R_X5Y145_SLICE_X7Y145_BO6;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_C3 = CLBLM_L_X10Y143_SLICE_X12Y143_DO6;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_C4 = CLBLM_L_X8Y147_SLICE_X11Y147_AQ;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_C5 = 1'b1;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_C6 = CLBLM_L_X12Y149_SLICE_X16Y149_CO6;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_D1 = 1'b1;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_D2 = CLBLM_L_X8Y148_SLICE_X10Y148_BQ;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_D3 = CLBLM_R_X5Y145_SLICE_X7Y145_BO6;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_D4 = CLBLM_L_X10Y148_SLICE_X12Y148_BO5;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_D5 = CLBLM_L_X8Y148_SLICE_X10Y148_A5Q;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_D6 = CLBLM_L_X12Y149_SLICE_X16Y149_CO6;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_SR = CLBLM_R_X7Y148_SLICE_X9Y148_DO6;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_A1 = CLBLM_R_X3Y148_SLICE_X2Y148_B5Q;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_A3 = CLBLM_R_X11Y151_SLICE_X15Y151_AQ;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_A4 = CLBLM_R_X5Y151_SLICE_X6Y151_BQ;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_A5 = CLBLM_L_X10Y151_SLICE_X13Y151_DO6;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_A6 = CLBLM_R_X11Y151_SLICE_X15Y151_CO6;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_AX = CLBLM_R_X11Y151_SLICE_X15Y151_CO5;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_C1 = CLBLM_R_X11Y146_SLICE_X14Y146_BO6;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_B1 = CLBLM_R_X3Y148_SLICE_X2Y148_B5Q;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_B2 = CLBLM_R_X11Y151_SLICE_X15Y151_BQ;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_B3 = CLBLM_L_X8Y146_SLICE_X10Y146_A5Q;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_B4 = CLBLM_L_X10Y151_SLICE_X13Y151_CO6;
  assign CLBLL_L_X4Y154_SLICE_X4Y154_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y154_SLICE_X4Y154_A2 = CLBLL_L_X4Y149_SLICE_X5Y149_AQ;
  assign CLBLL_L_X4Y154_SLICE_X4Y154_A3 = CLBLL_L_X4Y154_SLICE_X4Y154_AQ;
  assign CLBLL_L_X4Y154_SLICE_X4Y154_A4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y154_SLICE_X4Y154_A5 = CLBLM_R_X3Y151_SLICE_X3Y151_C5Q;
  assign CLBLL_L_X4Y154_SLICE_X4Y154_A6 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_C3 = 1'b1;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_D3 = 1'b1;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_D4 = 1'b1;
  assign CLBLL_L_X4Y154_SLICE_X4Y154_B1 = CLBLM_R_X3Y153_SLICE_X3Y153_A5Q;
  assign CLBLL_L_X4Y154_SLICE_X4Y154_B2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y154_SLICE_X4Y154_B3 = CLBLL_L_X4Y153_SLICE_X4Y153_CQ;
  assign CLBLL_L_X4Y154_SLICE_X4Y154_B4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y154_SLICE_X4Y154_B5 = CLBLM_R_X3Y150_SLICE_X2Y150_CO5;
  assign CLBLL_L_X4Y154_SLICE_X4Y154_B6 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_A3 = CLBLM_R_X7Y141_SLICE_X9Y141_AQ;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_A4 = CLBLM_L_X8Y148_SLICE_X11Y148_C5Q;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_A6 = CLBLM_R_X3Y148_SLICE_X2Y148_D5Q;
  assign CLBLL_L_X4Y154_SLICE_X4Y154_C1 = 1'b1;
  assign CLBLL_L_X4Y154_SLICE_X4Y154_C2 = 1'b1;
  assign CLBLL_L_X4Y154_SLICE_X4Y154_C3 = 1'b1;
  assign CLBLL_L_X4Y154_SLICE_X4Y154_C4 = 1'b1;
  assign CLBLL_L_X4Y154_SLICE_X4Y154_C5 = 1'b1;
  assign CLBLL_L_X4Y154_SLICE_X4Y154_C6 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_B3 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_B4 = 1'b1;
  assign CLBLL_L_X4Y154_SLICE_X4Y154_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_B6 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_C1 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_C2 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_C3 = 1'b1;
  assign CLBLL_L_X4Y154_SLICE_X4Y154_D1 = 1'b1;
  assign CLBLL_L_X4Y154_SLICE_X4Y154_D2 = 1'b1;
  assign CLBLL_L_X4Y154_SLICE_X4Y154_D3 = 1'b1;
  assign CLBLL_L_X4Y154_SLICE_X4Y154_D4 = 1'b1;
  assign CLBLL_L_X4Y154_SLICE_X4Y154_D5 = 1'b1;
  assign CLBLL_L_X4Y154_SLICE_X4Y154_D6 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_D1 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_D2 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_D3 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_D4 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_D5 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_D6 = 1'b1;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_B1 = CLBLM_R_X3Y148_SLICE_X2Y148_B5Q;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_A1 = CLBLM_R_X5Y149_SLICE_X7Y149_DQ;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_A2 = CLBLM_L_X8Y142_SLICE_X11Y142_CQ;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_A3 = CLBLM_R_X7Y141_SLICE_X8Y141_AQ;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_A4 = CLBLL_L_X4Y140_SLICE_X5Y140_AQ;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_A6 = CLBLM_R_X7Y143_SLICE_X8Y143_BQ;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_C2 = CLBLM_R_X11Y151_SLICE_X15Y151_A5Q;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_C3 = CLBLM_L_X10Y150_SLICE_X13Y150_C5Q;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_C4 = CLBLM_L_X10Y151_SLICE_X13Y151_CO6;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_C5 = CLBLM_R_X11Y151_SLICE_X15Y151_BQ;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_B1 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_B2 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_B3 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_B4 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_B5 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_B6 = 1'b1;
  assign CLBLL_L_X4Y154_SLICE_X5Y154_A1 = 1'b1;
  assign CLBLL_L_X4Y154_SLICE_X5Y154_A2 = 1'b1;
  assign CLBLL_L_X4Y154_SLICE_X5Y154_A3 = 1'b1;
  assign CLBLL_L_X4Y154_SLICE_X5Y154_A4 = CLBLM_R_X5Y153_SLICE_X6Y153_BQ;
  assign CLBLL_L_X4Y154_SLICE_X5Y154_A5 = 1'b1;
  assign CLBLL_L_X4Y154_SLICE_X5Y154_A6 = CLBLL_L_X4Y148_SLICE_X5Y148_CQ;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_C1 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_C2 = 1'b1;
  assign CLBLL_L_X4Y154_SLICE_X5Y154_B1 = 1'b1;
  assign CLBLL_L_X4Y154_SLICE_X5Y154_B2 = 1'b1;
  assign CLBLL_L_X4Y154_SLICE_X5Y154_B3 = 1'b1;
  assign CLBLL_L_X4Y154_SLICE_X5Y154_B4 = 1'b1;
  assign CLBLL_L_X4Y154_SLICE_X5Y154_B5 = 1'b1;
  assign CLBLL_L_X4Y154_SLICE_X5Y154_B6 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_D3 = CLBLM_L_X12Y151_SLICE_X16Y151_AQ;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_C6 = 1'b1;
  assign CLBLL_L_X4Y154_SLICE_X5Y154_C1 = 1'b1;
  assign CLBLL_L_X4Y154_SLICE_X5Y154_C2 = 1'b1;
  assign CLBLL_L_X4Y154_SLICE_X5Y154_C3 = 1'b1;
  assign CLBLL_L_X4Y154_SLICE_X5Y154_C4 = 1'b1;
  assign CLBLL_L_X4Y154_SLICE_X5Y154_C5 = 1'b1;
  assign CLBLL_L_X4Y154_SLICE_X5Y154_C6 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_D4 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_D1 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_D2 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_D3 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_D4 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_D5 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_D6 = 1'b1;
  assign CLBLL_L_X4Y154_SLICE_X5Y154_D1 = 1'b1;
  assign CLBLL_L_X4Y154_SLICE_X5Y154_D2 = 1'b1;
  assign CLBLL_L_X4Y154_SLICE_X5Y154_D3 = 1'b1;
  assign CLBLL_L_X4Y154_SLICE_X5Y154_D4 = 1'b1;
  assign CLBLL_L_X4Y154_SLICE_X5Y154_D5 = 1'b1;
  assign CLBLL_L_X4Y154_SLICE_X5Y154_D6 = 1'b1;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_B1 = CLBLM_L_X10Y153_SLICE_X12Y153_CQ;
  assign LIOI3_X0Y159_OLOGIC_X0Y160_D1 = CLBLL_L_X4Y145_SLICE_X5Y145_AQ;
  assign LIOI3_X0Y159_OLOGIC_X0Y160_T1 = 1'b1;
  assign LIOI3_X0Y159_OLOGIC_X0Y159_D1 = CLBLM_R_X3Y149_SLICE_X2Y149_CQ;
  assign LIOI3_X0Y159_OLOGIC_X0Y159_T1 = 1'b1;
  assign LIOB33_X0Y155_IOB_X0Y156_O = CLBLM_R_X7Y152_SLICE_X9Y152_BQ;
  assign LIOB33_X0Y155_IOB_X0Y155_O = CLBLM_L_X8Y150_SLICE_X11Y150_CQ;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_C1 = CLBLM_L_X8Y152_SLICE_X10Y152_D5Q;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_A1 = CLBLM_R_X5Y149_SLICE_X6Y149_D5Q;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_A2 = CLBLM_L_X8Y146_SLICE_X10Y146_CQ;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_A3 = CLBLM_L_X8Y148_SLICE_X11Y148_AQ;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_A4 = CLBLM_L_X8Y150_SLICE_X11Y150_B5Q;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_A5 = CLBLM_R_X11Y148_SLICE_X15Y148_AQ;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_T1 = 1'b1;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_B1 = CLBLM_L_X8Y151_SLICE_X10Y151_B5Q;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_B2 = CLBLM_L_X8Y152_SLICE_X10Y152_BQ;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_B4 = CLBLM_R_X7Y144_SLICE_X8Y144_A5Q;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_B5 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_B6 = 1'b1;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_C4 = CLBLM_R_X5Y148_SLICE_X6Y148_AO5;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_D1 = CLBLM_L_X12Y151_SLICE_X16Y151_CO5;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_C1 = CLBLL_L_X2Y149_SLICE_X0Y149_AQ;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_C2 = CLBLM_L_X10Y153_SLICE_X12Y153_AQ;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_C3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_C4 = CLBLM_L_X10Y150_SLICE_X13Y150_BQ;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_C5 = CLBLM_R_X7Y145_SLICE_X8Y145_C5Q;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_C6 = 1'b1;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_T1 = 1'b1;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_D1 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_D2 = CLBLM_L_X8Y143_SLICE_X11Y143_A5Q;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_D3 = CLBLM_L_X8Y148_SLICE_X11Y148_DQ;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_D4 = CLBLM_L_X8Y148_SLICE_X11Y148_BQ;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_D5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_D6 = CLBLM_R_X7Y148_SLICE_X8Y148_AQ;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_D1 = CLBLM_R_X11Y153_SLICE_X14Y153_AO5;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_A1 = 1'b1;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_A2 = 1'b1;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_A3 = CLBLM_R_X7Y151_SLICE_X9Y151_AQ;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_A4 = CLBLM_R_X5Y146_SLICE_X7Y146_CQ;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_A6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_T1 = 1'b1;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_B1 = CLBLM_R_X5Y154_SLICE_X7Y154_DQ;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_B2 = CLBLM_L_X8Y150_SLICE_X10Y150_AQ;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_B3 = CLBLM_L_X10Y145_SLICE_X12Y145_AO6;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_B4 = CLBLM_R_X7Y150_SLICE_X8Y150_D5Q;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_B5 = CLBLM_L_X8Y151_SLICE_X10Y151_DQ;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_B6 = 1'b1;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_BX = CLBLM_L_X8Y151_SLICE_X11Y151_BO6;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_C1 = CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_C2 = CLBLM_L_X10Y144_SLICE_X13Y144_CO6;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_C3 = CLBLL_L_X4Y149_SLICE_X4Y149_CQ;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_C4 = CLBLM_L_X8Y150_SLICE_X10Y150_A5Q;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_C5 = CLBLM_R_X11Y149_SLICE_X14Y149_AQ;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_C6 = 1'b1;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_D1 = CLBLL_L_X4Y141_SLICE_X5Y141_AQ;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_D2 = CLBLM_R_X3Y154_SLICE_X3Y154_AQ;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_D3 = CLBLM_R_X5Y151_SLICE_X6Y151_DQ;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_D4 = CLBLM_R_X7Y146_SLICE_X9Y146_AO5;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_D5 = 1'b1;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_D6 = CLBLM_L_X8Y148_SLICE_X10Y148_BO6;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_D3 = CLBLM_L_X8Y153_SLICE_X10Y153_BQ;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_D4 = 1'b1;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_SR = CLBLM_R_X7Y148_SLICE_X9Y148_AO5;
  assign LIOI3_X0Y155_OLOGIC_X0Y156_T1 = 1'b1;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_D6 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_A1 = CLBLM_R_X11Y151_SLICE_X14Y151_DO6;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_A2 = CLBLM_R_X3Y150_SLICE_X3Y150_BQ;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_A3 = CLBLM_L_X12Y151_SLICE_X16Y151_AQ;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_A4 = CLBLM_L_X8Y153_SLICE_X10Y153_AQ;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_A5 = CLBLM_R_X7Y145_SLICE_X8Y145_B5Q;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_A6 = CLBLM_R_X11Y152_SLICE_X14Y152_AQ;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_B1 = CLBLM_L_X12Y151_SLICE_X16Y151_DO6;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_B2 = CLBLM_L_X8Y153_SLICE_X10Y153_AQ;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_B3 = CLBLM_R_X3Y150_SLICE_X3Y150_BQ;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_B4 = CLBLM_L_X12Y151_SLICE_X16Y151_BQ;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_B5 = CLBLM_R_X7Y145_SLICE_X8Y145_B5Q;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_B6 = CLBLM_L_X10Y152_SLICE_X13Y152_AQ;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_A1 = CLBLM_R_X7Y150_SLICE_X9Y150_CQ;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_A2 = CLBLM_L_X10Y146_SLICE_X12Y146_AO5;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_A3 = CLBLM_R_X7Y142_SLICE_X9Y142_AQ;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_A4 = CLBLM_L_X8Y149_SLICE_X11Y149_BQ;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_A6 = CLBLM_R_X7Y147_SLICE_X9Y147_CQ;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_C1 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_C2 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_AX = CLBLM_L_X8Y142_SLICE_X10Y142_BO6;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_D4 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_B1 = CLBLM_L_X10Y152_SLICE_X12Y152_BQ;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_B2 = CLBLM_R_X7Y142_SLICE_X9Y142_BQ;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_B3 = CLBLM_R_X5Y144_SLICE_X6Y144_DQ;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_B4 = CLBLL_L_X4Y142_SLICE_X4Y142_A5Q;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_B6 = CLBLM_R_X3Y148_SLICE_X2Y148_D5Q;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_D5 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_D6 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_C2 = CLBLM_R_X7Y142_SLICE_X9Y142_CQ;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_C3 = CLBLM_R_X7Y150_SLICE_X9Y150_B5Q;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_C4 = CLBLM_R_X7Y142_SLICE_X9Y142_BQ;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_C5 = CLBLM_L_X10Y143_SLICE_X12Y143_BO6;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_C6 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_D3 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_D4 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_A1 = CLBLM_R_X5Y150_SLICE_X7Y150_AQ;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_A3 = CLBLM_R_X11Y152_SLICE_X15Y152_AO6;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_A4 = CLBLM_R_X11Y152_SLICE_X14Y152_BO6;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_D1 = CLBLM_R_X5Y142_SLICE_X6Y142_C5Q;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_D2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_D3 = CLBLM_R_X7Y142_SLICE_X9Y142_DQ;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_D4 = CLBLM_R_X7Y142_SLICE_X9Y142_AQ;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_D5 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_D6 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_A5 = CLBLM_R_X11Y150_SLICE_X14Y150_AQ;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_A6 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_B1 = CLBLM_L_X10Y153_SLICE_X12Y153_DO6;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_B2 = CLBLM_L_X8Y153_SLICE_X10Y153_AQ;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_B3 = CLBLM_R_X11Y151_SLICE_X14Y151_AQ;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_A1 = CLBLM_R_X7Y142_SLICE_X8Y142_B5Q;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_A2 = CLBLM_R_X7Y142_SLICE_X8Y142_BQ;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_A3 = CLBLM_R_X7Y148_SLICE_X8Y148_DO6;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_A4 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_A5 = CLBLM_R_X7Y142_SLICE_X8Y142_A5Q;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_A6 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_C1 = CLBLM_L_X12Y151_SLICE_X16Y151_AQ;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_C2 = CLBLM_R_X11Y152_SLICE_X14Y152_AQ;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_C3 = CLBLM_L_X10Y153_SLICE_X12Y153_DO6;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_B1 = CLBLM_R_X7Y142_SLICE_X8Y142_B5Q;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_B2 = CLBLM_R_X7Y142_SLICE_X8Y142_BQ;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_B3 = CLBLM_R_X7Y148_SLICE_X8Y148_DO6;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_B4 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_B5 = CLBLM_R_X7Y142_SLICE_X8Y142_A5Q;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_B6 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_D1 = CLBLM_L_X12Y151_SLICE_X16Y151_AQ;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_D2 = CLBLM_L_X10Y152_SLICE_X12Y152_BQ;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_C1 = CLBLM_R_X7Y142_SLICE_X9Y142_AQ;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_C2 = CLBLM_R_X5Y142_SLICE_X6Y142_AQ;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_C3 = CLBLM_L_X10Y149_SLICE_X12Y149_A5Q;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_C4 = CLBLM_R_X11Y146_SLICE_X15Y146_AQ;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_C5 = CLBLM_R_X5Y146_SLICE_X7Y146_AQ;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_C6 = CLBLM_R_X5Y144_SLICE_X7Y144_BQ;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_D3 = CLBLM_R_X11Y152_SLICE_X14Y152_AQ;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_D4 = CLBLM_L_X10Y152_SLICE_X13Y152_AQ;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_D5 = CLBLM_R_X11Y151_SLICE_X14Y151_DO6;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_D6 = CLBLM_L_X12Y151_SLICE_X16Y151_BQ;
  assign LIOI3_X0Y155_OLOGIC_X0Y155_T1 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_D1 = CLBLM_L_X10Y149_SLICE_X12Y149_A5Q;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_D2 = CLBLM_R_X5Y142_SLICE_X6Y142_AQ;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_D3 = CLBLM_R_X7Y142_SLICE_X9Y142_AQ;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_D4 = CLBLM_R_X11Y146_SLICE_X15Y146_AQ;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_D5 = CLBLM_R_X5Y146_SLICE_X7Y146_AQ;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_D6 = CLBLM_R_X5Y144_SLICE_X7Y144_BQ;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_C2 = CLBLM_R_X5Y142_SLICE_X7Y142_BQ;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_C3 = CLBLM_L_X8Y151_SLICE_X10Y151_CO5;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_C4 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_C5 = CLBLM_R_X5Y151_SLICE_X7Y151_BO5;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_B1 = CLBLM_L_X10Y145_SLICE_X13Y145_CO6;
  assign LIOB33_X0Y157_IOB_X0Y158_O = RIOB33_X105Y133_IOB_X1Y134_I;
  assign LIOB33_X0Y157_IOB_X0Y157_O = CLBLM_R_X7Y153_SLICE_X9Y153_CQ;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_C6 = 1'b1;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_B2 = CLBLM_R_X11Y147_SLICE_X14Y147_BO6;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_D1 = CLBLM_R_X3Y152_SLICE_X2Y152_BQ;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_A1 = CLBLM_R_X3Y148_SLICE_X2Y148_D5Q;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_A2 = CLBLM_L_X8Y145_SLICE_X10Y145_BQ;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_A3 = CLBLM_L_X8Y149_SLICE_X11Y149_AQ;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_A5 = CLBLM_R_X5Y144_SLICE_X6Y144_DQ;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_A6 = CLBLM_R_X7Y151_SLICE_X9Y151_CQ;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_D2 = CLBLM_L_X8Y152_SLICE_X11Y152_CO6;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_B1 = CLBLL_L_X4Y149_SLICE_X5Y149_CQ;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_B2 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_B3 = CLBLM_L_X8Y147_SLICE_X10Y147_AQ;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_B4 = CLBLM_L_X8Y149_SLICE_X11Y149_CQ;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_B6 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_D3 = CLBLM_R_X7Y151_SLICE_X9Y151_DQ;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_D4 = CLBLM_L_X8Y151_SLICE_X10Y151_DQ;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_C2 = CLBLL_L_X2Y151_SLICE_X1Y151_BQ;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_C3 = CLBLM_L_X8Y147_SLICE_X11Y147_AQ;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_C4 = 1'b1;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_C5 = CLBLM_R_X7Y151_SLICE_X9Y151_CQ;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_C6 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_D5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_D6 = CLBLM_R_X7Y147_SLICE_X8Y147_AQ;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_D1 = 1'b1;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_D2 = CLBLM_L_X8Y149_SLICE_X10Y149_CO6;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_D3 = CLBLM_L_X8Y150_SLICE_X10Y150_AQ;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_D4 = CLBLM_R_X7Y149_SLICE_X9Y149_BO6;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_D5 = CLBLM_L_X10Y145_SLICE_X12Y145_AO6;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_D6 = CLBLM_R_X11Y143_SLICE_X14Y143_CO5;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_A1 = 1'b1;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_A3 = CLBLM_R_X7Y149_SLICE_X9Y149_DQ;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_A4 = 1'b1;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_A5 = CLBLM_R_X5Y144_SLICE_X7Y144_CQ;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_A6 = 1'b1;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_B1 = 1'b1;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_B2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_B3 = CLBLM_R_X7Y146_SLICE_X9Y146_BQ;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_B4 = 1'b1;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_B5 = CLBLL_L_X2Y147_SLICE_X1Y147_AQ;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_B6 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_A1 = CLBLM_R_X5Y143_SLICE_X6Y143_CQ;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_C1 = CLBLM_L_X8Y150_SLICE_X11Y150_BQ;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_C2 = CLBLM_L_X10Y148_SLICE_X12Y148_BO5;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_C3 = CLBLM_R_X7Y149_SLICE_X9Y149_CQ;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_C4 = CLBLM_L_X8Y148_SLICE_X10Y148_CO6;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_C5 = CLBLM_L_X10Y144_SLICE_X12Y144_AO6;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_C6 = CLBLM_R_X5Y150_SLICE_X7Y150_A5Q;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_A2 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_A3 = 1'b1;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_A4 = CLBLM_L_X8Y146_SLICE_X11Y146_A5Q;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_D1 = CLBLM_L_X8Y146_SLICE_X10Y146_C5Q;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_D2 = CLBLM_L_X10Y144_SLICE_X12Y144_AO6;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_D3 = CLBLM_L_X10Y148_SLICE_X12Y148_BO5;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_D4 = CLBLM_L_X8Y148_SLICE_X10Y148_CO6;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_D5 = CLBLM_L_X8Y149_SLICE_X10Y149_B5Q;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_D6 = CLBLL_L_X4Y150_SLICE_X4Y150_AQ;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_A6 = CLBLM_R_X7Y144_SLICE_X9Y144_AQ;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_SR = CLBLM_R_X11Y148_SLICE_X14Y148_DO6;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_C4 = CLBLM_R_X7Y153_SLICE_X8Y153_DO5;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_C5 = CLBLM_R_X7Y154_SLICE_X9Y154_AO6;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_B1 = CLBLM_R_X5Y153_SLICE_X6Y153_AQ;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_C6 = CLBLL_L_X4Y154_SLICE_X4Y154_BO6;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_B2 = CLBLM_R_X7Y151_SLICE_X8Y151_BQ;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_A1 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_A2 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_A3 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_A4 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_B3 = CLBLM_R_X5Y153_SLICE_X7Y153_AQ;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_A5 = 1'b1;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_SR = CLBLM_R_X11Y148_SLICE_X14Y148_DO6;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_A6 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_B4 = CLBLM_R_X3Y148_SLICE_X2Y148_D5Q;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_B1 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_B2 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_B3 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_B4 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_B5 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_B6 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_B6 = CLBLM_R_X5Y144_SLICE_X6Y144_DQ;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_A1 = CLBLM_L_X8Y142_SLICE_X10Y142_CQ;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_A2 = CLBLM_R_X3Y147_SLICE_X3Y147_BQ;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_A3 = CLBLM_R_X7Y143_SLICE_X9Y143_AQ;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_A4 = CLBLM_R_X5Y144_SLICE_X6Y144_CQ;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_A6 = CLBLM_R_X5Y141_SLICE_X7Y141_A5Q;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_C1 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_C2 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_C3 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_B1 = CLBLM_R_X7Y144_SLICE_X8Y144_BO6;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_B2 = CLBLM_R_X7Y143_SLICE_X9Y143_BQ;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_B4 = CLBLL_L_X2Y148_SLICE_X0Y148_B5Q;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_B5 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_B6 = CLBLM_L_X8Y143_SLICE_X10Y143_BQ;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_D1 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_D2 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_C2 = CLBLM_R_X7Y143_SLICE_X9Y143_CQ;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_C3 = CLBLL_L_X4Y144_SLICE_X5Y144_B5Q;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_C4 = CLBLM_R_X7Y143_SLICE_X9Y143_BQ;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_C5 = CLBLM_R_X7Y144_SLICE_X8Y144_BO6;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_C6 = CLBLL_L_X2Y148_SLICE_X0Y148_B5Q;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_D3 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_D4 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_A1 = CLBLM_L_X10Y145_SLICE_X13Y145_CO6;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_A2 = CLBLM_R_X3Y151_SLICE_X3Y151_D5Q;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_A3 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_A4 = CLBLM_L_X10Y148_SLICE_X13Y148_CO6;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_D2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_D1 = CLBLM_L_X10Y142_SLICE_X13Y142_AQ;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_D2 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_D3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_D4 = CLBLM_R_X7Y143_SLICE_X9Y143_BQ;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_D5 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_D6 = CLBLM_R_X5Y148_SLICE_X6Y148_BQ;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_C3 = CLBLM_L_X10Y150_SLICE_X13Y150_A5Q;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_A6 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_C4 = CLBLM_R_X3Y151_SLICE_X3Y151_AQ;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_B1 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_B2 = 1'b1;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_D5 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_A2 = CLBLM_R_X7Y142_SLICE_X9Y142_BQ;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_A3 = CLBLM_R_X7Y143_SLICE_X8Y143_AQ;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_A4 = CLBLL_L_X2Y144_SLICE_X1Y144_AQ;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_D6 = CLBLM_R_X3Y151_SLICE_X3Y151_BQ;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_A5 = CLBLM_R_X5Y144_SLICE_X6Y144_CQ;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_A6 = CLBLM_R_X3Y147_SLICE_X3Y147_BQ;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_C5 = CLBLM_R_X5Y147_SLICE_X7Y147_BQ;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_C6 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_B2 = CLBLM_R_X7Y143_SLICE_X8Y143_BQ;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_B3 = CLBLM_R_X7Y142_SLICE_X8Y142_AQ;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_B4 = CLBLM_R_X7Y150_SLICE_X8Y150_C5Q;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_B5 = CLBLM_R_X7Y141_SLICE_X9Y141_AQ;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_B6 = CLBLM_L_X10Y143_SLICE_X12Y143_BO6;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_D1 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_D2 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_C1 = CLBLM_L_X10Y143_SLICE_X12Y143_AO6;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_C2 = CLBLM_R_X7Y143_SLICE_X8Y143_CQ;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_C3 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_SR = CLBLL_L_X2Y147_SLICE_X1Y147_BO6;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_C4 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_C5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_C6 = CLBLM_R_X5Y143_SLICE_X6Y143_BQ;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_D3 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_D4 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_D6 = 1'b1;
  assign LIOB33_X0Y159_IOB_X0Y160_O = CLBLL_L_X4Y145_SLICE_X5Y145_AQ;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_D1 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_D2 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_D3 = CLBLM_R_X7Y143_SLICE_X8Y143_DQ;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_D4 = CLBLM_R_X3Y144_SLICE_X2Y144_A5Q;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_D5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_D6 = CLBLM_L_X10Y143_SLICE_X12Y143_BO5;
  assign LIOB33_X0Y159_IOB_X0Y159_O = CLBLM_R_X3Y149_SLICE_X2Y149_CQ;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_D3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_D4 = CLBLM_R_X5Y152_SLICE_X6Y152_DQ;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_D5 = CLBLM_R_X5Y152_SLICE_X7Y152_D5Q;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_D6 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_A1 = CLBLM_L_X8Y150_SLICE_X11Y150_B5Q;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_A2 = CLBLM_R_X5Y149_SLICE_X6Y149_D5Q;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_A3 = CLBLM_L_X8Y150_SLICE_X11Y150_AQ;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_A4 = CLBLM_R_X5Y151_SLICE_X7Y151_AQ;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_A5 = CLBLM_L_X8Y147_SLICE_X10Y147_A5Q;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_B6 = CLBLM_R_X5Y152_SLICE_X6Y152_B5Q;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_B1 = CLBLM_L_X8Y152_SLICE_X11Y152_A5Q;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_B2 = CLBLM_R_X7Y151_SLICE_X8Y151_BQ;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_B3 = CLBLM_R_X7Y153_SLICE_X9Y153_CQ;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_B5 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_B6 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_C1 = CLBLM_L_X8Y149_SLICE_X10Y149_B5Q;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_C2 = CLBLM_R_X3Y154_SLICE_X3Y154_AQ;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_C3 = CLBLM_R_X7Y154_SLICE_X8Y154_CQ;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_C4 = CLBLM_L_X8Y151_SLICE_X11Y151_CO6;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_C5 = CLBLM_L_X8Y150_SLICE_X11Y150_DO6;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_C6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_D1 = CLBLM_L_X8Y154_SLICE_X10Y154_AQ;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_D2 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_D3 = CLBLM_R_X7Y146_SLICE_X9Y146_DO6;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_D4 = CLBLM_L_X10Y146_SLICE_X13Y146_AQ;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_D5 = CLBLM_R_X5Y145_SLICE_X7Y145_AQ;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_D6 = CLBLM_R_X7Y152_SLICE_X8Y152_CQ;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_A1 = CLBLM_L_X8Y142_SLICE_X10Y142_A5Q;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_A1 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_A2 = CLBLM_L_X8Y145_SLICE_X10Y145_AQ;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_A3 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_A5 = CLBLM_R_X3Y153_SLICE_X3Y153_AQ;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_A6 = 1'b1;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_C4 = CLBLM_R_X5Y152_SLICE_X6Y152_B5Q;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_C5 = CLBLM_R_X5Y152_SLICE_X7Y152_DQ;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign LIOI3_X0Y161_OLOGIC_X0Y162_D1 = CLBLM_R_X3Y153_SLICE_X3Y153_CO6;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_B1 = CLBLM_L_X10Y143_SLICE_X12Y143_BO5;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_B2 = CLBLM_R_X7Y148_SLICE_X8Y148_CO6;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_B3 = CLBLM_L_X8Y152_SLICE_X10Y152_AQ;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_B4 = CLBLM_R_X5Y150_SLICE_X7Y150_DO6;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_B5 = CLBLM_L_X8Y146_SLICE_X11Y146_CO6;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_B6 = CLBLM_L_X8Y150_SLICE_X10Y150_CO6;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_C6 = CLBLM_L_X8Y150_SLICE_X11Y150_BQ;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_A5 = CLBLM_R_X5Y144_SLICE_X6Y144_DQ;
  assign LIOI3_X0Y161_OLOGIC_X0Y162_T1 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_C1 = CLBLM_L_X12Y149_SLICE_X16Y149_CO6;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_C2 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_C3 = CLBLM_L_X10Y143_SLICE_X12Y143_BO6;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_C4 = CLBLM_L_X8Y152_SLICE_X10Y152_CQ;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_C5 = CLBLM_R_X7Y146_SLICE_X8Y146_AO6;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_C6 = CLBLM_L_X8Y149_SLICE_X10Y149_BQ;
  assign LIOI3_X0Y101_OLOGIC_X0Y102_D1 = CLBLM_R_X5Y140_SLICE_X7Y140_BQ;
  assign LIOI3_X0Y161_OLOGIC_X0Y161_D1 = CLBLM_R_X5Y151_SLICE_X6Y151_CQ;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign LIOI3_X0Y101_OLOGIC_X0Y102_T1 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_D1 = CLBLM_R_X7Y149_SLICE_X9Y149_DO6;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_D2 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_D3 = CLBLM_L_X8Y149_SLICE_X10Y149_DO6;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_D4 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_D5 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_D6 = 1'b1;
  assign LIOI3_X0Y161_OLOGIC_X0Y161_T1 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_B1 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_SR = CLBLM_R_X11Y148_SLICE_X15Y148_CO6;
  assign LIOI3_X0Y101_OLOGIC_X0Y101_D1 = CLBLM_R_X3Y142_SLICE_X2Y142_B5Q;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_B2 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y63_OLOGIC_X0Y64_D1 = CLBLL_L_X4Y140_SLICE_X5Y140_BO6;
  assign LIOI3_X0Y101_OLOGIC_X0Y101_T1 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_B5 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y63_OLOGIC_X0Y64_T1 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_A1 = CLBLM_R_X7Y142_SLICE_X9Y142_DQ;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_A2 = CLBLL_L_X2Y148_SLICE_X0Y148_B5Q;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_A3 = CLBLM_R_X7Y144_SLICE_X9Y144_AQ;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_A4 = CLBLM_R_X7Y152_SLICE_X8Y152_BQ;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_A5 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_AX = CLBLM_R_X7Y151_SLICE_X8Y151_DO6;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_B1 = CLBLM_L_X8Y143_SLICE_X11Y143_CQ;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_B2 = CLBLM_R_X7Y144_SLICE_X9Y144_BQ;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_B3 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_B4 = CLBLM_L_X8Y148_SLICE_X11Y148_B5Q;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_C4 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_B6 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_C5 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_C1 = CLBLM_R_X7Y142_SLICE_X9Y142_D5Q;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_C2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_C3 = CLBLM_L_X10Y149_SLICE_X13Y149_AQ;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_C4 = CLBLM_L_X10Y147_SLICE_X12Y147_CQ;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_C6 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_C5 = CLBLM_R_X7Y152_SLICE_X8Y152_BQ;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_C6 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_D1 = CLBLM_R_X3Y150_SLICE_X3Y150_BQ;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_D2 = CLBLM_R_X11Y147_SLICE_X15Y147_AQ;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_D3 = CLBLM_R_X7Y146_SLICE_X9Y146_B5Q;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_D4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_D5 = CLBLM_L_X8Y143_SLICE_X10Y143_DQ;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_D6 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_A1 = CLBLM_R_X5Y150_SLICE_X6Y150_CQ;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_A3 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_A4 = CLBLM_L_X8Y144_SLICE_X10Y144_AQ;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_A5 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_A6 = 1'b1;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_C5 = CLBLM_R_X3Y152_SLICE_X2Y152_BQ;
  assign LIOB33_X0Y161_IOB_X0Y161_O = CLBLM_R_X5Y151_SLICE_X6Y151_CQ;
  assign LIOB33_X0Y161_IOB_X0Y162_O = CLBLM_R_X3Y153_SLICE_X3Y153_CO6;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_B1 = CLBLM_R_X3Y152_SLICE_X3Y152_AQ;
  assign CLBLL_L_X2Y143_SLICE_X0Y143_A1 = 1'b1;
  assign CLBLL_L_X2Y143_SLICE_X0Y143_A2 = 1'b1;
  assign CLBLL_L_X2Y143_SLICE_X0Y143_A3 = 1'b1;
  assign CLBLL_L_X2Y143_SLICE_X0Y143_A4 = 1'b1;
  assign CLBLL_L_X2Y143_SLICE_X0Y143_A5 = 1'b1;
  assign CLBLL_L_X2Y143_SLICE_X0Y143_A6 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_B2 = CLBLM_R_X7Y152_SLICE_X8Y152_BQ;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_B3 = CLBLM_R_X3Y144_SLICE_X3Y144_CQ;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_B4 = CLBLL_L_X4Y151_SLICE_X5Y151_AQ;
  assign CLBLL_L_X2Y143_SLICE_X0Y143_B1 = 1'b1;
  assign CLBLL_L_X2Y143_SLICE_X0Y143_B2 = 1'b1;
  assign CLBLL_L_X2Y143_SLICE_X0Y143_B3 = 1'b1;
  assign CLBLL_L_X2Y143_SLICE_X0Y143_B4 = 1'b1;
  assign CLBLL_L_X2Y143_SLICE_X0Y143_B5 = 1'b1;
  assign CLBLL_L_X2Y143_SLICE_X0Y143_B6 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_BX = CLBLM_L_X8Y142_SLICE_X10Y142_DO5;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_C1 = CLBLM_R_X7Y144_SLICE_X8Y144_BQ;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_A2 = CLBLM_R_X3Y144_SLICE_X3Y144_CQ;
  assign CLBLL_L_X2Y143_SLICE_X0Y143_C1 = 1'b1;
  assign CLBLL_L_X2Y143_SLICE_X0Y143_C2 = 1'b1;
  assign CLBLL_L_X2Y143_SLICE_X0Y143_C3 = 1'b1;
  assign CLBLL_L_X2Y143_SLICE_X0Y143_C4 = 1'b1;
  assign CLBLL_L_X2Y143_SLICE_X0Y143_C5 = 1'b1;
  assign CLBLL_L_X2Y143_SLICE_X0Y143_C6 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_A4 = CLBLM_R_X5Y143_SLICE_X6Y143_BQ;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_D1 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_D2 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_D3 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_D4 = CLBLM_R_X7Y143_SLICE_X9Y143_CQ;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_D5 = 1'b1;
  assign CLBLL_L_X2Y143_SLICE_X0Y143_D1 = 1'b1;
  assign CLBLL_L_X2Y143_SLICE_X0Y143_D2 = 1'b1;
  assign CLBLL_L_X2Y143_SLICE_X0Y143_D3 = 1'b1;
  assign CLBLL_L_X2Y143_SLICE_X0Y143_D4 = 1'b1;
  assign CLBLL_L_X2Y143_SLICE_X0Y143_D5 = 1'b1;
  assign CLBLL_L_X2Y143_SLICE_X0Y143_D6 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_SR = CLBLM_R_X11Y148_SLICE_X15Y148_AO6;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_B2 = CLBLM_R_X7Y143_SLICE_X9Y143_BQ;
  assign CLBLL_L_X2Y143_SLICE_X1Y143_A1 = CLBLM_R_X3Y148_SLICE_X2Y148_D5Q;
  assign CLBLL_L_X2Y143_SLICE_X1Y143_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X2Y143_SLICE_X1Y143_A3 = CLBLL_L_X2Y143_SLICE_X1Y143_AQ;
  assign CLBLL_L_X2Y143_SLICE_X1Y143_A4 = CLBLM_R_X3Y150_SLICE_X3Y150_BQ;
  assign CLBLL_L_X2Y143_SLICE_X1Y143_A5 = CLBLM_R_X5Y144_SLICE_X6Y144_DQ;
  assign CLBLL_L_X2Y143_SLICE_X1Y143_A6 = CLBLL_L_X4Y148_SLICE_X4Y148_A5Q;
  assign CLBLL_L_X2Y143_SLICE_X1Y143_B1 = CLBLM_R_X7Y152_SLICE_X8Y152_BQ;
  assign CLBLL_L_X2Y143_SLICE_X1Y143_B2 = 1'b1;
  assign CLBLL_L_X2Y143_SLICE_X1Y143_B3 = 1'b1;
  assign CLBLL_L_X2Y143_SLICE_X1Y143_B4 = CLBLL_L_X4Y143_SLICE_X4Y143_DQ;
  assign CLBLL_L_X2Y143_SLICE_X1Y143_B5 = CLBLL_L_X4Y144_SLICE_X5Y144_D5Q;
  assign CLBLL_L_X2Y143_SLICE_X1Y143_B6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign RIOI3_X105Y145_ILOGIC_X1Y146_D = RIOB33_X105Y145_IOB_X1Y146_I;
  assign RIOI3_X105Y145_ILOGIC_X1Y145_D = RIOB33_X105Y145_IOB_X1Y145_I;
  assign CLBLL_L_X2Y143_SLICE_X1Y143_C1 = LIOB33_X0Y57_IOB_X0Y58_I;
  assign CLBLL_L_X2Y143_SLICE_X1Y143_C2 = CLBLL_L_X2Y143_SLICE_X1Y143_CQ;
  assign CLBLL_L_X2Y143_SLICE_X1Y143_C3 = CLBLL_L_X2Y143_SLICE_X1Y143_DQ;
  assign CLBLL_L_X2Y143_SLICE_X1Y143_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X2Y143_SLICE_X1Y143_C5 = 1'b1;
  assign CLBLL_L_X2Y143_SLICE_X1Y143_C6 = 1'b1;
  assign CLBLL_L_X2Y143_SLICE_X1Y143_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y63_D = LIOB33_X0Y63_IOB_X0Y63_I;
  assign CLBLL_L_X2Y143_SLICE_X1Y143_D1 = CLBLL_L_X2Y144_SLICE_X1Y144_AQ;
  assign CLBLL_L_X2Y143_SLICE_X1Y143_D2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X2Y143_SLICE_X1Y143_D3 = CLBLL_L_X2Y143_SLICE_X1Y143_DQ;
  assign CLBLL_L_X2Y143_SLICE_X1Y143_D4 = 1'b1;
  assign CLBLL_L_X2Y143_SLICE_X1Y143_D5 = CLBLM_L_X10Y143_SLICE_X12Y143_BO5;
  assign CLBLL_L_X2Y143_SLICE_X1Y143_D6 = CLBLM_R_X3Y144_SLICE_X3Y144_BQ;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_A1 = CLBLM_R_X7Y149_SLICE_X9Y149_CQ;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_A3 = 1'b1;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_A4 = CLBLM_R_X5Y141_SLICE_X7Y141_A5Q;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_A5 = 1'b1;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_A6 = 1'b1;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_B1 = CLBLM_R_X7Y151_SLICE_X8Y151_CQ;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_B2 = CLBLM_L_X8Y153_SLICE_X11Y153_BQ;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_B3 = CLBLM_L_X8Y150_SLICE_X11Y150_BQ;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_B4 = CLBLM_R_X5Y154_SLICE_X7Y154_DQ;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_B6 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_C4 = 1'b1;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_C1 = CLBLM_L_X8Y148_SLICE_X10Y148_AQ;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_C2 = CLBLM_L_X8Y151_SLICE_X11Y151_DO6;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_C3 = CLBLM_L_X8Y140_SLICE_X10Y140_A5Q;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_C4 = CLBLM_R_X7Y151_SLICE_X9Y151_DQ;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_C5 = CLBLM_L_X8Y151_SLICE_X11Y151_BO5;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_C6 = CLBLM_R_X5Y151_SLICE_X6Y151_DQ;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_C5 = CLBLM_R_X7Y143_SLICE_X9Y143_CQ;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_C6 = 1'b1;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_D1 = CLBLM_R_X7Y148_SLICE_X8Y148_AQ;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_D2 = 1'b1;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_D3 = CLBLM_R_X7Y154_SLICE_X8Y154_CQ;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_D4 = CLBLM_R_X5Y148_SLICE_X6Y148_B5Q;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_D5 = CLBLM_L_X8Y151_SLICE_X10Y151_DQ;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_D6 = 1'b1;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_SR = CLBLM_R_X11Y150_SLICE_X14Y150_DO6;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_A1 = CLBLL_L_X4Y148_SLICE_X4Y148_AQ;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_A2 = CLBLM_L_X10Y152_SLICE_X12Y152_AQ;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_A3 = CLBLM_L_X8Y151_SLICE_X10Y151_AQ;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_A4 = CLBLM_R_X3Y147_SLICE_X3Y147_BQ;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_A5 = CLBLM_R_X5Y144_SLICE_X6Y144_CQ;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_B1 = 1'b1;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_B2 = CLBLM_L_X8Y146_SLICE_X10Y146_C5Q;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_B3 = CLBLM_R_X7Y148_SLICE_X9Y148_C5Q;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_B5 = CLBLM_R_X11Y151_SLICE_X14Y151_AQ;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_B6 = 1'b1;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_C2 = CLBLM_R_X5Y153_SLICE_X6Y153_AQ;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_C3 = CLBLM_R_X7Y143_SLICE_X9Y143_BQ;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_C4 = CLBLL_L_X4Y150_SLICE_X5Y150_CQ;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_C5 = CLBLM_R_X3Y151_SLICE_X3Y151_AQ;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_C6 = 1'b1;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_D1 = CLBLM_R_X3Y152_SLICE_X2Y152_BQ;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_D2 = CLBLM_L_X8Y146_SLICE_X10Y146_A5Q;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_D3 = CLBLM_L_X8Y151_SLICE_X10Y151_DQ;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_D4 = CLBLM_L_X8Y152_SLICE_X11Y152_CO6;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_D5 = 1'b1;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_D6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_C3 = 1'b1;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_A1 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_C4 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_C5 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_A1 = CLBLM_L_X10Y143_SLICE_X12Y143_BO5;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_A2 = 1'b1;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_A3 = CLBLM_R_X7Y145_SLICE_X9Y145_AQ;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_A4 = CLBLM_R_X7Y145_SLICE_X9Y145_CQ;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_A5 = CLBLM_R_X7Y145_SLICE_X8Y145_AQ;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_B1 = CLBLM_R_X7Y153_SLICE_X8Y153_AQ;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_B2 = CLBLM_R_X7Y145_SLICE_X9Y145_BQ;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_B3 = CLBLM_R_X7Y145_SLICE_X9Y145_AQ;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_B4 = CLBLM_R_X5Y149_SLICE_X7Y149_DQ;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_B5 = CLBLM_L_X8Y142_SLICE_X11Y142_CQ;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_B6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_C1 = CLBLM_L_X8Y150_SLICE_X11Y150_B5Q;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_C2 = CLBLM_R_X7Y145_SLICE_X9Y145_CQ;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_C3 = CLBLM_R_X3Y146_SLICE_X3Y146_AQ;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_C5 = CLBLM_R_X5Y149_SLICE_X6Y149_D5Q;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_C6 = CLBLM_L_X8Y145_SLICE_X10Y145_AQ;
  assign LIOB33_X0Y163_IOB_X0Y163_O = CLBLM_R_X5Y159_SLICE_X6Y159_AO6;
  assign LIOB33_X0Y163_IOB_X0Y164_O = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_D1 = CLBLM_R_X5Y145_SLICE_X6Y145_AQ;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_D2 = CLBLM_L_X10Y146_SLICE_X12Y146_BO6;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_D3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_D4 = CLBLM_R_X7Y149_SLICE_X9Y149_CO6;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_D5 = CLBLM_R_X7Y147_SLICE_X9Y147_DO6;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_D6 = CLBLM_L_X8Y145_SLICE_X10Y145_BO6;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_A1 = CLBLM_R_X7Y145_SLICE_X8Y145_B5Q;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_A2 = CLBLM_R_X5Y144_SLICE_X6Y144_CQ;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_A3 = CLBLM_R_X7Y145_SLICE_X8Y145_AQ;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_A4 = CLBLM_L_X8Y142_SLICE_X10Y142_CQ;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_A6 = CLBLM_R_X3Y147_SLICE_X3Y147_BQ;
  assign CLBLL_L_X2Y144_SLICE_X0Y144_A1 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X0Y144_A2 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X0Y144_A3 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X0Y144_A4 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X0Y144_A5 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X0Y144_A6 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X0Y144_AX = CLBLM_R_X3Y144_SLICE_X2Y144_BO6;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X2Y144_SLICE_X0Y144_B1 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X0Y144_B2 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X0Y144_B3 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X0Y144_B4 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X0Y144_B5 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X0Y144_B6 = 1'b1;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_C2 = CLBLM_R_X3Y143_SLICE_X2Y143_CQ;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_C3 = CLBLM_R_X7Y145_SLICE_X8Y145_DQ;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_C4 = CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  assign CLBLL_L_X2Y144_SLICE_X0Y144_C1 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X0Y144_C2 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X0Y144_C3 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X0Y144_C4 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X0Y144_C5 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X0Y144_C6 = 1'b1;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_C5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_C6 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X0Y144_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_D1 = CLBLM_R_X7Y143_SLICE_X8Y143_AQ;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_D2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_D3 = CLBLM_R_X7Y145_SLICE_X8Y145_DQ;
  assign CLBLL_L_X2Y144_SLICE_X0Y144_D1 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X0Y144_D2 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X0Y144_D3 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X0Y144_D4 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X0Y144_D5 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X0Y144_D6 = 1'b1;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_D4 = CLBLM_L_X10Y143_SLICE_X12Y143_BO6;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_D5 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X0Y144_SR = CLBLM_R_X7Y144_SLICE_X8Y144_DO6;
  assign CLBLL_L_X2Y144_SLICE_X1Y144_A1 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X1Y144_A2 = CLBLM_R_X5Y142_SLICE_X7Y142_B5Q;
  assign CLBLL_L_X2Y144_SLICE_X1Y144_A3 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X1Y144_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X2Y144_SLICE_X1Y144_A5 = CLBLM_R_X3Y145_SLICE_X2Y145_DQ;
  assign CLBLL_L_X2Y144_SLICE_X1Y144_A6 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_C5 = CLBLL_L_X4Y143_SLICE_X5Y143_CQ;
  assign CLBLL_L_X2Y144_SLICE_X1Y144_B1 = LIOB33_X0Y63_IOB_X0Y63_I;
  assign CLBLL_L_X2Y144_SLICE_X1Y144_B2 = CLBLM_R_X3Y144_SLICE_X2Y144_AQ;
  assign CLBLL_L_X2Y144_SLICE_X1Y144_B3 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X1Y144_B4 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X1Y144_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X2Y144_SLICE_X1Y144_B6 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_C6 = CLBLM_R_X3Y147_SLICE_X3Y147_BQ;
  assign CLBLL_L_X2Y144_SLICE_X1Y144_C1 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X1Y144_C2 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X1Y144_C3 = CLBLM_R_X5Y144_SLICE_X7Y144_CQ;
  assign CLBLL_L_X2Y144_SLICE_X1Y144_C4 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X1Y144_C5 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X1Y144_C6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X2Y144_SLICE_X1Y144_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y144_SLICE_X1Y144_D1 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X1Y144_D2 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X1Y144_D3 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X1Y144_D4 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X1Y144_D5 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X1Y144_D6 = 1'b1;
  assign CLBLL_L_X2Y144_SLICE_X1Y144_SR = CLBLL_L_X2Y144_SLICE_X1Y144_CO6;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_A1 = CLBLM_L_X10Y145_SLICE_X13Y145_CO6;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_A2 = CLBLM_L_X8Y140_SLICE_X10Y140_A5Q;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_A3 = CLBLL_L_X4Y152_SLICE_X4Y152_AQ;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_A5 = CLBLM_L_X10Y148_SLICE_X13Y148_CO6;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_A6 = 1'b1;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_B1 = CLBLM_L_X8Y152_SLICE_X11Y152_DO6;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_B2 = CLBLL_L_X2Y148_SLICE_X0Y148_A5Q;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_B3 = CLBLL_L_X4Y144_SLICE_X5Y144_C5Q;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_B5 = CLBLM_L_X8Y153_SLICE_X11Y153_CO6;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_B6 = 1'b1;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_C1 = CLBLM_L_X8Y154_SLICE_X10Y154_AQ;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_C2 = CLBLM_R_X3Y154_SLICE_X3Y154_AQ;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_C3 = CLBLM_L_X8Y153_SLICE_X11Y153_BQ;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_C4 = CLBLM_R_X5Y154_SLICE_X7Y154_DQ;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_C5 = CLBLM_R_X7Y154_SLICE_X8Y154_CQ;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_C6 = CLBLM_R_X7Y152_SLICE_X8Y152_CQ;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_D1 = CLBLM_L_X8Y153_SLICE_X10Y153_AQ;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_D2 = CLBLM_R_X3Y150_SLICE_X3Y150_BQ;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_D3 = CLBLM_L_X10Y153_SLICE_X12Y153_BQ;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_D4 = CLBLM_L_X8Y153_SLICE_X10Y153_BQ;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_D5 = CLBLM_R_X7Y145_SLICE_X8Y145_B5Q;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_D6 = CLBLM_L_X8Y152_SLICE_X11Y152_B5Q;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_A2 = CLBLM_R_X3Y147_SLICE_X3Y147_BQ;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_A3 = CLBLM_L_X8Y152_SLICE_X10Y152_AQ;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_A4 = CLBLM_R_X11Y150_SLICE_X14Y150_AQ;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_A5 = CLBLM_L_X10Y146_SLICE_X12Y146_AQ;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_A6 = CLBLM_R_X5Y144_SLICE_X6Y144_CQ;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_B1 = CLBLM_L_X8Y146_SLICE_X10Y146_BQ;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_B2 = CLBLM_R_X3Y147_SLICE_X3Y147_BQ;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_B3 = CLBLL_L_X4Y145_SLICE_X4Y145_AQ;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_B5 = CLBLM_R_X5Y144_SLICE_X6Y144_CQ;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_B6 = CLBLM_L_X8Y152_SLICE_X10Y152_BQ;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_C2 = CLBLM_R_X5Y144_SLICE_X6Y144_DQ;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_C3 = CLBLM_R_X3Y148_SLICE_X2Y148_D5Q;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_C4 = CLBLM_L_X8Y151_SLICE_X11Y151_A5Q;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_C5 = CLBLM_L_X8Y152_SLICE_X10Y152_CQ;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_C6 = CLBLM_R_X5Y147_SLICE_X7Y147_CQ;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_D1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_D2 = CLBLL_L_X4Y149_SLICE_X4Y149_CQ;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_D3 = CLBLM_R_X7Y152_SLICE_X9Y152_CQ;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_D4 = CLBLM_L_X8Y146_SLICE_X10Y146_C5Q;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_D5 = 1'b1;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_D6 = 1'b1;
  assign LIOB33_X0Y165_IOB_X0Y166_O = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign LIOB33_X0Y165_IOB_X0Y165_O = LIOB33_X0Y57_IOB_X0Y57_I;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_A2 = CLBLM_R_X3Y150_SLICE_X2Y150_DQ;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_A3 = CLBLL_L_X4Y144_SLICE_X5Y144_DQ;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_A4 = CLBLM_R_X5Y150_SLICE_X6Y150_DQ;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_A5 = CLBLM_L_X8Y144_SLICE_X10Y144_A5Q;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_A6 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_B1 = CLBLM_R_X7Y144_SLICE_X9Y144_DQ;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_B2 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_B3 = CLBLL_L_X2Y149_SLICE_X0Y149_AQ;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_B4 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_B6 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_C1 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_C2 = CLBLL_L_X4Y146_SLICE_X4Y146_DQ;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_C3 = CLBLL_L_X2Y143_SLICE_X1Y143_DQ;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_C4 = CLBLM_L_X10Y143_SLICE_X12Y143_DO5;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_C5 = CLBLM_L_X8Y142_SLICE_X10Y142_BO5;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_C6 = CLBLM_L_X8Y147_SLICE_X10Y147_DO6;
  assign LIOI3_X0Y165_OLOGIC_X0Y166_D1 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y165_OLOGIC_X0Y166_T1 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_D1 = CLBLM_R_X5Y150_SLICE_X6Y150_DQ;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_D2 = CLBLM_R_X5Y146_SLICE_X6Y146_AQ;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_D3 = CLBLM_R_X3Y150_SLICE_X2Y150_DQ;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_D4 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_D5 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_D6 = CLBLM_L_X8Y146_SLICE_X11Y146_AQ;
  assign LIOI3_X0Y103_OLOGIC_X0Y104_D1 = CLBLM_R_X7Y144_SLICE_X9Y144_C5Q;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_SR = CLBLM_R_X11Y148_SLICE_X14Y148_CO6;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_D1 = CLBLL_L_X2Y148_SLICE_X1Y148_BO6;
  assign LIOI3_X0Y165_OLOGIC_X0Y165_D1 = LIOB33_X0Y57_IOB_X0Y57_I;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_A1 = CLBLM_R_X11Y149_SLICE_X14Y149_AQ;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_A2 = CLBLM_R_X5Y147_SLICE_X7Y147_A5Q;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_A1 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_A2 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_A3 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_A4 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_A5 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_A6 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_A3 = CLBLM_R_X5Y147_SLICE_X7Y147_BQ;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_A4 = CLBLM_L_X8Y150_SLICE_X10Y150_A5Q;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_A5 = CLBLM_L_X10Y143_SLICE_X13Y143_AO6;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_B1 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_B2 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_B3 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_B4 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_B5 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_B6 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_AX = CLBLM_R_X3Y144_SLICE_X3Y144_CQ;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_B1 = CLBLM_R_X7Y146_SLICE_X8Y146_DO6;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_B2 = CLBLM_R_X5Y147_SLICE_X7Y147_C5Q;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_C1 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_C2 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_C3 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_C4 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_C5 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_C6 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_BX = CLBLM_L_X8Y144_SLICE_X10Y144_A5Q;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_C1 = CLBLM_R_X7Y147_SLICE_X8Y147_AQ;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_C2 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_C3 = CLBLM_L_X10Y143_SLICE_X12Y143_BO5;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_C4 = CLBLM_L_X10Y143_SLICE_X12Y143_AO6;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_C5 = CLBLM_R_X7Y147_SLICE_X8Y147_CQ;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_C6 = CLBLM_L_X12Y149_SLICE_X16Y149_CO6;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_CE = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_D1 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_D2 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_D3 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_D4 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_D5 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X0Y145_D6 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_D1 = CLBLM_L_X8Y145_SLICE_X10Y145_CO5;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_D2 = CLBLM_L_X8Y142_SLICE_X10Y142_BO5;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_D3 = CLBLM_R_X7Y149_SLICE_X8Y149_DQ;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_D4 = CLBLM_R_X7Y146_SLICE_X8Y146_AO5;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_D5 = CLBLM_R_X5Y147_SLICE_X7Y147_B5Q;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_D6 = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_T1 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_A1 = CLBLL_L_X2Y147_SLICE_X1Y147_A5Q;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_A2 = CLBLM_R_X5Y147_SLICE_X6Y147_BQ;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_A3 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_A4 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_A6 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_B1 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_B2 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_B3 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_B4 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_B5 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_B6 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_C1 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_C2 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_C3 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_C4 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_C5 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_C6 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_D1 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_D2 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_D3 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_D4 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_D5 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_D6 = 1'b1;
  assign CLBLL_L_X2Y145_SLICE_X1Y145_SR = CLBLL_L_X2Y146_SLICE_X1Y146_BO6;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_D1 = CLBLL_L_X2Y146_SLICE_X1Y146_CO6;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_A1 = CLBLM_R_X3Y150_SLICE_X2Y150_CO5;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_A3 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_A4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_A5 = CLBLM_L_X12Y151_SLICE_X16Y151_BQ;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_A6 = 1'b1;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_B1 = 1'b1;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_B2 = CLBLM_L_X8Y153_SLICE_X11Y153_BQ;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_B3 = CLBLM_L_X10Y153_SLICE_X12Y153_BQ;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_B5 = CLBLM_R_X3Y152_SLICE_X2Y152_BQ;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_B6 = 1'b1;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_C1 = CLBLM_R_X11Y152_SLICE_X14Y152_DO6;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_C2 = CLBLM_L_X10Y152_SLICE_X12Y152_CQ;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_C3 = CLBLM_R_X7Y145_SLICE_X8Y145_B5Q;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_C4 = CLBLM_R_X3Y150_SLICE_X3Y150_BQ;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_C5 = CLBLM_L_X8Y153_SLICE_X10Y153_AQ;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_C6 = CLBLM_L_X8Y152_SLICE_X11Y152_BQ;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_D1 = 1'b1;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_D2 = 1'b1;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_D3 = 1'b1;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_D4 = 1'b1;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_D5 = 1'b1;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_D6 = 1'b1;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_A1 = CLBLM_L_X8Y153_SLICE_X10Y153_DO6;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_A2 = CLBLM_L_X8Y152_SLICE_X11Y152_BQ;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_A3 = CLBLM_L_X8Y153_SLICE_X10Y153_AQ;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_A4 = CLBLM_L_X8Y153_SLICE_X10Y153_DO5;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_A6 = CLBLM_R_X7Y143_SLICE_X9Y143_CQ;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_B1 = CLBLM_R_X7Y145_SLICE_X8Y145_B5Q;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_B2 = CLBLM_L_X8Y153_SLICE_X10Y153_BQ;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_B3 = CLBLM_L_X8Y153_SLICE_X10Y153_AQ;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_B5 = CLBLM_L_X8Y147_SLICE_X10Y147_BQ;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_B6 = CLBLM_R_X3Y150_SLICE_X3Y150_BQ;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_C1 = CLBLM_L_X8Y150_SLICE_X10Y150_AQ;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_C2 = CLBLM_L_X8Y153_SLICE_X10Y153_CQ;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_C3 = CLBLM_R_X7Y153_SLICE_X8Y153_BO6;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_C5 = 1'b1;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_C6 = CLBLM_R_X7Y154_SLICE_X9Y154_BO6;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_D1 = CLBLM_R_X11Y152_SLICE_X14Y152_DO6;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_D2 = CLBLM_R_X3Y150_SLICE_X3Y150_BQ;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_D3 = CLBLM_L_X8Y153_SLICE_X10Y153_AQ;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_D4 = CLBLM_L_X10Y152_SLICE_X12Y152_CQ;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_D5 = CLBLM_R_X7Y145_SLICE_X8Y145_B5Q;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_D6 = 1'b1;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_C4 = 1'b1;
  assign RIOI3_X105Y147_ILOGIC_X1Y148_D = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_C5 = 1'b1;
  assign RIOI3_X105Y147_ILOGIC_X1Y147_D = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_C6 = 1'b1;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_SR = CLBLM_R_X11Y150_SLICE_X14Y150_DO6;
  assign LIOB33_X0Y167_IOB_X0Y168_O = RIOB33_X105Y101_IOB_X1Y101_I;
  assign LIOB33_X0Y167_IOB_X0Y167_O = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_A1 = CLBLM_L_X8Y149_SLICE_X11Y149_BQ;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_A2 = CLBLM_L_X10Y147_SLICE_X12Y147_BQ;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_A3 = CLBLM_R_X7Y147_SLICE_X9Y147_AQ;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_A4 = CLBLM_R_X7Y145_SLICE_X9Y145_BQ;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_A5 = CLBLL_L_X4Y146_SLICE_X5Y146_DO6;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_D2 = 1'b1;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_B1 = 1'b1;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_B2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_B3 = CLBLM_R_X7Y144_SLICE_X8Y144_BQ;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_B4 = CLBLL_L_X4Y151_SLICE_X5Y151_AQ;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_B5 = CLBLM_L_X10Y149_SLICE_X12Y149_A5Q;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_B6 = 1'b1;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_C1 = CLBLL_L_X4Y143_SLICE_X5Y143_DQ;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_C2 = CLBLM_R_X7Y147_SLICE_X9Y147_CQ;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_C3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_C4 = CLBLM_R_X5Y147_SLICE_X7Y147_CQ;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_C5 = CLBLL_L_X4Y147_SLICE_X5Y147_CQ;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_C6 = 1'b1;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_D5 = 1'b1;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_D6 = 1'b1;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_D1 = CLBLM_R_X5Y148_SLICE_X6Y148_AQ;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_D2 = CLBLM_L_X10Y142_SLICE_X12Y142_CO6;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_D3 = CLBLL_L_X4Y147_SLICE_X5Y147_AQ;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_D4 = CLBLM_R_X11Y147_SLICE_X14Y147_AQ;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_D5 = CLBLM_R_X3Y146_SLICE_X3Y146_AQ;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_D6 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_A1 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_A2 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_A3 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_A4 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_A5 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_A6 = 1'b1;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_A1 = CLBLM_R_X5Y149_SLICE_X6Y149_D5Q;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_A2 = CLBLM_L_X8Y150_SLICE_X11Y150_B5Q;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_A3 = CLBLM_R_X7Y147_SLICE_X8Y147_AQ;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_B1 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_B2 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_B3 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_B4 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_B5 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_B6 = 1'b1;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_A4 = CLBLM_R_X5Y142_SLICE_X7Y142_C5Q;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_A6 = CLBLL_L_X2Y148_SLICE_X1Y148_A5Q;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_C1 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_C2 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_C3 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_C4 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_C5 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_C6 = 1'b1;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_B4 = CLBLM_R_X11Y145_SLICE_X15Y145_BO5;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_B5 = 1'b1;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_B6 = CLBLM_R_X3Y153_SLICE_X3Y153_A5Q;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_C1 = CLBLM_R_X5Y144_SLICE_X6Y144_CQ;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_C2 = CLBLM_R_X7Y147_SLICE_X8Y147_CQ;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_C3 = CLBLM_R_X7Y141_SLICE_X8Y141_AQ;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_C4 = CLBLL_L_X2Y148_SLICE_X1Y148_AQ;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_D1 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_D2 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_D3 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_D4 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_D5 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X0Y146_D6 = 1'b1;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_D1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_D2 = CLBLM_R_X11Y151_SLICE_X15Y151_A5Q;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_D3 = CLBLM_R_X5Y147_SLICE_X7Y147_B5Q;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_D4 = CLBLM_R_X5Y144_SLICE_X7Y144_CQ;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_D5 = CLBLM_L_X8Y148_SLICE_X11Y148_DQ;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_D6 = 1'b1;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_B4 = CLBLM_R_X5Y140_SLICE_X7Y140_AQ;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_C2 = CLBLM_R_X7Y150_SLICE_X9Y150_BQ;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_A3 = CLBLM_L_X10Y147_SLICE_X13Y147_AQ;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_C3 = CLBLM_R_X5Y152_SLICE_X7Y152_AQ;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_A2 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_A3 = CLBLM_R_X3Y154_SLICE_X3Y154_AQ;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_A4 = CLBLL_L_X2Y149_SLICE_X1Y149_AQ;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_A5 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_A6 = 1'b1;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_C4 = CLBLM_R_X5Y152_SLICE_X6Y152_AQ;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_C5 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_B2 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_B3 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_B4 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_B5 = CLBLM_R_X3Y151_SLICE_X3Y151_AQ;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_B6 = 1'b1;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_C6 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_C1 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_C2 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_C3 = CLBLM_R_X5Y149_SLICE_X7Y149_BQ;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_C4 = CLBLM_R_X3Y147_SLICE_X2Y147_CQ;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_C5 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_C6 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_D1 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_D2 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_D3 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_D4 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_D5 = 1'b1;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_D6 = 1'b1;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_C3 = CLBLM_L_X8Y144_SLICE_X10Y144_B5Q;
  assign CLBLL_L_X2Y146_SLICE_X1Y146_SR = CLBLM_R_X7Y144_SLICE_X8Y144_DO6;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_A1 = 1'b1;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_A2 = 1'b1;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_A3 = 1'b1;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_A4 = 1'b1;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_A5 = 1'b1;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_A6 = 1'b1;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_D1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_B1 = 1'b1;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_B2 = 1'b1;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_B3 = 1'b1;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_B4 = 1'b1;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_B5 = 1'b1;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_B6 = 1'b1;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_D2 = CLBLM_L_X8Y144_SLICE_X10Y144_B5Q;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_D3 = CLBLM_R_X7Y145_SLICE_X8Y145_B5Q;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_C1 = 1'b1;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_C2 = 1'b1;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_C3 = 1'b1;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_C4 = 1'b1;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_C5 = 1'b1;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_C6 = 1'b1;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_D4 = CLBLM_R_X5Y151_SLICE_X6Y151_CQ;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_D5 = CLBLM_R_X7Y149_SLICE_X9Y149_CQ;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_D6 = 1'b1;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_D1 = 1'b1;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_D2 = 1'b1;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_D3 = 1'b1;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_D4 = 1'b1;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_D5 = 1'b1;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_D6 = 1'b1;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_A1 = CLBLM_R_X7Y154_SLICE_X8Y154_CQ;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_A2 = CLBLM_R_X11Y151_SLICE_X15Y151_BQ;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_A3 = CLBLM_L_X8Y154_SLICE_X10Y154_AQ;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_A5 = CLBLM_R_X3Y152_SLICE_X2Y152_BQ;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_A6 = CLBLM_R_X7Y154_SLICE_X8Y154_DO5;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_B1 = CLBLM_R_X3Y151_SLICE_X3Y151_C5Q;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_B2 = CLBLM_R_X7Y153_SLICE_X8Y153_DO5;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_B3 = CLBLM_R_X7Y151_SLICE_X9Y151_AQ;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_B4 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_B5 = CLBLL_L_X4Y154_SLICE_X4Y154_AQ;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_B6 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_C1 = 1'b1;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_C2 = 1'b1;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_C3 = 1'b1;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_C4 = 1'b1;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_C5 = 1'b1;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_C6 = 1'b1;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_A1 = 1'b1;
  assign LIOB33_X0Y169_IOB_X0Y169_O = RIOB33_X105Y117_IOB_X1Y117_I;
  assign LIOB33_X0Y169_IOB_X0Y170_O = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_A3 = CLBLM_R_X7Y152_SLICE_X8Y152_AQ;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_D1 = 1'b1;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_D2 = 1'b1;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_D3 = 1'b1;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_D4 = 1'b1;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_D5 = 1'b1;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_D6 = 1'b1;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_A4 = CLBLM_L_X8Y152_SLICE_X10Y152_CQ;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_A5 = CLBLM_L_X10Y143_SLICE_X12Y143_BO6;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_A6 = CLBLM_L_X8Y146_SLICE_X10Y146_BQ;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_T1 = 1'b1;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_C5 = CLBLM_R_X5Y144_SLICE_X7Y144_AQ;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_B1 = 1'b1;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_C6 = CLBLM_L_X10Y143_SLICE_X12Y143_AO6;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_B2 = CLBLM_R_X7Y152_SLICE_X8Y152_BQ;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_B3 = CLBLM_R_X7Y151_SLICE_X8Y151_CQ;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_SR = CLBLM_R_X11Y150_SLICE_X14Y150_DO6;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_B4 = CLBLL_L_X2Y148_SLICE_X0Y148_B5Q;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_A1 = CLBLM_L_X8Y146_SLICE_X10Y146_CQ;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_A2 = CLBLM_L_X10Y147_SLICE_X13Y147_A5Q;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_A3 = CLBLM_R_X7Y148_SLICE_X9Y148_AQ;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_A4 = CLBLM_R_X5Y146_SLICE_X7Y146_BQ;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_A6 = 1'b1;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_B6 = 1'b1;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_B1 = CLBLM_L_X8Y147_SLICE_X11Y147_AQ;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_B2 = CLBLM_R_X3Y148_SLICE_X2Y148_C5Q;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_B3 = CLBLL_L_X4Y147_SLICE_X5Y147_AQ;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_B4 = CLBLL_L_X4Y151_SLICE_X5Y151_AQ;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_B6 = 1'b1;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_C1 = CLBLM_R_X7Y149_SLICE_X9Y149_BQ;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_C2 = CLBLM_R_X3Y149_SLICE_X3Y149_DQ;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_C3 = CLBLL_L_X2Y146_SLICE_X1Y146_A5Q;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_C5 = CLBLM_R_X5Y150_SLICE_X7Y150_AQ;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_C6 = 1'b1;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_D1 = 1'b1;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_D2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_D3 = 1'b1;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_D4 = 1'b1;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_D5 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_A2 = CLBLM_L_X10Y146_SLICE_X12Y146_AQ;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_A3 = CLBLM_R_X7Y144_SLICE_X9Y144_AQ;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_A4 = CLBLM_R_X7Y152_SLICE_X9Y152_DQ;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_A5 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_A6 = 1'b1;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_D2 = CLBLM_L_X8Y153_SLICE_X11Y153_BQ;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_D6 = CLBLL_L_X4Y151_SLICE_X5Y151_AQ;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_A1 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_B2 = CLBLL_L_X4Y144_SLICE_X5Y144_D5Q;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_B3 = CLBLM_L_X10Y147_SLICE_X12Y147_C5Q;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_B4 = CLBLL_L_X4Y153_SLICE_X5Y153_BQ;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_B5 = CLBLM_R_X3Y144_SLICE_X3Y144_A5Q;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_B6 = 1'b1;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_A2 = 1'b1;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_A3 = 1'b1;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_D5 = CLBLL_L_X4Y146_SLICE_X4Y146_BQ;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_C1 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_C2 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_C3 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_C4 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_C5 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_C6 = 1'b1;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_D6 = CLBLM_R_X3Y152_SLICE_X2Y152_BQ;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_B1 = CLBLM_R_X11Y149_SLICE_X14Y149_AQ;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_B2 = CLBLM_R_X3Y147_SLICE_X2Y147_C5Q;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_B3 = CLBLM_L_X10Y144_SLICE_X13Y144_CO6;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_B4 = CLBLM_L_X8Y150_SLICE_X10Y150_A5Q;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_B5 = CLBLM_R_X7Y148_SLICE_X9Y148_AQ;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_D1 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_D2 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_D3 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_D4 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_D5 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X0Y147_D6 = 1'b1;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_C4 = CLBLM_L_X8Y146_SLICE_X11Y146_A5Q;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_C6 = CLBLM_R_X5Y149_SLICE_X7Y149_C5Q;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_D1 = CLBLM_R_X3Y148_SLICE_X3Y148_CO5;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_D2 = 1'b1;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_D3 = CLBLL_L_X4Y148_SLICE_X4Y148_BO5;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_D4 = CLBLM_L_X10Y151_SLICE_X12Y151_BO6;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_D5 = CLBLM_R_X7Y152_SLICE_X8Y152_DO6;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_D6 = CLBLM_L_X10Y143_SLICE_X12Y143_AO5;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_SR = CLBLM_R_X11Y148_SLICE_X15Y148_BO6;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_A2 = CLBLM_R_X5Y147_SLICE_X6Y147_DQ;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_A3 = CLBLM_R_X3Y146_SLICE_X3Y146_C5Q;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_A4 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_A5 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_A6 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_B2 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_B3 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_B4 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_B5 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_B6 = CLBLM_R_X3Y144_SLICE_X3Y144_CQ;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_C1 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_C2 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_C3 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_C4 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_C5 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_C6 = 1'b1;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_D3 = CLBLM_L_X8Y153_SLICE_X10Y153_CQ;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_D4 = CLBLM_R_X7Y149_SLICE_X9Y149_AO5;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y167_OLOGIC_X0Y168_D1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_D5 = CLBLM_R_X7Y153_SLICE_X9Y153_BQ;
  assign LIOB33_X0Y179_IOB_X0Y180_O = RIOB33_X105Y127_IOB_X1Y127_I;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_D1 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_D2 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_D3 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_D4 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_D5 = 1'b1;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_D6 = 1'b1;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_D6 = CLBLM_R_X7Y153_SLICE_X9Y153_AQ;
  assign LIOB33_X0Y179_IOB_X0Y179_O = RIOB33_X105Y125_IOB_X1Y126_I;
  assign CLBLL_L_X2Y147_SLICE_X1Y147_SR = CLBLL_L_X2Y147_SLICE_X1Y147_BO6;
  assign LIOI3_X0Y105_OLOGIC_X0Y106_D1 = CLBLL_L_X4Y147_SLICE_X5Y147_DQ;
  assign LIOI3_X0Y167_OLOGIC_X0Y168_T1 = 1'b1;
  assign LIOI3_X0Y167_OLOGIC_X0Y167_D1 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign LIOI3_X0Y105_OLOGIC_X0Y106_T1 = 1'b1;
  assign RIOI3_X105Y151_OLOGIC_X1Y152_D1 = 1'b1;
  assign LIOI3_X0Y167_OLOGIC_X0Y167_T1 = 1'b1;
  assign LIOI3_X0Y105_OLOGIC_X0Y105_D1 = CLBLM_R_X5Y144_SLICE_X6Y144_B5Q;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_B5 = 1'b1;
  assign RIOI3_X105Y151_OLOGIC_X1Y152_T1 = 1'b1;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_B6 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_D1 = CLBLL_L_X4Y153_SLICE_X4Y153_A5Q;
  assign LIOI3_X0Y105_OLOGIC_X0Y105_T1 = 1'b1;
  assign RIOI3_X105Y151_OLOGIC_X1Y151_D1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_T1 = 1'b1;
  assign RIOI3_X105Y151_OLOGIC_X1Y151_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_D1 = CLBLM_R_X3Y146_SLICE_X2Y146_CQ;
  assign LIOB33_X0Y171_IOB_X0Y172_O = RIOB33_X105Y119_IOB_X1Y120_I;
  assign LIOB33_X0Y171_IOB_X0Y171_O = RIOB33_X105Y119_IOB_X1Y119_I;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_T1 = 1'b1;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_C4 = 1'b1;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_C5 = 1'b1;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_C6 = 1'b1;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_A1 = CLBLM_R_X7Y151_SLICE_X9Y151_CQ;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_A2 = CLBLM_R_X7Y152_SLICE_X8Y152_BQ;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_A3 = CLBLM_R_X7Y145_SLICE_X8Y145_AQ;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_A4 = CLBLL_L_X2Y151_SLICE_X1Y151_BQ;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_A6 = 1'b1;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_AX = CLBLM_R_X5Y148_SLICE_X6Y148_AQ;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_B1 = CLBLM_R_X7Y148_SLICE_X8Y148_BO5;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_B2 = CLBLM_L_X10Y143_SLICE_X12Y143_DO6;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_B3 = CLBLL_L_X4Y146_SLICE_X4Y146_AQ;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_B4 = CLBLL_L_X2Y149_SLICE_X1Y149_A5Q;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_B5 = CLBLM_R_X5Y152_SLICE_X7Y152_CQ;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_B6 = 1'b1;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_BX = CLBLM_R_X3Y152_SLICE_X2Y152_BQ;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_C1 = CLBLM_R_X7Y149_SLICE_X8Y149_AQ;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_C2 = CLBLM_R_X3Y147_SLICE_X3Y147_AQ;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_C3 = CLBLM_L_X8Y149_SLICE_X10Y149_A5Q;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_C4 = CLBLM_R_X7Y150_SLICE_X8Y150_DQ;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_C5 = CLBLM_R_X7Y143_SLICE_X9Y143_AQ;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_C6 = 1'b1;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_CE = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_CX = CLBLM_L_X8Y149_SLICE_X10Y149_A5Q;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_A1 = CLBLM_L_X8Y153_SLICE_X10Y153_AQ;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_A2 = CLBLM_R_X3Y148_SLICE_X3Y148_DO6;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_A3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_A4 = CLBLM_R_X3Y149_SLICE_X3Y149_DQ;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_A5 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_A6 = 1'b1;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_D1 = CLBLM_R_X7Y152_SLICE_X8Y152_AQ;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_D2 = CLBLM_L_X10Y142_SLICE_X12Y142_CO6;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_D3 = CLBLM_R_X7Y148_SLICE_X8Y148_BO5;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_B1 = CLBLM_R_X3Y150_SLICE_X2Y150_B5Q;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_B2 = CLBLM_L_X10Y150_SLICE_X12Y150_AQ;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_B3 = CLBLL_L_X2Y147_SLICE_X0Y147_AQ;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_B5 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_B6 = 1'b1;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_A1 = CLBLM_R_X7Y150_SLICE_X8Y150_DQ;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_A2 = CLBLM_R_X7Y150_SLICE_X8Y150_CQ;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_A3 = CLBLM_R_X7Y149_SLICE_X8Y149_AQ;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_C1 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_C2 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_C3 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_C4 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_C5 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_C6 = 1'b1;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_A5 = CLBLM_R_X3Y146_SLICE_X3Y146_CQ;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_B1 = CLBLM_L_X10Y143_SLICE_X12Y143_AO6;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_B2 = 1'b1;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_B4 = CLBLL_L_X4Y151_SLICE_X5Y151_AQ;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_D1 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_D2 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_D3 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_D4 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_D5 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X0Y148_D6 = 1'b1;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_C1 = CLBLM_R_X5Y142_SLICE_X7Y142_BQ;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_C2 = CLBLM_R_X3Y151_SLICE_X3Y151_BQ;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_C3 = 1'b1;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_C4 = CLBLM_L_X12Y149_SLICE_X16Y149_BQ;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_C5 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_A1 = CLBLM_R_X5Y149_SLICE_X6Y149_D5Q;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_C6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_D1 = CLBLM_R_X7Y143_SLICE_X8Y143_AQ;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_D2 = CLBLM_R_X7Y149_SLICE_X8Y149_CQ;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_D3 = CLBLM_R_X7Y149_SLICE_X8Y149_DQ;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_D4 = CLBLM_L_X10Y143_SLICE_X12Y143_BO5;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_D6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_D5 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_A1 = CLBLL_L_X4Y149_SLICE_X4Y149_C5Q;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_A3 = CLBLL_L_X4Y148_SLICE_X5Y148_BQ;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_A4 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_A5 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_A6 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_B1 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_B2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_B3 = CLBLM_R_X3Y146_SLICE_X2Y146_C5Q;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_B4 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_B5 = CLBLM_R_X3Y148_SLICE_X2Y148_BQ;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_B6 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_C1 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_C2 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_C3 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_C4 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_C5 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_C6 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_B2 = CLBLM_L_X8Y149_SLICE_X11Y149_BQ;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_D1 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_D2 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_D3 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_D4 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_D5 = 1'b1;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_D6 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_B3 = CLBLM_R_X7Y142_SLICE_X8Y142_DO6;
  assign CLBLL_L_X2Y148_SLICE_X1Y148_SR = CLBLL_L_X2Y146_SLICE_X1Y146_BO6;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_B6 = CLBLM_L_X8Y148_SLICE_X11Y148_B5Q;
  assign LIOB33_X0Y173_IOB_X0Y174_O = RIOB33_X105Y121_IOB_X1Y122_I;
  assign LIOB33_X0Y173_IOB_X0Y173_O = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_C3 = CLBLL_L_X2Y148_SLICE_X0Y148_B5Q;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_C4 = CLBLL_L_X4Y144_SLICE_X4Y144_DO6;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_C2 = CLBLM_R_X7Y152_SLICE_X8Y152_CQ;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_C3 = CLBLM_R_X7Y154_SLICE_X8Y154_DO6;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_A1 = CLBLM_L_X8Y150_SLICE_X11Y150_B5Q;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_A2 = CLBLM_L_X8Y143_SLICE_X11Y143_CQ;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_A3 = CLBLM_R_X7Y150_SLICE_X9Y150_AQ;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_A4 = CLBLM_R_X5Y149_SLICE_X6Y149_D5Q;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_A6 = CLBLM_R_X5Y151_SLICE_X7Y151_AQ;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_C4 = CLBLM_R_X5Y152_SLICE_X6Y152_AQ;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_B1 = CLBLL_L_X4Y150_SLICE_X4Y150_AQ;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_B2 = CLBLM_R_X7Y150_SLICE_X9Y150_DQ;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_B3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_B4 = CLBLL_L_X4Y151_SLICE_X5Y151_BQ;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_B6 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_A1 = CLBLM_R_X5Y143_SLICE_X7Y143_DQ;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_A2 = CLBLM_R_X5Y140_SLICE_X7Y140_BQ;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_A3 = CLBLM_R_X5Y140_SLICE_X7Y140_AQ;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_A4 = CLBLM_R_X11Y145_SLICE_X15Y145_BO5;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_A6 = 1'b1;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_C2 = CLBLM_L_X8Y146_SLICE_X10Y146_AQ;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_C3 = CLBLM_R_X7Y144_SLICE_X9Y144_B5Q;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_A1 = CLBLM_R_X3Y150_SLICE_X2Y150_B5Q;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_A2 = 1'b1;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_A3 = CLBLM_L_X10Y150_SLICE_X12Y150_CQ;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_A4 = CLBLM_R_X3Y151_SLICE_X2Y151_A5Q;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_A5 = CLBLM_R_X7Y148_SLICE_X9Y148_AQ;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_B3 = CLBLM_R_X5Y140_SLICE_X7Y140_AQ;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_B4 = RIOB33_X105Y123_IOB_X1Y123_I;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_B5 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_B1 = 1'b1;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_B2 = 1'b1;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_B3 = 1'b1;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_B4 = 1'b1;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_B5 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_C6 = 1'b1;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_B6 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_C1 = 1'b1;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_C1 = 1'b1;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_C2 = 1'b1;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_C3 = 1'b1;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_C4 = 1'b1;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_C5 = 1'b1;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_C6 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_D1 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_D2 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_D3 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_D4 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_D5 = 1'b1;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_D1 = 1'b1;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_D2 = 1'b1;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_D3 = 1'b1;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_D4 = 1'b1;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_D5 = 1'b1;
  assign CLBLL_L_X2Y149_SLICE_X0Y149_D6 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_A1 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_A2 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_A3 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_A4 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_A5 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_A6 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_B1 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_B2 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_B3 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_B4 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_B5 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_B6 = 1'b1;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_D1 = 1'b1;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_D2 = CLBLM_R_X7Y154_SLICE_X8Y154_BQ;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_C1 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_C2 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_C3 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_C4 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_C5 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_C6 = 1'b1;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_D3 = CLBLM_R_X3Y148_SLICE_X2Y148_C5Q;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_D4 = CLBLM_R_X7Y150_SLICE_X8Y150_BQ;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_D5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_D6 = 1'b1;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_A1 = CLBLM_R_X5Y149_SLICE_X7Y149_BQ;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_A2 = CLBLL_L_X2Y144_SLICE_X1Y144_BQ;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_A3 = CLBLM_R_X7Y148_SLICE_X9Y148_AQ;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_A5 = CLBLM_L_X10Y150_SLICE_X12Y150_CQ;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_A6 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_D1 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_D2 = 1'b1;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_B1 = CLBLL_L_X4Y152_SLICE_X5Y152_CQ;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_B2 = CLBLL_L_X2Y149_SLICE_X1Y149_BQ;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_B3 = CLBLL_L_X2Y149_SLICE_X1Y149_CQ;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_B4 = CLBLL_L_X2Y149_SLICE_X1Y149_DQ;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_B5 = CLBLM_R_X3Y150_SLICE_X2Y150_DQ;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_B6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_D3 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_D4 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_D5 = 1'b1;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_C1 = CLBLL_L_X2Y149_SLICE_X1Y149_BQ;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_C2 = CLBLL_L_X4Y152_SLICE_X5Y152_CQ;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_C3 = CLBLL_L_X2Y149_SLICE_X1Y149_DQ;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_C5 = CLBLM_R_X5Y142_SLICE_X7Y142_C5Q;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_C6 = CLBLL_L_X2Y149_SLICE_X1Y149_CQ;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_C1 = CLBLM_R_X7Y152_SLICE_X9Y152_AQ;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_C2 = CLBLM_R_X5Y144_SLICE_X6Y144_D5Q;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_C3 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_D1 = CLBLL_L_X2Y149_SLICE_X1Y149_BQ;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_D2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_D3 = CLBLL_L_X2Y149_SLICE_X1Y149_DQ;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_D4 = CLBLL_L_X2Y147_SLICE_X0Y147_B5Q;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_D5 = CLBLL_L_X4Y152_SLICE_X5Y152_CQ;
  assign CLBLL_L_X2Y149_SLICE_X1Y149_D6 = CLBLL_L_X2Y149_SLICE_X1Y149_CQ;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_C4 = CLBLM_L_X8Y148_SLICE_X11Y148_CQ;
  assign LIOB33_X0Y175_IOB_X0Y176_O = RIOB33_X105Y115_IOB_X1Y116_I;
  assign LIOB33_X0Y175_IOB_X0Y175_O = RIOB33_X105Y123_IOB_X1Y123_I;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_C2 = CLBLM_L_X8Y148_SLICE_X10Y148_BO5;
  assign LIOI3_X0Y171_OLOGIC_X0Y172_D1 = RIOB33_X105Y119_IOB_X1Y120_I;
  assign RIOI3_SING_X105Y100_ILOGIC_X1Y100_D = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign LIOI3_X0Y171_OLOGIC_X0Y172_T1 = 1'b1;
  assign LIOI3_X0Y109_OLOGIC_X0Y110_D1 = CLBLM_R_X5Y143_SLICE_X6Y143_DQ;
  assign LIOI3_X0Y171_OLOGIC_X0Y171_D1 = RIOB33_X105Y119_IOB_X1Y119_I;
  assign LIOI3_X0Y109_OLOGIC_X0Y110_T1 = 1'b1;
  assign RIOI3_X105Y153_OLOGIC_X1Y154_D1 = 1'b1;
  assign LIOI3_X0Y171_OLOGIC_X0Y171_T1 = 1'b1;
  assign LIOI3_X0Y109_OLOGIC_X0Y109_D1 = CLBLL_L_X2Y153_SLICE_X1Y153_AQ;
  assign RIOI3_X105Y153_OLOGIC_X1Y154_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_D1 = CLBLM_R_X3Y144_SLICE_X3Y144_A5Q;
  assign RIOB33_X105Y185_IOB_X1Y186_O = CLBLM_R_X7Y154_SLICE_X9Y154_CO6;
  assign LIOI3_X0Y109_OLOGIC_X0Y109_T1 = 1'b1;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_C5 = CLBLM_L_X10Y146_SLICE_X12Y146_CO5;
  assign RIOB33_X105Y185_IOB_X1Y185_O = CLBLM_L_X8Y154_SLICE_X10Y154_BO6;
  assign RIOI3_X105Y153_OLOGIC_X1Y153_D1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_T1 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_A1 = CLBLM_R_X3Y148_SLICE_X2Y148_DQ;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_A2 = CLBLM_R_X7Y146_SLICE_X8Y146_BQ;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_A3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_A4 = CLBLM_R_X7Y153_SLICE_X8Y153_DO6;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_A5 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_A6 = CLBLM_L_X10Y150_SLICE_X12Y150_CQ;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_D1 = CLBLM_R_X7Y150_SLICE_X9Y150_B5Q;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_B1 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_B2 = CLBLM_R_X5Y149_SLICE_X7Y149_D5Q;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_B4 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_B5 = CLBLM_L_X8Y146_SLICE_X10Y146_AQ;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_B6 = CLBLM_R_X5Y153_SLICE_X7Y153_CO6;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_T1 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_A1 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_A2 = CLBLL_L_X4Y153_SLICE_X4Y153_AQ;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_A3 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_A4 = CLBLM_R_X7Y141_SLICE_X9Y141_AQ;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_A1 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_A2 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_A3 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_A4 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_A5 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_A6 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_A6 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_B1 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_B1 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_B2 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_B3 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_B4 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_B5 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_B6 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_B3 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_B4 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_B6 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_C1 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_C2 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_C3 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_C4 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_C5 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_C6 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_C3 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_C4 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_C5 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_C6 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_D1 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_D2 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_D1 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_D2 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_D3 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_D4 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_D5 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X0Y150_D6 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_D3 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_D4 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_A1 = CLBLM_R_X5Y143_SLICE_X7Y143_CQ;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_A2 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_A3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_A4 = CLBLM_R_X5Y141_SLICE_X6Y141_BO6;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_A5 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_A6 = CLBLM_R_X5Y153_SLICE_X7Y153_CO6;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_C1 = CLBLM_R_X5Y152_SLICE_X7Y152_BQ;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_C2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_B1 = CLBLL_L_X4Y147_SLICE_X4Y147_D5Q;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_B2 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_B3 = CLBLL_L_X4Y150_SLICE_X4Y150_AQ;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_B4 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_B6 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_D1 = CLBLM_R_X7Y151_SLICE_X8Y151_C5Q;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_D2 = CLBLM_R_X7Y151_SLICE_X8Y151_AQ;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_C1 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_C2 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_C3 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_C4 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_C5 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_A1 = CLBLM_R_X3Y152_SLICE_X2Y152_AQ;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_A2 = CLBLM_L_X8Y146_SLICE_X10Y146_AQ;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_A3 = CLBLL_L_X2Y150_SLICE_X1Y150_AQ;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_A4 = CLBLM_R_X7Y150_SLICE_X9Y150_CQ;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_A5 = CLBLM_R_X3Y148_SLICE_X2Y148_DQ;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_C6 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_AX = CLBLL_L_X2Y150_SLICE_X1Y150_DO6;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_B2 = CLBLM_R_X3Y153_SLICE_X3Y153_CQ;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_B3 = CLBLL_L_X4Y144_SLICE_X5Y144_C5Q;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_D3 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_D4 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_D5 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_D6 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_B4 = CLBLM_R_X3Y151_SLICE_X3Y151_CQ;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_B5 = LIOB33_X0Y61_IOB_X0Y61_I;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_B6 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_D1 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_C1 = CLBLL_L_X2Y147_SLICE_X0Y147_BQ;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_C2 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_C3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_C4 = CLBLM_R_X3Y151_SLICE_X3Y151_CQ;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_C5 = CLBLM_R_X7Y153_SLICE_X9Y153_AQ;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_C6 = 1'b1;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign LIOB33_X0Y177_IOB_X0Y177_O = RIOB33_X105Y123_IOB_X1Y124_I;
  assign LIOB33_X0Y177_IOB_X0Y178_O = RIOB33_X105Y125_IOB_X1Y125_I;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_D1 = CLBLM_R_X3Y145_SLICE_X2Y145_DQ;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_D2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_D3 = CLBLL_L_X4Y151_SLICE_X5Y151_DQ;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_D4 = CLBLM_R_X3Y143_SLICE_X2Y143_AQ;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_D5 = CLBLM_R_X3Y147_SLICE_X2Y147_C5Q;
  assign CLBLL_L_X2Y150_SLICE_X1Y150_D6 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_B3 = CLBLM_R_X11Y143_SLICE_X14Y143_CO5;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_B4 = CLBLM_R_X11Y145_SLICE_X14Y145_BO6;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_B6 = CLBLM_R_X11Y148_SLICE_X14Y148_CQ;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_B5 = CLBLM_R_X11Y144_SLICE_X14Y144_AO6;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_C1 = CLBLM_L_X12Y151_SLICE_X16Y151_AQ;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_C2 = CLBLM_L_X10Y151_SLICE_X13Y151_CO6;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_C3 = CLBLM_R_X11Y151_SLICE_X15Y151_BQ;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_B6 = CLBLM_L_X10Y142_SLICE_X13Y142_BO6;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_C5 = CLBLM_L_X8Y146_SLICE_X10Y146_A5Q;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_C6 = 1'b1;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign RIOI3_SING_X105Y149_ILOGIC_X1Y149_D = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_A1 = CLBLM_R_X3Y148_SLICE_X2Y148_B5Q;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_A3 = CLBLM_R_X7Y152_SLICE_X9Y152_AQ;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_A4 = CLBLM_R_X3Y152_SLICE_X3Y152_AQ;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_A5 = CLBLM_L_X10Y151_SLICE_X12Y151_AO6;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_A6 = 1'b1;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_B1 = CLBLM_L_X8Y142_SLICE_X10Y142_AQ;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_B2 = CLBLM_R_X7Y152_SLICE_X9Y152_BQ;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_B3 = CLBLM_R_X5Y152_SLICE_X6Y152_C5Q;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_B4 = CLBLM_R_X7Y154_SLICE_X8Y154_BQ;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_B5 = CLBLM_R_X7Y155_SLICE_X8Y155_AQ;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_B6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_D1 = 1'b1;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_D2 = 1'b1;
  assign CLBLL_L_X2Y151_SLICE_X0Y151_A1 = 1'b1;
  assign CLBLL_L_X2Y151_SLICE_X0Y151_A2 = 1'b1;
  assign CLBLL_L_X2Y151_SLICE_X0Y151_A3 = 1'b1;
  assign CLBLL_L_X2Y151_SLICE_X0Y151_A4 = 1'b1;
  assign CLBLL_L_X2Y151_SLICE_X0Y151_A5 = 1'b1;
  assign CLBLL_L_X2Y151_SLICE_X0Y151_A6 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_A1 = CLBLM_R_X5Y143_SLICE_X7Y143_BQ;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_A2 = CLBLM_R_X5Y149_SLICE_X7Y149_CQ;
  assign CLBLL_L_X2Y151_SLICE_X0Y151_B1 = 1'b1;
  assign CLBLL_L_X2Y151_SLICE_X0Y151_B2 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_B3 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_B4 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_B5 = CLBLM_R_X5Y142_SLICE_X6Y142_AQ;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_B6 = 1'b1;
  assign CLBLL_L_X2Y151_SLICE_X0Y151_B3 = 1'b1;
  assign CLBLL_L_X2Y151_SLICE_X0Y151_B4 = 1'b1;
  assign CLBLL_L_X2Y151_SLICE_X0Y151_B5 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_C1 = CLBLM_R_X5Y141_SLICE_X7Y141_AQ;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_C2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X2Y151_SLICE_X0Y151_B6 = 1'b1;
  assign CLBLL_L_X2Y151_SLICE_X0Y151_C1 = 1'b1;
  assign CLBLL_L_X2Y151_SLICE_X0Y151_C2 = 1'b1;
  assign CLBLL_L_X2Y151_SLICE_X0Y151_C3 = 1'b1;
  assign CLBLL_L_X2Y151_SLICE_X0Y151_C4 = 1'b1;
  assign CLBLL_L_X2Y151_SLICE_X0Y151_C5 = 1'b1;
  assign CLBLL_L_X2Y151_SLICE_X0Y151_C6 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_C3 = CLBLM_R_X3Y144_SLICE_X3Y144_AQ;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_C4 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_C5 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_C6 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y151_SLICE_X0Y151_D1 = 1'b1;
  assign CLBLL_L_X2Y151_SLICE_X0Y151_D2 = 1'b1;
  assign CLBLL_L_X2Y151_SLICE_X0Y151_D3 = 1'b1;
  assign CLBLL_L_X2Y151_SLICE_X0Y151_D4 = 1'b1;
  assign CLBLL_L_X2Y151_SLICE_X0Y151_D5 = 1'b1;
  assign CLBLL_L_X2Y151_SLICE_X0Y151_D6 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_SR = CLBLL_L_X4Y151_SLICE_X4Y151_CO6;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_D2 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_D4 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_D5 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_D6 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_A1 = CLBLM_L_X8Y142_SLICE_X10Y142_DO6;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_A2 = CLBLM_R_X7Y143_SLICE_X9Y143_BQ;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_A3 = CLBLM_R_X5Y142_SLICE_X6Y142_AQ;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_A4 = CLBLM_L_X8Y149_SLICE_X11Y149_BQ;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_A6 = CLBLL_L_X4Y144_SLICE_X5Y144_CQ;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_B1 = CLBLM_R_X5Y144_SLICE_X6Y144_B5Q;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_B2 = CLBLM_R_X5Y142_SLICE_X6Y142_BQ;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_B3 = CLBLM_R_X11Y145_SLICE_X15Y145_BO5;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_B4 = CLBLM_R_X5Y143_SLICE_X6Y143_AQ;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_B5 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_B6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_D1 = CLBLM_R_X7Y149_SLICE_X8Y149_BQ;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_D2 = CLBLM_L_X8Y152_SLICE_X11Y152_AQ;
  assign CLBLL_L_X2Y151_SLICE_X1Y151_A1 = CLBLM_R_X3Y151_SLICE_X2Y151_CO6;
  assign CLBLL_L_X2Y151_SLICE_X1Y151_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_C3 = CLBLL_L_X4Y142_SLICE_X5Y142_BQ;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_C4 = CLBLL_L_X4Y141_SLICE_X5Y141_A5Q;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_C5 = CLBLL_L_X4Y143_SLICE_X4Y143_BQ;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_C6 = 1'b1;
  assign CLBLL_L_X2Y151_SLICE_X1Y151_A3 = LIOB33_X0Y55_IOB_X0Y55_I;
  assign CLBLL_L_X2Y151_SLICE_X1Y151_A4 = CLBLM_R_X3Y151_SLICE_X2Y151_AQ;
  assign CLBLL_L_X2Y151_SLICE_X1Y151_A5 = CLBLM_R_X5Y149_SLICE_X7Y149_CQ;
  assign CLBLL_L_X2Y151_SLICE_X1Y151_A6 = CLBLL_L_X2Y151_SLICE_X1Y151_AQ;
  assign CLBLL_L_X2Y151_SLICE_X1Y151_B1 = CLBLM_R_X3Y144_SLICE_X3Y144_CQ;
  assign CLBLL_L_X2Y151_SLICE_X1Y151_B2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X2Y151_SLICE_X1Y151_B3 = CLBLM_R_X5Y144_SLICE_X7Y144_CQ;
  assign CLBLL_L_X2Y151_SLICE_X1Y151_B4 = CLBLM_R_X7Y144_SLICE_X9Y144_AQ;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_D1 = CLBLM_L_X8Y142_SLICE_X11Y142_CQ;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_D2 = CLBLM_R_X5Y149_SLICE_X7Y149_DQ;
  assign CLBLL_L_X2Y151_SLICE_X1Y151_B5 = CLBLM_R_X3Y152_SLICE_X3Y152_AQ;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_D4 = CLBLM_R_X5Y142_SLICE_X6Y142_DQ;
  assign CLBLL_L_X2Y151_SLICE_X1Y151_B6 = CLBLL_L_X2Y149_SLICE_X1Y149_CQ;
  assign CLBLL_L_X2Y151_SLICE_X1Y151_C1 = CLBLM_R_X3Y151_SLICE_X2Y151_AQ;
  assign CLBLL_L_X2Y151_SLICE_X1Y151_C2 = CLBLM_R_X3Y151_SLICE_X2Y151_A5Q;
  assign CLBLL_L_X2Y151_SLICE_X1Y151_C3 = CLBLM_R_X3Y147_SLICE_X3Y147_B5Q;
  assign CLBLL_L_X2Y151_SLICE_X1Y151_C4 = CLBLM_R_X3Y151_SLICE_X3Y151_DQ;
  assign CLBLL_L_X2Y151_SLICE_X1Y151_C5 = CLBLL_L_X2Y151_SLICE_X1Y151_AQ;
  assign CLBLL_L_X2Y151_SLICE_X1Y151_C6 = LIOB33_X0Y55_IOB_X0Y55_I;
  assign CLBLL_L_X2Y151_SLICE_X1Y151_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_D5 = CLBLL_L_X4Y145_SLICE_X4Y145_A5Q;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_D6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_B4 = CLBLM_L_X10Y144_SLICE_X13Y144_AO6;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_B5 = CLBLM_R_X3Y142_SLICE_X2Y142_BQ;
  assign CLBLL_L_X2Y151_SLICE_X1Y151_D1 = 1'b1;
  assign CLBLL_L_X2Y151_SLICE_X1Y151_D2 = 1'b1;
  assign CLBLL_L_X2Y151_SLICE_X1Y151_D3 = 1'b1;
  assign CLBLL_L_X2Y151_SLICE_X1Y151_D4 = 1'b1;
  assign CLBLL_L_X2Y151_SLICE_X1Y151_D5 = 1'b1;
  assign CLBLL_L_X2Y151_SLICE_X1Y151_D6 = 1'b1;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_C3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_C4 = CLBLM_R_X7Y155_SLICE_X9Y155_AO5;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_C5 = CLBLM_R_X7Y153_SLICE_X9Y153_CQ;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I0 = LIOB33_X0Y77_IOB_X0Y78_I;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I1 = 1'b1;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_C6 = CLBLM_R_X7Y152_SLICE_X9Y152_BQ;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_B2 = CLBLM_R_X11Y151_SLICE_X14Y151_BQ;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_B3 = 1'b1;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_B4 = CLBLM_L_X10Y151_SLICE_X13Y151_BO5;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_B6 = CLBLM_L_X10Y147_SLICE_X13Y147_B5Q;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_D1 = CLBLM_R_X7Y153_SLICE_X9Y153_BQ;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_C1 = CLBLM_L_X10Y149_SLICE_X12Y149_AQ;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_D2 = CLBLM_L_X8Y153_SLICE_X10Y153_CQ;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_D3 = CLBLM_R_X7Y153_SLICE_X8Y153_DO6;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_D4 = CLBLM_L_X10Y151_SLICE_X12Y151_CO6;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_D5 = CLBLM_R_X7Y153_SLICE_X9Y153_AQ;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_D6 = 1'b1;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_C6 = CLBLM_L_X10Y149_SLICE_X12Y149_BQ;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign RIOI3_X105Y197_OLOGIC_X1Y198_D1 = CLBLM_R_X11Y149_SLICE_X14Y149_CO6;
  assign RIOI3_SING_X105Y150_OLOGIC_X1Y150_D1 = 1'b1;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_A1 = 1'b1;
  assign RIOI3_SING_X105Y150_OLOGIC_X1Y150_T1 = 1'b1;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_A2 = CLBLM_L_X8Y153_SLICE_X10Y153_BQ;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_A3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_A4 = 1'b1;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_D1 = 1'b1;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_A5 = 1'b1;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_D2 = 1'b1;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_A6 = 1'b1;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_D3 = CLBLM_L_X10Y153_SLICE_X12Y153_DO6;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_D4 = CLBLM_R_X11Y151_SLICE_X14Y151_AQ;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_D5 = CLBLM_R_X11Y152_SLICE_X14Y152_A5Q;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_D6 = CLBLM_L_X10Y152_SLICE_X12Y152_AQ;
  assign RIOI3_X105Y197_OLOGIC_X1Y198_T1 = 1'b1;
  assign LIOB33_X0Y181_IOB_X0Y182_O = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_B2 = CLBLM_R_X11Y149_SLICE_X15Y149_BQ;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_A1 = CLBLM_R_X7Y153_SLICE_X9Y153_DO6;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_A2 = CLBLM_R_X7Y153_SLICE_X8Y153_BO6;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_A3 = CLBLM_R_X7Y153_SLICE_X9Y153_AQ;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_A4 = CLBLM_R_X7Y154_SLICE_X9Y154_BO6;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_A6 = CLBLM_R_X3Y151_SLICE_X3Y151_DQ;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_AX = CLBLM_L_X8Y153_SLICE_X11Y153_AO6;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_B4 = CLBLM_L_X10Y150_SLICE_X12Y150_CQ;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_B1 = CLBLM_R_X7Y152_SLICE_X9Y152_DQ;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_B2 = CLBLM_R_X7Y154_SLICE_X9Y154_BO6;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_B4 = CLBLM_L_X8Y153_SLICE_X10Y153_CQ;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_B5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_A1 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_A2 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_A3 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_A4 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_A5 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_A6 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_A1 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_A3 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_B1 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_B2 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_B3 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_B4 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_B1 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_B5 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_B6 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_A6 = CLBLM_R_X5Y145_SLICE_X7Y145_A5Q;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_C1 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_C2 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_C3 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_C4 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_C5 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_C6 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_B3 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_B4 = CLBLM_L_X8Y144_SLICE_X11Y144_AQ;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_B6 = CLBLL_L_X2Y145_SLICE_X1Y145_AQ;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_C2 = CLBLM_L_X8Y144_SLICE_X10Y144_AQ;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_C3 = CLBLM_R_X3Y143_SLICE_X2Y143_DQ;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_D1 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_D2 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_D3 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_D4 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_D5 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X0Y152_D6 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_D1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_D2 = CLBLM_R_X5Y149_SLICE_X7Y149_DQ;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_D3 = CLBLM_R_X5Y143_SLICE_X7Y143_DQ;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_D4 = CLBLM_R_X5Y141_SLICE_X7Y141_AQ;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_D5 = CLBLM_L_X8Y142_SLICE_X11Y142_CQ;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_D6 = CLBLL_L_X4Y153_SLICE_X5Y153_BQ;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_B1 = CLBLM_R_X7Y152_SLICE_X9Y152_DQ;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_A1 = CLBLM_R_X5Y153_SLICE_X7Y153_A5Q;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_A2 = CLBLM_L_X8Y142_SLICE_X11Y142_CQ;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_A3 = CLBLM_R_X5Y143_SLICE_X6Y143_AQ;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_A4 = CLBLM_R_X5Y151_SLICE_X6Y151_DQ;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_A6 = CLBLM_R_X5Y149_SLICE_X7Y149_DQ;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_C1 = CLBLM_R_X7Y149_SLICE_X9Y149_DQ;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_C2 = CLBLM_R_X3Y151_SLICE_X3Y151_C5Q;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_C3 = CLBLL_L_X4Y154_SLICE_X4Y154_AQ;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_B1 = CLBLL_L_X4Y148_SLICE_X5Y148_B5Q;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_B2 = CLBLM_R_X5Y143_SLICE_X6Y143_BQ;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_B3 = CLBLL_L_X4Y142_SLICE_X4Y142_AQ;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_B5 = CLBLM_L_X8Y150_SLICE_X11Y150_B5Q;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_B6 = CLBLM_R_X5Y149_SLICE_X6Y149_D5Q;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_A1 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_A2 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_A3 = CLBLL_L_X4Y145_SLICE_X5Y145_BQ;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_A4 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_A5 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_C2 = CLBLM_R_X5Y143_SLICE_X6Y143_CQ;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_C3 = CLBLL_L_X4Y144_SLICE_X4Y144_AQ;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_A6 = CLBLL_L_X2Y150_SLICE_X1Y150_A5Q;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_B1 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_B2 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_B3 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_B4 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_B5 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_B6 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_C4 = CLBLM_R_X5Y144_SLICE_X6Y144_CQ;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_C1 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_C2 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_C3 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_C4 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_C5 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_D5 = CLBLM_R_X7Y147_SLICE_X8Y147_DQ;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_C6 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_D6 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_D4 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_D1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_D2 = CLBLL_L_X4Y144_SLICE_X4Y144_AQ;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_D3 = CLBLM_R_X3Y145_SLICE_X2Y145_CQ;
  assign RIOI3_X105Y155_OLOGIC_X1Y155_T1 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_D1 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_D2 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_D3 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_D4 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_D5 = 1'b1;
  assign CLBLL_L_X2Y152_SLICE_X1Y152_D6 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_D1 = CLBLM_R_X5Y159_SLICE_X6Y159_AO6;
  assign RIOI3_X105Y189_OLOGIC_X1Y190_D1 = CLBLM_R_X11Y153_SLICE_X14Y153_AO6;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_D1 = CLBLM_R_X3Y150_SLICE_X2Y150_CO5;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_T1 = 1'b1;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_D2 = CLBLM_R_X7Y153_SLICE_X9Y153_A5Q;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_D3 = CLBLM_R_X7Y152_SLICE_X9Y152_DQ;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_D4 = CLBLM_R_X7Y154_SLICE_X8Y154_AQ;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_D5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_D6 = 1'b1;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_SR = CLBLM_R_X5Y153_SLICE_X7Y153_DO6;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE0 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE1 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE0 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE1 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S0 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S1 = 1'b1;
  assign LIOB33_X0Y63_IOB_X0Y64_O = CLBLL_L_X4Y140_SLICE_X5Y140_BO6;
  assign LIOI3_X0Y51_ILOGIC_X0Y52_D = LIOB33_X0Y51_IOB_X0Y52_I;
  assign LIOI3_X0Y51_ILOGIC_X0Y51_D = LIOB33_X0Y51_IOB_X0Y51_I;
  assign RIOI3_SING_X105Y199_OLOGIC_X1Y199_D1 = CLBLM_R_X11Y149_SLICE_X14Y149_AQ;
  assign RIOB33_X105Y151_IOB_X1Y152_O = 1'b1;
  assign RIOB33_X105Y151_IOB_X1Y151_O = 1'b1;
  assign RIOI3_SING_X105Y199_OLOGIC_X1Y199_T1 = 1'b1;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_A1 = CLBLM_R_X7Y153_SLICE_X8Y153_DO5;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_A2 = CLBLM_R_X3Y151_SLICE_X3Y151_C5Q;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_A3 = CLBLL_L_X4Y154_SLICE_X4Y154_AQ;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_A4 = CLBLM_R_X7Y151_SLICE_X9Y151_AQ;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_A5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_A6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y58_D = LIOB33_X0Y57_IOB_X0Y58_I;
  assign LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y57_D = LIOB33_X0Y57_IOB_X0Y57_I;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_A1 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_A2 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_A3 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_A4 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_A5 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_A6 = 1'b1;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_B1 = CLBLM_R_X7Y153_SLICE_X8Y153_DO6;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_B2 = CLBLM_L_X8Y153_SLICE_X10Y153_CQ;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_B3 = CLBLM_R_X7Y153_SLICE_X9Y153_BQ;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_B1 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_B2 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_A3 = CLBLM_L_X10Y143_SLICE_X12Y143_AQ;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_A4 = CLBLM_R_X5Y144_SLICE_X7Y144_AQ;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_A6 = CLBLL_L_X4Y146_SLICE_X5Y146_A5Q;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_B3 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_B4 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_B5 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_B6 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_A2 = CLBLM_L_X8Y150_SLICE_X11Y150_B5Q;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_C1 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_C2 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_C3 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_C4 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_C5 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_C6 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_B1 = CLBLM_R_X7Y142_SLICE_X8Y142_CO6;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_C2 = CLBLM_R_X5Y144_SLICE_X7Y144_CQ;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_B4 = CLBLM_R_X3Y149_SLICE_X2Y149_A5Q;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_C5 = CLBLM_L_X8Y149_SLICE_X10Y149_B5Q;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_C6 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_D1 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_D2 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_D3 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_D4 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_D5 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_D6 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_D1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_D2 = CLBLM_R_X5Y144_SLICE_X7Y144_AQ;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_D3 = CLBLM_R_X5Y144_SLICE_X7Y144_DQ;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_D4 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_D5 = CLBLM_L_X10Y143_SLICE_X12Y143_BO5;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_D6 = CLBLM_R_X7Y143_SLICE_X9Y143_AQ;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_A6 = CLBLM_R_X3Y153_SLICE_X3Y153_A5Q;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_B1 = CLBLM_R_X7Y154_SLICE_X8Y154_BQ;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_B2 = CLBLL_L_X4Y149_SLICE_X4Y149_D5Q;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_B3 = CLBLM_R_X5Y152_SLICE_X6Y152_C5Q;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_A1 = CLBLM_R_X3Y148_SLICE_X2Y148_D5Q;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_A2 = CLBLM_R_X5Y144_SLICE_X6Y144_DQ;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_A3 = CLBLM_R_X5Y144_SLICE_X6Y144_AQ;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_A4 = CLBLM_L_X8Y147_SLICE_X10Y147_B5Q;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_A6 = CLBLM_R_X3Y146_SLICE_X3Y146_CQ;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_C1 = CLBLM_R_X7Y154_SLICE_X8Y154_DO5;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_C2 = CLBLM_R_X7Y154_SLICE_X8Y154_CQ;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_C3 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_B1 = CLBLL_L_X4Y150_SLICE_X5Y150_C5Q;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_A1 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_A2 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_B4 = CLBLM_L_X8Y143_SLICE_X11Y143_BQ;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_B5 = RIOB33_X105Y119_IOB_X1Y119_I;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_B6 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_A3 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_A4 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_A5 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_A6 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_AX = CLBLM_R_X3Y153_SLICE_X2Y153_AO6;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_B1 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_B2 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_B3 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_B4 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_C6 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_B5 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_B6 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_C5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_C1 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_C2 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_C3 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_C4 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_C5 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_C6 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_D2 = CLBLM_R_X7Y150_SLICE_X9Y150_B5Q;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_D3 = CLBLM_L_X10Y150_SLICE_X13Y150_A5Q;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_D4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_D6 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_D5 = CLBLM_R_X5Y153_SLICE_X7Y153_A5Q;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_D1 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_D1 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_D2 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_D3 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_D4 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_D5 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_D6 = 1'b1;
  assign LIOB33_X0Y65_IOB_X0Y66_O = CLBLM_R_X7Y152_SLICE_X9Y152_DQ;
  assign LIOB33_X0Y65_IOB_X0Y65_O = CLBLL_L_X4Y140_SLICE_X5Y140_CO6;
  assign RIOI3_X105Y135_ILOGIC_X1Y135_D = RIOB33_X105Y135_IOB_X1Y135_I;
  assign RIOB33_X105Y153_IOB_X1Y154_O = 1'b1;
  assign RIOB33_X105Y153_IOB_X1Y153_O = 1'b1;
  assign LIOB33_X0Y185_IOB_X0Y186_O = RIOB33_X105Y119_IOB_X1Y120_I;
  assign LIOB33_X0Y185_IOB_X0Y185_O = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_A1 = 1'b1;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_A2 = 1'b1;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_B1 = CLBLM_R_X3Y147_SLICE_X3Y147_B5Q;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_A3 = CLBLM_R_X7Y154_SLICE_X8Y154_BQ;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_A4 = 1'b1;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_A5 = CLBLM_R_X7Y155_SLICE_X8Y155_AQ;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_A6 = 1'b1;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_B2 = CLBLM_R_X5Y144_SLICE_X6Y144_CQ;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_B1 = 1'b1;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_B2 = 1'b1;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_B3 = CLBLM_L_X10Y147_SLICE_X13Y147_DQ;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_B3 = 1'b1;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_B4 = 1'b1;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_B5 = 1'b1;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_B6 = 1'b1;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_A1 = CLBLM_R_X5Y145_SLICE_X6Y145_DQ;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_A2 = 1'b1;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_A3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_A4 = CLBLL_L_X2Y144_SLICE_X1Y144_A5Q;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_A5 = 1'b1;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_A6 = 1'b1;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_C1 = 1'b1;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_C2 = 1'b1;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_C3 = 1'b1;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_B1 = CLBLM_L_X8Y150_SLICE_X10Y150_A5Q;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_B2 = CLBLL_L_X4Y151_SLICE_X4Y151_AQ;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_B3 = CLBLM_R_X5Y142_SLICE_X7Y142_BQ;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_B4 = CLBLM_R_X11Y149_SLICE_X14Y149_AQ;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_B5 = CLBLM_L_X10Y143_SLICE_X13Y143_AO6;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_B6 = 1'b1;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_D1 = 1'b1;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_D2 = 1'b1;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_C1 = CLBLM_L_X8Y148_SLICE_X10Y148_CO5;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_C2 = CLBLM_R_X5Y142_SLICE_X7Y142_B5Q;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_C3 = CLBLM_R_X5Y145_SLICE_X7Y145_BO6;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_C4 = CLBLL_L_X4Y142_SLICE_X4Y142_CO5;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_C5 = CLBLM_R_X5Y145_SLICE_X7Y145_DO6;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_C6 = CLBLM_R_X5Y151_SLICE_X7Y151_DO6;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_D3 = 1'b1;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_D4 = 1'b1;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_A2 = CLBLM_R_X7Y155_SLICE_X8Y155_BQ;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_A3 = CLBLM_R_X7Y155_SLICE_X8Y155_AQ;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_A4 = CLBLM_R_X5Y150_SLICE_X6Y150_AQ;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_A5 = CLBLM_R_X7Y154_SLICE_X8Y154_BQ;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_D1 = CLBLM_R_X5Y145_SLICE_X6Y145_DQ;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_D2 = CLBLM_L_X8Y142_SLICE_X10Y142_BO5;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_D3 = CLBLM_L_X8Y145_SLICE_X10Y145_CO5;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_D4 = CLBLM_R_X5Y145_SLICE_X7Y145_A5Q;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_D5 = CLBLM_R_X5Y145_SLICE_X7Y145_BO5;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_D6 = 1'b1;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_A6 = CLBLM_R_X5Y152_SLICE_X6Y152_C5Q;
  assign CLBLM_R_X5Y145_SLICE_X7Y145_SR = CLBLL_L_X4Y151_SLICE_X4Y151_CO6;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_B1 = CLBLM_L_X8Y146_SLICE_X11Y146_A5Q;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_B2 = CLBLM_R_X7Y155_SLICE_X8Y155_BQ;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_B3 = CLBLM_R_X7Y155_SLICE_X8Y155_AQ;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_A1 = CLBLM_R_X3Y147_SLICE_X3Y147_BQ;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_A2 = CLBLL_L_X2Y147_SLICE_X1Y147_A5Q;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_A3 = CLBLM_R_X5Y145_SLICE_X6Y145_AQ;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_A4 = CLBLM_R_X5Y153_SLICE_X6Y153_BQ;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_A6 = CLBLM_R_X5Y144_SLICE_X6Y144_CQ;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_C1 = 1'b1;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_C2 = 1'b1;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_C3 = 1'b1;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_B1 = CLBLM_R_X5Y146_SLICE_X7Y146_B5Q;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_B2 = 1'b1;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_B4 = CLBLM_R_X3Y145_SLICE_X2Y145_C5Q;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_B5 = CLBLM_R_X11Y146_SLICE_X14Y146_AQ;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_B6 = 1'b1;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_D1 = 1'b1;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_D2 = 1'b1;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_C2 = CLBLM_R_X5Y145_SLICE_X6Y145_CQ;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_C3 = CLBLM_R_X3Y149_SLICE_X3Y149_CQ;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_C4 = CLBLM_R_X5Y142_SLICE_X6Y142_CQ;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_C5 = 1'b1;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_C6 = CLBLM_L_X10Y143_SLICE_X12Y143_AO6;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_D3 = 1'b1;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_D4 = 1'b1;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_D5 = 1'b1;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_D6 = 1'b1;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_D1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_D2 = 1'b1;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_D3 = CLBLM_R_X5Y145_SLICE_X6Y145_DQ;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_D4 = CLBLM_L_X10Y143_SLICE_X12Y143_BO5;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_D5 = CLBLL_L_X4Y145_SLICE_X4Y145_A5Q;
  assign CLBLM_R_X5Y145_SLICE_X6Y145_D6 = CLBLM_R_X5Y145_SLICE_X6Y145_AQ;
  assign LIOI3_X0Y175_OLOGIC_X0Y176_D1 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign LIOI3_X0Y175_OLOGIC_X0Y176_T1 = 1'b1;
  assign LIOI3_X0Y115_OLOGIC_X0Y116_D1 = CLBLM_R_X5Y152_SLICE_X6Y152_CQ;
  assign LIOI3_X0Y175_OLOGIC_X0Y175_D1 = RIOB33_X105Y123_IOB_X1Y123_I;
  assign LIOI3_X0Y115_OLOGIC_X0Y116_T1 = 1'b1;
  assign RIOI3_X105Y159_OLOGIC_X1Y160_D1 = 1'b1;
  assign LIOI3_X0Y175_OLOGIC_X0Y175_T1 = 1'b1;
  assign LIOI3_X0Y115_OLOGIC_X0Y115_D1 = CLBLM_R_X3Y151_SLICE_X3Y151_CQ;
  assign RIOI3_X105Y159_OLOGIC_X1Y160_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_D1 = CLBLM_R_X3Y150_SLICE_X3Y150_BQ;
  assign LIOI3_X0Y115_OLOGIC_X0Y115_T1 = 1'b1;
  assign RIOI3_X105Y159_OLOGIC_X1Y159_D1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_T1 = 1'b1;
  assign RIOI3_X105Y159_OLOGIC_X1Y159_T1 = 1'b1;
  assign RIOB33_X105Y155_IOB_X1Y156_O = 1'b1;
  assign RIOB33_X105Y155_IOB_X1Y155_O = 1'b1;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_D1 = CLBLM_L_X10Y150_SLICE_X12Y150_CQ;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_T1 = 1'b1;
  assign LIOB33_X0Y187_IOB_X0Y188_O = CLBLM_R_X3Y150_SLICE_X3Y150_BQ;
  assign LIOB33_X0Y187_IOB_X0Y187_O = CLBLM_L_X10Y150_SLICE_X12Y150_CQ;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_A1 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_A2 = CLBLM_L_X8Y143_SLICE_X11Y143_A5Q;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_A3 = CLBLM_R_X5Y146_SLICE_X7Y146_AQ;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_A4 = CLBLM_R_X5Y147_SLICE_X6Y147_BQ;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_A6 = CLBLM_L_X8Y149_SLICE_X11Y149_BQ;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_B1 = CLBLM_R_X3Y152_SLICE_X3Y152_AQ;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_B2 = CLBLM_R_X5Y147_SLICE_X7Y147_A5Q;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_B4 = CLBLM_R_X5Y146_SLICE_X6Y146_B5Q;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_B5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_B6 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_C2 = CLBLM_R_X5Y146_SLICE_X7Y146_CQ;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_C3 = CLBLM_R_X3Y148_SLICE_X3Y148_A5Q;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_C4 = CLBLM_R_X3Y142_SLICE_X3Y142_BQ;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_C5 = CLBLM_R_X5Y149_SLICE_X6Y149_D5Q;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_C6 = CLBLM_L_X8Y150_SLICE_X11Y150_B5Q;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_D1 = CLBLM_R_X11Y145_SLICE_X15Y145_BO5;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_D2 = CLBLL_L_X4Y146_SLICE_X4Y146_DQ;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_D3 = CLBLM_R_X5Y146_SLICE_X7Y146_DQ;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_D4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_D5 = CLBLM_R_X3Y146_SLICE_X3Y146_DQ;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_D6 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_A1 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_A2 = CLBLM_R_X3Y145_SLICE_X2Y145_CQ;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_A3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_A4 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_A5 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_A6 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_B1 = CLBLM_L_X10Y153_SLICE_X13Y153_AQ;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_B2 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_B3 = CLBLL_L_X4Y146_SLICE_X5Y146_BQ;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_B4 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_B6 = 1'b1;
  assign LIOI3_X0Y53_ILOGIC_X0Y54_D = LIOB33_X0Y53_IOB_X0Y54_I;
  assign LIOI3_X0Y53_ILOGIC_X0Y53_D = LIOB33_X0Y53_IOB_X0Y53_I;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_C1 = CLBLM_R_X5Y145_SLICE_X7Y145_BO6;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_C2 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_C3 = CLBLM_R_X5Y146_SLICE_X6Y146_BQ;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_C4 = CLBLM_L_X10Y143_SLICE_X12Y143_DO5;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_C5 = CLBLM_R_X5Y147_SLICE_X6Y147_CQ;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_C6 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_D1 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_D2 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_D3 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_D4 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_D5 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_D6 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_SR = CLBLM_R_X11Y148_SLICE_X14Y148_CO6;
  assign RIOB33_X105Y157_IOB_X1Y158_O = 1'b1;
  assign RIOB33_X105Y157_IOB_X1Y157_O = 1'b1;
  assign LIOB33_X0Y189_IOB_X0Y190_O = CLBLM_R_X7Y155_SLICE_X9Y155_AO6;
  assign LIOB33_X0Y189_IOB_X0Y189_O = CLBLM_R_X3Y149_SLICE_X3Y149_DQ;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_D1 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_B1 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_C3 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_C4 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_B4 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_C5 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_C6 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_B6 = 1'b1;
  assign LIOI3_X0Y61_ILOGIC_X0Y62_D = LIOB33_X0Y61_IOB_X0Y62_I;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_T1 = 1'b1;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_A1 = 1'b1;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_A2 = CLBLM_R_X7Y151_SLICE_X9Y151_DQ;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_A3 = CLBLM_R_X5Y143_SLICE_X7Y143_AQ;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_A4 = 1'b1;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_A6 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_D1 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_D2 = 1'b1;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_B1 = 1'b1;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_B2 = CLBLM_R_X5Y147_SLICE_X6Y147_B5Q;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_B3 = CLBLM_R_X5Y149_SLICE_X6Y149_AQ;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_B4 = 1'b1;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_B6 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_C6 = 1'b1;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_C2 = CLBLM_R_X3Y148_SLICE_X3Y148_A5Q;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_C3 = CLBLM_R_X7Y148_SLICE_X9Y148_CQ;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_C4 = 1'b1;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_C5 = 1'b1;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_C6 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_D5 = 1'b1;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_D6 = 1'b1;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_D1 = 1'b1;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_D2 = CLBLM_L_X8Y151_SLICE_X10Y151_B5Q;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_D3 = CLBLM_R_X5Y140_SLICE_X7Y140_B5Q;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_D4 = 1'b1;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_D5 = 1'b1;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_D6 = 1'b1;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_SR = CLBLM_R_X11Y148_SLICE_X15Y148_BO6;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_A1 = CLBLM_R_X7Y150_SLICE_X9Y150_CQ;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_A2 = CLBLM_R_X5Y151_SLICE_X6Y151_AQ;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_A3 = CLBLM_R_X5Y147_SLICE_X6Y147_AQ;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_A4 = CLBLM_R_X11Y144_SLICE_X14Y144_AQ;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_A5 = CLBLM_L_X8Y146_SLICE_X10Y146_AQ;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_B1 = CLBLM_R_X5Y149_SLICE_X7Y149_C5Q;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_B2 = 1'b1;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_B4 = CLBLM_R_X5Y150_SLICE_X7Y150_A5Q;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_B5 = CLBLM_R_X5Y147_SLICE_X6Y147_CQ;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_B6 = 1'b1;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_B4 = CLBLM_L_X10Y150_SLICE_X12Y150_CQ;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_C1 = CLBLM_R_X5Y142_SLICE_X6Y142_BQ;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_C2 = CLBLM_R_X5Y147_SLICE_X6Y147_CQ;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_C3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_C4 = CLBLM_L_X10Y143_SLICE_X12Y143_AO6;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_C5 = 1'b1;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_C6 = CLBLL_L_X4Y149_SLICE_X5Y149_AQ;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_B5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_B6 = CLBLM_R_X7Y153_SLICE_X9Y153_AQ;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_D1 = CLBLM_L_X8Y142_SLICE_X11Y142_CQ;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_D2 = CLBLL_L_X4Y144_SLICE_X5Y144_DQ;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_D3 = CLBLM_R_X5Y147_SLICE_X6Y147_DQ;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_D4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_D5 = CLBLM_R_X5Y149_SLICE_X7Y149_DQ;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_D6 = CLBLL_L_X2Y146_SLICE_X1Y146_A5Q;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_B1 = CLBLM_R_X11Y149_SLICE_X14Y149_AQ;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_B2 = CLBLM_R_X5Y151_SLICE_X6Y151_BQ;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_B3 = CLBLM_R_X11Y145_SLICE_X14Y145_BQ;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_C1 = CLBLM_R_X7Y154_SLICE_X8Y154_AQ;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_B4 = CLBLM_R_X11Y142_SLICE_X14Y142_DO6;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_C2 = CLBLM_R_X7Y152_SLICE_X9Y152_DQ;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_B5 = CLBLM_L_X8Y150_SLICE_X10Y150_A5Q;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_C3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_B6 = 1'b1;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_C4 = CLBLM_R_X7Y154_SLICE_X9Y154_AO5;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_C5 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_C6 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_B4 = CLBLM_R_X3Y150_SLICE_X3Y150_BQ;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_C1 = CLBLM_L_X10Y142_SLICE_X13Y142_BO6;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_B5 = CLBLM_R_X7Y145_SLICE_X8Y145_B5Q;
  assign LIOB33_X0Y183_IOB_X0Y184_O = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_C2 = CLBLM_L_X10Y146_SLICE_X12Y146_CO6;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_B6 = CLBLM_R_X11Y152_SLICE_X14Y152_A5Q;
  assign LIOB33_X0Y183_IOB_X0Y183_O = RIOB33_X105Y129_IOB_X1Y130_I;
  assign RIOB33_X105Y159_IOB_X1Y159_O = 1'b1;
  assign RIOB33_X105Y159_IOB_X1Y160_O = 1'b1;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_C3 = CLBLM_R_X11Y146_SLICE_X15Y146_CO6;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_C4 = CLBLM_R_X11Y144_SLICE_X14Y144_CO6;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_C5 = CLBLM_R_X11Y147_SLICE_X15Y147_DO6;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_C6 = CLBLM_L_X10Y146_SLICE_X13Y146_DO6;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_D1 = 1'b1;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_D2 = 1'b1;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_D3 = 1'b1;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_D4 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_C4 = CLBLM_R_X11Y152_SLICE_X14Y152_A5Q;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_D5 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_C5 = CLBLM_R_X11Y151_SLICE_X14Y151_AQ;
  assign LIOB33_X0Y191_IOB_X0Y191_O = CLBLL_L_X4Y145_SLICE_X4Y145_BO6;
  assign LIOB33_X0Y191_IOB_X0Y192_O = CLBLL_L_X4Y154_SLICE_X4Y154_AO5;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_D6 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_C6 = CLBLM_L_X10Y152_SLICE_X12Y152_AQ;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_A1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_A2 = CLBLM_R_X7Y153_SLICE_X9Y153_DO5;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_A3 = CLBLM_R_X3Y150_SLICE_X2Y150_CO5;
  assign LIOI3_X0Y177_OLOGIC_X0Y178_D1 = RIOB33_X105Y125_IOB_X1Y125_I;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_SR = CLBLM_R_X11Y148_SLICE_X15Y148_AO6;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_A5 = CLBLM_R_X3Y151_SLICE_X3Y151_BQ;
  assign LIOI3_X0Y177_OLOGIC_X0Y178_T1 = 1'b1;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_D1 = CLBLM_R_X11Y147_SLICE_X15Y147_AQ;
  assign LIOI3_X0Y177_OLOGIC_X0Y177_D1 = RIOB33_X105Y123_IOB_X1Y124_I;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_T1 = 1'b1;
  assign RIOI3_X105Y161_OLOGIC_X1Y162_D1 = CLBLM_L_X10Y150_SLICE_X13Y150_C5Q;
  assign LIOI3_X0Y177_OLOGIC_X0Y177_T1 = 1'b1;
  assign LIOI3_X0Y117_OLOGIC_X0Y117_D1 = CLBLM_R_X7Y144_SLICE_X9Y144_B5Q;
  assign RIOI3_X105Y161_OLOGIC_X1Y162_T1 = 1'b1;
  assign LIOI3_X0Y117_OLOGIC_X0Y117_T1 = 1'b1;
  assign RIOI3_X105Y161_OLOGIC_X1Y161_D1 = CLBLM_L_X8Y153_SLICE_X11Y153_AO5;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_B4 = CLBLM_R_X7Y155_SLICE_X8Y155_BQ;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_A1 = CLBLM_L_X10Y150_SLICE_X13Y150_CQ;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_A2 = CLBLM_R_X7Y149_SLICE_X8Y149_CQ;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_A3 = CLBLM_R_X5Y150_SLICE_X6Y150_AQ;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_A4 = CLBLM_R_X5Y146_SLICE_X7Y146_BQ;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_A5 = CLBLM_R_X5Y143_SLICE_X7Y143_AQ;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_A6 = CLBLM_R_X7Y147_SLICE_X9Y147_BQ;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_B5 = CLBLM_R_X7Y155_SLICE_X8Y155_AQ;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_AX = CLBLM_R_X5Y148_SLICE_X6Y148_AO6;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_B6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_B1 = CLBLM_R_X11Y149_SLICE_X14Y149_AQ;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_B2 = CLBLM_L_X8Y150_SLICE_X10Y150_A5Q;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_B3 = CLBLM_R_X5Y145_SLICE_X7Y145_BO6;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_B4 = CLBLL_L_X4Y144_SLICE_X5Y144_D5Q;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_B5 = CLBLM_L_X10Y144_SLICE_X13Y144_CO6;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_B6 = CLBLM_R_X7Y148_SLICE_X9Y148_CQ;
  assign RIOI3_X105Y161_OLOGIC_X1Y161_T1 = 1'b1;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_C1 = CLBLL_L_X4Y145_SLICE_X5Y145_AO6;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_C2 = CLBLM_L_X8Y146_SLICE_X11Y146_BO6;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_C3 = CLBLM_L_X10Y143_SLICE_X12Y143_BO5;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_C4 = CLBLM_R_X3Y149_SLICE_X3Y149_BQ;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_C5 = CLBLM_R_X5Y148_SLICE_X7Y148_DO6;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_C6 = CLBLM_R_X5Y148_SLICE_X7Y148_BO6;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_D1 = 1'b1;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_D2 = 1'b1;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_D3 = CLBLM_R_X7Y149_SLICE_X8Y149_BQ;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_D4 = CLBLM_R_X5Y149_SLICE_X6Y149_CQ;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_D5 = CLBLM_L_X8Y142_SLICE_X10Y142_BO5;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_D6 = CLBLM_L_X10Y143_SLICE_X12Y143_AO5;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_SR = CLBLL_L_X4Y151_SLICE_X4Y151_CO6;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_A1 = CLBLL_L_X4Y148_SLICE_X4Y148_BO5;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_A3 = CLBLL_L_X4Y149_SLICE_X4Y149_AQ;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_A4 = CLBLL_L_X4Y148_SLICE_X5Y148_AQ;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_A5 = CLBLL_L_X4Y148_SLICE_X5Y148_BQ;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_A6 = 1'b1;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_C4 = CLBLM_R_X7Y151_SLICE_X8Y151_AQ;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_AX = CLBLM_R_X3Y150_SLICE_X2Y150_CO6;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_B1 = CLBLL_L_X2Y150_SLICE_X1Y150_AQ;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_B2 = 1'b1;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_B3 = CLBLL_L_X4Y147_SLICE_X5Y147_DQ;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_B4 = 1'b1;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_B6 = 1'b1;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_C5 = CLBLM_R_X3Y152_SLICE_X2Y152_BQ;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_C6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_C1 = CLBLL_L_X4Y147_SLICE_X4Y147_C5Q;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_C2 = CLBLM_R_X7Y145_SLICE_X8Y145_B5Q;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_C3 = CLBLM_R_X5Y151_SLICE_X6Y151_BQ;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_C4 = CLBLM_L_X10Y150_SLICE_X12Y150_AQ;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_C5 = CLBLL_L_X4Y149_SLICE_X4Y149_D5Q;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_C6 = 1'b1;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_D1 = 1'b1;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_D2 = 1'b1;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_D3 = 1'b1;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_D4 = 1'b1;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_D5 = 1'b1;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_D6 = 1'b1;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_SR = CLBLL_L_X4Y145_SLICE_X5Y145_BO6;
  assign RIOB33_X105Y161_IOB_X1Y162_O = CLBLM_L_X10Y150_SLICE_X13Y150_C5Q;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_D1 = CLBLM_L_X8Y153_SLICE_X11Y153_BQ;
  assign RIOB33_X105Y161_IOB_X1Y161_O = CLBLM_L_X8Y153_SLICE_X11Y153_AO5;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_D2 = CLBLM_R_X7Y154_SLICE_X8Y154_CQ;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_D3 = CLBLM_L_X8Y154_SLICE_X10Y154_AQ;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_D4 = CLBLM_R_X3Y154_SLICE_X3Y154_AQ;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_D5 = CLBLM_R_X5Y154_SLICE_X7Y154_DQ;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_D6 = 1'b1;
  assign LIOB33_X0Y193_IOB_X0Y194_O = RIOB33_X105Y103_IOB_X1Y103_I;
  assign LIOB33_X0Y193_IOB_X0Y193_O = CLBLL_L_X2Y166_SLICE_X0Y166_AO6;
  assign LIOI3_X0Y55_ILOGIC_X0Y56_D = LIOB33_X0Y55_IOB_X0Y56_I;
  assign LIOI3_X0Y55_ILOGIC_X0Y55_D = LIOB33_X0Y55_IOB_X0Y55_I;
  assign RIOI3_X105Y101_ILOGIC_X1Y102_D = RIOB33_X105Y101_IOB_X1Y102_I;
  assign RIOI3_X105Y101_ILOGIC_X1Y101_D = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_A1 = CLBLM_L_X8Y142_SLICE_X10Y142_C5Q;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_A2 = CLBLM_R_X5Y149_SLICE_X6Y149_D5Q;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_A3 = CLBLM_R_X5Y149_SLICE_X7Y149_AQ;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_A4 = CLBLM_R_X3Y150_SLICE_X3Y150_CQ;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_A6 = CLBLM_L_X8Y150_SLICE_X11Y150_B5Q;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_B1 = CLBLM_R_X7Y145_SLICE_X8Y145_CQ;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_B2 = CLBLM_R_X5Y152_SLICE_X6Y152_A5Q;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_B4 = CLBLM_R_X7Y150_SLICE_X8Y150_CQ;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_B5 = CLBLM_R_X7Y144_SLICE_X9Y144_DQ;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_B6 = 1'b1;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_C1 = CLBLM_L_X8Y149_SLICE_X10Y149_AQ;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_C2 = CLBLM_R_X5Y147_SLICE_X7Y147_A5Q;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_C3 = CLBLL_L_X4Y151_SLICE_X5Y151_CQ;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_C5 = CLBLM_R_X3Y151_SLICE_X3Y151_AQ;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_C6 = 1'b1;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_D1 = CLBLM_L_X8Y142_SLICE_X11Y142_CQ;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_D2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_D3 = CLBLM_R_X5Y140_SLICE_X7Y140_B5Q;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_D4 = CLBLM_R_X7Y152_SLICE_X9Y152_C5Q;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_D5 = CLBLM_R_X5Y149_SLICE_X7Y149_AQ;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_D6 = 1'b1;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_A1 = CLBLL_L_X4Y148_SLICE_X5Y148_B5Q;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_A2 = CLBLM_R_X7Y147_SLICE_X8Y147_D5Q;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_A3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_A4 = CLBLM_L_X8Y149_SLICE_X11Y149_CQ;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_A5 = CLBLM_R_X5Y150_SLICE_X6Y150_CQ;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_A6 = 1'b1;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_B5 = CLBLM_L_X8Y144_SLICE_X10Y144_B5Q;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_B6 = 1'b1;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_B1 = CLBLM_L_X10Y150_SLICE_X12Y150_AQ;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_B2 = CLBLM_L_X8Y148_SLICE_X11Y148_DQ;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_B3 = CLBLL_L_X4Y149_SLICE_X4Y149_D5Q;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_B5 = CLBLM_R_X5Y148_SLICE_X6Y148_CO5;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_B6 = CLBLL_L_X4Y152_SLICE_X5Y152_B5Q;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_C1 = CLBLL_L_X4Y147_SLICE_X5Y147_BQ;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_C2 = CLBLM_R_X5Y149_SLICE_X6Y149_CQ;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_C3 = 1'b1;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_C4 = CLBLM_L_X10Y143_SLICE_X12Y143_BO5;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_C5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_C6 = CLBLM_R_X5Y143_SLICE_X6Y143_CQ;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_D1 = CLBLL_L_X4Y150_SLICE_X5Y150_BQ;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_D2 = CLBLM_R_X5Y152_SLICE_X6Y152_DQ;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_D3 = CLBLL_L_X4Y146_SLICE_X5Y146_B5Q;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_D4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_D5 = CLBLM_L_X8Y150_SLICE_X11Y150_B5Q;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_D6 = 1'b1;
  assign RIOB33_X105Y163_IOB_X1Y163_O = CLBLM_L_X10Y149_SLICE_X12Y149_BQ;
  assign RIOB33_X105Y163_IOB_X1Y164_O = CLBLM_R_X11Y151_SLICE_X15Y151_A5Q;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_C3 = CLBLM_R_X7Y146_SLICE_X9Y146_B5Q;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_C4 = CLBLM_L_X8Y150_SLICE_X10Y150_A5Q;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_C5 = CLBLM_R_X11Y142_SLICE_X14Y142_BO5;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_B1 = CLBLM_R_X7Y143_SLICE_X9Y143_DQ;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_C6 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_B2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign LIOB33_X0Y195_IOB_X0Y196_O = CLBLL_L_X4Y154_SLICE_X5Y154_AO6;
  assign LIOB33_X0Y195_IOB_X0Y195_O = CLBLL_L_X2Y152_SLICE_X1Y152_AO6;
  assign LIOI3_X0Y111_OLOGIC_X0Y112_D1 = CLBLM_R_X3Y145_SLICE_X2Y145_B5Q;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_D4 = CLBLM_L_X8Y144_SLICE_X10Y144_B5Q;
  assign LIOI3_X0Y111_OLOGIC_X0Y112_T1 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_B5 = CLBLM_R_X7Y144_SLICE_X9Y144_AQ;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_B6 = CLBLM_R_X5Y144_SLICE_X7Y144_CQ;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_C2 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_C3 = CLBLM_R_X7Y143_SLICE_X8Y143_DQ;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_C4 = CLBLM_L_X8Y145_SLICE_X10Y145_CO5;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_C5 = CLBLM_L_X8Y142_SLICE_X10Y142_BO5;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_D1 = CLBLM_R_X3Y145_SLICE_X2Y145_CQ;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_C6 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_B2 = CLBLM_L_X8Y147_SLICE_X10Y147_B5Q;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_A1 = CLBLM_R_X5Y152_SLICE_X7Y152_CQ;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_A2 = 1'b1;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_A3 = CLBLL_L_X4Y150_SLICE_X5Y150_DQ;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_A4 = 1'b1;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_A6 = 1'b1;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_B1 = CLBLM_R_X5Y150_SLICE_X6Y150_DQ;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_B2 = CLBLM_R_X7Y151_SLICE_X9Y151_DQ;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_B3 = CLBLM_L_X8Y151_SLICE_X10Y151_DQ;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_B4 = CLBLM_L_X8Y152_SLICE_X11Y152_CO6;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_B5 = CLBLM_R_X5Y151_SLICE_X6Y151_DQ;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_B6 = 1'b1;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_C1 = CLBLM_R_X5Y152_SLICE_X7Y152_AQ;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_C2 = CLBLM_R_X7Y150_SLICE_X8Y150_BQ;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_C3 = CLBLM_R_X7Y148_SLICE_X9Y148_BQ;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_C4 = CLBLL_L_X4Y147_SLICE_X4Y147_CQ;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_C5 = CLBLL_L_X4Y149_SLICE_X4Y149_B5Q;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_C6 = CLBLM_R_X5Y150_SLICE_X6Y150_BQ;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_T1 = 1'b1;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_D1 = CLBLM_L_X10Y143_SLICE_X12Y143_AO5;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_D2 = CLBLM_R_X5Y154_SLICE_X7Y154_CQ;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_D3 = 1'b1;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_D4 = CLBLM_L_X8Y142_SLICE_X10Y142_BO5;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_D5 = 1'b1;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_D6 = CLBLL_L_X4Y151_SLICE_X5Y151_BQ;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_SR = CLBLM_R_X11Y148_SLICE_X15Y148_CO6;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_A1 = CLBLM_L_X10Y147_SLICE_X13Y147_BQ;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_A2 = CLBLM_R_X5Y153_SLICE_X6Y153_AQ;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_A3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_A4 = CLBLM_R_X5Y152_SLICE_X6Y152_A5Q;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_A5 = CLBLL_L_X2Y148_SLICE_X0Y148_AQ;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_A6 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_D6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign LIOI3_X0Y179_OLOGIC_X0Y180_D1 = RIOB33_X105Y127_IOB_X1Y127_I;
  assign RIOB33_X105Y165_IOB_X1Y165_O = CLBLM_R_X3Y153_SLICE_X2Y153_AO5;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_B1 = CLBLL_L_X4Y153_SLICE_X5Y153_BQ;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_B2 = CLBLM_R_X7Y146_SLICE_X9Y146_BQ;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_B4 = 1'b1;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_B5 = 1'b1;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_B6 = CLBLM_R_X5Y154_SLICE_X7Y154_CQ;
  assign RIOB33_X105Y165_IOB_X1Y166_O = CLBLM_L_X10Y153_SLICE_X13Y153_AQ;
  assign LIOI3_X0Y179_OLOGIC_X0Y180_T1 = 1'b1;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_C2 = CLBLM_R_X7Y145_SLICE_X9Y145_DQ;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_C2 = 1'b1;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_C3 = CLBLM_L_X8Y152_SLICE_X10Y152_DQ;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_C4 = CLBLL_L_X4Y150_SLICE_X5Y150_AQ;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_C5 = CLBLM_R_X5Y144_SLICE_X6Y144_BQ;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_C6 = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_D1 = CLBLL_L_X4Y149_SLICE_X4Y149_D5Q;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign LIOI3_X0Y179_OLOGIC_X0Y179_D1 = RIOB33_X105Y125_IOB_X1Y126_I;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_T1 = 1'b1;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_D1 = 1'b1;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_D2 = CLBLM_R_X7Y145_SLICE_X8Y145_CQ;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_D3 = CLBLM_R_X5Y150_SLICE_X7Y150_BO5;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_D4 = CLBLM_R_X5Y150_SLICE_X6Y150_DQ;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_D5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_D6 = CLBLM_R_X3Y152_SLICE_X2Y152_BQ;
  assign LIOI3_X0Y179_OLOGIC_X0Y179_T1 = 1'b1;
  assign RIOI3_X105Y165_OLOGIC_X1Y166_D1 = CLBLM_L_X10Y153_SLICE_X13Y153_AQ;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_D1 = CLBLM_L_X8Y146_SLICE_X10Y146_AQ;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_C3 = 1'b1;
  assign RIOI3_X105Y165_OLOGIC_X1Y166_T1 = 1'b1;
  assign LIOB33_X0Y197_IOB_X0Y198_O = 1'b1;
  assign LIOB33_X0Y197_IOB_X0Y197_O = CLBLM_R_X3Y153_SLICE_X3Y153_BO5;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_T1 = 1'b1;
  assign RIOI3_X105Y165_OLOGIC_X1Y165_D1 = CLBLM_R_X3Y153_SLICE_X2Y153_AO5;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_C4 = 1'b1;
  assign RIOI3_X105Y165_OLOGIC_X1Y165_T1 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_C5 = 1'b1;
  assign LIOI3_X0Y173_OLOGIC_X0Y174_D1 = RIOB33_X105Y121_IOB_X1Y122_I;
  assign LIOI3_X0Y59_ILOGIC_X0Y60_D = LIOB33_X0Y59_IOB_X0Y60_I;
  assign LIOI3_X0Y59_ILOGIC_X0Y59_D = LIOB33_X0Y59_IOB_X0Y59_I;
  assign RIOI3_X105Y103_ILOGIC_X1Y104_D = RIOB33_X105Y103_IOB_X1Y104_I;
  assign RIOI3_X105Y103_ILOGIC_X1Y103_D = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_A1 = 1'b1;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_A2 = CLBLL_L_X4Y148_SLICE_X4Y148_BQ;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_A3 = CLBLM_R_X5Y152_SLICE_X6Y152_C5Q;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_A5 = 1'b1;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_A6 = 1'b1;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_B1 = CLBLM_R_X7Y143_SLICE_X9Y143_CQ;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_B2 = CLBLM_R_X3Y151_SLICE_X3Y151_BQ;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_B3 = CLBLL_L_X4Y153_SLICE_X5Y153_BQ;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_B4 = CLBLL_L_X4Y151_SLICE_X5Y151_AQ;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_B5 = CLBLM_R_X7Y143_SLICE_X9Y143_BQ;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_B6 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_A1 = CLBLM_R_X3Y141_SLICE_X3Y141_DO6;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_A2 = CLBLL_L_X4Y142_SLICE_X5Y142_AQ;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_A3 = CLBLM_R_X7Y150_SLICE_X9Y150_B5Q;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_A4 = CLBLM_R_X3Y142_SLICE_X3Y142_BQ;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_A5 = CLBLM_L_X10Y142_SLICE_X12Y142_AQ;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_A6 = CLBLL_L_X4Y141_SLICE_X5Y141_BO5;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_C2 = CLBLM_L_X8Y152_SLICE_X11Y152_CO6;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_C3 = CLBLM_R_X7Y151_SLICE_X9Y151_DQ;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_B1 = CLBLL_L_X4Y141_SLICE_X5Y141_BO5;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_B2 = CLBLL_L_X4Y142_SLICE_X5Y142_AQ;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_B3 = CLBLM_R_X3Y142_SLICE_X3Y142_BQ;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_B4 = CLBLM_R_X5Y142_SLICE_X6Y142_C5Q;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_B5 = CLBLM_R_X3Y141_SLICE_X2Y141_BO6;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_B6 = CLBLM_L_X10Y142_SLICE_X12Y142_AQ;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_D1 = CLBLM_L_X10Y143_SLICE_X12Y143_AO6;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_C1 = CLBLM_R_X3Y141_SLICE_X2Y141_BO6;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_C2 = CLBLL_L_X4Y142_SLICE_X5Y142_AQ;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_C3 = CLBLM_R_X5Y142_SLICE_X6Y142_C5Q;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_C4 = CLBLL_L_X4Y141_SLICE_X5Y141_BO5;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_C5 = CLBLM_R_X5Y144_SLICE_X6Y144_D5Q;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_C6 = CLBLM_R_X3Y142_SLICE_X3Y142_BQ;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_D3 = CLBLM_L_X10Y143_SLICE_X12Y143_BO5;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_D4 = CLBLL_L_X4Y150_SLICE_X5Y150_AQ;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_A1 = CLBLM_R_X3Y148_SLICE_X2Y148_B5Q;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_A3 = CLBLM_R_X5Y151_SLICE_X6Y151_AQ;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_A4 = CLBLM_R_X5Y149_SLICE_X6Y149_BQ;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_A5 = CLBLM_R_X7Y150_SLICE_X8Y150_AQ;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_A6 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_D1 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_D2 = CLBLL_L_X4Y142_SLICE_X5Y142_AQ;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_D3 = CLBLM_R_X5Y142_SLICE_X6Y142_C5Q;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_D4 = CLBLL_L_X4Y143_SLICE_X4Y143_CQ;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_D5 = CLBLM_L_X10Y142_SLICE_X12Y142_AQ;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_D6 = CLBLM_R_X3Y142_SLICE_X3Y142_BQ;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_B1 = CLBLM_R_X7Y152_SLICE_X9Y152_D5Q;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_B2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_B3 = RIOB33_X105Y123_IOB_X1Y124_I;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_B4 = CLBLM_R_X11Y151_SLICE_X15Y151_AQ;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_B5 = CLBLM_R_X5Y153_SLICE_X7Y153_AQ;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_A2 = CLBLL_L_X2Y153_SLICE_X1Y153_AQ;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_A3 = CLBLM_R_X3Y145_SLICE_X2Y145_C5Q;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_A4 = CLBLM_R_X5Y143_SLICE_X6Y143_DQ;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_A5 = CLBLM_R_X3Y146_SLICE_X2Y146_CQ;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_A6 = 1'b1;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_C1 = CLBLL_L_X4Y144_SLICE_X4Y144_BO6;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_C2 = CLBLM_R_X5Y150_SLICE_X7Y150_CO6;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_C3 = CLBLM_R_X7Y145_SLICE_X9Y145_DQ;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_B1 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_B2 = CLBLM_R_X3Y146_SLICE_X2Y146_BQ;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_B3 = CLBLL_L_X4Y143_SLICE_X5Y143_C5Q;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_B4 = CLBLM_R_X3Y145_SLICE_X2Y145_CQ;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_B5 = CLBLM_R_X3Y145_SLICE_X2Y145_B5Q;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_B6 = CLBLM_R_X3Y141_SLICE_X2Y141_AO5;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_D1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_D2 = CLBLM_R_X5Y151_SLICE_X7Y151_CO6;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_C1 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_C2 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_C3 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_C4 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_C5 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_C6 = 1'b1;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_D3 = CLBLM_L_X8Y151_SLICE_X10Y151_DQ;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_D4 = CLBLM_R_X5Y151_SLICE_X6Y151_A5Q;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_D5 = 1'b1;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_D6 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_D1 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_D2 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_D3 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_D4 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_D5 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_D6 = 1'b1;
  assign LIOI3_X0Y173_OLOGIC_X0Y173_T1 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_C4 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_C5 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_C6 = 1'b1;
  assign RIOB33_X105Y169_IOB_X1Y170_O = CLBLM_R_X7Y153_SLICE_X9Y153_CQ;
  assign RIOB33_X105Y169_IOB_X1Y169_O = CLBLM_R_X7Y152_SLICE_X9Y152_BQ;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_A1 = CLBLL_L_X4Y152_SLICE_X5Y152_B5Q;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_A2 = 1'b1;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_A3 = CLBLM_R_X5Y153_SLICE_X6Y153_AQ;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_A4 = CLBLM_L_X8Y149_SLICE_X10Y149_BQ;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_A5 = 1'b1;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_B1 = CLBLM_R_X5Y144_SLICE_X6Y144_DQ;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_B2 = CLBLM_R_X5Y152_SLICE_X7Y152_BQ;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_B3 = CLBLM_R_X7Y150_SLICE_X9Y150_C5Q;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_B4 = CLBLM_R_X5Y151_SLICE_X7Y151_A5Q;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_B5 = CLBLM_R_X3Y148_SLICE_X2Y148_D5Q;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_B6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_A2 = LIOB33_X0Y53_IOB_X0Y54_I;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_A3 = CLBLM_R_X3Y142_SLICE_X3Y142_AQ;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_A4 = CLBLM_R_X3Y143_SLICE_X3Y143_DO6;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_A5 = CLBLM_R_X3Y143_SLICE_X3Y143_CO5;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_A6 = CLBLL_L_X4Y142_SLICE_X5Y142_CQ;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_C2 = CLBLM_R_X5Y152_SLICE_X7Y152_CQ;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_C3 = CLBLM_R_X5Y152_SLICE_X7Y152_BQ;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_B2 = CLBLM_R_X5Y144_SLICE_X6Y144_D5Q;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_B3 = CLBLM_R_X3Y141_SLICE_X3Y141_BO6;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_B4 = CLBLM_R_X3Y142_SLICE_X3Y142_DO6;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_B5 = CLBLM_L_X8Y148_SLICE_X11Y148_CQ;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_B6 = CLBLL_L_X4Y142_SLICE_X4Y142_DO6;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_D1 = CLBLM_R_X3Y147_SLICE_X3Y147_AQ;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_C1 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_C2 = CLBLM_R_X3Y142_SLICE_X3Y142_CQ;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_C3 = CLBLM_R_X3Y145_SLICE_X3Y145_CQ;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_C4 = CLBLM_R_X3Y143_SLICE_X3Y143_CO6;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_C5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_C6 = LIOB33_X0Y53_IOB_X0Y54_I;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_D3 = CLBLM_R_X7Y143_SLICE_X9Y143_CQ;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_D4 = CLBLL_L_X4Y152_SLICE_X5Y152_BQ;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_A1 = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_A2 = CLBLM_R_X7Y152_SLICE_X8Y152_CQ;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_A3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_A4 = CLBLL_L_X4Y150_SLICE_X5Y150_D5Q;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_A5 = CLBLM_R_X3Y150_SLICE_X2Y150_AQ;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_D1 = CLBLL_L_X4Y142_SLICE_X5Y142_AQ;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_D2 = CLBLM_R_X5Y144_SLICE_X6Y144_D5Q;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_D3 = CLBLM_R_X3Y142_SLICE_X3Y142_BQ;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_D4 = CLBLL_L_X4Y143_SLICE_X4Y143_CQ;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_D5 = CLBLM_L_X10Y142_SLICE_X12Y142_AQ;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_D6 = CLBLM_R_X5Y142_SLICE_X6Y142_C5Q;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_A6 = 1'b1;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_B1 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_B2 = CLBLM_R_X5Y152_SLICE_X6Y152_BQ;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_B3 = CLBLL_L_X2Y150_SLICE_X1Y150_A5Q;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_A2 = CLBLM_R_X3Y145_SLICE_X3Y145_A5Q;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_A3 = CLBLM_R_X3Y142_SLICE_X2Y142_AQ;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_A4 = CLBLM_L_X8Y146_SLICE_X10Y146_AQ;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_A5 = CLBLM_R_X7Y150_SLICE_X9Y150_CQ;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_A6 = CLBLM_R_X3Y142_SLICE_X3Y142_CQ;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_C3 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_C5 = CLBLL_L_X4Y153_SLICE_X4Y153_BQ;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_AX = CLBLM_R_X3Y142_SLICE_X2Y142_CO6;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_C6 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_B2 = CLBLL_L_X4Y143_SLICE_X5Y143_C5Q;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_B3 = CLBLM_R_X5Y153_SLICE_X6Y153_DQ;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_B4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_B5 = CLBLM_R_X3Y142_SLICE_X3Y142_AQ;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_B6 = 1'b1;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_D1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_D2 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_C1 = CLBLM_R_X5Y145_SLICE_X7Y145_A5Q;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_C2 = LIOB33_X0Y59_IOB_X0Y60_I;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_C3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_C4 = CLBLM_R_X3Y142_SLICE_X2Y142_A5Q;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_C5 = CLBLM_R_X3Y143_SLICE_X2Y143_DQ;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_C6 = 1'b1;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_D3 = CLBLM_R_X5Y152_SLICE_X6Y152_DQ;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_D4 = CLBLM_R_X7Y153_SLICE_X8Y153_AQ;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_D5 = CLBLM_R_X5Y152_SLICE_X6Y152_BQ;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_D6 = CLBLM_L_X8Y143_SLICE_X11Y143_A5Q;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_A5 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_D1 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_D2 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_D3 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_D4 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_D5 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_D6 = 1'b1;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_C4 = 1'b1;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_C5 = 1'b1;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_C6 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_B3 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_B4 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_B5 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_B6 = 1'b1;
  assign LIOI3_X0Y183_OLOGIC_X0Y184_D1 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign LIOI3_X0Y183_OLOGIC_X0Y184_T1 = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_D1 = CLBLM_R_X7Y152_SLICE_X9Y152_DQ;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_C1 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_C2 = 1'b1;
  assign LIOI3_X0Y183_OLOGIC_X0Y183_D1 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_T1 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_C3 = 1'b1;
  assign RIOI3_X105Y167_OLOGIC_X1Y168_D1 = CLBLM_L_X8Y150_SLICE_X11Y150_CQ;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_C4 = 1'b1;
  assign LIOI3_X0Y183_OLOGIC_X0Y183_T1 = 1'b1;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_D5 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_C5 = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_D1 = CLBLM_R_X3Y149_SLICE_X2Y149_CQ;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_D6 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_C6 = 1'b1;
  assign RIOI3_X105Y167_OLOGIC_X1Y168_T1 = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_T1 = 1'b1;
  assign RIOI3_X105Y167_OLOGIC_X1Y167_D1 = CLBLM_L_X8Y152_SLICE_X10Y152_DQ;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_D1 = CLBLL_L_X4Y143_SLICE_X5Y143_C5Q;
  assign RIOI3_X105Y167_OLOGIC_X1Y167_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_D1 = CLBLM_R_X3Y145_SLICE_X2Y145_C5Q;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_T1 = 1'b1;
  assign RIOB33_X105Y171_IOB_X1Y172_O = CLBLL_L_X4Y145_SLICE_X5Y145_AQ;
  assign RIOB33_X105Y171_IOB_X1Y171_O = CLBLM_R_X7Y153_SLICE_X8Y153_CO5;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_D5 = 1'b1;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_A2 = 1'b1;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_A3 = 1'b1;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_A4 = CLBLM_L_X8Y151_SLICE_X11Y151_A5Q;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_A5 = CLBLM_R_X7Y155_SLICE_X8Y155_BQ;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_A6 = 1'b1;
  assign LIOB33_SING_X0Y149_IOB_X0Y149_O = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_B1 = CLBLM_R_X7Y150_SLICE_X9Y150_C5Q;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_B2 = CLBLL_L_X4Y153_SLICE_X5Y153_CO6;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_B3 = CLBLM_R_X7Y149_SLICE_X9Y149_DQ;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_B4 = CLBLM_L_X10Y150_SLICE_X12Y150_CQ;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_B5 = CLBLM_R_X7Y144_SLICE_X9Y144_B5Q;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_B6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_B5 = CLBLM_R_X7Y154_SLICE_X8Y154_BQ;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_B6 = CLBLM_R_X5Y152_SLICE_X6Y152_C5Q;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_A1 = CLBLM_R_X3Y143_SLICE_X3Y143_BO5;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_A2 = CLBLM_R_X3Y145_SLICE_X3Y145_BQ;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_A3 = CLBLM_R_X3Y143_SLICE_X3Y143_AQ;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_A5 = CLBLL_L_X2Y143_SLICE_X1Y143_BQ;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_A6 = CLBLM_R_X3Y145_SLICE_X3Y145_CQ;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_C1 = CLBLM_R_X3Y150_SLICE_X2Y150_CO5;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_C2 = CLBLM_L_X10Y150_SLICE_X12Y150_CQ;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_C3 = CLBLL_L_X4Y154_SLICE_X4Y154_AQ;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_B1 = LIOB33_X0Y53_IOB_X0Y54_I;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_B2 = CLBLM_R_X3Y143_SLICE_X3Y143_CO6;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_B3 = CLBLM_R_X3Y142_SLICE_X3Y142_CQ;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_B4 = CLBLM_R_X3Y143_SLICE_X2Y143_BQ;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_B6 = 1'b1;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_D1 = 1'b1;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_C1 = CLBLM_R_X3Y142_SLICE_X3Y142_AQ;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_C2 = CLBLM_R_X3Y145_SLICE_X3Y145_BQ;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_C3 = 1'b1;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_C4 = CLBLM_R_X3Y145_SLICE_X3Y145_CQ;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_C5 = CLBLM_R_X3Y143_SLICE_X3Y143_AQ;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_C6 = 1'b1;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_D3 = 1'b1;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_D4 = 1'b1;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_A1 = CLBLM_R_X5Y153_SLICE_X6Y153_CQ;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_A2 = CLBLL_L_X2Y148_SLICE_X0Y148_B5Q;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_A3 = CLBLM_R_X5Y153_SLICE_X6Y153_AQ;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_A4 = CLBLM_R_X3Y152_SLICE_X2Y152_DO6;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_A5 = 1'b1;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_D1 = CLBLM_R_X3Y142_SLICE_X3Y142_AQ;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_D2 = CLBLM_R_X3Y142_SLICE_X3Y142_CQ;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_D3 = CLBLM_R_X3Y145_SLICE_X3Y145_BQ;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_D4 = CLBLM_R_X3Y145_SLICE_X3Y145_CQ;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_D5 = CLBLM_R_X3Y143_SLICE_X3Y143_AQ;
  assign CLBLM_R_X3Y143_SLICE_X3Y143_D6 = CLBLM_R_X3Y143_SLICE_X2Y143_BQ;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_B1 = CLBLM_R_X5Y152_SLICE_X7Y152_DQ;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_B2 = CLBLM_R_X5Y153_SLICE_X6Y153_BQ;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_B3 = CLBLM_R_X5Y153_SLICE_X6Y153_CQ;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_B4 = CLBLM_R_X7Y152_SLICE_X9Y152_D5Q;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_A2 = CLBLM_R_X3Y143_SLICE_X2Y143_DQ;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_A3 = CLBLM_R_X3Y142_SLICE_X2Y142_A5Q;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_A4 = CLBLL_L_X2Y150_SLICE_X1Y150_DO5;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_A5 = CLBLM_R_X5Y149_SLICE_X6Y149_BQ;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_A6 = LIOB33_X0Y59_IOB_X0Y60_I;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_C1 = CLBLM_R_X5Y153_SLICE_X6Y153_BQ;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_C2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_C3 = 1'b1;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_B1 = LIOB33_X0Y53_IOB_X0Y54_I;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_B2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_B3 = CLBLM_R_X3Y143_SLICE_X3Y143_CO6;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_B4 = CLBLM_L_X8Y143_SLICE_X11Y143_DQ;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_B5 = CLBLM_R_X3Y143_SLICE_X2Y143_BQ;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_B6 = CLBLM_R_X3Y142_SLICE_X3Y142_CQ;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_D1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_D2 = CLBLM_L_X10Y143_SLICE_X12Y143_BO6;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_C1 = CLBLM_R_X3Y143_SLICE_X2Y143_BQ;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_C2 = CLBLM_R_X3Y143_SLICE_X2Y143_CQ;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_C3 = CLBLL_L_X4Y154_SLICE_X4Y154_AQ;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_C4 = CLBLM_R_X3Y142_SLICE_X3Y142_CQ;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_C5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_C6 = CLBLM_R_X3Y143_SLICE_X3Y143_CO6;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_D3 = CLBLM_R_X5Y153_SLICE_X6Y153_DQ;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_D4 = CLBLM_R_X7Y154_SLICE_X8Y154_AQ;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_D5 = 1'b1;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_D6 = CLBLM_R_X3Y152_SLICE_X2Y152_CQ;
  assign LIOI3_X0Y61_ILOGIC_X0Y61_D = LIOB33_X0Y61_IOB_X0Y61_I;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_D1 = CLBLL_L_X4Y141_SLICE_X5Y141_AQ;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_D2 = 1'b1;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_D3 = CLBLM_R_X3Y143_SLICE_X2Y143_DQ;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_D4 = 1'b1;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_D5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y143_SLICE_X2Y143_D6 = LIOB33_X0Y59_IOB_X0Y60_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y106_D = RIOB33_X105Y105_IOB_X1Y106_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y105_D = RIOB33_X105Y105_IOB_X1Y105_I;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_D = RIOB33_X105Y113_IOB_X1Y113_I;
  assign RIOB33_X105Y173_IOB_X1Y174_O = CLBLM_R_X5Y159_SLICE_X6Y159_AO6;
  assign RIOB33_X105Y173_IOB_X1Y173_O = CLBLM_R_X5Y151_SLICE_X6Y151_CQ;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_A1 = 1'b1;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_A2 = CLBLM_R_X5Y154_SLICE_X7Y154_BQ;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_A3 = CLBLM_R_X5Y154_SLICE_X7Y154_AQ;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_A4 = CLBLM_R_X7Y149_SLICE_X8Y149_BQ;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_A5 = CLBLL_L_X4Y152_SLICE_X5Y152_C5Q;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_B1 = CLBLM_R_X7Y153_SLICE_X9Y153_BQ;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_B2 = CLBLM_R_X5Y154_SLICE_X7Y154_BQ;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_B3 = CLBLM_R_X5Y154_SLICE_X7Y154_AQ;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_B4 = 1'b1;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_B5 = CLBLL_L_X4Y152_SLICE_X5Y152_C5Q;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_B6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_A1 = CLBLM_R_X3Y147_SLICE_X3Y147_DO6;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_A3 = CLBLM_R_X3Y145_SLICE_X3Y145_DQ;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_A4 = CLBLM_R_X5Y144_SLICE_X6Y144_AQ;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_A5 = CLBLL_L_X2Y148_SLICE_X0Y148_AQ;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_A6 = 1'b1;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_C1 = CLBLM_L_X8Y152_SLICE_X11Y152_BQ;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_C2 = CLBLM_R_X5Y154_SLICE_X7Y154_CQ;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_C3 = 1'b1;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_B1 = CLBLM_R_X7Y144_SLICE_X9Y144_D5Q;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_B2 = CLBLM_R_X3Y144_SLICE_X3Y144_BQ;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_B4 = CLBLM_R_X5Y144_SLICE_X6Y144_CQ;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_B5 = CLBLL_L_X2Y146_SLICE_X1Y146_AQ;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_B6 = CLBLM_R_X3Y147_SLICE_X3Y147_BQ;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_D1 = CLBLM_R_X3Y154_SLICE_X3Y154_AQ;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_C1 = CLBLM_R_X3Y145_SLICE_X3Y145_AQ;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_C2 = CLBLM_R_X3Y144_SLICE_X3Y144_CQ;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_C3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_C4 = CLBLL_L_X4Y144_SLICE_X4Y144_DO6;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_C5 = CLBLL_L_X2Y148_SLICE_X0Y148_B5Q;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_C6 = CLBLM_R_X5Y144_SLICE_X7Y144_CQ;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_D3 = CLBLM_R_X5Y154_SLICE_X7Y154_DQ;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_D4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_A1 = CLBLL_L_X2Y150_SLICE_X1Y150_AQ;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_A2 = CLBLM_L_X8Y153_SLICE_X10Y153_CQ;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_A3 = CLBLM_R_X5Y154_SLICE_X6Y154_AQ;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_A4 = 1'b1;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_D1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_D2 = CLBLM_R_X3Y143_SLICE_X3Y143_AQ;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_D3 = CLBLM_R_X3Y144_SLICE_X3Y144_DQ;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_D4 = CLBLL_L_X2Y153_SLICE_X1Y153_AQ;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_D5 = CLBLL_L_X4Y152_SLICE_X5Y152_C5Q;
  assign CLBLM_R_X3Y144_SLICE_X3Y144_D6 = 1'b1;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_A6 = CLBLM_L_X10Y143_SLICE_X12Y143_AO6;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_B1 = 1'b1;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_B2 = 1'b1;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_B3 = 1'b1;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_B4 = 1'b1;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_A1 = 1'b1;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_A3 = 1'b1;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_A4 = CLBLM_R_X3Y144_SLICE_X3Y144_BQ;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_A5 = CLBLM_L_X8Y142_SLICE_X11Y142_CQ;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_A6 = 1'b1;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_C1 = 1'b1;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_C2 = 1'b1;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_C3 = 1'b1;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_B1 = CLBLM_R_X3Y146_SLICE_X2Y146_CQ;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_B2 = CLBLM_R_X3Y142_SLICE_X2Y142_BQ;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_B4 = CLBLM_R_X3Y145_SLICE_X2Y145_BQ;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_B5 = CLBLL_L_X4Y143_SLICE_X5Y143_C5Q;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_B6 = 1'b1;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_D1 = 1'b1;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_D2 = 1'b1;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_D3 = 1'b1;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_C1 = CLBLM_R_X5Y148_SLICE_X7Y148_AO6;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_C2 = CLBLM_R_X7Y144_SLICE_X9Y144_CQ;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_C3 = CLBLL_L_X2Y147_SLICE_X0Y147_B5Q;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_C4 = CLBLM_R_X5Y142_SLICE_X7Y142_AO5;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_C5 = CLBLL_L_X2Y147_SLICE_X0Y147_AQ;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_C6 = 1'b1;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_D4 = 1'b1;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_D5 = 1'b1;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_D6 = 1'b1;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_C1 = CLBLM_R_X5Y142_SLICE_X7Y142_C5Q;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_C2 = CLBLM_L_X8Y144_SLICE_X10Y144_B5Q;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_D1 = 1'b1;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_D2 = 1'b1;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_D3 = 1'b1;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_D4 = 1'b1;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_D5 = 1'b1;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_D6 = 1'b1;
  assign CLBLM_R_X3Y144_SLICE_X2Y144_SR = CLBLM_R_X3Y146_SLICE_X2Y146_DO6;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_C5 = CLBLM_L_X8Y144_SLICE_X11Y144_A5Q;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_C2 = CLBLM_L_X10Y141_SLICE_X12Y141_AO6;
  assign LIOI3_X0Y173_OLOGIC_X0Y174_T1 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_C3 = CLBLM_R_X7Y151_SLICE_X9Y151_BQ;
  assign RIOB33_X105Y175_IOB_X1Y176_O = CLBLL_L_X2Y151_SLICE_X1Y151_CO6;
  assign RIOB33_X105Y175_IOB_X1Y175_O = CLBLM_R_X3Y153_SLICE_X3Y153_CO6;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_B2 = CLBLM_R_X7Y149_SLICE_X8Y149_AQ;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_B3 = CLBLM_R_X3Y149_SLICE_X3Y149_CQ;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_B4 = CLBLM_R_X7Y143_SLICE_X8Y143_CQ;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_B5 = CLBLM_R_X5Y149_SLICE_X7Y149_B5Q;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_B6 = 1'b1;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_C1 = CLBLM_R_X7Y144_SLICE_X9Y144_D5Q;
  assign LIOI3_X0Y185_OLOGIC_X0Y186_D1 = RIOB33_X105Y119_IOB_X1Y120_I;
  assign LIOI3_X0Y185_OLOGIC_X0Y186_T1 = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_D1 = CLBLM_R_X5Y144_SLICE_X6Y144_CQ;
  assign LIOI3_X0Y185_OLOGIC_X0Y185_D1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_T1 = 1'b1;
  assign RIOI3_X105Y171_OLOGIC_X1Y172_D1 = CLBLL_L_X4Y145_SLICE_X5Y145_AQ;
  assign LIOI3_X0Y65_OLOGIC_X0Y66_D1 = CLBLM_R_X7Y152_SLICE_X9Y152_DQ;
  assign LIOI3_X0Y185_OLOGIC_X0Y185_T1 = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_D1 = CLBLM_R_X5Y144_SLICE_X6Y144_DQ;
  assign RIOI3_X105Y171_OLOGIC_X1Y172_T1 = 1'b1;
  assign LIOI3_X0Y65_OLOGIC_X0Y66_T1 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_A1 = CLBLM_R_X3Y146_SLICE_X3Y146_BQ;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_A3 = CLBLM_R_X3Y146_SLICE_X3Y146_AQ;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_A4 = CLBLL_L_X4Y150_SLICE_X5Y150_CQ;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_A5 = CLBLL_L_X4Y141_SLICE_X4Y141_AQ;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_A6 = 1'b1;
  assign LIOI3_X0Y65_OLOGIC_X0Y65_D1 = CLBLL_L_X4Y140_SLICE_X5Y140_CO6;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_T1 = 1'b1;
  assign RIOI3_X105Y171_OLOGIC_X1Y171_D1 = CLBLM_R_X7Y153_SLICE_X8Y153_CO5;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_B1 = CLBLM_R_X3Y145_SLICE_X3Y145_CQ;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_B2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_B3 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_B4 = CLBLM_R_X3Y143_SLICE_X3Y143_BO6;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_B5 = CLBLM_R_X11Y147_SLICE_X14Y147_AQ;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_B6 = CLBLM_R_X3Y145_SLICE_X3Y145_BQ;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_D1 = CLBLM_R_X3Y150_SLICE_X3Y150_AQ;
  assign LIOI3_X0Y65_OLOGIC_X0Y65_T1 = 1'b1;
  assign RIOI3_X105Y171_OLOGIC_X1Y171_T1 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_C1 = CLBLM_R_X3Y143_SLICE_X3Y143_BO6;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_C2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_C3 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_C4 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_C5 = CLBLM_R_X3Y145_SLICE_X3Y145_CQ;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_C6 = CLBLM_R_X3Y151_SLICE_X2Y151_BQ;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_T1 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_D1 = CLBLM_R_X3Y147_SLICE_X2Y147_AQ;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_D2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_D3 = CLBLM_R_X3Y145_SLICE_X3Y145_DQ;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_D4 = CLBLM_R_X5Y149_SLICE_X7Y149_DQ;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_D5 = CLBLL_L_X2Y145_SLICE_X1Y145_A5Q;
  assign CLBLM_R_X3Y145_SLICE_X3Y145_D6 = CLBLM_L_X8Y142_SLICE_X11Y142_CQ;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_D6 = CLBLM_R_X7Y151_SLICE_X8Y151_BQ;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_D1 = CLBLM_R_X3Y149_SLICE_X2Y149_CQ;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_A1 = CLBLM_R_X3Y146_SLICE_X2Y146_B5Q;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_A2 = CLBLM_R_X3Y148_SLICE_X2Y148_D5Q;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_A3 = CLBLM_R_X5Y144_SLICE_X6Y144_DQ;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_A5 = CLBLM_R_X3Y144_SLICE_X2Y144_AQ;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_A6 = CLBLM_R_X3Y145_SLICE_X2Y145_AQ;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_T1 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_B1 = CLBLM_R_X3Y146_SLICE_X2Y146_CQ;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_B2 = CLBLL_L_X4Y148_SLICE_X4Y148_A5Q;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_B3 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_B4 = CLBLL_L_X4Y148_SLICE_X5Y148_CQ;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_B6 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_C2 = CLBLM_R_X3Y145_SLICE_X2Y145_B5Q;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_C3 = CLBLM_R_X5Y146_SLICE_X6Y146_AQ;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_C4 = CLBLM_R_X5Y144_SLICE_X6Y144_D5Q;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_C5 = CLBLL_L_X2Y145_SLICE_X1Y145_A5Q;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_C6 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_D1 = CLBLM_R_X3Y143_SLICE_X2Y143_AQ;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_D2 = 1'b1;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_D3 = CLBLM_R_X3Y145_SLICE_X2Y145_DQ;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_D4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_D5 = CLBLM_R_X3Y146_SLICE_X2Y146_B5Q;
  assign CLBLM_R_X3Y145_SLICE_X2Y145_D6 = CLBLL_L_X2Y153_SLICE_X1Y153_AQ;
  assign RIOB33_X105Y177_IOB_X1Y178_O = CLBLM_R_X3Y150_SLICE_X3Y150_BQ;
  assign RIOB33_X105Y177_IOB_X1Y177_O = CLBLM_L_X10Y142_SLICE_X12Y142_AQ;
  assign LIOI3_X0Y173_OLOGIC_X0Y173_D1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign RIOI3_X105Y109_ILOGIC_X1Y110_D = RIOB33_X105Y109_IOB_X1Y110_I;
  assign RIOI3_X105Y109_ILOGIC_X1Y109_D = RIOB33_X105Y109_IOB_X1Y109_I;
  assign RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y138_D = RIOB33_X105Y137_IOB_X1Y138_I;
  assign RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y137_D = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_A1 = CLBLM_R_X3Y146_SLICE_X3Y146_CQ;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_A2 = 1'b1;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_A3 = CLBLM_R_X3Y146_SLICE_X3Y146_AQ;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_A4 = CLBLM_R_X7Y142_SLICE_X9Y142_D5Q;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_A6 = CLBLM_R_X3Y147_SLICE_X3Y147_CO6;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_B1 = CLBLM_R_X7Y150_SLICE_X9Y150_CQ;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_B2 = CLBLM_R_X3Y146_SLICE_X3Y146_BQ;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_B3 = CLBLL_L_X2Y144_SLICE_X0Y144_AQ;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_B4 = CLBLM_L_X8Y146_SLICE_X10Y146_AQ;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_B6 = CLBLM_R_X3Y148_SLICE_X2Y148_CQ;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_C1 = CLBLM_R_X5Y143_SLICE_X6Y143_DQ;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_C2 = CLBLM_R_X5Y149_SLICE_X6Y149_AQ;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_C3 = CLBLM_R_X3Y145_SLICE_X3Y145_BQ;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_C5 = CLBLL_L_X4Y143_SLICE_X5Y143_C5Q;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_C6 = 1'b1;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_D1 = CLBLL_L_X2Y144_SLICE_X1Y144_A5Q;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_D2 = CLBLM_L_X8Y142_SLICE_X11Y142_CQ;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_D3 = CLBLM_R_X3Y146_SLICE_X3Y146_DQ;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_D4 = CLBLM_R_X5Y149_SLICE_X7Y149_DQ;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_D5 = CLBLM_R_X3Y147_SLICE_X2Y147_CQ;
  assign CLBLM_R_X3Y146_SLICE_X3Y146_D6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_A2 = CLBLM_R_X5Y144_SLICE_X6Y144_DQ;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_A3 = CLBLM_R_X3Y146_SLICE_X2Y146_AQ;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_A4 = CLBLM_R_X3Y148_SLICE_X2Y148_D5Q;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_A5 = CLBLL_L_X2Y144_SLICE_X0Y144_AQ;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_A6 = CLBLM_R_X3Y151_SLICE_X3Y151_AQ;
  assign LIOB33_X0Y139_IOB_X0Y139_O = CLBLL_L_X2Y148_SLICE_X0Y148_AQ;
  assign LIOB33_X0Y139_IOB_X0Y140_O = CLBLL_L_X2Y147_SLICE_X0Y147_BQ;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_B1 = LIOB33_X0Y59_IOB_X0Y59_I;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_B2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_B3 = CLBLM_R_X3Y146_SLICE_X2Y146_AQ;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_B4 = CLBLM_R_X3Y147_SLICE_X2Y147_BQ;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_B5 = CLBLL_L_X4Y143_SLICE_X5Y143_C5Q;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_B6 = 1'b1;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_C1 = CLBLM_R_X3Y145_SLICE_X2Y145_C5Q;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_C2 = CLBLM_R_X3Y145_SLICE_X3Y145_A5Q;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_C3 = CLBLM_R_X3Y150_SLICE_X2Y150_B5Q;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_C5 = RIOB33_X105Y121_IOB_X1Y122_I;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_C6 = 1'b1;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_D1 = CLBLL_L_X4Y150_SLICE_X5Y150_CQ;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_D2 = 1'b1;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_D3 = 1'b1;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_D4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_D5 = 1'b1;
  assign CLBLM_R_X3Y146_SLICE_X2Y146_D6 = 1'b1;
  assign RIOB33_X105Y179_IOB_X1Y180_O = CLBLM_L_X10Y150_SLICE_X12Y150_CQ;
  assign RIOB33_X105Y179_IOB_X1Y179_O = CLBLM_R_X3Y149_SLICE_X3Y149_DQ;
  assign CLBLL_L_X2Y166_SLICE_X0Y166_A1 = 1'b1;
  assign CLBLL_L_X2Y166_SLICE_X0Y166_A2 = 1'b1;
  assign CLBLL_L_X2Y166_SLICE_X0Y166_A3 = 1'b1;
  assign CLBLL_L_X2Y166_SLICE_X0Y166_A4 = 1'b1;
  assign CLBLL_L_X2Y166_SLICE_X0Y166_A5 = CLBLM_R_X11Y143_SLICE_X14Y143_AQ;
  assign CLBLL_L_X2Y166_SLICE_X0Y166_A6 = 1'b1;
  assign CLBLL_L_X2Y166_SLICE_X0Y166_B1 = 1'b1;
  assign CLBLL_L_X2Y166_SLICE_X0Y166_B2 = 1'b1;
  assign CLBLL_L_X2Y166_SLICE_X0Y166_B3 = 1'b1;
  assign CLBLL_L_X2Y166_SLICE_X0Y166_B4 = 1'b1;
  assign CLBLL_L_X2Y166_SLICE_X0Y166_B5 = 1'b1;
  assign CLBLL_L_X2Y166_SLICE_X0Y166_B6 = 1'b1;
  assign CLBLL_L_X2Y166_SLICE_X0Y166_C1 = 1'b1;
  assign CLBLL_L_X2Y166_SLICE_X0Y166_C2 = 1'b1;
  assign CLBLL_L_X2Y166_SLICE_X0Y166_C3 = 1'b1;
  assign CLBLL_L_X2Y166_SLICE_X0Y166_C4 = 1'b1;
  assign CLBLL_L_X2Y166_SLICE_X0Y166_C5 = 1'b1;
  assign CLBLL_L_X2Y166_SLICE_X0Y166_C6 = 1'b1;
  assign CLBLL_L_X2Y166_SLICE_X0Y166_D1 = 1'b1;
  assign CLBLL_L_X2Y166_SLICE_X0Y166_D2 = 1'b1;
  assign CLBLL_L_X2Y166_SLICE_X0Y166_D3 = 1'b1;
  assign CLBLL_L_X2Y166_SLICE_X0Y166_D4 = 1'b1;
  assign CLBLL_L_X2Y166_SLICE_X0Y166_D5 = 1'b1;
  assign CLBLL_L_X2Y166_SLICE_X0Y166_D6 = 1'b1;
  assign RIOI3_X105Y189_OLOGIC_X1Y190_T1 = 1'b1;
  assign CLBLL_L_X2Y166_SLICE_X1Y166_A1 = 1'b1;
  assign CLBLL_L_X2Y166_SLICE_X1Y166_A2 = 1'b1;
  assign CLBLL_L_X2Y166_SLICE_X1Y166_A3 = 1'b1;
  assign CLBLL_L_X2Y166_SLICE_X1Y166_A4 = 1'b1;
  assign CLBLL_L_X2Y166_SLICE_X1Y166_A5 = 1'b1;
  assign CLBLL_L_X2Y166_SLICE_X1Y166_A6 = 1'b1;
  assign CLBLL_L_X2Y166_SLICE_X1Y166_B1 = 1'b1;
  assign CLBLL_L_X2Y166_SLICE_X1Y166_B2 = 1'b1;
  assign CLBLL_L_X2Y166_SLICE_X1Y166_B3 = 1'b1;
  assign CLBLL_L_X2Y166_SLICE_X1Y166_B4 = 1'b1;
  assign CLBLL_L_X2Y166_SLICE_X1Y166_B5 = 1'b1;
  assign CLBLL_L_X2Y166_SLICE_X1Y166_B6 = 1'b1;
  assign CLBLL_L_X2Y166_SLICE_X1Y166_C1 = 1'b1;
  assign CLBLL_L_X2Y166_SLICE_X1Y166_C2 = 1'b1;
  assign CLBLL_L_X2Y166_SLICE_X1Y166_C3 = 1'b1;
  assign CLBLL_L_X2Y166_SLICE_X1Y166_C4 = 1'b1;
  assign CLBLL_L_X2Y166_SLICE_X1Y166_C5 = 1'b1;
  assign CLBLL_L_X2Y166_SLICE_X1Y166_C6 = 1'b1;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_A1 = CLBLL_L_X2Y147_SLICE_X0Y147_BQ;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_A2 = CLBLL_L_X4Y148_SLICE_X4Y148_CO6;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_A3 = CLBLM_R_X3Y146_SLICE_X3Y146_CQ;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_A5 = CLBLM_R_X3Y147_SLICE_X3Y147_CO5;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_A6 = CLBLM_R_X3Y147_SLICE_X3Y147_AQ;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_AX = CLBLM_R_X3Y147_SLICE_X2Y147_DO5;
  assign CLBLL_L_X2Y166_SLICE_X1Y166_D1 = 1'b1;
  assign CLBLL_L_X2Y166_SLICE_X1Y166_D2 = 1'b1;
  assign CLBLL_L_X2Y166_SLICE_X1Y166_D3 = 1'b1;
  assign CLBLL_L_X2Y166_SLICE_X1Y166_D4 = 1'b1;
  assign CLBLL_L_X2Y166_SLICE_X1Y166_D5 = 1'b1;
  assign CLBLL_L_X2Y166_SLICE_X1Y166_D6 = 1'b1;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_B5 = CLBLM_R_X5Y147_SLICE_X6Y147_AQ;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_B6 = 1'b1;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_C1 = CLBLM_R_X3Y148_SLICE_X2Y148_AQ;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_C2 = CLBLL_L_X4Y147_SLICE_X4Y147_BQ;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_C3 = CLBLL_L_X4Y148_SLICE_X4Y148_CO6;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_C4 = CLBLM_R_X3Y147_SLICE_X3Y147_AQ;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_C5 = CLBLM_R_X3Y146_SLICE_X3Y146_AQ;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_C6 = 1'b1;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_D1 = CLBLM_R_X3Y147_SLICE_X2Y147_AQ;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_D2 = CLBLM_R_X3Y147_SLICE_X2Y147_BQ;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_D3 = CLBLM_R_X3Y147_SLICE_X3Y147_A5Q;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_D4 = CLBLM_R_X3Y150_SLICE_X3Y150_BQ;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_D5 = CLBLM_R_X3Y144_SLICE_X3Y144_AQ;
  assign CLBLM_R_X3Y147_SLICE_X3Y147_D6 = CLBLM_R_X5Y153_SLICE_X7Y153_BO6;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_A1 = CLBLM_R_X3Y147_SLICE_X2Y147_DO6;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_A2 = CLBLM_R_X3Y147_SLICE_X2Y147_BQ;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_A3 = CLBLM_R_X3Y147_SLICE_X2Y147_AQ;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_A4 = CLBLM_R_X5Y153_SLICE_X7Y153_BO6;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_A5 = CLBLM_R_X7Y144_SLICE_X8Y144_BQ;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_B1 = CLBLM_R_X3Y147_SLICE_X3Y147_A5Q;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_B2 = CLBLM_R_X3Y147_SLICE_X2Y147_BQ;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_B4 = CLBLM_R_X3Y150_SLICE_X3Y150_BQ;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_B5 = CLBLM_R_X3Y146_SLICE_X2Y146_C5Q;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_B6 = CLBLM_R_X5Y153_SLICE_X7Y153_BO6;
  assign LIOI3_X0Y189_OLOGIC_X0Y190_D1 = CLBLM_R_X7Y155_SLICE_X9Y155_AO6;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_C1 = CLBLM_R_X3Y151_SLICE_X2Y151_AQ;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_C2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_C3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_C4 = CLBLM_R_X5Y147_SLICE_X7Y147_AQ;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_C5 = CLBLM_R_X3Y146_SLICE_X3Y146_DQ;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_C6 = 1'b1;
  assign LIOI3_X0Y189_OLOGIC_X0Y190_T1 = 1'b1;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_D1 = CLBLM_L_X8Y142_SLICE_X11Y142_CQ;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_D1 = CLBLM_R_X11Y147_SLICE_X15Y147_AQ;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_D2 = CLBLM_R_X3Y147_SLICE_X3Y147_A5Q;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_D3 = CLBLM_R_X3Y150_SLICE_X3Y150_BQ;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_D4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_D5 = CLBLM_R_X5Y153_SLICE_X7Y153_BO6;
  assign CLBLM_R_X3Y147_SLICE_X2Y147_D6 = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_T1 = 1'b1;
  assign LIOI3_X0Y189_OLOGIC_X0Y189_D1 = CLBLM_R_X3Y149_SLICE_X3Y149_DQ;
  assign RIOI3_X105Y173_OLOGIC_X1Y174_D1 = CLBLM_R_X5Y159_SLICE_X6Y159_AO6;
  assign LIOI3_X0Y189_OLOGIC_X0Y189_T1 = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_D1 = CLBLM_L_X8Y150_SLICE_X11Y150_B5Q;
  assign RIOB33_X105Y181_IOB_X1Y182_O = CLBLM_R_X7Y153_SLICE_X8Y153_DO6;
  assign RIOB33_X105Y181_IOB_X1Y181_O = CLBLM_R_X7Y155_SLICE_X9Y155_AO6;
  assign RIOI3_X105Y173_OLOGIC_X1Y174_T1 = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_T1 = 1'b1;
  assign RIOI3_X105Y173_OLOGIC_X1Y173_D1 = CLBLM_R_X5Y151_SLICE_X6Y151_CQ;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_D1 = CLBLL_L_X4Y142_SLICE_X4Y142_BO5;
  assign RIOI3_X105Y173_OLOGIC_X1Y173_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_D1 = CLBLM_R_X11Y151_SLICE_X15Y151_A5Q;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_D1 = CLBLL_L_X2Y75_SLICE_X0Y75_AO6;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_D1 = CLBLM_L_X10Y149_SLICE_X12Y149_BQ;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_T1 = 1'b1;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_C6 = 1'b1;
  assign RIOI3_X105Y111_ILOGIC_X1Y112_D = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_A1 = 1'b1;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_A2 = CLBLM_R_X5Y150_SLICE_X6Y150_BQ;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_A3 = CLBLM_R_X5Y144_SLICE_X6Y144_C5Q;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_A4 = 1'b1;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_A6 = 1'b1;
  assign RIOI3_X105Y111_ILOGIC_X1Y111_D = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_B1 = CLBLM_R_X3Y144_SLICE_X3Y144_AQ;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_B2 = CLBLM_R_X3Y150_SLICE_X3Y150_BQ;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_B3 = CLBLM_R_X3Y147_SLICE_X2Y147_AQ;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_B4 = CLBLM_R_X3Y147_SLICE_X2Y147_BQ;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_B5 = CLBLM_R_X3Y147_SLICE_X3Y147_A5Q;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_B6 = 1'b1;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_C1 = CLBLL_L_X4Y147_SLICE_X4Y147_BQ;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_C2 = CLBLM_R_X3Y147_SLICE_X3Y147_AQ;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_C3 = CLBLM_R_X3Y146_SLICE_X3Y146_AQ;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_C4 = CLBLM_R_X3Y146_SLICE_X3Y146_CQ;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_C5 = CLBLL_L_X4Y148_SLICE_X4Y148_CO6;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_C6 = 1'b1;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_D5 = 1'b1;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_D1 = CLBLM_R_X7Y147_SLICE_X9Y147_AQ;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_D2 = CLBLM_L_X8Y149_SLICE_X11Y149_BQ;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_D3 = CLBLL_L_X4Y147_SLICE_X5Y147_CQ;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_D4 = CLBLM_R_X7Y142_SLICE_X8Y142_DO6;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_D5 = CLBLL_L_X2Y148_SLICE_X0Y148_A5Q;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_D6 = CLBLL_L_X4Y143_SLICE_X5Y143_AQ;
  assign CLBLM_R_X3Y148_SLICE_X3Y148_SR = CLBLM_R_X3Y146_SLICE_X2Y146_DO6;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_A1 = CLBLM_R_X3Y148_SLICE_X3Y148_CO6;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_A3 = CLBLM_R_X3Y148_SLICE_X2Y148_AQ;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_A4 = 1'b1;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_A5 = CLBLL_L_X2Y149_SLICE_X1Y149_DQ;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_A6 = CLBLM_R_X3Y146_SLICE_X3Y146_CQ;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_D6 = 1'b1;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_B2 = CLBLL_L_X4Y152_SLICE_X4Y152_CQ;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_B3 = CLBLM_R_X3Y147_SLICE_X3Y147_A5Q;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_B4 = CLBLM_R_X3Y149_SLICE_X2Y149_A5Q;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_B5 = CLBLM_R_X3Y142_SLICE_X2Y142_B5Q;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_B6 = 1'b1;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_C1 = CLBLM_R_X3Y150_SLICE_X3Y150_AQ;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_C2 = CLBLM_R_X3Y148_SLICE_X2Y148_AQ;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_C3 = 1'b1;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_C4 = CLBLM_R_X11Y146_SLICE_X14Y146_BO6;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_C5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_C6 = 1'b1;
  assign RIOB33_X105Y183_IOB_X1Y183_O = 1'b0;
  assign RIOB33_X105Y183_IOB_X1Y184_O = CLBLL_L_X4Y154_SLICE_X5Y154_AO6;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_D1 = CLBLM_R_X3Y144_SLICE_X3Y144_D5Q;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_D2 = CLBLL_L_X4Y147_SLICE_X4Y147_BQ;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_D3 = 1'b1;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_D4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_D5 = CLBLM_R_X5Y144_SLICE_X6Y144_DQ;
  assign CLBLM_R_X3Y148_SLICE_X2Y148_D6 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_A1 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_A2 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_A3 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_A4 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_A5 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_A6 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_B1 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_B2 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_B3 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_B4 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_B5 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_B6 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_C1 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_C2 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_C3 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_C4 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_C5 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_C6 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_D1 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_D2 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_D3 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_D4 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_D5 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_D6 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_A1 = CLBLM_L_X8Y144_SLICE_X11Y144_A5Q;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_A2 = CLBLM_R_X11Y146_SLICE_X14Y146_AQ;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_A3 = CLBLM_R_X7Y146_SLICE_X9Y146_B5Q;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_A4 = CLBLM_R_X7Y144_SLICE_X8Y144_AQ;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_A5 = CLBLM_R_X5Y142_SLICE_X7Y142_C5Q;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_A6 = CLBLM_L_X8Y144_SLICE_X10Y144_B5Q;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_B1 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_B2 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_B3 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_B4 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_B5 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_B6 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_C1 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_C2 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_C3 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_C4 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_C5 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_C6 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_D1 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_D2 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_D3 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_D4 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_D5 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_D6 = 1'b1;
  assign CLBLM_R_X5Y159_SLICE_X7Y159_A1 = 1'b1;
  assign CLBLM_R_X5Y159_SLICE_X7Y159_A2 = 1'b1;
  assign CLBLM_R_X5Y159_SLICE_X7Y159_A3 = 1'b1;
  assign CLBLM_R_X5Y159_SLICE_X7Y159_A4 = 1'b1;
  assign CLBLM_R_X5Y159_SLICE_X7Y159_A5 = 1'b1;
  assign CLBLM_R_X5Y159_SLICE_X7Y159_A6 = 1'b1;
  assign CLBLM_R_X5Y159_SLICE_X7Y159_B1 = 1'b1;
  assign CLBLM_R_X5Y159_SLICE_X7Y159_B2 = 1'b1;
  assign CLBLM_R_X5Y159_SLICE_X7Y159_B3 = 1'b1;
  assign CLBLM_R_X5Y159_SLICE_X7Y159_B4 = 1'b1;
  assign CLBLM_R_X5Y159_SLICE_X7Y159_B5 = 1'b1;
  assign CLBLM_R_X5Y159_SLICE_X7Y159_B6 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_A6 = CLBLM_R_X11Y145_SLICE_X15Y145_BO5;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_A1 = CLBLM_R_X3Y152_SLICE_X3Y152_DO6;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_A2 = CLBLM_R_X5Y153_SLICE_X7Y153_BO6;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_A3 = CLBLM_R_X3Y149_SLICE_X3Y149_AQ;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_A4 = CLBLL_L_X4Y147_SLICE_X4Y147_AQ;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_A6 = 1'b1;
  assign CLBLM_R_X5Y159_SLICE_X7Y159_C1 = 1'b1;
  assign CLBLM_R_X5Y159_SLICE_X7Y159_C2 = 1'b1;
  assign CLBLM_R_X5Y159_SLICE_X7Y159_C3 = 1'b1;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_B1 = CLBLM_R_X5Y144_SLICE_X6Y144_CQ;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_B2 = CLBLM_R_X3Y149_SLICE_X3Y149_BQ;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_B3 = CLBLM_R_X3Y148_SLICE_X3Y148_AQ;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_B4 = CLBLM_R_X5Y148_SLICE_X7Y148_AQ;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_B5 = CLBLM_R_X3Y147_SLICE_X3Y147_BQ;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_B6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y159_SLICE_X7Y159_D1 = 1'b1;
  assign CLBLM_R_X5Y159_SLICE_X7Y159_D2 = 1'b1;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_C2 = CLBLL_L_X4Y147_SLICE_X5Y147_B5Q;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_C3 = CLBLM_R_X7Y150_SLICE_X9Y150_CQ;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_C4 = CLBLM_L_X8Y146_SLICE_X10Y146_AQ;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_C5 = CLBLM_R_X3Y149_SLICE_X3Y149_CQ;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_C6 = CLBLM_R_X3Y149_SLICE_X3Y149_AQ;
  assign CLBLM_R_X5Y159_SLICE_X7Y159_D4 = 1'b1;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y159_SLICE_X6Y159_A1 = CLBLM_R_X7Y145_SLICE_X9Y145_DQ;
  assign CLBLM_R_X5Y159_SLICE_X6Y159_A2 = 1'b1;
  assign CLBLM_R_X5Y159_SLICE_X6Y159_A3 = 1'b1;
  assign CLBLM_R_X5Y159_SLICE_X6Y159_A4 = CLBLM_L_X8Y152_SLICE_X10Y152_DQ;
  assign CLBLM_R_X5Y159_SLICE_X6Y159_A5 = 1'b1;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_D1 = CLBLL_L_X4Y147_SLICE_X4Y147_AQ;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_D2 = CLBLM_R_X3Y150_SLICE_X3Y150_DO6;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_D3 = 1'b1;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_D4 = 1'b1;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_D5 = CLBLM_R_X7Y143_SLICE_X8Y143_DQ;
  assign CLBLM_R_X3Y149_SLICE_X3Y149_D6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y159_SLICE_X6Y159_A6 = 1'b1;
  assign CLBLM_R_X5Y159_SLICE_X6Y159_B1 = 1'b1;
  assign CLBLM_R_X5Y159_SLICE_X6Y159_B2 = 1'b1;
  assign CLBLM_R_X5Y159_SLICE_X6Y159_B3 = 1'b1;
  assign CLBLM_R_X5Y159_SLICE_X6Y159_B4 = 1'b1;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_A2 = CLBLM_R_X5Y150_SLICE_X6Y150_A5Q;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_A3 = CLBLM_R_X3Y149_SLICE_X2Y149_AQ;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_A4 = CLBLM_L_X8Y152_SLICE_X10Y152_DQ;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_A5 = CLBLM_R_X7Y153_SLICE_X9Y153_A5Q;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_A6 = 1'b1;
  assign CLBLM_R_X5Y159_SLICE_X6Y159_C1 = 1'b1;
  assign CLBLM_R_X5Y159_SLICE_X6Y159_C2 = 1'b1;
  assign CLBLM_R_X5Y159_SLICE_X6Y159_C3 = 1'b1;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_B1 = CLBLL_L_X2Y149_SLICE_X1Y149_CQ;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_B2 = CLBLM_R_X7Y150_SLICE_X8Y150_D5Q;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_B4 = 1'b1;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_B5 = CLBLL_L_X2Y149_SLICE_X1Y149_BQ;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_B6 = CLBLL_L_X2Y149_SLICE_X1Y149_DQ;
  assign CLBLM_R_X5Y159_SLICE_X6Y159_D1 = 1'b1;
  assign CLBLM_R_X5Y159_SLICE_X6Y159_D2 = 1'b1;
  assign CLBLM_R_X5Y159_SLICE_X6Y159_D3 = 1'b1;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_C2 = CLBLM_R_X3Y147_SLICE_X3Y147_B5Q;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_C3 = CLBLL_L_X2Y149_SLICE_X1Y149_BQ;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_C4 = CLBLL_L_X2Y149_SLICE_X1Y149_DQ;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_C5 = CLBLL_L_X2Y149_SLICE_X1Y149_CQ;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_C6 = 1'b1;
  assign CLBLM_R_X5Y159_SLICE_X6Y159_D4 = 1'b1;
  assign CLBLM_R_X5Y159_SLICE_X6Y159_D5 = 1'b1;
  assign CLBLM_R_X5Y159_SLICE_X6Y159_D6 = 1'b1;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_D1 = 1'b1;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_D2 = 1'b1;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_D3 = CLBLM_R_X5Y149_SLICE_X6Y149_A5Q;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_D4 = CLBLM_R_X5Y151_SLICE_X6Y151_B5Q;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_D5 = 1'b1;
  assign CLBLM_R_X3Y149_SLICE_X2Y149_D6 = 1'b1;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_A1 = 1'b1;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_A2 = 1'b1;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_A3 = 1'b1;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_A4 = 1'b1;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_A5 = 1'b1;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_A6 = 1'b1;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_B1 = 1'b1;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_B2 = 1'b1;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_B3 = 1'b1;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_B4 = 1'b1;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_B5 = 1'b1;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_B6 = 1'b1;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_C1 = 1'b1;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_C2 = 1'b1;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_C3 = 1'b1;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_C4 = 1'b1;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_C5 = 1'b1;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_C6 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_CE = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_D1 = 1'b1;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_D2 = 1'b1;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_D3 = 1'b1;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_D4 = 1'b1;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_D5 = 1'b1;
  assign CLBLM_L_X12Y144_SLICE_X17Y144_D6 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_A1 = CLBLM_R_X11Y142_SLICE_X14Y142_DO6;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_A2 = RIOB33_X105Y143_IOB_X1Y144_I;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_A3 = CLBLM_R_X11Y149_SLICE_X14Y149_AQ;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_A4 = CLBLM_L_X8Y150_SLICE_X10Y150_A5Q;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_A5 = CLBLM_R_X11Y148_SLICE_X14Y148_DQ;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_A6 = 1'b1;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_B1 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_B2 = CLBLM_L_X12Y145_SLICE_X17Y145_BO6;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_B3 = CLBLM_L_X12Y145_SLICE_X17Y145_AO6;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_B4 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_B5 = CLBLM_R_X7Y149_SLICE_X9Y149_BQ;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_B6 = CLBLM_R_X11Y144_SLICE_X14Y144_AQ;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_C1 = CLBLM_L_X12Y144_SLICE_X16Y144_AO6;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_C2 = CLBLM_L_X12Y145_SLICE_X16Y145_BO6;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_C3 = CLBLM_R_X11Y145_SLICE_X15Y145_BO5;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_C4 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_C5 = CLBLM_R_X11Y144_SLICE_X15Y144_AO5;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_C6 = CLBLM_R_X11Y143_SLICE_X15Y143_DO6;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_A6 = 1'b1;
  assign LIOI3_X0Y191_OLOGIC_X0Y192_D1 = CLBLL_L_X4Y154_SLICE_X4Y154_AO5;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_D1 = CLBLM_L_X12Y146_SLICE_X16Y146_AO6;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_D2 = CLBLM_L_X12Y144_SLICE_X16Y144_AO6;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_D3 = CLBLM_R_X11Y144_SLICE_X15Y144_AO5;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_D4 = CLBLM_R_X11Y145_SLICE_X15Y145_BO5;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_D5 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_L_X12Y144_SLICE_X16Y144_D6 = CLBLM_R_X11Y143_SLICE_X15Y143_DO6;
  assign LIOI3_X0Y191_OLOGIC_X0Y192_T1 = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_D1 = CLBLM_R_X3Y149_SLICE_X2Y149_BQ;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_D3 = 1'b1;
  assign LIOI3_X0Y191_OLOGIC_X0Y191_D1 = CLBLL_L_X4Y145_SLICE_X4Y145_BO6;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_T1 = 1'b1;
  assign RIOI3_X105Y175_OLOGIC_X1Y176_D1 = CLBLL_L_X2Y151_SLICE_X1Y151_CO6;
  assign LIOI3_X0Y191_OLOGIC_X0Y191_T1 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_B3 = CLBLM_R_X5Y145_SLICE_X7Y145_BO6;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_D1 = CLBLM_R_X3Y149_SLICE_X2Y149_CQ;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_B4 = CLBLM_R_X7Y148_SLICE_X8Y148_BO6;
  assign RIOI3_X105Y175_OLOGIC_X1Y176_T1 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_B5 = CLBLM_R_X7Y146_SLICE_X8Y146_CO6;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_D4 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_B6 = CLBLL_L_X4Y142_SLICE_X5Y142_DO6;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_T1 = 1'b1;
  assign RIOI3_X105Y175_OLOGIC_X1Y175_D1 = CLBLM_R_X3Y153_SLICE_X3Y153_CO6;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_D1 = CLBLM_R_X3Y144_SLICE_X2Y144_CO6;
  assign RIOI3_X105Y175_OLOGIC_X1Y175_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_T1 = 1'b1;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_D5 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_D1 = CLBLM_R_X7Y153_SLICE_X8Y153_DO6;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_D1 = CLBLL_L_X2Y150_SLICE_X1Y150_DO5;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_D1 = CLBLM_R_X103Y178_SLICE_X163Y178_AO6;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_D6 = 1'b1;
  assign LIOB33_X0Y101_IOB_X0Y102_O = CLBLM_R_X5Y140_SLICE_X7Y140_BQ;
  assign LIOB33_X0Y101_IOB_X0Y101_O = CLBLM_R_X3Y142_SLICE_X2Y142_B5Q;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_T1 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_A1 = CLBLL_L_X4Y150_SLICE_X4Y150_CO6;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_A2 = 1'b1;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_A3 = CLBLM_R_X3Y150_SLICE_X3Y150_CQ;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_A4 = CLBLL_L_X4Y149_SLICE_X4Y149_BQ;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_A5 = 1'b1;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign RIOB33_X105Y167_IOB_X1Y168_O = CLBLM_L_X8Y150_SLICE_X11Y150_CQ;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_B1 = CLBLL_L_X4Y150_SLICE_X4Y150_CO6;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_B2 = CLBLM_R_X3Y152_SLICE_X2Y152_BQ;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_B3 = CLBLM_R_X3Y150_SLICE_X3Y150_CQ;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_B4 = CLBLM_L_X10Y148_SLICE_X12Y148_AQ;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_B5 = CLBLM_R_X3Y152_SLICE_X2Y152_AQ;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_B6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign RIOB33_X105Y187_IOB_X1Y187_O = CLBLM_R_X103Y178_SLICE_X163Y178_AO6;
  assign RIOB33_X105Y187_IOB_X1Y188_O = CLBLM_R_X7Y153_SLICE_X8Y153_DO6;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_C1 = CLBLM_R_X5Y148_SLICE_X6Y148_BQ;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_C2 = CLBLM_R_X7Y152_SLICE_X8Y152_BQ;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_C3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_C4 = CLBLM_R_X7Y144_SLICE_X9Y144_AQ;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_C5 = 1'b1;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_C6 = CLBLL_L_X4Y150_SLICE_X4Y150_AO5;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign RIOB33_X105Y167_IOB_X1Y167_O = CLBLM_L_X8Y152_SLICE_X10Y152_DQ;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_D1 = CLBLM_R_X3Y152_SLICE_X2Y152_AQ;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_D2 = CLBLM_R_X3Y150_SLICE_X3Y150_CQ;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_D3 = 1'b1;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_D4 = CLBLL_L_X4Y150_SLICE_X4Y150_CO6;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_D5 = 1'b1;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_D6 = CLBLM_R_X3Y152_SLICE_X2Y152_BQ;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_A1 = CLBLM_L_X8Y153_SLICE_X11Y153_BQ;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_A2 = CLBLM_R_X3Y150_SLICE_X2Y150_BQ;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_A3 = CLBLM_R_X11Y150_SLICE_X14Y150_CO6;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_A4 = CLBLM_L_X8Y148_SLICE_X10Y148_DO6;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_A5 = 1'b1;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_B1 = CLBLM_R_X5Y152_SLICE_X6Y152_CQ;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_B2 = CLBLL_L_X4Y154_SLICE_X4Y154_AQ;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_B3 = CLBLM_R_X3Y150_SLICE_X2Y150_AQ;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_B5 = CLBLM_R_X3Y148_SLICE_X3Y148_AQ;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_B6 = 1'b1;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_C1 = CLBLM_R_X3Y150_SLICE_X2Y150_BQ;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_C2 = CLBLL_L_X4Y153_SLICE_X4Y153_A5Q;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_C3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_C4 = CLBLL_L_X2Y150_SLICE_X1Y150_BO5;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_C5 = CLBLL_L_X2Y150_SLICE_X1Y150_CQ;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_C6 = 1'b1;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_D1 = CLBLM_R_X5Y150_SLICE_X7Y150_BO6;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_D2 = 1'b1;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_D3 = CLBLM_R_X3Y150_SLICE_X2Y150_DQ;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_D4 = CLBLM_R_X3Y144_SLICE_X3Y144_A5Q;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_D5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_D6 = CLBLM_R_X3Y152_SLICE_X2Y152_BQ;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_A1 = 1'b1;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_A2 = CLBLM_R_X13Y145_SLICE_X18Y145_AO6;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_A3 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_A4 = CLBLM_R_X11Y145_SLICE_X14Y145_CQ;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_A5 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_A6 = CLBLM_R_X11Y145_SLICE_X14Y145_DQ;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_B1 = CLBLM_R_X11Y146_SLICE_X15Y146_BO5;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_B2 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_B3 = CLBLM_L_X10Y145_SLICE_X12Y145_AQ;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_B4 = CLBLM_R_X11Y145_SLICE_X15Y145_AQ;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_B5 = 1'b1;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_B6 = RIOB33_X105Y137_IOB_X1Y138_I;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_B5 = CLBLM_R_X7Y153_SLICE_X9Y153_BQ;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_C1 = CLBLM_R_X11Y145_SLICE_X15Y145_BO5;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_C2 = 1'b1;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_C3 = 1'b1;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_C4 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_C5 = CLBLM_L_X12Y145_SLICE_X16Y145_AO6;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_C6 = CLBLM_R_X7Y145_SLICE_X9Y145_BQ;
  assign RIOI3_X105Y115_ILOGIC_X1Y116_D = RIOB33_X105Y115_IOB_X1Y116_I;
  assign RIOI3_X105Y115_ILOGIC_X1Y115_D = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_D1 = 1'b1;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_D2 = 1'b1;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_D3 = 1'b1;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_D4 = 1'b1;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_D5 = 1'b1;
  assign CLBLM_L_X12Y145_SLICE_X17Y145_D6 = 1'b1;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_B6 = CLBLM_R_X5Y149_SLICE_X7Y149_DQ;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_A1 = CLBLM_R_X11Y145_SLICE_X14Y145_DQ;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_A2 = CLBLM_L_X8Y150_SLICE_X10Y150_A5Q;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_A3 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_A4 = CLBLM_R_X11Y142_SLICE_X14Y142_DO6;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_A5 = CLBLM_R_X11Y149_SLICE_X14Y149_AQ;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_A6 = 1'b1;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_B1 = CLBLM_R_X11Y149_SLICE_X14Y149_AQ;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_B2 = CLBLM_R_X11Y145_SLICE_X14Y145_CQ;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_B3 = CLBLM_R_X11Y142_SLICE_X14Y142_BO6;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_B4 = CLBLM_L_X8Y150_SLICE_X10Y150_A5Q;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_B5 = CLBLM_L_X10Y147_SLICE_X12Y147_AQ;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_B6 = CLBLM_R_X11Y142_SLICE_X14Y142_DO6;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_C1 = CLBLM_R_X11Y142_SLICE_X14Y142_BO6;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_C2 = CLBLM_R_X7Y146_SLICE_X9Y146_B5Q;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_C3 = CLBLM_R_X11Y149_SLICE_X14Y149_AQ;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_C4 = CLBLL_L_X4Y144_SLICE_X5Y144_BQ;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_C5 = CLBLM_L_X10Y147_SLICE_X13Y147_AQ;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_C6 = CLBLM_L_X8Y150_SLICE_X10Y150_A5Q;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_A1 = CLBLM_L_X10Y153_SLICE_X12Y153_DO6;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_D1 = CLBLM_R_X11Y145_SLICE_X15Y145_BO5;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_D2 = CLBLM_L_X12Y145_SLICE_X16Y145_AO6;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_D3 = RIOB33_X105Y137_IOB_X1Y138_I;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_D4 = CLBLM_R_X3Y145_SLICE_X3Y145_DQ;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_D5 = 1'b1;
  assign CLBLM_L_X12Y145_SLICE_X16Y145_D6 = 1'b1;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_A2 = CLBLM_L_X8Y149_SLICE_X11Y149_B5Q;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_A3 = CLBLM_R_X11Y151_SLICE_X14Y151_AQ;
  assign LIOB33_X0Y141_IOB_X0Y142_O = CLBLM_R_X3Y149_SLICE_X2Y149_CQ;
  assign LIOB33_X0Y141_IOB_X0Y141_O = CLBLL_L_X2Y150_SLICE_X1Y150_C5Q;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_A4 = CLBLM_L_X10Y151_SLICE_X12Y151_DO6;
  assign LIOB33_X0Y103_IOB_X0Y104_O = CLBLM_R_X7Y144_SLICE_X9Y144_C5Q;
  assign LIOB33_X0Y103_IOB_X0Y103_O = CLBLL_L_X4Y150_SLICE_X5Y150_DQ;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_C1 = CLBLM_R_X5Y152_SLICE_X6Y152_C5Q;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_A5 = CLBLM_L_X10Y152_SLICE_X13Y152_CO5;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_C2 = CLBLM_L_X8Y149_SLICE_X10Y149_BQ;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign RIOB33_X105Y189_IOB_X1Y190_O = CLBLM_R_X11Y153_SLICE_X14Y153_AO6;
  assign RIOB33_X105Y189_IOB_X1Y189_O = CLBLM_R_X103Y178_SLICE_X163Y178_AO6;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_A1 = CLBLL_L_X4Y151_SLICE_X4Y151_BO5;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_A2 = CLBLM_R_X5Y148_SLICE_X6Y148_B5Q;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_A3 = CLBLM_R_X3Y151_SLICE_X3Y151_AQ;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_A5 = CLBLL_L_X2Y148_SLICE_X0Y148_B5Q;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_A6 = CLBLM_R_X3Y150_SLICE_X3Y150_AQ;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_B1 = CLBLL_L_X4Y151_SLICE_X4Y151_BO6;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_B2 = CLBLM_R_X3Y151_SLICE_X3Y151_BQ;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_B3 = CLBLL_L_X2Y148_SLICE_X0Y148_B5Q;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_B4 = CLBLL_L_X4Y143_SLICE_X5Y143_AQ;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_B5 = CLBLM_R_X3Y150_SLICE_X3Y150_AQ;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_B6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_C2 = CLBLM_R_X7Y144_SLICE_X9Y144_AQ;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_C3 = CLBLM_R_X5Y145_SLICE_X6Y145_B5Q;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_C4 = CLBLM_R_X7Y153_SLICE_X8Y153_DO5;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_C5 = CLBLL_L_X4Y154_SLICE_X4Y154_AQ;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_C6 = 1'b1;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_D1 = CLBLM_R_X3Y147_SLICE_X3Y147_BQ;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_D2 = CLBLL_L_X4Y147_SLICE_X5Y147_B5Q;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_D3 = CLBLM_R_X3Y151_SLICE_X2Y151_DO6;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_D4 = CLBLM_L_X12Y149_SLICE_X16Y149_CO6;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_D5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_D6 = 1'b1;
  assign RIOI3_X105Y153_OLOGIC_X1Y153_T1 = 1'b1;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_A1 = 1'b1;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_A2 = CLBLM_R_X5Y150_SLICE_X6Y150_A5Q;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_A3 = CLBLM_R_X3Y151_SLICE_X2Y151_AQ;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_A4 = CLBLL_L_X2Y151_SLICE_X1Y151_AQ;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_A6 = CLBLM_R_X3Y151_SLICE_X2Y151_CO6;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_AX = CLBLM_R_X3Y151_SLICE_X2Y151_CO5;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_B1 = CLBLM_R_X3Y143_SLICE_X2Y143_AQ;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_B2 = CLBLL_L_X4Y149_SLICE_X5Y149_CQ;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_B3 = CLBLM_R_X3Y145_SLICE_X2Y145_DQ;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_B4 = CLBLM_R_X7Y152_SLICE_X9Y152_BQ;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_B5 = CLBLM_R_X3Y148_SLICE_X2Y148_C5Q;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_B6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_C1 = CLBLM_R_X7Y152_SLICE_X8Y152_AQ;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_C2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_C3 = CLBLM_R_X3Y147_SLICE_X3Y147_B5Q;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_C4 = CLBLM_R_X3Y151_SLICE_X2Y151_A5Q;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_C5 = CLBLM_R_X3Y151_SLICE_X3Y151_DQ;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_C6 = 1'b1;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_D1 = LIOB33_X0Y55_IOB_X0Y55_I;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_D2 = CLBLM_R_X3Y151_SLICE_X2Y151_AQ;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_D3 = CLBLM_R_X3Y147_SLICE_X3Y147_B5Q;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_D4 = CLBLM_R_X3Y151_SLICE_X2Y151_A5Q;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_D5 = CLBLM_R_X3Y151_SLICE_X3Y151_DQ;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_D6 = CLBLL_L_X2Y151_SLICE_X1Y151_AQ;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_A1 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_A2 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_A3 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_A4 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_A5 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_A6 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_B1 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_B2 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_B3 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_B4 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_B5 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_B6 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_C1 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_C2 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_C3 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_C4 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_C5 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_C6 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_D1 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_D2 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_D3 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_D4 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_D5 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_D6 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_A1 = CLBLM_R_X11Y149_SLICE_X14Y149_AQ;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_A2 = CLBLM_R_X11Y148_SLICE_X14Y148_BQ;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_A3 = CLBLM_R_X11Y142_SLICE_X14Y142_BO6;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_A4 = CLBLM_L_X12Y149_SLICE_X16Y149_BQ;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_A5 = CLBLM_L_X8Y150_SLICE_X10Y150_A5Q;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_A6 = CLBLM_R_X11Y142_SLICE_X14Y142_DO6;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_B1 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_B2 = CLBLM_R_X7Y149_SLICE_X9Y149_BQ;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_B3 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_B4 = CLBLM_R_X11Y146_SLICE_X15Y146_CO5;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_B5 = CLBLM_R_X11Y142_SLICE_X14Y142_CO5;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_B6 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_C1 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_C2 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_C3 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_C4 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_C5 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_C6 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_D1 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_D2 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_D3 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_D4 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_D5 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_D6 = 1'b1;
  assign LIOB33_X0Y105_IOB_X0Y106_O = CLBLL_L_X4Y147_SLICE_X5Y147_DQ;
  assign LIOB33_X0Y105_IOB_X0Y105_O = CLBLM_R_X5Y144_SLICE_X6Y144_B5Q;
  assign CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_CE = 1'b1;
  assign RIOB33_X105Y191_IOB_X1Y192_O = CLBLM_L_X12Y151_SLICE_X16Y151_CO6;
  assign RIOB33_X105Y191_IOB_X1Y191_O = CLBLM_R_X11Y149_SLICE_X14Y149_AO6;
  assign LIOI3_X0Y195_OLOGIC_X0Y196_D1 = CLBLL_L_X4Y154_SLICE_X5Y154_AO6;
  assign LIOI3_X0Y195_OLOGIC_X0Y196_T1 = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_D1 = CLBLM_R_X3Y149_SLICE_X2Y149_BQ;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_A1 = CLBLL_L_X4Y149_SLICE_X4Y149_B5Q;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_A2 = CLBLL_L_X2Y150_SLICE_X1Y150_A5Q;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_A3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_A4 = CLBLL_L_X4Y145_SLICE_X5Y145_BQ;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_A5 = CLBLM_R_X3Y152_SLICE_X3Y152_CO6;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_A6 = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_T1 = 1'b1;
  assign LIOI3_X0Y195_OLOGIC_X0Y195_D1 = CLBLL_L_X2Y152_SLICE_X1Y152_AO6;
  assign RIOI3_X105Y177_OLOGIC_X1Y178_D1 = CLBLM_R_X3Y150_SLICE_X3Y150_BQ;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_B1 = CLBLM_R_X5Y153_SLICE_X7Y153_BO6;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_B2 = CLBLM_R_X3Y148_SLICE_X3Y148_BO5;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_B3 = CLBLL_L_X4Y150_SLICE_X5Y150_D5Q;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_B4 = CLBLM_R_X3Y150_SLICE_X3Y150_BQ;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_B5 = CLBLM_R_X3Y153_SLICE_X3Y153_AQ;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_B6 = CLBLM_R_X3Y153_SLICE_X3Y153_BQ;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_D1 = CLBLM_R_X3Y142_SLICE_X2Y142_CO5;
  assign LIOI3_X0Y195_OLOGIC_X0Y195_T1 = 1'b1;
  assign RIOI3_X105Y177_OLOGIC_X1Y178_T1 = 1'b1;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_C1 = CLBLM_R_X3Y150_SLICE_X3Y150_AQ;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_C2 = CLBLM_R_X7Y144_SLICE_X9Y144_AQ;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_C3 = CLBLM_R_X7Y152_SLICE_X8Y152_BQ;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_C4 = CLBLM_R_X3Y152_SLICE_X3Y152_AQ;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_C5 = CLBLL_L_X2Y148_SLICE_X0Y148_B5Q;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_C6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_T1 = 1'b1;
  assign RIOI3_X105Y177_OLOGIC_X1Y177_D1 = CLBLM_L_X10Y142_SLICE_X12Y142_AQ;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_D1 = CLBLM_R_X3Y153_SLICE_X3Y153_AQ;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_D2 = CLBLM_R_X3Y148_SLICE_X3Y148_BO5;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_D3 = CLBLM_R_X3Y153_SLICE_X3Y153_BQ;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_D4 = CLBLL_L_X4Y150_SLICE_X5Y150_D5Q;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_D5 = 1'b1;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_D6 = CLBLM_R_X3Y150_SLICE_X3Y150_BQ;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_D1 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign RIOI3_X105Y177_OLOGIC_X1Y177_T1 = 1'b1;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_A1 = CLBLM_R_X7Y152_SLICE_X8Y152_BQ;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_A2 = CLBLL_L_X4Y152_SLICE_X4Y152_DQ;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_A3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_A4 = CLBLL_L_X4Y150_SLICE_X4Y150_AO5;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_A5 = 1'b1;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_A6 = CLBLM_R_X7Y144_SLICE_X9Y144_AQ;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_T1 = 1'b1;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_B1 = CLBLM_R_X5Y152_SLICE_X7Y152_DQ;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_B2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_B3 = CLBLM_R_X3Y152_SLICE_X2Y152_AQ;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_B4 = CLBLL_L_X4Y150_SLICE_X4Y150_CO6;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_B5 = 1'b1;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_B6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_D1 = CLBLM_R_X7Y153_SLICE_X9Y153_CQ;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_C1 = CLBLM_R_X3Y148_SLICE_X2Y148_D5Q;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_C2 = CLBLM_R_X3Y152_SLICE_X2Y152_CQ;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_C3 = CLBLM_R_X7Y152_SLICE_X8Y152_BQ;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_C5 = CLBLM_R_X5Y144_SLICE_X6Y144_DQ;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_C6 = CLBLL_L_X2Y144_SLICE_X1Y144_B5Q;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_T1 = 1'b1;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_D1 = CLBLM_R_X5Y151_SLICE_X7Y151_BO6;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_D2 = CLBLL_L_X4Y150_SLICE_X4Y150_AO5;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_D3 = CLBLM_R_X7Y152_SLICE_X8Y152_BQ;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_D4 = CLBLL_L_X4Y150_SLICE_X5Y150_CQ;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_D5 = 1'b1;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_D6 = CLBLM_R_X7Y144_SLICE_X9Y144_AQ;
  assign LIOB33_X0Y107_IOB_X0Y108_O = CLBLL_L_X4Y143_SLICE_X5Y143_C5Q;
  assign LIOB33_X0Y107_IOB_X0Y107_O = CLBLM_R_X3Y145_SLICE_X2Y145_C5Q;
  assign RIOI3_X105Y117_ILOGIC_X1Y118_D = RIOB33_X105Y117_IOB_X1Y118_I;
  assign RIOI3_X105Y117_ILOGIC_X1Y117_D = RIOB33_X105Y117_IOB_X1Y117_I;
  assign RIOB33_X105Y193_IOB_X1Y194_O = CLBLM_L_X12Y151_SLICE_X16Y151_CO5;
  assign RIOB33_X105Y193_IOB_X1Y193_O = CLBLM_R_X11Y153_SLICE_X14Y153_AO5;
  assign CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_I = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLM_R_X5Y159_SLICE_X7Y159_C4 = 1'b1;
  assign CLBLM_R_X5Y159_SLICE_X7Y159_C5 = 1'b1;
  assign CLBLM_R_X5Y159_SLICE_X7Y159_C6 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_A2 = CLBLM_R_X3Y148_SLICE_X3Y148_BO6;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_A3 = CLBLM_R_X3Y153_SLICE_X3Y153_AQ;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_A4 = CLBLM_R_X5Y153_SLICE_X7Y153_BO6;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_A5 = CLBLM_R_X3Y153_SLICE_X3Y153_BQ;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_A6 = CLBLM_L_X8Y151_SLICE_X10Y151_BQ;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_AX = CLBLM_R_X3Y153_SLICE_X3Y153_BO6;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_B1 = CLBLM_R_X3Y143_SLICE_X2Y143_AQ;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_B2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_B4 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_B5 = CLBLM_R_X3Y150_SLICE_X2Y150_CO5;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_B6 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_BX = CLBLM_R_X3Y153_SLICE_X3Y153_CO5;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_C1 = CLBLM_R_X3Y153_SLICE_X3Y153_BQ;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_C2 = CLBLM_R_X3Y148_SLICE_X3Y148_BO6;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_C3 = CLBLM_R_X5Y153_SLICE_X7Y153_BO6;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_C5 = CLBLL_L_X4Y153_SLICE_X5Y153_AQ;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_C6 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_CX = CLBLM_R_X7Y153_SLICE_X8Y153_BO5;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_D1 = CLBLM_R_X3Y153_SLICE_X3Y153_BQ;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_D2 = CLBLM_R_X3Y148_SLICE_X3Y148_BO5;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_D3 = CLBLM_R_X3Y150_SLICE_X3Y150_BQ;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_D4 = CLBLM_R_X3Y149_SLICE_X3Y149_AQ;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_D5 = CLBLM_R_X3Y153_SLICE_X3Y153_AQ;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_D6 = CLBLL_L_X4Y150_SLICE_X5Y150_D5Q;
  assign LIOI3_X0Y155_OLOGIC_X0Y155_D1 = CLBLM_L_X8Y150_SLICE_X11Y150_CQ;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_A2 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_A3 = CLBLM_R_X3Y153_SLICE_X2Y153_AQ;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_A4 = CLBLM_R_X3Y151_SLICE_X3Y151_D5Q;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_A5 = CLBLM_R_X5Y143_SLICE_X6Y143_DQ;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_A6 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_AX = CLBLM_R_X3Y152_SLICE_X2Y152_CQ;
  assign CLBLM_R_X5Y159_SLICE_X7Y159_D3 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_B1 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_B2 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_B3 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_B4 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_B5 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_B6 = 1'b1;
  assign CLBLM_R_X5Y159_SLICE_X7Y159_D5 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_C1 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_C2 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_C3 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_C4 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_C5 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_C6 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_CE = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y159_SLICE_X7Y159_D6 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_D1 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_D2 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_D3 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_D4 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_D5 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_D6 = 1'b1;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_C4 = 1'b1;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_C5 = 1'b1;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_C6 = 1'b1;
  assign LIOB33_X0Y109_IOB_X0Y110_O = CLBLM_R_X5Y143_SLICE_X6Y143_DQ;
  assign LIOB33_X0Y109_IOB_X0Y109_O = CLBLL_L_X2Y153_SLICE_X1Y153_AQ;
  assign CLBLM_R_X5Y159_SLICE_X6Y159_B5 = 1'b1;
  assign CLBLM_R_X5Y159_SLICE_X6Y159_B6 = 1'b1;
  assign RIOB33_X105Y195_IOB_X1Y196_O = CLBLM_R_X11Y150_SLICE_X14Y150_BO6;
  assign RIOB33_X105Y195_IOB_X1Y195_O = CLBLM_R_X11Y149_SLICE_X14Y149_BO6;
  assign CLBLM_R_X5Y159_SLICE_X6Y159_C4 = 1'b1;
  assign CLBLM_R_X5Y159_SLICE_X6Y159_C5 = 1'b1;
  assign CLBLM_R_X5Y159_SLICE_X6Y159_C6 = 1'b1;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_A1 = 1'b1;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_A2 = CLBLM_R_X7Y142_SLICE_X9Y142_CQ;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_A1 = 1'b1;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_A2 = CLBLM_L_X8Y153_SLICE_X11Y153_BQ;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_A3 = CLBLM_R_X3Y154_SLICE_X3Y154_AQ;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_A4 = CLBLM_R_X3Y152_SLICE_X2Y152_BQ;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_A5 = CLBLL_L_X2Y151_SLICE_X1Y151_AQ;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_B1 = 1'b1;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_B2 = 1'b1;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_B3 = 1'b1;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_B4 = 1'b1;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_B5 = 1'b1;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_B6 = 1'b1;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_C1 = 1'b1;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_C2 = 1'b1;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_C3 = 1'b1;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_C4 = 1'b1;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_C5 = 1'b1;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_C6 = 1'b1;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_A3 = 1'b1;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_D1 = 1'b1;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_D2 = 1'b1;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_D3 = 1'b1;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_D4 = 1'b1;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_D5 = 1'b1;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_D6 = 1'b1;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_B1 = CLBLM_R_X11Y149_SLICE_X14Y149_AQ;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_B2 = CLBLM_L_X12Y143_SLICE_X16Y143_AO6;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_A1 = 1'b1;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_A2 = 1'b1;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_A3 = 1'b1;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_A4 = 1'b1;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_A5 = 1'b1;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_A6 = 1'b1;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_B3 = CLBLM_R_X7Y149_SLICE_X9Y149_C5Q;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_B1 = 1'b1;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_B2 = 1'b1;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_B3 = 1'b1;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_B4 = 1'b1;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_B5 = 1'b1;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_B6 = 1'b1;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_B6 = 1'b1;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_C1 = 1'b1;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_C2 = 1'b1;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_C3 = 1'b1;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_C4 = 1'b1;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_C5 = 1'b1;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_C6 = 1'b1;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_D1 = 1'b1;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_D2 = 1'b1;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_D3 = 1'b1;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_D4 = 1'b1;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_D5 = 1'b1;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_D6 = 1'b1;
  assign LIOI3_X0Y197_OLOGIC_X0Y198_D1 = 1'b1;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_A1 = 1'b1;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_A2 = 1'b1;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_A3 = 1'b1;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_A4 = 1'b1;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_A5 = 1'b1;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_A6 = 1'b1;
  assign LIOI3_X0Y197_OLOGIC_X0Y198_T1 = 1'b1;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_B1 = 1'b1;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_B2 = 1'b1;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_B3 = 1'b1;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_B4 = 1'b1;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_B5 = 1'b1;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_B6 = 1'b1;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_B6 = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_D1 = CLBLM_L_X8Y153_SLICE_X10Y153_AQ;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_C1 = 1'b1;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_C2 = 1'b1;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_C3 = 1'b1;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_C4 = 1'b1;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_C5 = 1'b1;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_C6 = 1'b1;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_C5 = CLBLM_R_X11Y145_SLICE_X14Y145_BO5;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_C6 = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_T1 = 1'b1;
  assign LIOI3_X0Y197_OLOGIC_X0Y197_D1 = CLBLM_R_X3Y153_SLICE_X3Y153_BO5;
  assign RIOI3_X105Y179_OLOGIC_X1Y180_D1 = CLBLM_L_X10Y150_SLICE_X12Y150_CQ;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_CE = LIOB33_X0Y61_IOB_X0Y62_I;
  assign LIOI3_X0Y197_OLOGIC_X0Y197_T1 = 1'b1;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_D1 = 1'b1;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_D2 = 1'b1;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_D3 = 1'b1;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_D4 = 1'b1;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_D5 = 1'b1;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_D6 = 1'b1;
  assign LIOB33_X0Y111_IOB_X0Y111_O = CLBLM_R_X3Y145_SLICE_X2Y145_CQ;
  assign LIOB33_X0Y111_IOB_X0Y112_O = CLBLM_R_X3Y145_SLICE_X2Y145_B5Q;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_D1 = CLBLM_R_X3Y149_SLICE_X2Y149_BQ;
  assign RIOI3_X105Y179_OLOGIC_X1Y180_T1 = 1'b1;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_A1 = CLBLM_R_X11Y148_SLICE_X14Y148_AO6;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_A2 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_A3 = CLBLM_R_X11Y149_SLICE_X15Y149_BQ;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_A4 = CLBLM_L_X10Y147_SLICE_X13Y147_AQ;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_A5 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_T1 = 1'b1;
  assign RIOI3_X105Y179_OLOGIC_X1Y179_D1 = CLBLM_R_X3Y149_SLICE_X3Y149_DQ;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_B1 = CLBLM_R_X11Y145_SLICE_X15Y145_BO5;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_B2 = CLBLM_L_X12Y149_SLICE_X16Y149_BQ;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_B3 = CLBLL_L_X4Y149_SLICE_X5Y149_DQ;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_B4 = 1'b1;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_B5 = CLBLM_L_X10Y149_SLICE_X12Y149_AQ;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_B6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_D1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign RIOI3_X105Y179_OLOGIC_X1Y179_T1 = 1'b1;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_C1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_C2 = CLBLM_L_X12Y149_SLICE_X16Y149_AQ;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_C3 = 1'b1;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_C4 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_C5 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_C6 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_T1 = 1'b1;
  assign RIOB33_X105Y197_IOB_X1Y198_O = CLBLM_R_X11Y149_SLICE_X14Y149_CO6;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOB33_X105Y197_IOB_X1Y197_O = CLBLM_R_X11Y150_SLICE_X14Y150_BO5;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_D1 = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_D1 = CLBLM_R_X11Y149_SLICE_X15Y149_BQ;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_D2 = 1'b1;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_D3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_D4 = 1'b1;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_D5 = CLBLM_R_X11Y148_SLICE_X14Y148_AO6;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_D6 = 1'b1;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_A5 = CLBLM_R_X7Y147_SLICE_X9Y147_AQ;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_T1 = 1'b1;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_B2 = CLBLM_R_X7Y147_SLICE_X8Y147_BQ;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_B3 = CLBLM_R_X5Y147_SLICE_X6Y147_DQ;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_C5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_C6 = CLBLM_R_X3Y147_SLICE_X3Y147_BQ;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_C4 = CLBLM_L_X10Y150_SLICE_X12Y150_CQ;
  assign RIOI3_X105Y121_ILOGIC_X1Y122_D = RIOB33_X105Y121_IOB_X1Y122_I;
  assign RIOI3_X105Y121_ILOGIC_X1Y121_D = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_C5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_C6 = 1'b1;
  assign LIOB33_X0Y113_IOB_X0Y114_O = CLBLL_L_X4Y153_SLICE_X4Y153_A5Q;
  assign LIOB33_X0Y113_IOB_X0Y113_O = CLBLM_R_X3Y146_SLICE_X2Y146_CQ;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign LIOB33_X0Y181_IOB_X0Y181_O = RIOB33_X105Y127_IOB_X1Y128_I;
  assign LIOB33_SING_X0Y100_IOB_X0Y100_O = CLBLM_R_X3Y149_SLICE_X2Y149_AQ;
  assign LIOI3_X0Y103_OLOGIC_X0Y104_T1 = 1'b1;
  assign LIOI3_X0Y103_OLOGIC_X0Y103_D1 = CLBLL_L_X4Y150_SLICE_X5Y150_DQ;
  assign LIOB33_X0Y115_IOB_X0Y116_O = CLBLM_R_X5Y152_SLICE_X6Y152_CQ;
  assign LIOB33_X0Y115_IOB_X0Y115_O = CLBLM_R_X3Y151_SLICE_X3Y151_CQ;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_A1 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_A2 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_A3 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_A4 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_A5 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_A6 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_B1 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_B2 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_B3 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_B4 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_B5 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_B6 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_A1 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_A2 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_C3 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_C4 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_C5 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_C6 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_A3 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_A4 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_A5 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_A6 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_B1 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_B2 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_B3 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_B4 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_B5 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_B6 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_D1 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_D5 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_D6 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_D2 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_C1 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_C2 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_C3 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_C4 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_C5 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_C6 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_A1 = CLBLM_L_X12Y151_SLICE_X16Y151_AQ;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_A3 = CLBLM_L_X10Y151_SLICE_X12Y151_DO6;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_A4 = CLBLM_L_X10Y152_SLICE_X13Y152_CO5;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_A5 = CLBLM_L_X10Y151_SLICE_X12Y151_AQ;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_A6 = CLBLM_R_X11Y151_SLICE_X14Y151_DO6;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_D1 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_D2 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_D3 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_D4 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_D5 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_D6 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_B6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_B1 = CLBLM_L_X12Y151_SLICE_X16Y151_DO6;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_B2 = CLBLM_L_X12Y151_SLICE_X16Y151_BQ;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_B3 = CLBLM_R_X11Y148_SLICE_X15Y148_AQ;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_B4 = CLBLM_L_X10Y152_SLICE_X13Y152_CO5;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_B5 = CLBLM_L_X10Y151_SLICE_X12Y151_DO6;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_A1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_A2 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_C4 = CLBLM_R_X3Y151_SLICE_X3Y151_D5Q;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_C5 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_C6 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_A3 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_A4 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_A5 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_A6 = CLBLM_R_X5Y141_SLICE_X6Y141_AQ;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_C2 = CLBLM_L_X10Y145_SLICE_X12Y145_BO6;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_B1 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_B2 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_B3 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_B4 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_B5 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_B6 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_D1 = CLBLM_R_X11Y152_SLICE_X14Y152_AQ;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_D2 = CLBLM_L_X10Y152_SLICE_X12Y152_BQ;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_C1 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_C2 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_C3 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_C4 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_C5 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_C6 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_D5 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_D6 = CLBLM_R_X11Y151_SLICE_X14Y151_DO6;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_D1 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_D2 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_D3 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_D4 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_D5 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_D6 = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_D1 = CLBLL_L_X2Y147_SLICE_X0Y147_BQ;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_T1 = 1'b1;
  assign RIOI3_X105Y183_OLOGIC_X1Y184_D1 = CLBLL_L_X4Y154_SLICE_X5Y154_AO6;
  assign CLBLM_R_X13Y145_SLICE_X19Y145_A1 = 1'b1;
  assign CLBLM_R_X13Y145_SLICE_X19Y145_A2 = 1'b1;
  assign CLBLM_R_X13Y145_SLICE_X19Y145_A3 = 1'b1;
  assign CLBLM_R_X13Y145_SLICE_X19Y145_A4 = 1'b1;
  assign CLBLM_R_X13Y145_SLICE_X19Y145_A5 = 1'b1;
  assign CLBLM_R_X13Y145_SLICE_X19Y145_A6 = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_D1 = CLBLL_L_X2Y148_SLICE_X0Y148_AQ;
  assign RIOI3_X105Y183_OLOGIC_X1Y184_T1 = 1'b1;
  assign CLBLM_R_X13Y145_SLICE_X19Y145_B1 = 1'b1;
  assign CLBLM_R_X13Y145_SLICE_X19Y145_B2 = 1'b1;
  assign CLBLM_R_X13Y145_SLICE_X19Y145_B3 = 1'b1;
  assign CLBLM_R_X13Y145_SLICE_X19Y145_B4 = 1'b1;
  assign CLBLM_R_X13Y145_SLICE_X19Y145_B5 = 1'b1;
  assign CLBLM_R_X13Y145_SLICE_X19Y145_B6 = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_T1 = 1'b1;
  assign CLBLM_R_X13Y145_SLICE_X19Y145_C1 = 1'b1;
  assign CLBLM_R_X13Y145_SLICE_X19Y145_C2 = 1'b1;
  assign CLBLM_R_X13Y145_SLICE_X19Y145_C3 = 1'b1;
  assign CLBLM_R_X13Y145_SLICE_X19Y145_C4 = 1'b1;
  assign CLBLM_R_X13Y145_SLICE_X19Y145_C5 = 1'b1;
  assign CLBLM_R_X13Y145_SLICE_X19Y145_C6 = 1'b1;
  assign LIOB33_SING_X0Y150_IOB_X0Y150_O = CLBLL_L_X4Y142_SLICE_X4Y142_DO5;
  assign RIOI3_X105Y183_OLOGIC_X1Y183_D1 = 1'b0;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_D1 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign RIOI3_X105Y183_OLOGIC_X1Y183_T1 = 1'b1;
  assign CLBLM_R_X13Y145_SLICE_X19Y145_D1 = 1'b1;
  assign CLBLM_R_X13Y145_SLICE_X19Y145_D2 = 1'b1;
  assign CLBLM_R_X13Y145_SLICE_X19Y145_D3 = 1'b1;
  assign CLBLM_R_X13Y145_SLICE_X19Y145_D4 = 1'b1;
  assign CLBLM_R_X13Y145_SLICE_X19Y145_D5 = 1'b1;
  assign CLBLM_R_X13Y145_SLICE_X19Y145_D6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_T1 = 1'b1;
  assign CLBLM_R_X13Y145_SLICE_X18Y145_A1 = CLBLM_R_X11Y148_SLICE_X14Y148_DQ;
  assign CLBLM_R_X13Y145_SLICE_X18Y145_A2 = 1'b1;
  assign CLBLM_R_X13Y145_SLICE_X18Y145_A3 = CLBLM_R_X11Y148_SLICE_X14Y148_BQ;
  assign CLBLM_R_X13Y145_SLICE_X18Y145_A4 = RIOB33_X105Y143_IOB_X1Y144_I;
  assign CLBLM_R_X13Y145_SLICE_X18Y145_A5 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_R_X13Y145_SLICE_X18Y145_A6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_D1 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLM_R_X13Y145_SLICE_X18Y145_B1 = 1'b1;
  assign CLBLM_R_X13Y145_SLICE_X18Y145_B2 = 1'b1;
  assign CLBLM_R_X13Y145_SLICE_X18Y145_B3 = 1'b1;
  assign CLBLM_R_X13Y145_SLICE_X18Y145_B4 = 1'b1;
  assign CLBLM_R_X13Y145_SLICE_X18Y145_B5 = 1'b1;
  assign CLBLM_R_X13Y145_SLICE_X18Y145_B6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_T1 = 1'b1;
  assign CLBLM_R_X13Y145_SLICE_X18Y145_C1 = 1'b1;
  assign CLBLM_R_X13Y145_SLICE_X18Y145_C2 = 1'b1;
  assign CLBLM_R_X13Y145_SLICE_X18Y145_C3 = 1'b1;
  assign CLBLM_R_X13Y145_SLICE_X18Y145_C4 = 1'b1;
  assign CLBLM_R_X13Y145_SLICE_X18Y145_C5 = 1'b1;
  assign CLBLM_R_X13Y145_SLICE_X18Y145_C6 = 1'b1;
  assign CLBLM_R_X13Y145_SLICE_X18Y145_D1 = 1'b1;
  assign CLBLM_R_X13Y145_SLICE_X18Y145_D2 = 1'b1;
  assign CLBLM_R_X13Y145_SLICE_X18Y145_D3 = 1'b1;
  assign CLBLM_R_X13Y145_SLICE_X18Y145_D4 = 1'b1;
  assign CLBLM_R_X13Y145_SLICE_X18Y145_D5 = 1'b1;
  assign CLBLM_R_X13Y145_SLICE_X18Y145_D6 = 1'b1;
  assign LIOB33_X0Y117_IOB_X0Y118_O = CLBLM_R_X11Y147_SLICE_X15Y147_AQ;
  assign LIOB33_X0Y117_IOB_X0Y117_O = CLBLM_R_X7Y144_SLICE_X9Y144_B5Q;
  assign LIOB33_SING_X0Y199_IOB_X0Y199_O = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_A1 = CLBLM_L_X8Y142_SLICE_X11Y142_CQ;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_A3 = CLBLM_L_X10Y142_SLICE_X13Y142_AQ;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_A4 = CLBLM_R_X5Y149_SLICE_X7Y149_DQ;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_A5 = CLBLM_R_X3Y144_SLICE_X2Y144_A5Q;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_A6 = CLBLM_L_X10Y147_SLICE_X13Y147_CQ;
  assign RIOI3_X105Y197_OLOGIC_X1Y197_D1 = CLBLM_R_X11Y150_SLICE_X14Y150_BO5;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_B1 = CLBLM_L_X8Y144_SLICE_X11Y144_A5Q;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_B2 = CLBLM_L_X8Y144_SLICE_X10Y144_B5Q;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_B3 = CLBLM_R_X11Y146_SLICE_X14Y146_AQ;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_B4 = CLBLM_R_X7Y144_SLICE_X8Y144_AQ;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_B5 = CLBLM_R_X5Y142_SLICE_X7Y142_C5Q;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_B6 = CLBLM_R_X7Y146_SLICE_X9Y146_B5Q;
  assign LIOI3_X0Y77_ILOGIC_X0Y78_D = LIOB33_X0Y77_IOB_X0Y78_I;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_C1 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_C2 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_C3 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_C4 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_C5 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_C6 = 1'b1;
  assign RIOI3_X105Y123_ILOGIC_X1Y124_D = RIOB33_X105Y123_IOB_X1Y124_I;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_X105Y123_ILOGIC_X1Y123_D = RIOB33_X105Y123_IOB_X1Y123_I;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_D1 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_D2 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_D3 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_D4 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_D5 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_D6 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_A1 = CLBLM_L_X8Y144_SLICE_X11Y144_A5Q;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_A2 = CLBLM_R_X7Y144_SLICE_X8Y144_AQ;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_A3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_A4 = CLBLM_L_X8Y144_SLICE_X10Y144_B5Q;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_A5 = CLBLM_R_X3Y141_SLICE_X3Y141_AO6;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_A6 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_B1 = CLBLM_L_X8Y144_SLICE_X11Y144_A5Q;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_B2 = CLBLM_R_X5Y142_SLICE_X7Y142_C5Q;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_B3 = CLBLM_R_X7Y146_SLICE_X9Y146_B5Q;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_B4 = CLBLM_R_X7Y144_SLICE_X8Y144_AQ;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_B5 = CLBLM_R_X11Y146_SLICE_X14Y146_AQ;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_B6 = CLBLM_L_X8Y144_SLICE_X10Y144_B5Q;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_C3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_C1 = CLBLM_R_X11Y146_SLICE_X14Y146_AQ;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_C2 = CLBLM_R_X7Y146_SLICE_X9Y146_B5Q;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_C3 = CLBLM_L_X8Y150_SLICE_X10Y150_A5Q;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_C4 = CLBLM_L_X10Y142_SLICE_X12Y142_AO5;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_C5 = CLBLM_R_X11Y149_SLICE_X14Y149_AQ;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_C6 = CLBLM_R_X5Y142_SLICE_X7Y142_C5Q;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_D = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_D = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_D1 = CLBLM_R_X11Y146_SLICE_X14Y146_AQ;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_D2 = CLBLM_R_X7Y144_SLICE_X8Y144_AQ;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_D3 = CLBLM_L_X8Y144_SLICE_X10Y144_B5Q;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_D4 = CLBLM_R_X7Y146_SLICE_X9Y146_B5Q;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_D5 = CLBLM_L_X8Y144_SLICE_X11Y144_A5Q;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_D6 = CLBLM_R_X5Y142_SLICE_X7Y142_C5Q;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign LIOI3_X0Y165_OLOGIC_X0Y165_T1 = 1'b1;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_D3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_D4 = CLBLM_R_X7Y154_SLICE_X8Y154_CQ;
  assign LIOB33_X0Y119_IOB_X0Y120_O = CLBLM_R_X3Y150_SLICE_X3Y150_AQ;
  assign LIOB33_X0Y119_IOB_X0Y119_O = CLBLM_R_X3Y149_SLICE_X2Y149_CQ;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_B2 = CLBLM_R_X11Y143_SLICE_X14Y143_CO6;
  assign RIOI3_X105Y141_ILOGIC_X1Y142_D = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_C1 = CLBLM_L_X8Y150_SLICE_X11Y150_AQ;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_C2 = CLBLM_L_X10Y150_SLICE_X12Y150_CQ;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_C3 = CLBLM_L_X10Y143_SLICE_X12Y143_CO6;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_B3 = CLBLM_R_X11Y149_SLICE_X14Y149_AQ;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_A1 = CLBLM_R_X5Y142_SLICE_X7Y142_C5Q;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_A2 = CLBLM_R_X7Y144_SLICE_X8Y144_AQ;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_A3 = CLBLM_L_X8Y144_SLICE_X10Y144_B5Q;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_A4 = CLBLM_R_X11Y146_SLICE_X14Y146_AQ;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_A5 = CLBLM_L_X8Y144_SLICE_X11Y144_A5Q;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_A6 = CLBLM_R_X7Y146_SLICE_X9Y146_B5Q;
  assign RIOI3_X105Y141_ILOGIC_X1Y141_D = RIOB33_X105Y141_IOB_X1Y141_I;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_B1 = CLBLM_R_X11Y142_SLICE_X14Y142_DO6;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_B2 = CLBLM_L_X8Y144_SLICE_X10Y144_CO6;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_B3 = CLBLM_R_X11Y142_SLICE_X14Y142_BO5;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_B4 = LIOB33_X0Y53_IOB_X0Y53_I;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_B5 = CLBLM_L_X10Y143_SLICE_X12Y143_AQ;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_B6 = CLBLM_R_X11Y142_SLICE_X14Y142_CO6;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_C1 = CLBLM_R_X5Y142_SLICE_X6Y142_DQ;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_C2 = LIOB33_X0Y51_IOB_X0Y52_I;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_C3 = CLBLM_R_X11Y145_SLICE_X15Y145_BO5;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_C4 = CLBLM_L_X10Y146_SLICE_X13Y146_BO6;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_C5 = CLBLM_L_X10Y146_SLICE_X13Y146_BO5;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_C6 = CLBLM_R_X11Y142_SLICE_X14Y142_CO5;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_B4 = CLBLM_R_X11Y146_SLICE_X14Y146_AQ;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_D1 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_D2 = CLBLM_R_X11Y142_SLICE_X14Y142_CO6;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_D3 = LIOB33_X0Y51_IOB_X0Y51_I;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_D4 = CLBLM_R_X11Y142_SLICE_X14Y142_DO6;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_D5 = CLBLM_R_X11Y142_SLICE_X14Y142_BO5;
  assign CLBLM_L_X10Y143_SLICE_X13Y143_D6 = CLBLM_L_X10Y148_SLICE_X13Y148_BO6;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_A1 = CLBLM_L_X10Y142_SLICE_X12Y142_BO6;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_A2 = CLBLM_L_X8Y150_SLICE_X10Y150_A5Q;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_A3 = CLBLM_R_X11Y149_SLICE_X14Y149_AQ;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_A4 = CLBLM_L_X12Y149_SLICE_X16Y149_CO6;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_A5 = 1'b1;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_A6 = 1'b1;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_AX = CLBLM_L_X8Y143_SLICE_X11Y143_AQ;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_B1 = CLBLM_L_X8Y150_SLICE_X10Y150_A5Q;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_B2 = CLBLM_L_X12Y149_SLICE_X16Y149_CO6;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_B3 = CLBLM_R_X11Y149_SLICE_X14Y149_AQ;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_B4 = CLBLM_L_X8Y142_SLICE_X11Y142_DO6;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_B5 = 1'b1;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_B6 = 1'b1;
  assign CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_CE = 1'b1;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_C1 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_C2 = CLBLM_L_X8Y142_SLICE_X11Y142_AQ;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_C3 = CLBLM_L_X10Y149_SLICE_X12Y149_B5Q;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_C4 = CLBLM_L_X8Y142_SLICE_X11Y142_BQ;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_C5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_C6 = 1'b1;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_CE = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_D3 = 1'b1;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_B6 = 1'b1;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_D4 = CLBLM_L_X8Y146_SLICE_X10Y146_A5Q;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_D1 = CLBLM_R_X11Y149_SLICE_X14Y149_AQ;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_D2 = 1'b1;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_D3 = CLBLM_L_X8Y142_SLICE_X11Y142_DO6;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_D4 = CLBLM_L_X8Y150_SLICE_X10Y150_A5Q;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_D5 = CLBLM_L_X10Y142_SLICE_X12Y142_BO6;
  assign CLBLM_L_X10Y143_SLICE_X12Y143_D6 = 1'b1;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_D6 = 1'b1;
  assign LIOB33_X0Y121_IOB_X0Y122_O = CLBLL_L_X4Y149_SLICE_X4Y149_D5Q;
  assign LIOB33_X0Y121_IOB_X0Y121_O = CLBLM_L_X8Y146_SLICE_X10Y146_AQ;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_A5 = CLBLM_L_X10Y145_SLICE_X12Y145_AO6;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_A6 = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_D1 = CLBLM_R_X3Y149_SLICE_X2Y149_CQ;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_A1 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_A2 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_A3 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_A4 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_A5 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_A6 = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_T1 = 1'b1;
  assign RIOI3_X105Y185_OLOGIC_X1Y186_D1 = CLBLM_R_X7Y154_SLICE_X9Y154_CO6;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_B1 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_B2 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_B3 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_B4 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_B5 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_B6 = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_D1 = CLBLL_L_X2Y150_SLICE_X1Y150_C5Q;
  assign RIOI3_X105Y185_OLOGIC_X1Y186_T1 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_C1 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_C2 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_C3 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_C4 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_C5 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_C6 = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_T1 = 1'b1;
  assign RIOI3_X105Y185_OLOGIC_X1Y185_D1 = CLBLM_L_X8Y154_SLICE_X10Y154_BO6;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_D1 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_D2 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_D3 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_D4 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_D5 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_D6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_D1 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign RIOI3_X105Y185_OLOGIC_X1Y185_T1 = 1'b1;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_B6 = CLBLM_R_X11Y146_SLICE_X14Y146_CO6;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_D1 = CLBLL_L_X2Y166_SLICE_X0Y166_AO6;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_A1 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_A2 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_A3 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_A5 = CLBLM_L_X8Y150_SLICE_X11Y150_B5Q;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_A6 = 1'b1;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_C1 = CLBLM_L_X10Y142_SLICE_X13Y142_BO6;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_T1 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_B1 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_B2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_B3 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_B4 = CLBLL_L_X4Y150_SLICE_X4Y150_AQ;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_B5 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_B6 = CLBLM_R_X5Y153_SLICE_X7Y153_CO6;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_A1 = CLBLM_L_X8Y144_SLICE_X10Y144_B5Q;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_A2 = CLBLM_R_X7Y144_SLICE_X8Y144_AQ;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_A6 = CLBLM_L_X8Y144_SLICE_X10Y144_CO6;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_A3 = CLBLM_R_X11Y146_SLICE_X14Y146_AQ;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_C1 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_C2 = CLBLM_R_X5Y153_SLICE_X7Y153_CO6;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_C3 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_C4 = CLBLL_L_X4Y147_SLICE_X4Y147_D5Q;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_C5 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_C6 = CLBLL_L_X4Y150_SLICE_X4Y150_AQ;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_A5 = CLBLM_L_X8Y144_SLICE_X11Y144_A5Q;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_B5 = CLBLM_L_X12Y144_SLICE_X16Y144_AO5;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_B6 = CLBLM_R_X11Y143_SLICE_X15Y143_DO6;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_B1 = CLBLM_R_X11Y144_SLICE_X15Y144_AO5;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_B2 = CLBLM_R_X11Y144_SLICE_X15Y144_CO6;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_B3 = CLBLM_R_X11Y145_SLICE_X15Y145_BO5;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_C2 = CLBLM_R_X11Y146_SLICE_X14Y146_AQ;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_D1 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_D2 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_D3 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_D4 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_D5 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_D6 = 1'b1;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_C1 = CLBLM_R_X5Y142_SLICE_X7Y142_C5Q;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_SR = CLBLL_L_X4Y145_SLICE_X5Y145_CO6;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_C4 = CLBLM_L_X8Y144_SLICE_X11Y144_A5Q;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_C5 = CLBLM_R_X7Y146_SLICE_X9Y146_B5Q;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_C6 = CLBLM_R_X7Y144_SLICE_X8Y144_AQ;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_D1 = CLBLM_R_X11Y145_SLICE_X15Y145_BO5;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_D2 = CLBLM_L_X8Y143_SLICE_X10Y143_DQ;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_D3 = CLBLM_L_X10Y143_SLICE_X13Y143_DO6;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_D4 = CLBLM_R_X11Y144_SLICE_X15Y144_AO5;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_D5 = CLBLM_R_X11Y143_SLICE_X15Y143_DO6;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_D6 = CLBLM_R_X11Y144_SLICE_X15Y144_CO6;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_A1 = CLBLM_L_X10Y142_SLICE_X12Y142_DO6;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_A2 = CLBLM_L_X12Y143_SLICE_X16Y143_AO6;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_A3 = CLBLM_R_X11Y149_SLICE_X14Y149_AQ;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_A4 = CLBLM_R_X7Y142_SLICE_X9Y142_DQ;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_A5 = CLBLM_L_X8Y150_SLICE_X10Y150_A5Q;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_A6 = 1'b1;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_B1 = CLBLM_L_X10Y142_SLICE_X12Y142_DO6;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_B2 = CLBLM_R_X7Y142_SLICE_X9Y142_A5Q;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_B3 = CLBLM_L_X10Y144_SLICE_X13Y144_AO6;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_B4 = CLBLM_R_X11Y149_SLICE_X14Y149_AQ;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_B5 = CLBLM_L_X8Y150_SLICE_X10Y150_A5Q;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_B6 = CLBLL_L_X4Y144_SLICE_X5Y144_DQ;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_C1 = CLBLM_L_X8Y150_SLICE_X10Y150_A5Q;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_C2 = CLBLM_L_X10Y148_SLICE_X12Y148_AQ;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_C3 = CLBLM_L_X10Y142_SLICE_X12Y142_DO6;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_C4 = CLBLM_R_X3Y144_SLICE_X3Y144_DQ;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_C5 = CLBLM_R_X11Y149_SLICE_X14Y149_AQ;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_C6 = CLBLM_R_X11Y142_SLICE_X14Y142_BO6;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_A5 = 1'b1;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_A6 = CLBLL_L_X4Y148_SLICE_X5Y148_DQ;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_D1 = CLBLM_L_X10Y144_SLICE_X12Y144_AO5;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_D2 = CLBLM_L_X10Y143_SLICE_X13Y143_CO6;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_D3 = CLBLM_L_X10Y144_SLICE_X13Y144_BO6;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_D4 = CLBLM_L_X10Y144_SLICE_X12Y144_CO6;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_D5 = CLBLM_R_X11Y143_SLICE_X14Y143_CO5;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_D6 = CLBLM_L_X10Y142_SLICE_X13Y142_BO6;
  assign CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_I = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_B6 = 1'b1;
  assign RIOI3_X105Y125_ILOGIC_X1Y126_D = RIOB33_X105Y125_IOB_X1Y126_I;
  assign RIOI3_X105Y125_ILOGIC_X1Y125_D = RIOB33_X105Y125_IOB_X1Y125_I;
  assign LIOB33_X0Y123_IOB_X0Y124_O = CLBLM_R_X7Y152_SLICE_X9Y152_DQ;
  assign LIOB33_X0Y123_IOB_X0Y123_O = CLBLM_R_X3Y149_SLICE_X2Y149_CQ;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_C1 = CLBLM_R_X5Y145_SLICE_X7Y145_BO6;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_C2 = CLBLM_L_X8Y150_SLICE_X10Y150_A5Q;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_C3 = CLBLM_R_X11Y149_SLICE_X14Y149_AQ;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_C5 = CLBLM_L_X10Y144_SLICE_X13Y144_CO6;
  assign RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y120_D = RIOB33_X105Y119_IOB_X1Y120_I;
  assign RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_D = RIOB33_X105Y119_IOB_X1Y119_I;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_A1 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_A2 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_A3 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_A4 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_A5 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_A6 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_AX = CLBLM_R_X3Y141_SLICE_X2Y141_AO6;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_B1 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_B2 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_B3 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_B4 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_B5 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_B6 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_C1 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_C2 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_C3 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_C4 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_C5 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_C6 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_D1 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_D2 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_D3 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_D4 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_D5 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_D6 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_SR = CLBLM_R_X11Y148_SLICE_X15Y148_CO6;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_A1 = CLBLM_R_X5Y143_SLICE_X6Y143_D5Q;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_A2 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_A3 = CLBLL_L_X4Y140_SLICE_X5Y140_AQ;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_A5 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_A6 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_B1 = LIOB33_X0Y57_IOB_X0Y58_I;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_B2 = CLBLM_R_X3Y142_SLICE_X3Y142_BQ;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_B3 = CLBLL_L_X4Y142_SLICE_X5Y142_AQ;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_B4 = CLBLL_L_X4Y142_SLICE_X5Y142_A5Q;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_B5 = CLBLL_L_X2Y143_SLICE_X1Y143_CQ;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_B6 = 1'b1;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_A1 = CLBLM_R_X11Y145_SLICE_X14Y145_BO5;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_C1 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_C2 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_C3 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_C4 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_C5 = CLBLM_R_X3Y152_SLICE_X3Y152_AQ;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_C6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_A3 = CLBLM_L_X8Y144_SLICE_X10Y144_BQ;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_A4 = CLBLM_R_X5Y145_SLICE_X6Y145_BQ;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_B2 = CLBLL_L_X4Y141_SLICE_X5Y141_AQ;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_B3 = CLBLM_L_X10Y145_SLICE_X12Y145_AO6;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_A5 = CLBLM_L_X10Y144_SLICE_X13Y144_AO6;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_A6 = 1'b1;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_B6 = 1'b1;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_B1 = CLBLM_L_X10Y147_SLICE_X13Y147_B5Q;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_D1 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_D2 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_D3 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_D4 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_D5 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_D6 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_SR = CLBLL_L_X4Y145_SLICE_X5Y145_BO6;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_C1 = CLBLM_L_X8Y145_SLICE_X11Y145_AO6;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_C2 = CLBLM_L_X10Y146_SLICE_X13Y146_CO6;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_C3 = CLBLM_L_X10Y145_SLICE_X12Y145_DO6;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_C4 = CLBLM_R_X11Y143_SLICE_X14Y143_CO5;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_C5 = CLBLM_R_X11Y145_SLICE_X14Y145_CO6;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_C6 = CLBLM_R_X7Y146_SLICE_X8Y146_BO6;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_D1 = CLBLM_R_X7Y147_SLICE_X9Y147_DO5;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_D2 = CLBLM_L_X10Y142_SLICE_X13Y142_BO6;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_D3 = CLBLM_L_X10Y144_SLICE_X13Y144_DO6;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_D4 = CLBLM_R_X11Y143_SLICE_X14Y143_CO5;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_D5 = CLBLM_L_X10Y145_SLICE_X13Y145_BO5;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_D6 = CLBLM_R_X11Y145_SLICE_X14Y145_AO5;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_A1 = CLBLM_L_X10Y142_SLICE_X12Y142_DO6;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_A2 = 1'b1;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_A3 = CLBLM_R_X5Y146_SLICE_X6Y146_AQ;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_A4 = CLBLM_L_X8Y150_SLICE_X10Y150_A5Q;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_A5 = CLBLM_R_X11Y149_SLICE_X14Y149_AQ;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_A6 = 1'b1;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_AX = CLBLM_R_X7Y148_SLICE_X9Y148_BQ;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_B1 = CLBLM_L_X10Y148_SLICE_X12Y148_CO6;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_B2 = CLBLM_L_X8Y145_SLICE_X11Y145_BO6;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_B3 = CLBLM_L_X8Y145_SLICE_X10Y145_CO6;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_B4 = CLBLM_L_X10Y144_SLICE_X12Y144_DO6;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_B5 = CLBLM_L_X10Y145_SLICE_X12Y145_CO6;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_B6 = CLBLM_L_X10Y145_SLICE_X12Y145_AO5;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_C1 = CLBLM_L_X10Y143_SLICE_X12Y143_AO6;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_C2 = 1'b1;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_C3 = CLBLM_L_X10Y146_SLICE_X12Y146_DO6;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_C4 = CLBLM_L_X8Y148_SLICE_X10Y148_CO6;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_C5 = CLBLM_R_X7Y145_SLICE_X9Y145_CQ;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_C6 = CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_CE = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_D1 = CLBLM_L_X10Y143_SLICE_X12Y143_DO5;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_D2 = 1'b1;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_D3 = CLBLM_L_X10Y143_SLICE_X12Y143_DO6;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_D4 = CLBLM_L_X8Y141_SLICE_X10Y141_CQ;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_D5 = CLBLM_R_X5Y153_SLICE_X6Y153_DQ;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_D6 = CLBLM_L_X10Y148_SLICE_X12Y148_BO6;
  assign LIOB33_X0Y125_IOB_X0Y126_O = CLBLM_R_X5Y144_SLICE_X6Y144_CQ;
  assign LIOB33_X0Y125_IOB_X0Y125_O = CLBLM_R_X5Y144_SLICE_X6Y144_DQ;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_C4 = CLBLM_R_X7Y151_SLICE_X8Y151_DO5;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_A1 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_A2 = CLBLL_L_X2Y148_SLICE_X0Y148_BQ;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_A3 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_A5 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_A6 = 1'b1;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_C5 = 1'b1;
  assign RIOI3_X105Y191_OLOGIC_X1Y192_T1 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_AX = CLBLL_L_X4Y142_SLICE_X4Y142_CO6;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_B1 = LIOB33_X0Y57_IOB_X0Y58_I;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_B2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_B3 = CLBLL_L_X4Y143_SLICE_X4Y143_AQ;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_B4 = CLBLL_L_X2Y143_SLICE_X1Y143_CQ;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_B5 = CLBLL_L_X4Y142_SLICE_X5Y142_A5Q;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_B6 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_C2 = CLBLM_L_X10Y143_SLICE_X12Y143_AO5;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_C3 = CLBLL_L_X4Y143_SLICE_X4Y143_DQ;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_C4 = CLBLM_L_X10Y143_SLICE_X12Y143_BO6;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_C5 = CLBLL_L_X2Y143_SLICE_X1Y143_AQ;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_C6 = 1'b1;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_C6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_A1 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_A2 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_A3 = LIOB33_X0Y55_IOB_X0Y56_I;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_A4 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_D4 = CLBLM_L_X10Y142_SLICE_X12Y142_AQ;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_D5 = CLBLL_L_X4Y142_SLICE_X5Y142_BQ;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_D6 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_A5 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_A6 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_D1 = CLBLL_L_X4Y142_SLICE_X5Y142_AQ;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_D2 = CLBLM_R_X3Y142_SLICE_X3Y142_BQ;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_D3 = CLBLL_L_X4Y141_SLICE_X5Y141_BO5;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_B1 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_B2 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_B3 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_B4 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_B5 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_B6 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_SR = CLBLL_L_X4Y141_SLICE_X5Y141_CO6;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_C1 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_C2 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_C3 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_C4 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_C5 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_C6 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_B6 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_D1 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_D2 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_D3 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_D4 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_D5 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_D6 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_A1 = CLBLM_L_X10Y142_SLICE_X12Y142_AQ;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_A2 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_A3 = CLBLL_L_X4Y141_SLICE_X5Y141_BO6;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_A5 = CLBLM_L_X10Y147_SLICE_X13Y147_A5Q;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_A6 = CLBLM_R_X3Y141_SLICE_X3Y141_CO6;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_AX = CLBLL_L_X4Y142_SLICE_X4Y142_BO6;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_B1 = LIOB33_X0Y57_IOB_X0Y58_I;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_B2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_B3 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_B4 = CLBLL_L_X2Y143_SLICE_X1Y143_CQ;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_B5 = CLBLM_R_X5Y143_SLICE_X6Y143_AQ;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_B6 = CLBLL_L_X4Y142_SLICE_X5Y142_A5Q;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_C1 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_C2 = CLBLL_L_X4Y142_SLICE_X5Y142_CQ;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_C3 = CLBLM_L_X10Y150_SLICE_X13Y150_B5Q;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_C4 = CLBLM_L_X10Y143_SLICE_X12Y143_AO6;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_C5 = CLBLL_L_X4Y143_SLICE_X4Y143_BQ;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_C6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_A1 = 1'b1;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_A3 = 1'b1;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_A4 = CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_A5 = 1'b1;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_A6 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_A1 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_A2 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_A3 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_A4 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_D4 = CLBLL_L_X4Y143_SLICE_X5Y143_BQ;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_D5 = CLBLM_L_X10Y143_SLICE_X12Y143_BO6;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_D6 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_A5 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_A6 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_D1 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_D2 = CLBLL_L_X4Y142_SLICE_X5Y142_CQ;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_D3 = CLBLM_L_X10Y143_SLICE_X12Y143_AO5;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_B1 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_B2 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_B3 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_B4 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_B5 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_B6 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_C1 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_C2 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_C3 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_C4 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_C5 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_C6 = 1'b1;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_D1 = CLBLM_R_X3Y146_SLICE_X3Y146_C5Q;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_D2 = CLBLM_R_X11Y142_SLICE_X14Y142_BO6;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_D3 = CLBLM_L_X8Y152_SLICE_X11Y152_AQ;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_D4 = CLBLM_R_X7Y146_SLICE_X9Y146_B5Q;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_D5 = CLBLM_R_X11Y149_SLICE_X14Y149_AQ;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_D6 = CLBLM_L_X8Y150_SLICE_X10Y150_A5Q;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_D1 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_D2 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_D3 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_D4 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_D5 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_D6 = 1'b1;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_A1 = CLBLM_L_X10Y149_SLICE_X12Y149_A5Q;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_A2 = CLBLM_L_X10Y147_SLICE_X12Y147_B5Q;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_A3 = CLBLM_L_X8Y149_SLICE_X11Y149_BQ;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_A4 = CLBLM_R_X5Y146_SLICE_X7Y146_AQ;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_A5 = CLBLM_R_X11Y146_SLICE_X15Y146_AQ;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_A6 = 1'b1;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_AX = CLBLM_R_X11Y145_SLICE_X15Y145_AO6;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_B1 = CLBLL_L_X4Y147_SLICE_X4Y147_BQ;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_B2 = CLBLL_L_X4Y150_SLICE_X5Y150_BQ;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_B3 = CLBLM_L_X10Y148_SLICE_X13Y148_AQ;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_B4 = CLBLM_L_X10Y147_SLICE_X12Y147_CQ;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_B5 = CLBLM_L_X10Y142_SLICE_X12Y142_CO6;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_B6 = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_T1 = 1'b1;
  assign RIOI3_X105Y189_OLOGIC_X1Y189_D1 = CLBLM_R_X103Y178_SLICE_X163Y178_AO6;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_C1 = CLBLM_R_X5Y142_SLICE_X6Y142_BQ;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_C2 = 1'b1;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_C3 = CLBLM_R_X5Y146_SLICE_X7Y146_DQ;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_C4 = CLBLM_R_X11Y144_SLICE_X15Y144_CO6;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_C5 = 1'b1;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_C6 = 1'b1;
  assign RIOI3_X105Y189_OLOGIC_X1Y189_T1 = 1'b1;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_D1 = CLBLM_L_X10Y142_SLICE_X12Y142_CO6;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_D2 = CLBLM_L_X10Y147_SLICE_X12Y147_CQ;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_D3 = CLBLM_R_X11Y143_SLICE_X14Y143_CO5;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_D4 = CLBLM_R_X11Y144_SLICE_X15Y144_CO6;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_D5 = CLBLM_R_X7Y146_SLICE_X9Y146_B5Q;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_D6 = CLBLM_L_X10Y150_SLICE_X13Y150_A5Q;
  assign LIOB33_X0Y127_IOB_X0Y127_O = CLBLM_L_X8Y150_SLICE_X11Y150_B5Q;
  assign LIOB33_X0Y127_IOB_X0Y128_O = CLBLM_L_X8Y142_SLICE_X11Y142_CQ;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_SR = CLBLM_R_X11Y148_SLICE_X14Y148_DO6;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_D6 = 1'b1;
  assign LIOI3_X0Y153_OLOGIC_X0Y154_D1 = CLBLM_L_X8Y152_SLICE_X10Y152_DQ;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_A2 = CLBLM_R_X7Y150_SLICE_X8Y150_C5Q;
  assign LIOI3_X0Y153_OLOGIC_X0Y154_T1 = 1'b1;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_A2 = CLBLL_L_X2Y147_SLICE_X1Y147_AQ;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_A3 = CLBLL_L_X4Y143_SLICE_X4Y143_AQ;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_A4 = CLBLM_R_X5Y149_SLICE_X6Y149_D5Q;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_A5 = CLBLM_L_X8Y149_SLICE_X11Y149_BQ;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_A6 = CLBLM_L_X8Y150_SLICE_X11Y150_B5Q;
  assign LIOI3_X0Y153_OLOGIC_X0Y153_D1 = CLBLM_L_X10Y153_SLICE_X13Y153_AQ;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_B1 = CLBLL_L_X2Y144_SLICE_X1Y144_BQ;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_B2 = CLBLL_L_X4Y143_SLICE_X4Y143_BQ;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_B4 = CLBLM_R_X5Y149_SLICE_X6Y149_D5Q;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_B5 = CLBLL_L_X4Y150_SLICE_X4Y150_AQ;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_B6 = CLBLM_L_X8Y150_SLICE_X11Y150_B5Q;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_C1 = CLBLL_L_X4Y142_SLICE_X5Y142_AQ;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_C2 = CLBLM_L_X10Y142_SLICE_X12Y142_AQ;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_C3 = CLBLL_L_X4Y147_SLICE_X4Y147_CQ;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_C4 = CLBLM_R_X3Y142_SLICE_X3Y142_BQ;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_C5 = CLBLM_R_X7Y150_SLICE_X9Y150_B5Q;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_C6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_D1 = 1'b1;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_D2 = CLBLL_L_X4Y143_SLICE_X4Y143_AQ;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_D3 = CLBLL_L_X4Y143_SLICE_X4Y143_DQ;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_D4 = CLBLM_L_X10Y143_SLICE_X12Y143_AO6;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_D5 = CLBLL_L_X4Y143_SLICE_X5Y143_BQ;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_D6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign RIOI3_X105Y127_ILOGIC_X1Y128_D = RIOB33_X105Y127_IOB_X1Y128_I;
  assign RIOI3_X105Y127_ILOGIC_X1Y127_D = RIOB33_X105Y127_IOB_X1Y127_I;
  assign LIOI3_X0Y153_OLOGIC_X0Y153_T1 = 1'b1;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_A1 = CLBLM_R_X5Y143_SLICE_X7Y143_DQ;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_A2 = CLBLM_R_X5Y142_SLICE_X6Y142_CQ;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_A3 = CLBLL_L_X4Y143_SLICE_X5Y143_AQ;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_A5 = CLBLM_L_X8Y149_SLICE_X11Y149_BQ;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_A6 = CLBLM_R_X7Y142_SLICE_X8Y142_DO6;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_B1 = CLBLL_L_X2Y145_SLICE_X1Y145_AQ;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_B2 = CLBLL_L_X4Y143_SLICE_X5Y143_BQ;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_B3 = CLBLM_R_X3Y148_SLICE_X2Y148_D5Q;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_B5 = CLBLM_R_X5Y144_SLICE_X6Y144_DQ;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_B6 = CLBLM_R_X5Y150_SLICE_X7Y150_A5Q;
  assign RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y132_D = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_C1 = CLBLM_R_X11Y143_SLICE_X14Y143_AQ;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_C2 = CLBLL_L_X2Y153_SLICE_X1Y153_AQ;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_C3 = CLBLM_L_X8Y140_SLICE_X10Y140_AQ;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_C5 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_C6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y131_D = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_A2 = CLBLL_L_X4Y147_SLICE_X4Y147_D5Q;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_A3 = CLBLM_R_X5Y145_SLICE_X7Y145_AQ;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_A4 = CLBLM_L_X8Y147_SLICE_X11Y147_BO6;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_A5 = CLBLM_R_X11Y147_SLICE_X14Y147_BO6;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_D1 = CLBLM_R_X5Y143_SLICE_X6Y143_D5Q;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_D2 = CLBLM_L_X8Y143_SLICE_X11Y143_A5Q;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_D3 = CLBLL_L_X4Y143_SLICE_X5Y143_DQ;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_D4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_D5 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_D6 = CLBLL_L_X2Y149_SLICE_X1Y149_BQ;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_A6 = 1'b1;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_B1 = CLBLM_R_X7Y147_SLICE_X8Y147_CQ;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_B2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_B3 = CLBLL_L_X4Y144_SLICE_X5Y144_BQ;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_B4 = 1'b1;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_B5 = CLBLM_L_X10Y150_SLICE_X13Y150_AQ;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_B6 = 1'b1;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_C1 = CLBLM_R_X5Y149_SLICE_X7Y149_DQ;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_C2 = CLBLM_L_X10Y147_SLICE_X13Y147_CQ;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_C3 = CLBLM_L_X8Y151_SLICE_X11Y151_AQ;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_C4 = CLBLM_L_X8Y147_SLICE_X10Y147_AQ;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_C5 = CLBLM_L_X8Y142_SLICE_X11Y142_CQ;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_C6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_X105Y155_OLOGIC_X1Y156_D1 = 1'b1;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_D1 = CLBLM_R_X5Y149_SLICE_X7Y149_DQ;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_D2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_D3 = CLBLM_L_X10Y147_SLICE_X13Y147_DQ;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_D4 = CLBLM_L_X8Y142_SLICE_X11Y142_CQ;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_D5 = CLBLM_L_X8Y151_SLICE_X11Y151_AQ;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_D6 = CLBLM_R_X3Y151_SLICE_X3Y151_D5Q;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_D6 = 1'b1;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_A1 = CLBLM_L_X10Y147_SLICE_X12Y147_B5Q;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_A2 = CLBLM_R_X11Y145_SLICE_X15Y145_BO5;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_A3 = CLBLM_L_X10Y147_SLICE_X12Y147_AQ;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_A4 = CLBLM_R_X7Y141_SLICE_X8Y141_AQ;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_A5 = 1'b1;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign LIOB33_X0Y129_IOB_X0Y130_O = CLBLM_R_X3Y149_SLICE_X2Y149_BQ;
  assign LIOB33_X0Y129_IOB_X0Y129_O = CLBLM_R_X3Y149_SLICE_X2Y149_CQ;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_B1 = CLBLM_L_X10Y148_SLICE_X12Y148_A5Q;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_B2 = CLBLM_L_X10Y147_SLICE_X12Y147_BQ;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_B3 = CLBLM_R_X3Y151_SLICE_X3Y151_C5Q;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_B5 = CLBLM_L_X8Y148_SLICE_X10Y148_BQ;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_B6 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_C3 = CLBLM_R_X11Y151_SLICE_X14Y151_BQ;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_C1 = CLBLM_L_X10Y150_SLICE_X13Y150_A5Q;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_C2 = 1'b1;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_C3 = CLBLL_L_X4Y148_SLICE_X4Y148_AQ;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_C5 = CLBLM_R_X11Y148_SLICE_X14Y148_DQ;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_C6 = 1'b1;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_D1 = CLBLM_R_X7Y146_SLICE_X9Y146_B5Q;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_D2 = CLBLM_R_X11Y144_SLICE_X15Y144_CO6;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_D3 = CLBLM_R_X7Y147_SLICE_X8Y147_BQ;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_D4 = CLBLM_R_X11Y143_SLICE_X14Y143_CO5;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_D5 = CLBLM_L_X10Y150_SLICE_X13Y150_AQ;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_D6 = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y156_T1 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_D3 = CLBLM_R_X7Y152_SLICE_X9Y152_AQ;
  assign RIOI3_X105Y155_OLOGIC_X1Y155_D1 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_D4 = CLBLM_L_X10Y151_SLICE_X13Y151_CO6;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_A1 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_A2 = CLBLL_L_X2Y153_SLICE_X1Y153_AQ;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_A3 = CLBLM_R_X5Y143_SLICE_X6Y143_DQ;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_A4 = CLBLM_R_X3Y144_SLICE_X3Y144_DQ;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_A5 = CLBLM_R_X3Y146_SLICE_X3Y146_C5Q;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_A6 = CLBLL_L_X4Y144_SLICE_X4Y144_CO6;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_AX = CLBLM_L_X10Y150_SLICE_X12Y150_DO5;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_B1 = CLBLM_R_X3Y145_SLICE_X3Y145_AQ;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_B2 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_B3 = CLBLM_R_X7Y143_SLICE_X9Y143_DQ;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_B4 = CLBLL_L_X2Y143_SLICE_X1Y143_BQ;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_B5 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_B6 = CLBLL_L_X4Y147_SLICE_X5Y147_C5Q;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_C1 = CLBLM_R_X7Y142_SLICE_X9Y142_A5Q;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_C2 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_C3 = CLBLM_R_X3Y146_SLICE_X2Y146_BQ;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_C4 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_C5 = CLBLM_R_X3Y145_SLICE_X2Y145_B5Q;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_C6 = CLBLL_L_X4Y144_SLICE_X5Y144_BQ;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_D1 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_D2 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_D3 = CLBLM_R_X3Y152_SLICE_X3Y152_AQ;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_D4 = CLBLM_R_X7Y144_SLICE_X9Y144_AQ;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_D5 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_D6 = CLBLM_R_X7Y152_SLICE_X8Y152_BQ;
  assign CLBLL_L_X4Y144_SLICE_X4Y144_SR = CLBLL_L_X4Y145_SLICE_X5Y145_CO6;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_A1 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_A2 = CLBLM_R_X5Y144_SLICE_X6Y144_AQ;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_A3 = CLBLL_L_X4Y144_SLICE_X5Y144_AQ;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_A4 = CLBLM_L_X10Y143_SLICE_X12Y143_BO6;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_A5 = CLBLM_R_X7Y142_SLICE_X9Y142_A5Q;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_B1 = CLBLM_R_X3Y145_SLICE_X2Y145_B5Q;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_B2 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_B3 = CLBLL_L_X4Y144_SLICE_X5Y144_CQ;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_B5 = CLBLL_L_X2Y149_SLICE_X1Y149_AQ;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_B6 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_C1 = CLBLM_R_X5Y142_SLICE_X7Y142_CQ;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_C2 = CLBLL_L_X4Y153_SLICE_X4Y153_A5Q;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_C3 = CLBLL_L_X4Y146_SLICE_X5Y146_A5Q;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_C5 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_C6 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_C1 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_A1 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_D1 = CLBLM_R_X3Y143_SLICE_X2Y143_BQ;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_D2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_D3 = 1'b1;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_D4 = CLBLL_L_X4Y152_SLICE_X5Y152_CQ;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_D5 = CLBLM_L_X8Y152_SLICE_X11Y152_A5Q;
  assign CLBLL_L_X4Y144_SLICE_X5Y144_D6 = 1'b1;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_A2 = 1'b1;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_A3 = CLBLM_L_X10Y143_SLICE_X12Y143_AO6;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_A4 = CLBLM_R_X5Y146_SLICE_X7Y146_CQ;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_A5 = CLBLM_L_X8Y148_SLICE_X11Y148_AQ;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_A6 = 1'b1;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_AX = CLBLM_L_X10Y150_SLICE_X13Y150_DO6;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_B1 = CLBLM_R_X11Y149_SLICE_X14Y149_AQ;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_B2 = CLBLM_L_X10Y147_SLICE_X13Y147_BQ;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_B3 = CLBLM_L_X10Y146_SLICE_X12Y146_AQ;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_B4 = CLBLM_L_X8Y150_SLICE_X10Y150_A5Q;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_B5 = CLBLM_L_X10Y143_SLICE_X13Y143_AO6;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_B6 = 1'b1;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_C1 = CLBLM_L_X10Y148_SLICE_X13Y148_AO6;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_C2 = CLBLM_L_X8Y149_SLICE_X11Y149_DO6;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_C3 = CLBLM_L_X10Y149_SLICE_X13Y149_DO6;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_C4 = CLBLM_L_X8Y145_SLICE_X10Y145_BO5;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_C5 = CLBLM_R_X11Y144_SLICE_X15Y144_BO6;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_C6 = CLBLM_R_X5Y148_SLICE_X7Y148_CO6;
  assign LIOB33_X0Y131_IOB_X0Y131_O = CLBLL_L_X2Y75_SLICE_X0Y75_AO6;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOB33_X0Y131_IOB_X0Y132_O = CLBLL_L_X4Y142_SLICE_X4Y142_BO5;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_D1 = CLBLM_L_X10Y147_SLICE_X12Y147_C5Q;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_D2 = CLBLM_L_X8Y150_SLICE_X10Y150_A5Q;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_D3 = CLBLM_L_X10Y144_SLICE_X13Y144_CO6;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_D4 = CLBLM_R_X11Y149_SLICE_X14Y149_AQ;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_D5 = CLBLM_L_X10Y150_SLICE_X13Y150_B5Q;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_D6 = CLBLM_L_X10Y143_SLICE_X13Y143_AO6;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_SR = CLBLM_R_X11Y148_SLICE_X15Y148_AO6;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_A2 = CLBLM_L_X8Y148_SLICE_X10Y148_BQ;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_A3 = 1'b1;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_A4 = CLBLM_L_X8Y147_SLICE_X10Y147_A5Q;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_A5 = 1'b1;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_A6 = 1'b1;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_B1 = CLBLM_L_X10Y144_SLICE_X13Y144_CO6;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_B2 = CLBLM_L_X8Y150_SLICE_X10Y150_A5Q;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_B3 = CLBLM_R_X7Y147_SLICE_X9Y147_C5Q;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_B4 = CLBLM_R_X5Y147_SLICE_X7Y147_CQ;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_B5 = CLBLM_R_X11Y149_SLICE_X14Y149_AQ;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_B6 = 1'b1;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_C1 = CLBLM_L_X10Y143_SLICE_X12Y143_BO6;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_C2 = CLBLM_R_X7Y151_SLICE_X8Y151_CQ;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_C3 = CLBLM_L_X10Y148_SLICE_X13Y148_DO6;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_C4 = CLBLM_L_X10Y144_SLICE_X12Y144_AO6;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_C5 = CLBLM_L_X10Y148_SLICE_X12Y148_DO6;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_C6 = CLBLM_L_X8Y149_SLICE_X11Y149_AQ;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_D1 = 1'b1;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_D2 = CLBLM_L_X10Y143_SLICE_X12Y143_BO5;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_D3 = CLBLM_L_X8Y152_SLICE_X10Y152_BQ;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_D4 = CLBLM_L_X10Y148_SLICE_X12Y148_A5Q;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_D5 = CLBLM_L_X10Y148_SLICE_X12Y148_BO5;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_D6 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_D3 = CLBLM_R_X7Y145_SLICE_X8Y145_B5Q;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_D4 = CLBLM_R_X3Y150_SLICE_X3Y150_BQ;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_SR = CLBLM_R_X11Y148_SLICE_X14Y148_CO6;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_D6 = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_D1 = CLBLM_R_X3Y149_SLICE_X2Y149_DO6;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_A1 = 1'b1;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_A2 = 1'b1;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_A3 = 1'b1;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_A4 = 1'b1;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_A5 = 1'b1;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_A6 = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_T1 = 1'b1;
  assign RIOI3_X105Y191_OLOGIC_X1Y192_D1 = CLBLM_L_X12Y151_SLICE_X16Y151_CO6;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_D4 = 1'b1;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_B1 = 1'b1;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_B2 = 1'b1;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_B3 = 1'b1;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_B4 = 1'b1;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_B5 = 1'b1;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_B6 = 1'b1;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_D5 = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_D1 = CLBLM_R_X5Y147_SLICE_X7Y147_DO6;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_D6 = 1'b1;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_C1 = 1'b1;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_C2 = 1'b1;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_C3 = 1'b1;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_C4 = 1'b1;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_C5 = 1'b1;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_C6 = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_T1 = 1'b1;
  assign RIOI3_X105Y191_OLOGIC_X1Y191_D1 = CLBLM_R_X11Y149_SLICE_X14Y149_AO6;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_D1 = 1'b1;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_D2 = 1'b1;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_D3 = 1'b1;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_D4 = 1'b1;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_D5 = 1'b1;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_D6 = 1'b1;
  assign RIOI3_X105Y191_OLOGIC_X1Y191_T1 = 1'b1;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_A1 = CLBLM_R_X11Y145_SLICE_X15Y145_BO5;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_A2 = CLBLM_L_X10Y147_SLICE_X13Y147_CQ;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_A3 = CLBLM_R_X11Y142_SLICE_X14Y142_AQ;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_A5 = CLBLM_R_X11Y146_SLICE_X15Y146_AQ;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_A6 = 1'b1;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_B1 = CLBLM_L_X8Y144_SLICE_X11Y144_A5Q;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_A1 = CLBLL_L_X2Y148_SLICE_X0Y148_B5Q;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_A3 = 1'b1;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_A4 = CLBLL_L_X2Y143_SLICE_X1Y143_CQ;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_A5 = 1'b1;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_A6 = 1'b1;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_B2 = CLBLM_R_X7Y144_SLICE_X8Y144_AQ;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_B3 = CLBLM_R_X5Y142_SLICE_X7Y142_C5Q;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_B4 = CLBLM_R_X11Y146_SLICE_X14Y146_AQ;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_B1 = CLBLM_L_X10Y142_SLICE_X12Y142_AQ;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_B2 = CLBLL_L_X4Y145_SLICE_X4Y145_CO6;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_B3 = CLBLL_L_X4Y144_SLICE_X4Y144_AO6;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_B4 = CLBLM_R_X3Y142_SLICE_X3Y142_BQ;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_B5 = CLBLL_L_X4Y142_SLICE_X5Y142_AQ;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_B6 = CLBLM_R_X3Y143_SLICE_X2Y143_CQ;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_C1 = CLBLM_R_X11Y149_SLICE_X14Y149_AQ;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_C2 = CLBLM_L_X8Y144_SLICE_X11Y144_A5Q;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_C1 = CLBLM_R_X3Y144_SLICE_X2Y144_BO5;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_C2 = 1'b1;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_C3 = CLBLM_R_X3Y145_SLICE_X2Y145_C5Q;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_C4 = CLBLM_R_X5Y145_SLICE_X6Y145_BQ;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_C5 = CLBLM_R_X3Y145_SLICE_X2Y145_CQ;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_C6 = CLBLL_L_X4Y147_SLICE_X5Y147_BQ;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_D1 = CLBLM_R_X5Y142_SLICE_X7Y142_C5Q;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_D5 = CLBLM_R_X7Y146_SLICE_X9Y146_B5Q;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_D6 = CLBLM_R_X7Y144_SLICE_X8Y144_AQ;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_D2 = CLBLM_R_X11Y146_SLICE_X14Y146_AQ;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_D3 = CLBLM_L_X8Y144_SLICE_X11Y144_A5Q;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_D1 = 1'b1;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_D2 = 1'b1;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_D3 = 1'b1;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_D4 = 1'b1;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_D5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_D6 = CLBLL_L_X4Y153_SLICE_X5Y153_BQ;
  assign CLBLL_L_X4Y145_SLICE_X4Y145_SR = CLBLL_L_X4Y145_SLICE_X4Y145_DO6;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_A1 = CLBLL_L_X4Y141_SLICE_X4Y141_AQ;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_A2 = CLBLM_L_X12Y149_SLICE_X16Y149_CO6;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_A3 = CLBLM_L_X10Y143_SLICE_X12Y143_BO6;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_A4 = CLBLM_R_X3Y145_SLICE_X2Y145_AQ;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_A5 = CLBLM_R_X7Y146_SLICE_X8Y146_AO6;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_A6 = 1'b1;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_AX = CLBLL_L_X4Y142_SLICE_X5Y142_AQ;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_B1 = 1'b1;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_B2 = CLBLM_R_X7Y150_SLICE_X8Y150_C5Q;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_B3 = 1'b1;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_B4 = 1'b1;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_B6 = 1'b1;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_B6 = CLBLM_R_X11Y147_SLICE_X14Y147_CO6;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_BX = CLBLM_R_X5Y144_SLICE_X6Y144_CQ;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_C1 = CLBLM_R_X7Y152_SLICE_X8Y152_BQ;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_C2 = 1'b1;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_C3 = 1'b1;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_C4 = 1'b1;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_C5 = 1'b1;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_C6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_CE = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOB33_X0Y133_IOB_X0Y134_O = CLBLM_R_X3Y149_SLICE_X2Y149_BQ;
  assign LIOB33_X0Y133_IOB_X0Y133_O = CLBLM_R_X3Y142_SLICE_X2Y142_CO5;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_D1 = 1'b1;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_D2 = 1'b1;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_D3 = 1'b1;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_D4 = 1'b1;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_D5 = 1'b1;
  assign CLBLL_L_X4Y145_SLICE_X5Y145_D6 = 1'b1;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_A1 = 1'b1;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_A3 = CLBLM_L_X8Y152_SLICE_X11Y152_AQ;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_A4 = 1'b1;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_A5 = 1'b1;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_A6 = 1'b1;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_AX = CLBLM_R_X7Y149_SLICE_X9Y149_AO6;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_B1 = CLBLM_R_X7Y148_SLICE_X9Y148_B5Q;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_B2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_B3 = 1'b1;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_B4 = CLBLM_R_X11Y149_SLICE_X15Y149_AQ;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_B5 = CLBLM_R_X3Y152_SLICE_X3Y152_A5Q;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_B6 = 1'b1;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_D4 = CLBLM_L_X10Y143_SLICE_X12Y143_DO6;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_C1 = CLBLM_L_X8Y150_SLICE_X10Y150_BO6;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_C2 = CLBLM_L_X10Y148_SLICE_X13Y148_AO5;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_C3 = CLBLM_L_X10Y147_SLICE_X12Y147_DO6;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_C4 = CLBLM_L_X8Y150_SLICE_X10Y150_DO6;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_C5 = CLBLM_L_X10Y148_SLICE_X13Y148_BO5;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_C6 = CLBLM_R_X11Y144_SLICE_X14Y144_BO6;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_D5 = CLBLM_L_X8Y149_SLICE_X10Y149_A5Q;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_D6 = CLBLM_R_X7Y147_SLICE_X8Y147_D5Q;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_D1 = CLBLM_L_X8Y150_SLICE_X10Y150_A5Q;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_D2 = 1'b1;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_D3 = CLBLM_L_X10Y143_SLICE_X13Y143_AO6;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_D4 = CLBLM_L_X10Y149_SLICE_X13Y149_A5Q;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_D5 = CLBLM_L_X10Y149_SLICE_X13Y149_AQ;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_D6 = CLBLM_R_X11Y149_SLICE_X14Y149_AQ;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_DX = CLBLL_L_X4Y149_SLICE_X4Y149_CQ;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_SR = CLBLM_R_X11Y148_SLICE_X15Y148_CO6;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_A1 = CLBLM_L_X10Y150_SLICE_X13Y150_C5Q;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_A2 = CLBLM_L_X10Y148_SLICE_X12Y148_A5Q;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_A3 = CLBLM_L_X10Y146_SLICE_X12Y146_AO6;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_A5 = 1'b1;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_A6 = 1'b1;
  assign RIOI3_X105Y129_ILOGIC_X1Y130_D = RIOB33_X105Y129_IOB_X1Y130_I;
  assign RIOI3_X105Y129_ILOGIC_X1Y129_D = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_B1 = CLBLM_R_X11Y151_SLICE_X15Y151_A5Q;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_B2 = CLBLM_L_X8Y148_SLICE_X11Y148_C5Q;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_B4 = CLBLM_L_X10Y150_SLICE_X13Y150_CQ;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_B5 = CLBLL_L_X4Y143_SLICE_X4Y143_CQ;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_B6 = 1'b1;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_C1 = CLBLM_L_X10Y143_SLICE_X12Y143_AO6;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_C2 = CLBLM_L_X10Y149_SLICE_X12Y149_CQ;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_C3 = 1'b1;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_C5 = CLBLM_L_X10Y149_SLICE_X13Y149_A5Q;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_C6 = CLBLM_L_X8Y150_SLICE_X11Y150_AQ;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_A4 = CLBLM_R_X7Y150_SLICE_X8Y150_AQ;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_D1 = CLBLM_L_X8Y149_SLICE_X11Y149_AQ;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_D2 = CLBLM_L_X10Y143_SLICE_X12Y143_AO6;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_D3 = CLBLM_L_X10Y149_SLICE_X12Y149_DQ;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_D4 = CLBLM_R_X5Y149_SLICE_X7Y149_AQ;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_D5 = 1'b1;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_D6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_A1 = RIOB33_X105Y127_IOB_X1Y127_I;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_A2 = RIOB33_X105Y125_IOB_X1Y125_I;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_A3 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_A4 = RIOB33_X105Y125_IOB_X1Y126_I;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_A5 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_A6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y144_D = RIOB33_X105Y143_IOB_X1Y144_I;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_B1 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_B2 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_B3 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_B4 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_B5 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_B6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y143_D = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_C1 = 1'b1;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_C4 = CLBLM_L_X8Y151_SLICE_X10Y151_DQ;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_C2 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_C3 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_C4 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_C5 = 1'b1;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_C5 = CLBLM_R_X5Y151_SLICE_X6Y151_DQ;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_C6 = 1'b1;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_C6 = CLBLM_R_X3Y152_SLICE_X2Y152_BQ;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_D1 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_D2 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_D3 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_D4 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_D5 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_D6 = 1'b1;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_B5 = CLBLM_R_X7Y149_SLICE_X8Y149_BQ;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_A1 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_A2 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_A3 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_A4 = 1'b1;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_B6 = CLBLM_R_X7Y150_SLICE_X9Y150_AQ;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_A1 = CLBLM_L_X10Y142_SLICE_X13Y142_AQ;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_A2 = CLBLM_R_X11Y143_SLICE_X14Y143_BO6;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_A3 = CLBLM_L_X12Y145_SLICE_X16Y145_AO6;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_A4 = CLBLM_R_X11Y143_SLICE_X15Y143_BO6;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_A5 = RIOB33_X105Y139_IOB_X1Y140_I;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_A6 = CLBLM_R_X11Y145_SLICE_X15Y145_BO5;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_A5 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_A6 = 1'b1;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_B1 = CLBLM_R_X11Y142_SLICE_X14Y142_DO6;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_B2 = CLBLM_R_X11Y142_SLICE_X14Y142_BO5;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_B3 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_B4 = CLBLM_R_X11Y142_SLICE_X14Y142_CO6;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_B5 = CLBLM_R_X11Y148_SLICE_X14Y148_AQ;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_B6 = CLBLM_L_X8Y144_SLICE_X10Y144_CO6;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_B2 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_B3 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_B5 = 1'b1;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_C1 = CLBLM_R_X11Y142_SLICE_X14Y142_CO6;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_C2 = CLBLM_R_X11Y142_SLICE_X14Y142_BO5;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_C3 = CLBLM_R_X11Y142_SLICE_X14Y142_DO6;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_C4 = CLBLM_L_X10Y148_SLICE_X13Y148_BO6;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_C5 = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_C6 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_C1 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_C2 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_C3 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_C4 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_C5 = 1'b1;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_D2 = 1'b1;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_D1 = CLBLM_R_X11Y142_SLICE_X14Y142_CO6;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_D2 = CLBLM_R_X11Y142_SLICE_X14Y142_BO5;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_D3 = 1'b1;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_D4 = CLBLM_L_X10Y148_SLICE_X13Y148_BO6;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_D5 = CLBLM_R_X11Y143_SLICE_X14Y143_CO6;
  assign CLBLM_R_X11Y143_SLICE_X15Y143_D6 = CLBLM_R_X11Y142_SLICE_X14Y142_BO6;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_D1 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_D2 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_D3 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_D4 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_D5 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_D6 = 1'b1;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_A1 = CLBLM_R_X11Y143_SLICE_X14Y143_DO6;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_D5 = CLBLM_L_X12Y149_SLICE_X16Y149_CO6;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_A2 = CLBLM_R_X7Y144_SLICE_X9Y144_CQ;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_A3 = CLBLM_L_X12Y144_SLICE_X16Y144_BO6;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_A5 = RIOB33_X105Y139_IOB_X1Y139_I;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_D6 = CLBLM_L_X8Y151_SLICE_X10Y151_AQ;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_A1 = CLBLM_L_X8Y146_SLICE_X10Y146_DQ;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_A2 = CLBLM_L_X10Y143_SLICE_X12Y143_BO6;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_A3 = CLBLL_L_X4Y146_SLICE_X4Y146_AQ;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_A5 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_A6 = CLBLM_R_X3Y146_SLICE_X2Y146_AQ;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_A6 = CLBLM_L_X10Y143_SLICE_X12Y143_AQ;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_B1 = CLBLM_L_X8Y150_SLICE_X10Y150_A5Q;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_B1 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_B2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_B3 = CLBLM_R_X3Y142_SLICE_X2Y142_BQ;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_B4 = CLBLL_L_X2Y148_SLICE_X0Y148_BQ;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_B5 = CLBLM_R_X3Y144_SLICE_X3Y144_D5Q;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_B6 = CLBLL_L_X4Y148_SLICE_X5Y148_CQ;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_B5 = CLBLM_R_X11Y149_SLICE_X15Y149_CQ;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_SR = CLBLL_L_X4Y145_SLICE_X5Y145_CO6;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_C2 = CLBLL_L_X4Y146_SLICE_X4Y146_CQ;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_C3 = CLBLM_R_X3Y149_SLICE_X2Y149_CQ;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_C4 = CLBLM_R_X5Y147_SLICE_X6Y147_AQ;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_C5 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_C6 = CLBLM_L_X10Y143_SLICE_X12Y143_AO6;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_C3 = CLBLM_R_X7Y146_SLICE_X9Y146_B5Q;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_C4 = CLBLM_R_X7Y144_SLICE_X8Y144_AQ;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_C6 = 1'b1;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_D1 = CLBLM_R_X11Y148_SLICE_X14Y148_AQ;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_D2 = RIOB33_X105Y139_IOB_X1Y140_I;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_D1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_D2 = CLBLM_R_X3Y146_SLICE_X3Y146_BQ;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_D3 = CLBLL_L_X4Y146_SLICE_X4Y146_DQ;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_D4 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_D5 = CLBLL_L_X4Y147_SLICE_X4Y147_DQ;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_D6 = CLBLM_L_X10Y143_SLICE_X12Y143_AO6;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_D3 = CLBLM_R_X11Y145_SLICE_X14Y145_AQ;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_D4 = RIOB33_X105Y141_IOB_X1Y141_I;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_D5 = 1'b1;
  assign CLBLM_R_X11Y143_SLICE_X14Y143_D6 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_A1 = CLBLM_R_X7Y148_SLICE_X9Y148_AQ;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_A2 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_A3 = CLBLL_L_X4Y144_SLICE_X5Y144_AQ;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_A5 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_A6 = 1'b1;
  assign LIOB33_X0Y135_IOB_X0Y136_O = CLBLM_L_X8Y153_SLICE_X10Y153_AQ;
  assign LIOB33_X0Y135_IOB_X0Y135_O = CLBLM_R_X3Y149_SLICE_X2Y149_BQ;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_B1 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_B2 = CLBLM_L_X8Y142_SLICE_X11Y142_BQ;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_B3 = CLBLL_L_X2Y146_SLICE_X1Y146_AQ;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_B4 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_B6 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_C2 = CLBLM_R_X7Y144_SLICE_X9Y144_AQ;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_C3 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_C4 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_C5 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_C6 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_D1 = CLBLM_R_X7Y142_SLICE_X8Y142_DO6;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_D2 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_D3 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_D4 = CLBLL_L_X4Y143_SLICE_X5Y143_AQ;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_D5 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_D6 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_SR = CLBLL_L_X4Y146_SLICE_X5Y146_CO6;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_A2 = CLBLM_L_X10Y145_SLICE_X12Y145_BO6;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_A3 = CLBLM_L_X10Y149_SLICE_X12Y149_DQ;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_A4 = CLBLM_L_X10Y149_SLICE_X13Y149_CO6;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_A5 = CLBLM_L_X8Y152_SLICE_X10Y152_D5Q;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_A6 = 1'b1;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_B6 = 1'b1;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_B2 = CLBLM_L_X10Y150_SLICE_X13Y150_BQ;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_B3 = CLBLM_R_X11Y150_SLICE_X15Y150_AQ;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_B4 = CLBLM_R_X11Y152_SLICE_X14Y152_AQ;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_B5 = CLBLM_R_X3Y148_SLICE_X2Y148_B5Q;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_B6 = CLBLM_L_X8Y146_SLICE_X10Y146_A5Q;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_BX = CLBLM_L_X10Y151_SLICE_X13Y151_BO6;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_A1 = 1'b1;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_A2 = 1'b1;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_A3 = 1'b1;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_C4 = CLBLM_L_X10Y149_SLICE_X12Y149_BQ;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_C5 = CLBLL_L_X4Y150_SLICE_X5Y150_CQ;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_C6 = 1'b1;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_A4 = 1'b1;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_A5 = 1'b1;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_A6 = 1'b1;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_C1 = CLBLM_L_X10Y149_SLICE_X13Y149_A5Q;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_C2 = CLBLM_R_X11Y151_SLICE_X14Y151_BQ;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_B1 = 1'b1;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_B2 = 1'b1;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_B3 = 1'b1;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_B4 = 1'b1;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_D2 = CLBLM_L_X10Y147_SLICE_X13Y147_B5Q;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_B5 = 1'b1;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_B6 = 1'b1;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_D5 = CLBLM_L_X10Y148_SLICE_X12Y148_AQ;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_D6 = 1'b1;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_D1 = CLBLM_L_X8Y154_SLICE_X10Y154_AQ;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_C1 = 1'b1;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_C2 = 1'b1;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_C3 = 1'b1;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_C4 = 1'b1;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_C5 = 1'b1;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_C6 = 1'b1;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_A2 = CLBLM_L_X10Y151_SLICE_X12Y151_BO6;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_A3 = CLBLM_R_X11Y151_SLICE_X14Y151_CO6;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_A4 = CLBLL_L_X4Y150_SLICE_X5Y150_BQ;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_A5 = CLBLM_L_X8Y145_SLICE_X11Y145_AQ;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_A6 = 1'b1;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_D1 = 1'b1;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_D2 = 1'b1;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_D3 = 1'b1;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_D4 = 1'b1;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_D5 = 1'b1;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_D6 = 1'b1;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_B6 = CLBLM_R_X11Y152_SLICE_X14Y152_A5Q;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_B2 = CLBLM_L_X10Y150_SLICE_X12Y150_BQ;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_B3 = CLBLM_R_X3Y148_SLICE_X2Y148_B5Q;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_B4 = CLBLM_L_X10Y150_SLICE_X12Y150_DO6;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_B5 = 1'b1;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_A1 = 1'b1;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_C5 = CLBLM_L_X10Y151_SLICE_X12Y151_CO6;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_C6 = 1'b1;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_A3 = CLBLM_R_X5Y142_SLICE_X6Y142_DQ;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_A4 = CLBLM_R_X7Y144_SLICE_X9Y144_A5Q;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_A5 = 1'b1;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_A6 = 1'b1;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_B1 = 1'b1;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_B2 = 1'b1;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_B3 = 1'b1;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_B4 = 1'b1;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_B5 = 1'b1;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_B6 = 1'b1;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_D1 = CLBLM_R_X11Y150_SLICE_X15Y150_AQ;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_D2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_C1 = 1'b1;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_C2 = 1'b1;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_C3 = 1'b1;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_C4 = 1'b1;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_C5 = 1'b1;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_C6 = 1'b1;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_D5 = CLBLM_L_X10Y150_SLICE_X13Y150_BQ;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_D1 = 1'b1;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_D2 = 1'b1;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_D3 = 1'b1;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_D4 = 1'b1;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_D5 = 1'b1;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_D6 = 1'b1;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_SR = CLBLM_R_X11Y148_SLICE_X15Y148_CO6;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_A1 = CLBLM_L_X8Y150_SLICE_X10Y150_A5Q;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_A2 = CLBLM_R_X11Y149_SLICE_X14Y149_AQ;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_A3 = CLBLM_R_X11Y143_SLICE_X14Y143_CO6;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_A4 = CLBLM_R_X11Y146_SLICE_X14Y146_AQ;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_A5 = CLBLM_R_X11Y149_SLICE_X15Y149_AQ;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_A6 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_B1 = CLBLM_L_X10Y144_SLICE_X12Y144_BO6;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_B2 = CLBLM_R_X11Y143_SLICE_X15Y143_AO6;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_B3 = CLBLM_L_X10Y142_SLICE_X13Y142_BO6;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_B4 = CLBLM_L_X12Y144_SLICE_X16Y144_CO6;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_B5 = CLBLM_R_X11Y143_SLICE_X14Y143_CO5;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_B6 = CLBLM_R_X11Y145_SLICE_X15Y145_CO6;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_C1 = CLBLM_R_X11Y146_SLICE_X14Y146_AQ;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_C2 = CLBLM_R_X7Y144_SLICE_X8Y144_AQ;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_C3 = CLBLM_L_X8Y144_SLICE_X11Y144_A5Q;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_C4 = CLBLM_L_X8Y144_SLICE_X10Y144_B5Q;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_C5 = CLBLM_R_X5Y142_SLICE_X7Y142_C5Q;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_C6 = CLBLM_L_X10Y148_SLICE_X13Y148_BO6;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_D1 = CLBLM_R_X11Y144_SLICE_X15Y144_CO6;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_D2 = CLBLM_R_X11Y143_SLICE_X15Y143_CO6;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_D3 = CLBLM_R_X11Y143_SLICE_X15Y143_DO6;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_D4 = CLBLM_R_X11Y144_SLICE_X15Y144_AO5;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_D5 = CLBLM_R_X11Y145_SLICE_X15Y145_BO5;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_D6 = CLBLM_R_X11Y142_SLICE_X14Y142_AQ;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_A1 = CLBLM_L_X12Y145_SLICE_X16Y145_AO6;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_A2 = CLBLM_L_X10Y143_SLICE_X13Y143_BO6;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_A1 = 1'b1;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_A3 = CLBLL_L_X4Y148_SLICE_X4Y148_CO5;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_A4 = CLBLM_R_X3Y147_SLICE_X3Y147_CO5;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_A5 = CLBLM_R_X5Y144_SLICE_X7Y144_BQ;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_A6 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_A3 = CLBLM_R_X11Y144_SLICE_X15Y144_AO6;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_A4 = RIOB33_X105Y139_IOB_X1Y139_I;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_A5 = CLBLM_L_X10Y147_SLICE_X13Y147_DQ;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_B1 = CLBLL_L_X4Y148_SLICE_X4Y148_CO6;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_B2 = CLBLL_L_X4Y147_SLICE_X4Y147_BQ;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_B4 = CLBLM_R_X3Y147_SLICE_X3Y147_AQ;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_B5 = CLBLM_R_X7Y145_SLICE_X8Y145_C5Q;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_B6 = CLBLM_R_X3Y146_SLICE_X3Y146_CQ;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_AX = CLBLM_R_X11Y142_SLICE_X14Y142_AQ;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_B1 = CLBLM_L_X12Y144_SLICE_X16Y144_DO6;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_B2 = CLBLM_L_X10Y145_SLICE_X13Y145_BO6;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_C2 = CLBLM_R_X5Y144_SLICE_X7Y144_CQ;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_C3 = CLBLL_L_X4Y143_SLICE_X5Y143_DQ;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_C4 = CLBLL_L_X2Y150_SLICE_X1Y150_C5Q;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_C5 = CLBLM_R_X5Y147_SLICE_X7Y147_C5Q;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_C6 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_C1 = CLBLM_R_X11Y142_SLICE_X14Y142_CO5;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_C2 = CLBLM_R_X11Y144_SLICE_X15Y144_AO5;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_C3 = CLBLM_R_X11Y145_SLICE_X15Y145_BO5;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_C4 = CLBLM_R_X11Y143_SLICE_X14Y143_BO5;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_C5 = CLBLM_L_X12Y145_SLICE_X16Y145_AO6;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_C6 = CLBLM_R_X11Y144_SLICE_X15Y144_CO6;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_D1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_D2 = CLBLM_R_X5Y145_SLICE_X6Y145_B5Q;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_D3 = CLBLL_L_X2Y148_SLICE_X1Y148_A5Q;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_D4 = CLBLL_L_X2Y144_SLICE_X1Y144_B5Q;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_D5 = CLBLM_R_X3Y147_SLICE_X2Y147_C5Q;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_D6 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_D1 = CLBLM_R_X3Y145_SLICE_X2Y145_BQ;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_D2 = CLBLM_R_X7Y150_SLICE_X8Y150_C5Q;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_D3 = CLBLM_R_X7Y146_SLICE_X9Y146_B5Q;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_D4 = CLBLM_L_X8Y150_SLICE_X10Y150_A5Q;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_D5 = CLBLM_R_X11Y149_SLICE_X14Y149_AQ;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_D6 = CLBLM_R_X11Y142_SLICE_X14Y142_BO6;
  assign LIOB33_X0Y137_IOB_X0Y138_O = CLBLM_R_X3Y144_SLICE_X3Y144_A5Q;
  assign LIOB33_X0Y137_IOB_X0Y137_O = CLBLM_R_X7Y150_SLICE_X9Y150_B5Q;
  assign LIOI3_X0Y151_OLOGIC_X0Y152_D1 = CLBLM_R_X3Y150_SLICE_X2Y150_B5Q;
  assign LIOI3_SING_X0Y50_ILOGIC_X0Y50_D = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign LIOI3_X0Y151_OLOGIC_X0Y152_T1 = 1'b1;
  assign RIOI3_X105Y195_OLOGIC_X1Y196_D1 = CLBLM_R_X11Y150_SLICE_X14Y150_BO6;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_A1 = CLBLL_L_X4Y150_SLICE_X5Y150_BQ;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_A2 = CLBLM_R_X5Y147_SLICE_X7Y147_AQ;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_A3 = CLBLL_L_X4Y147_SLICE_X5Y147_AQ;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_A5 = CLBLL_L_X4Y151_SLICE_X4Y151_AO5;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_A6 = CLBLM_R_X3Y146_SLICE_X3Y146_CQ;
  assign LIOI3_X0Y151_OLOGIC_X0Y151_D1 = CLBLM_R_X3Y149_SLICE_X2Y149_CQ;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_B2 = 1'b1;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_B1 = CLBLM_R_X3Y145_SLICE_X2Y145_CQ;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_B2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_B3 = CLBLM_R_X3Y147_SLICE_X3Y147_AQ;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_B4 = CLBLM_L_X8Y148_SLICE_X11Y148_AQ;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_B5 = CLBLL_L_X4Y147_SLICE_X5Y147_C5Q;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_B6 = 1'b1;
  assign RIOI3_X105Y195_OLOGIC_X1Y196_T1 = 1'b1;
  assign LIOI3_X0Y151_OLOGIC_X0Y151_T1 = 1'b1;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_C2 = CLBLM_R_X5Y146_SLICE_X6Y146_BQ;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_C3 = CLBLM_R_X3Y152_SLICE_X3Y152_AQ;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_C4 = CLBLM_R_X7Y148_SLICE_X9Y148_CQ;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_C5 = CLBLL_L_X4Y152_SLICE_X4Y152_CQ;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_C6 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_B5 = 1'b1;
  assign RIOI3_X105Y195_OLOGIC_X1Y195_D1 = CLBLM_R_X11Y149_SLICE_X14Y149_BO6;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_X105Y195_OLOGIC_X1Y195_T1 = 1'b1;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_D1 = CLBLM_R_X5Y153_SLICE_X6Y153_BQ;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_D2 = CLBLM_R_X3Y148_SLICE_X2Y148_CQ;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_D3 = CLBLL_L_X4Y147_SLICE_X5Y147_DQ;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_D4 = CLBLL_L_X4Y148_SLICE_X5Y148_CQ;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_D5 = CLBLM_R_X5Y154_SLICE_X7Y154_AQ;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_D6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_A1 = CLBLM_R_X3Y148_SLICE_X2Y148_B5Q;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_A2 = CLBLM_R_X3Y142_SLICE_X2Y142_A5Q;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_A3 = CLBLM_L_X10Y151_SLICE_X12Y151_AO6;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_A4 = CLBLM_R_X7Y152_SLICE_X9Y152_AQ;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_A6 = CLBLM_L_X10Y151_SLICE_X13Y151_AQ;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_C1 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_B1 = CLBLM_R_X7Y152_SLICE_X9Y152_AQ;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_B2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_B3 = CLBLM_L_X10Y151_SLICE_X13Y151_AQ;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_B4 = CLBLM_L_X10Y151_SLICE_X12Y151_AO6;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_B5 = CLBLM_L_X10Y151_SLICE_X12Y151_AQ;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_B6 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_C2 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_D1 = 1'b1;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_A1 = 1'b1;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_A2 = 1'b1;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_A3 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_C4 = CLBLM_L_X10Y151_SLICE_X13Y151_AQ;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_C5 = CLBLM_R_X7Y152_SLICE_X9Y152_AQ;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_C6 = CLBLM_L_X10Y152_SLICE_X13Y152_BQ;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_A4 = 1'b1;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_A5 = 1'b1;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_A6 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_C1 = CLBLM_R_X11Y151_SLICE_X15Y151_AQ;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_C2 = CLBLM_L_X10Y151_SLICE_X12Y151_AO5;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_B1 = 1'b1;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_B2 = 1'b1;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_B3 = 1'b1;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_B4 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_D2 = CLBLM_L_X10Y151_SLICE_X12Y151_AO6;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_B5 = 1'b1;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_B6 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_D5 = CLBLM_L_X10Y151_SLICE_X13Y151_AQ;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_D6 = CLBLM_L_X10Y152_SLICE_X13Y152_BQ;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_D1 = CLBLM_R_X11Y151_SLICE_X14Y151_BQ;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_C1 = 1'b1;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_C2 = 1'b1;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_C3 = 1'b1;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_C4 = 1'b1;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_C5 = 1'b1;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_C6 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_A1 = CLBLM_L_X8Y146_SLICE_X10Y146_A5Q;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_A2 = CLBLM_L_X10Y150_SLICE_X12Y150_A5Q;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_A3 = CLBLM_R_X11Y150_SLICE_X15Y150_AQ;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_A4 = CLBLM_L_X10Y150_SLICE_X12Y150_BQ;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_A5 = CLBLM_L_X10Y150_SLICE_X13Y150_BQ;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_AX = CLBLM_L_X8Y151_SLICE_X10Y151_CO6;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_A6 = 1'b1;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_D1 = 1'b1;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_D2 = 1'b1;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_D3 = 1'b1;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_D4 = 1'b1;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_D5 = 1'b1;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_D6 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_B1 = CLBLM_R_X3Y148_SLICE_X2Y148_B5Q;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_B2 = CLBLM_L_X10Y150_SLICE_X12Y150_A5Q;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_B3 = CLBLM_R_X11Y150_SLICE_X15Y150_AQ;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_B4 = CLBLM_L_X10Y150_SLICE_X12Y150_BQ;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_B5 = CLBLM_L_X10Y150_SLICE_X13Y150_BQ;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_B6 = CLBLM_L_X8Y146_SLICE_X10Y146_A5Q;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_A1 = CLBLM_L_X8Y142_SLICE_X10Y142_A5Q;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_C4 = CLBLM_R_X5Y149_SLICE_X7Y149_D5Q;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_C5 = CLBLM_R_X7Y153_SLICE_X8Y153_DO5;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_C6 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_A2 = CLBLM_L_X8Y142_SLICE_X11Y142_BQ;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_A3 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_A4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_A5 = 1'b1;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_B1 = 1'b1;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_B2 = CLBLM_L_X8Y141_SLICE_X10Y141_BQ;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_B3 = CLBLM_L_X10Y143_SLICE_X12Y143_AO6;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_B5 = CLBLM_R_X3Y142_SLICE_X2Y142_AQ;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_B6 = CLBLM_L_X8Y144_SLICE_X11Y144_A5Q;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_D1 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_D2 = 1'b1;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_C1 = 1'b1;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_C2 = CLBLM_L_X8Y141_SLICE_X10Y141_CQ;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_C3 = CLBLM_L_X10Y142_SLICE_X12Y142_AQ;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_C4 = CLBLM_L_X8Y143_SLICE_X10Y143_BQ;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_C5 = CLBLM_L_X10Y143_SLICE_X12Y143_AO6;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_C6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_D5 = 1'b1;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_SR = CLBLM_R_X11Y148_SLICE_X14Y148_CO6;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_D5 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_D6 = 1'b1;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_D1 = CLBLM_R_X7Y143_SLICE_X9Y143_BQ;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_D2 = 1'b1;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_D3 = 1'b1;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_D4 = 1'b1;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_D5 = 1'b1;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_D6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_SR = CLBLL_L_X4Y141_SLICE_X5Y141_CO6;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_A1 = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_A2 = CLBLM_L_X10Y145_SLICE_X12Y145_AQ;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_A3 = CLBLM_R_X11Y146_SLICE_X15Y146_CO5;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_A5 = CLBLM_R_X11Y142_SLICE_X14Y142_CO5;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_A6 = 1'b1;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_AX = CLBLM_L_X10Y146_SLICE_X13Y146_AQ;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_B1 = CLBLM_R_X11Y149_SLICE_X14Y149_AQ;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_B2 = CLBLM_L_X12Y149_SLICE_X16Y149_CO6;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_B3 = CLBLM_L_X8Y150_SLICE_X10Y150_A5Q;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_B4 = CLBLM_R_X11Y142_SLICE_X14Y142_BO6;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_B5 = CLBLM_R_X7Y146_SLICE_X9Y146_B5Q;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_B6 = 1'b1;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_C1 = CLBLM_L_X12Y143_SLICE_X16Y143_AO6;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_C2 = CLBLL_L_X4Y145_SLICE_X5Y145_BQ;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_C3 = CLBLM_R_X11Y149_SLICE_X14Y149_AQ;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_C4 = CLBLM_L_X8Y150_SLICE_X10Y150_A5Q;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_C5 = CLBLM_L_X8Y152_SLICE_X11Y152_A5Q;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_C6 = CLBLM_R_X11Y145_SLICE_X15Y145_BO6;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_CE = LIOB33_X0Y61_IOB_X0Y62_I;
  assign RIOI3_X105Y133_ILOGIC_X1Y134_D = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_X105Y133_ILOGIC_X1Y133_D = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_D1 = CLBLM_R_X11Y146_SLICE_X15Y146_CO5;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_D2 = CLBLM_R_X11Y144_SLICE_X14Y144_AQ;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_D3 = 1'b1;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_D4 = CLBLM_L_X12Y145_SLICE_X16Y145_CO6;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_D5 = 1'b1;
  assign CLBLM_R_X11Y145_SLICE_X15Y145_D6 = CLBLM_L_X10Y142_SLICE_X13Y142_BO6;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_A1 = CLBLM_R_X5Y149_SLICE_X6Y149_DQ;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_A3 = 1'b1;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_A4 = CLBLM_R_X3Y149_SLICE_X3Y149_BQ;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_A5 = 1'b1;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_A6 = 1'b1;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_A1 = CLBLM_R_X11Y144_SLICE_X14Y144_DO6;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_A2 = CLBLM_L_X10Y142_SLICE_X13Y142_BO6;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_A3 = CLBLM_R_X11Y146_SLICE_X15Y146_CO5;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_B1 = CLBLL_L_X4Y143_SLICE_X5Y143_AQ;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_B2 = CLBLM_R_X7Y142_SLICE_X8Y142_DO6;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_B3 = CLBLM_R_X7Y147_SLICE_X9Y147_AQ;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_B4 = CLBLL_L_X2Y148_SLICE_X0Y148_A5Q;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_B5 = CLBLL_L_X4Y148_SLICE_X5Y148_AQ;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_B6 = 1'b1;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_A5 = CLBLM_R_X11Y145_SLICE_X15Y145_AQ;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_A6 = 1'b1;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_BX = CLBLL_L_X2Y148_SLICE_X1Y148_BO5;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_AX = CLBLM_R_X3Y145_SLICE_X2Y145_AQ;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_C1 = CLBLL_L_X4Y147_SLICE_X5Y147_AQ;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_C2 = CLBLL_L_X4Y150_SLICE_X5Y150_BQ;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_C3 = CLBLM_R_X7Y149_SLICE_X8Y149_AQ;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_C4 = CLBLM_R_X7Y150_SLICE_X8Y150_AQ;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_C5 = CLBLM_R_X7Y150_SLICE_X8Y150_CQ;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_C6 = 1'b1;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_B4 = 1'b1;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_B5 = CLBLM_L_X8Y150_SLICE_X10Y150_A5Q;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_BX = CLBLM_R_X7Y147_SLICE_X9Y147_BQ;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_C1 = CLBLM_L_X10Y142_SLICE_X13Y142_BO6;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_C2 = CLBLM_R_X11Y145_SLICE_X15Y145_AO5;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_C3 = CLBLM_R_X11Y147_SLICE_X14Y147_AQ;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_C4 = CLBLM_L_X12Y145_SLICE_X16Y145_DO6;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_D1 = CLBLL_L_X4Y148_SLICE_X5Y148_AQ;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_D2 = CLBLM_L_X8Y149_SLICE_X11Y149_BQ;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_D3 = CLBLL_L_X4Y147_SLICE_X4Y147_DQ;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_D4 = CLBLL_L_X4Y149_SLICE_X4Y149_AQ;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_D5 = CLBLL_L_X4Y148_SLICE_X4Y148_BO5;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_D6 = CLBLL_L_X4Y148_SLICE_X5Y148_BQ;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_CX = CLBLM_R_X11Y147_SLICE_X14Y147_A5Q;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_SR = CLBLM_R_X5Y153_SLICE_X7Y153_DO6;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_D1 = CLBLM_R_X11Y142_SLICE_X14Y142_CO5;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_D2 = CLBLM_L_X12Y145_SLICE_X16Y145_AO6;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_D3 = 1'b1;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_D4 = RIOB33_X105Y141_IOB_X1Y141_I;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_D5 = 1'b1;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_D6 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X11Y145_SLICE_X14Y145_DX = CLBLM_R_X11Y145_SLICE_X14Y145_CQ;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_A1 = CLBLL_L_X4Y148_SLICE_X5Y148_AQ;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_A2 = CLBLM_L_X10Y149_SLICE_X12Y149_B5Q;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_A3 = CLBLM_R_X5Y147_SLICE_X6Y147_B5Q;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_A5 = CLBLM_L_X8Y149_SLICE_X11Y149_BQ;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_A6 = CLBLL_L_X4Y148_SLICE_X4Y148_BO5;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_B1 = CLBLM_R_X7Y145_SLICE_X8Y145_AQ;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_B2 = CLBLM_R_X5Y145_SLICE_X6Y145_BQ;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_B3 = CLBLM_R_X5Y144_SLICE_X6Y144_C5Q;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_B5 = CLBLL_L_X4Y148_SLICE_X4Y148_DO6;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_B6 = 1'b1;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_C2 = CLBLM_R_X7Y152_SLICE_X9Y152_C5Q;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_C3 = CLBLL_L_X4Y146_SLICE_X4Y146_BQ;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_C4 = CLBLM_R_X3Y144_SLICE_X3Y144_D5Q;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_C5 = CLBLL_L_X4Y148_SLICE_X5Y148_CQ;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_C6 = CLBLL_L_X2Y148_SLICE_X0Y148_BQ;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_D1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_D2 = 1'b1;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_D3 = CLBLM_R_X5Y149_SLICE_X6Y149_D5Q;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_D4 = CLBLM_R_X3Y143_SLICE_X2Y143_AQ;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_D5 = CLBLM_R_X3Y145_SLICE_X2Y145_DQ;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_D6 = CLBLM_L_X10Y147_SLICE_X13Y147_A5Q;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_A1 = CLBLM_L_X10Y152_SLICE_X13Y152_DO6;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_A2 = 1'b1;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_A3 = CLBLM_L_X10Y152_SLICE_X13Y152_AQ;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_A4 = CLBLM_R_X11Y152_SLICE_X15Y152_BO6;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_A6 = CLBLM_L_X10Y150_SLICE_X12Y150_A5Q;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_B1 = CLBLM_L_X10Y151_SLICE_X13Y151_BO5;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_B2 = CLBLM_L_X10Y152_SLICE_X13Y152_BQ;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_B3 = CLBLM_R_X11Y151_SLICE_X14Y151_BQ;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_B5 = CLBLM_L_X10Y152_SLICE_X12Y152_CQ;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_B6 = CLBLM_R_X3Y148_SLICE_X2Y148_B5Q;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_A1 = CLBLM_L_X8Y152_SLICE_X11Y152_B5Q;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_A2 = CLBLM_L_X8Y142_SLICE_X11Y142_BQ;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_A3 = CLBLM_L_X8Y142_SLICE_X11Y142_AQ;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_C4 = CLBLM_L_X8Y153_SLICE_X10Y153_AQ;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_C5 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_A5 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_D2 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_A6 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_C2 = CLBLM_R_X3Y150_SLICE_X3Y150_BQ;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_B1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_B2 = CLBLM_L_X8Y142_SLICE_X11Y142_BQ;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_B3 = CLBLM_L_X8Y142_SLICE_X11Y142_AQ;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_B5 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_B6 = CLBLL_L_X4Y142_SLICE_X4Y142_AQ;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_D1 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_C1 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_C2 = CLBLL_L_X4Y142_SLICE_X4Y142_A5Q;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_C3 = CLBLM_R_X5Y146_SLICE_X7Y146_DQ;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_C4 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_C5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_C6 = 1'b1;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_D4 = CLBLM_L_X10Y152_SLICE_X13Y152_CO6;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_A1 = CLBLM_L_X10Y152_SLICE_X12Y152_DO6;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_A2 = CLBLM_R_X5Y149_SLICE_X7Y149_D5Q;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_A3 = CLBLM_L_X10Y152_SLICE_X13Y152_CO5;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_A4 = CLBLM_L_X10Y152_SLICE_X12Y152_AQ;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_D1 = CLBLM_L_X8Y144_SLICE_X11Y144_A5Q;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_D2 = CLBLM_R_X7Y146_SLICE_X9Y146_B5Q;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_D3 = CLBLM_L_X8Y144_SLICE_X10Y144_B5Q;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_D4 = CLBLM_R_X11Y146_SLICE_X14Y146_AQ;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_D5 = CLBLM_R_X7Y144_SLICE_X8Y144_AQ;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_D6 = CLBLM_R_X5Y142_SLICE_X7Y142_C5Q;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_A6 = CLBLM_L_X10Y151_SLICE_X12Y151_DO6;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_B1 = CLBLM_R_X11Y152_SLICE_X14Y152_CO6;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_B2 = CLBLM_L_X10Y152_SLICE_X12Y152_BQ;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_B3 = CLBLM_L_X10Y152_SLICE_X13Y152_CO5;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_B4 = CLBLM_L_X10Y151_SLICE_X12Y151_DO6;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_A1 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_A2 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_A3 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_A4 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_A6 = 1'b1;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_C1 = CLBLM_R_X11Y152_SLICE_X15Y152_BO6;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_C2 = CLBLM_L_X10Y152_SLICE_X13Y152_CO6;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_AX = CLBLM_R_X5Y142_SLICE_X7Y142_AO6;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_C3 = CLBLM_R_X11Y152_SLICE_X14Y152_DO6;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_C3 = CLBLM_R_X7Y145_SLICE_X8Y145_B5Q;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_B1 = CLBLM_L_X8Y150_SLICE_X10Y150_A5Q;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_B2 = CLBLM_L_X8Y142_SLICE_X11Y142_DO6;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_B3 = CLBLM_R_X11Y149_SLICE_X14Y149_AQ;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_B4 = CLBLM_R_X3Y146_SLICE_X2Y146_BQ;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_B6 = 1'b1;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_D1 = CLBLM_R_X11Y151_SLICE_X14Y151_AQ;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_D2 = CLBLM_R_X11Y152_SLICE_X14Y152_A5Q;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_C2 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_C3 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_C4 = CLBLM_L_X8Y148_SLICE_X11Y148_BQ;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_C5 = CLBLM_R_X3Y142_SLICE_X2Y142_AQ;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_C6 = 1'b1;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_D3 = CLBLM_L_X10Y153_SLICE_X12Y153_BQ;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_D4 = CLBLM_L_X10Y153_SLICE_X12Y153_AQ;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_D5 = CLBLM_L_X8Y152_SLICE_X11Y152_B5Q;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_C6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_D1 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_D1 = CLBLM_L_X10Y149_SLICE_X12Y149_A5Q;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_D2 = CLBLM_R_X11Y146_SLICE_X15Y146_AQ;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_D3 = CLBLM_R_X5Y146_SLICE_X7Y146_AQ;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_D4 = CLBLM_R_X7Y142_SLICE_X9Y142_AQ;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_D5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_D6 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_SR = CLBLM_L_X8Y141_SLICE_X10Y141_DO6;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_A1 = CLBLM_L_X8Y149_SLICE_X11Y149_BQ;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_A2 = CLBLM_L_X8Y151_SLICE_X10Y151_BQ;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_A3 = CLBLM_R_X11Y146_SLICE_X15Y146_AQ;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_D2 = CLBLM_L_X12Y151_SLICE_X16Y151_BQ;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_A5 = CLBLM_L_X12Y149_SLICE_X16Y149_AQ;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_A6 = CLBLM_R_X5Y146_SLICE_X7Y146_AQ;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_D3 = 1'b1;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_B1 = CLBLM_R_X11Y148_SLICE_X14Y148_CQ;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_B2 = CLBLM_R_X11Y145_SLICE_X14Y145_BQ;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_B4 = RIOB33_X105Y145_IOB_X1Y145_I;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_B5 = CLBLM_R_X5Y151_SLICE_X6Y151_BQ;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_B6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_T1 = 1'b1;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_D5 = CLBLM_L_X10Y152_SLICE_X13Y152_AQ;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_C1 = RIOB33_X105Y145_IOB_X1Y145_I;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_C2 = CLBLM_R_X11Y149_SLICE_X14Y149_AQ;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_C3 = CLBLM_R_X11Y148_SLICE_X14Y148_CQ;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_C4 = CLBLM_L_X8Y150_SLICE_X10Y150_A5Q;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_D6 = CLBLM_L_X12Y151_SLICE_X16Y151_DO6;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_C5 = CLBLM_R_X11Y142_SLICE_X14Y142_DO6;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_C6 = 1'b1;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_D1 = CLBLM_R_X11Y146_SLICE_X14Y146_AO6;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_D2 = CLBLM_L_X10Y142_SLICE_X13Y142_BO6;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_D3 = CLBLM_L_X10Y146_SLICE_X12Y146_BO5;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_D4 = CLBLM_R_X11Y144_SLICE_X15Y144_DO6;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_A1 = CLBLM_R_X5Y151_SLICE_X6Y151_B5Q;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_A2 = CLBLL_L_X4Y149_SLICE_X4Y149_BQ;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_A3 = CLBLL_L_X4Y149_SLICE_X4Y149_AQ;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_A4 = CLBLM_L_X8Y149_SLICE_X11Y149_BQ;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_A5 = CLBLL_L_X4Y148_SLICE_X4Y148_BO6;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_D5 = CLBLM_R_X11Y143_SLICE_X14Y143_CO5;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_D6 = CLBLM_R_X11Y145_SLICE_X15Y145_DO6;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_A1 = 1'b1;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_B1 = CLBLL_L_X4Y147_SLICE_X4Y147_C5Q;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_B2 = CLBLL_L_X4Y151_SLICE_X4Y151_AQ;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_B3 = CLBLM_R_X3Y151_SLICE_X3Y151_BQ;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_B5 = CLBLM_L_X10Y150_SLICE_X13Y150_B5Q;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_B6 = 1'b1;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_A2 = CLBLM_L_X8Y144_SLICE_X10Y144_A5Q;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_A3 = 1'b1;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_A4 = CLBLM_L_X8Y147_SLICE_X11Y147_A5Q;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_C2 = CLBLM_R_X5Y148_SLICE_X7Y148_AQ;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_C3 = CLBLL_L_X4Y149_SLICE_X4Y149_DQ;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_C4 = CLBLM_L_X10Y150_SLICE_X12Y150_CQ;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_C5 = 1'b1;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_C6 = 1'b1;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_AX = CLBLM_R_X11Y145_SLICE_X14Y145_AO6;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_B1 = CLBLM_R_X11Y147_SLICE_X14Y147_DO6;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_B2 = CLBLM_R_X5Y145_SLICE_X7Y145_CO6;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_B3 = CLBLM_R_X11Y146_SLICE_X14Y146_DO6;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_B4 = CLBLM_R_X11Y143_SLICE_X14Y143_CO5;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_B5 = CLBLM_L_X8Y145_SLICE_X10Y145_DO6;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_D1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_D2 = CLBLL_L_X2Y148_SLICE_X1Y148_AQ;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_D3 = CLBLM_R_X3Y148_SLICE_X2Y148_D5Q;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_D4 = CLBLM_R_X5Y148_SLICE_X6Y148_CO6;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_D5 = CLBLL_L_X4Y149_SLICE_X4Y149_D5Q;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_D6 = 1'b1;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_C3 = CLBLM_R_X11Y147_SLICE_X15Y147_BO6;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_C4 = CLBLM_L_X12Y145_SLICE_X16Y145_AO5;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_C6 = CLBLM_R_X11Y144_SLICE_X14Y144_CO6;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_D1 = CLBLM_L_X12Y145_SLICE_X17Y145_CO6;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_D2 = CLBLM_L_X10Y142_SLICE_X13Y142_BO6;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_D3 = CLBLM_R_X7Y150_SLICE_X8Y150_DQ;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_D4 = CLBLM_L_X12Y146_SLICE_X16Y146_BO6;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_D5 = 1'b1;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_D6 = CLBLM_R_X11Y145_SLICE_X14Y145_BO5;
  assign LIOI3_SING_X0Y100_OLOGIC_X0Y100_D1 = CLBLM_R_X3Y149_SLICE_X2Y149_AQ;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_SR = CLBLM_R_X11Y148_SLICE_X15Y148_BO6;
  assign LIOI3_SING_X0Y100_OLOGIC_X0Y100_T1 = 1'b1;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_A1 = CLBLM_R_X5Y149_SLICE_X6Y149_DQ;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_A2 = CLBLM_L_X8Y146_SLICE_X10Y146_AQ;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_A3 = CLBLL_L_X4Y149_SLICE_X5Y149_AQ;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_A4 = CLBLL_L_X4Y146_SLICE_X5Y146_AQ;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_A6 = CLBLM_R_X7Y150_SLICE_X9Y150_CQ;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_B1 = CLBLL_L_X4Y148_SLICE_X5Y148_DQ;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_B2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_B3 = CLBLM_R_X3Y145_SLICE_X2Y145_DQ;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_B4 = CLBLM_R_X7Y150_SLICE_X8Y150_C5Q;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_B5 = CLBLL_L_X4Y146_SLICE_X4Y146_AQ;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_B6 = CLBLM_R_X3Y143_SLICE_X2Y143_AQ;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_C1 = CLBLL_L_X4Y149_SLICE_X5Y149_BQ;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_C2 = CLBLM_R_X5Y149_SLICE_X6Y149_A5Q;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_C3 = CLBLM_L_X10Y147_SLICE_X13Y147_AQ;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_C4 = CLBLM_R_X3Y143_SLICE_X2Y143_AQ;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_C5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_C6 = CLBLM_R_X3Y145_SLICE_X2Y145_DQ;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_D1 = CLBLL_L_X4Y146_SLICE_X5Y146_AQ;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_D2 = CLBLM_L_X8Y142_SLICE_X11Y142_CQ;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_D3 = CLBLM_R_X5Y149_SLICE_X7Y149_DQ;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_D4 = CLBLL_L_X4Y149_SLICE_X5Y149_DQ;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_D5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_D6 = CLBLM_R_X5Y152_SLICE_X6Y152_CQ;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_B6 = CLBLM_R_X7Y155_SLICE_X8Y155_AQ;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_A1 = CLBLM_R_X5Y148_SLICE_X6Y148_AO5;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_A2 = CLBLM_R_X11Y149_SLICE_X15Y149_AQ;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_A3 = CLBLM_L_X10Y153_SLICE_X13Y153_AQ;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_A5 = CLBLM_L_X8Y149_SLICE_X11Y149_BQ;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_A6 = CLBLM_L_X10Y153_SLICE_X12Y153_CQ;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_B1 = 1'b1;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_B2 = 1'b1;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_B3 = 1'b1;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_B4 = 1'b1;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_B5 = 1'b1;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_B6 = 1'b1;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_C2 = 1'b1;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_C3 = 1'b1;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_C4 = 1'b1;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_C5 = 1'b1;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_C6 = 1'b1;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_A2 = CLBLM_L_X8Y143_SLICE_X11Y143_BQ;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_A3 = CLBLM_L_X8Y143_SLICE_X11Y143_AQ;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_A4 = CLBLM_L_X10Y143_SLICE_X12Y143_AO6;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_A5 = CLBLM_L_X8Y148_SLICE_X10Y148_AQ;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_A6 = 1'b1;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_C5 = CLBLM_R_X7Y144_SLICE_X8Y144_A5Q;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_AX = CLBLM_L_X10Y143_SLICE_X12Y143_CO5;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_B1 = CLBLM_R_X5Y149_SLICE_X6Y149_D5Q;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_B2 = CLBLM_L_X8Y143_SLICE_X11Y143_BQ;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_D1 = 1'b1;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_D2 = 1'b1;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_B3 = CLBLM_L_X8Y145_SLICE_X11Y145_AQ;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_B4 = CLBLM_L_X8Y150_SLICE_X11Y150_B5Q;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_D5 = 1'b1;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_D6 = 1'b1;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_B6 = CLBLM_L_X8Y141_SLICE_X10Y141_CQ;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_C1 = CLBLM_L_X8Y142_SLICE_X11Y142_C5Q;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_C2 = CLBLM_L_X8Y143_SLICE_X11Y143_CQ;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_C3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_C4 = CLBLM_L_X8Y143_SLICE_X11Y143_A5Q;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_C5 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_C6 = CLBLM_R_X7Y146_SLICE_X8Y146_BQ;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_A1 = CLBLM_R_X7Y147_SLICE_X9Y147_C5Q;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_A2 = CLBLM_L_X10Y151_SLICE_X12Y151_DO6;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_A3 = CLBLM_L_X10Y153_SLICE_X12Y153_AQ;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_A4 = CLBLM_L_X10Y153_SLICE_X12Y153_DO5;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_A5 = CLBLM_L_X10Y152_SLICE_X13Y152_CO5;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_D1 = CLBLM_L_X10Y150_SLICE_X12Y150_BQ;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_D2 = CLBLM_L_X8Y142_SLICE_X11Y142_CQ;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_D3 = CLBLM_L_X8Y143_SLICE_X11Y143_DQ;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_D4 = CLBLM_L_X8Y142_SLICE_X10Y142_AQ;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_D5 = CLBLM_R_X5Y149_SLICE_X7Y149_DQ;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_B5 = CLBLM_L_X10Y152_SLICE_X13Y152_CO5;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_B6 = CLBLM_L_X8Y153_SLICE_X10Y153_BQ;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_D6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_B2 = CLBLM_L_X10Y153_SLICE_X12Y153_BQ;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_B3 = CLBLM_L_X10Y151_SLICE_X12Y151_DO6;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_A1 = CLBLM_L_X8Y147_SLICE_X10Y147_BQ;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_A2 = CLBLM_R_X7Y145_SLICE_X8Y145_BQ;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_C5 = CLBLM_L_X8Y149_SLICE_X11Y149_BQ;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_C6 = CLBLL_L_X4Y151_SLICE_X5Y151_A5Q;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_A3 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_A5 = CLBLM_R_X5Y144_SLICE_X6Y144_CQ;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_A6 = CLBLM_R_X3Y147_SLICE_X3Y147_BQ;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_C2 = CLBLM_L_X10Y153_SLICE_X12Y153_CQ;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_C3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_B1 = CLBLM_R_X7Y148_SLICE_X9Y148_B5Q;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_B2 = CLBLM_L_X8Y143_SLICE_X10Y143_BQ;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_B3 = CLBLM_R_X5Y144_SLICE_X6Y144_DQ;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_B5 = CLBLM_R_X7Y150_SLICE_X9Y150_CQ;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_B6 = CLBLM_L_X8Y146_SLICE_X10Y146_AQ;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_D1 = CLBLM_L_X10Y153_SLICE_X12Y153_BQ;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_D2 = CLBLM_L_X10Y153_SLICE_X12Y153_AQ;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_C1 = CLBLM_L_X8Y142_SLICE_X11Y142_C5Q;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_C2 = CLBLM_L_X8Y143_SLICE_X10Y143_CQ;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_C3 = CLBLM_L_X8Y146_SLICE_X10Y146_AQ;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_C4 = CLBLM_R_X7Y150_SLICE_X9Y150_CQ;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_C5 = CLBLM_R_X7Y145_SLICE_X8Y145_BQ;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_C6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_D5 = CLBLM_L_X8Y152_SLICE_X11Y152_B5Q;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_X105Y197_OLOGIC_X1Y197_T1 = 1'b1;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_D1 = CLBLM_L_X8Y146_SLICE_X11Y146_AQ;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_D2 = 1'b1;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_D3 = CLBLM_L_X8Y143_SLICE_X10Y143_DQ;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_D4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_D5 = CLBLM_L_X8Y143_SLICE_X11Y143_DQ;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_D6 = CLBLM_L_X8Y153_SLICE_X10Y153_BQ;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_D6 = CLBLM_R_X11Y145_SLICE_X15Y145_BO5;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_D1 = CLBLM_R_X7Y153_SLICE_X9Y153_CQ;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_T1 = 1'b1;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_A1 = CLBLM_L_X10Y148_SLICE_X13Y148_AQ;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_A2 = CLBLL_L_X4Y152_SLICE_X5Y152_B5Q;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_A3 = CLBLM_R_X11Y147_SLICE_X15Y147_AQ;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_A6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_D1 = CLBLM_R_X7Y152_SLICE_X9Y152_BQ;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_D2 = 1'b1;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_B1 = CLBLL_L_X4Y147_SLICE_X5Y147_BQ;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_B2 = CLBLM_R_X7Y146_SLICE_X9Y146_B5Q;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_B3 = CLBLM_R_X11Y142_SLICE_X14Y142_BO6;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_B4 = CLBLM_L_X8Y150_SLICE_X10Y150_A5Q;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_B5 = CLBLM_R_X3Y148_SLICE_X2Y148_C5Q;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_B6 = CLBLM_R_X11Y149_SLICE_X14Y149_AQ;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_D3 = 1'b1;
  assign LIOB33_X0Y143_IOB_X0Y143_O = CLBLL_L_X2Y150_SLICE_X1Y150_DO5;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_D4 = 1'b1;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_C1 = CLBLM_R_X11Y146_SLICE_X15Y146_CO5;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_C2 = CLBLM_R_X7Y146_SLICE_X9Y146_B5Q;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_C3 = CLBLM_L_X10Y142_SLICE_X13Y142_BO6;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_C4 = CLBLM_R_X11Y144_SLICE_X15Y144_CO6;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_C5 = CLBLM_L_X10Y147_SLICE_X13Y147_A5Q;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_C6 = CLBLM_R_X11Y145_SLICE_X14Y145_AQ;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_D5 = 1'b1;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_D6 = 1'b1;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_A1 = CLBLM_R_X7Y152_SLICE_X8Y152_BQ;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_A2 = CLBLM_R_X5Y144_SLICE_X7Y144_CQ;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_A3 = CLBLM_R_X3Y144_SLICE_X3Y144_CQ;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_A4 = CLBLM_R_X7Y144_SLICE_X9Y144_AQ;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_A5 = CLBLM_R_X3Y152_SLICE_X3Y152_AQ;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_A6 = 1'b1;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_D1 = 1'b1;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_D2 = CLBLM_R_X11Y147_SLICE_X14Y147_A5Q;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_AX = CLBLL_L_X4Y151_SLICE_X5Y151_DQ;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_D3 = CLBLM_L_X10Y145_SLICE_X12Y145_AO6;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_B1 = CLBLM_R_X7Y152_SLICE_X8Y152_BQ;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_B2 = CLBLL_L_X4Y150_SLICE_X5Y150_CQ;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_B3 = CLBLM_R_X7Y144_SLICE_X9Y144_AQ;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_B4 = CLBLM_R_X5Y151_SLICE_X7Y151_BO6;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_B6 = CLBLL_L_X4Y150_SLICE_X4Y150_AO5;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_A4 = CLBLM_L_X10Y149_SLICE_X12Y149_CQ;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_A6 = 1'b1;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_C1 = CLBLM_R_X5Y153_SLICE_X6Y153_AQ;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_C2 = CLBLL_L_X4Y153_SLICE_X5Y153_BQ;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_C3 = CLBLM_R_X3Y151_SLICE_X3Y151_AQ;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_C4 = CLBLL_L_X4Y150_SLICE_X5Y150_CQ;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_C5 = CLBLM_R_X3Y151_SLICE_X3Y151_BQ;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_C6 = CLBLM_R_X5Y151_SLICE_X7Y151_BO6;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_CE = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_B1 = CLBLM_L_X8Y144_SLICE_X11Y144_DO6;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_B2 = CLBLM_R_X7Y146_SLICE_X9Y146_CO6;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_B3 = CLBLM_R_X11Y147_SLICE_X15Y147_CO6;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_B4 = CLBLM_R_X11Y143_SLICE_X14Y143_CO5;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_B5 = CLBLM_R_X7Y149_SLICE_X9Y149_BO5;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_D1 = CLBLL_L_X2Y150_SLICE_X1Y150_C5Q;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_D2 = CLBLL_L_X4Y147_SLICE_X4Y147_C5Q;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_D3 = CLBLM_R_X3Y144_SLICE_X3Y144_A5Q;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_D4 = CLBLL_L_X2Y148_SLICE_X0Y148_AQ;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_D5 = CLBLM_L_X8Y153_SLICE_X10Y153_AQ;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_D6 = CLBLL_L_X2Y147_SLICE_X0Y147_BQ;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_C1 = CLBLM_L_X10Y147_SLICE_X12Y147_DO5;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_C2 = CLBLM_R_X11Y144_SLICE_X14Y144_CO6;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_C3 = CLBLM_R_X11Y145_SLICE_X14Y145_DO6;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_C4 = CLBLM_R_X11Y146_SLICE_X14Y146_AO5;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_C5 = CLBLM_L_X10Y142_SLICE_X13Y142_BO6;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_C6 = CLBLM_L_X10Y145_SLICE_X13Y145_AO5;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_D1 = CLBLM_R_X5Y145_SLICE_X7Y145_AQ;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_D2 = 1'b1;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_D3 = 1'b1;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_D4 = CLBLM_L_X10Y144_SLICE_X12Y144_AO6;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_D5 = 1'b1;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_D6 = 1'b1;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_A4 = CLBLM_R_X11Y148_SLICE_X14Y148_BO6;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_A5 = CLBLM_L_X10Y147_SLICE_X13Y147_A5Q;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_SR = CLBLM_R_X11Y148_SLICE_X15Y148_BO6;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_A1 = CLBLL_L_X4Y150_SLICE_X5Y150_AQ;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_A2 = CLBLM_R_X3Y149_SLICE_X2Y149_BQ;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_A3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_A4 = CLBLL_L_X4Y148_SLICE_X4Y148_BQ;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_A5 = CLBLM_R_X5Y149_SLICE_X6Y149_D5Q;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_A6 = CLBLM_L_X8Y150_SLICE_X11Y150_B5Q;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_B1 = 1'b1;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_B2 = CLBLL_L_X4Y150_SLICE_X5Y150_BQ;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_B3 = CLBLL_L_X4Y148_SLICE_X5Y148_AQ;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_B5 = CLBLL_L_X4Y151_SLICE_X4Y151_AO5;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_B6 = CLBLM_R_X3Y146_SLICE_X3Y146_CQ;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_C4 = 1'b1;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_AX = CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_C5 = CLBLM_L_X10Y147_SLICE_X12Y147_AQ;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_C1 = CLBLM_R_X5Y143_SLICE_X6Y143_DQ;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_C2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_C3 = CLBLL_L_X4Y150_SLICE_X4Y150_BO6;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_C4 = CLBLL_L_X4Y149_SLICE_X5Y149_BQ;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_C5 = CLBLL_L_X2Y148_SLICE_X0Y148_B5Q;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_C6 = 1'b1;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_C6 = 1'b1;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_B1 = CLBLM_L_X8Y152_SLICE_X11Y152_A5Q;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_B2 = CLBLM_R_X3Y148_SLICE_X2Y148_C5Q;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_B3 = 1'b1;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_D1 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign RIOI3_X105Y135_ILOGIC_X1Y136_D = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_D1 = CLBLM_R_X5Y150_SLICE_X6Y150_C5Q;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_D2 = CLBLM_R_X3Y152_SLICE_X3Y152_BO6;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_D3 = CLBLM_R_X5Y144_SLICE_X7Y144_DQ;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_D4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_D5 = 1'b1;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_D6 = 1'b1;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_B4 = CLBLM_L_X10Y150_SLICE_X13Y150_A5Q;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_T1 = 1'b1;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_B6 = CLBLM_L_X10Y150_SLICE_X13Y150_AQ;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_D1 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign LIOI3_X0Y103_OLOGIC_X0Y103_T1 = 1'b1;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_D2 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_A1 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_A2 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_A3 = CLBLM_L_X8Y142_SLICE_X10Y142_C5Q;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_A5 = CLBLM_R_X5Y147_SLICE_X7Y147_C5Q;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_A6 = 1'b1;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_D3 = CLBLM_R_X7Y149_SLICE_X8Y149_AQ;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_D4 = CLBLM_R_X3Y152_SLICE_X3Y152_A5Q;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_B1 = CLBLM_R_X5Y148_SLICE_X6Y148_B5Q;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_B2 = CLBLM_R_X7Y148_SLICE_X8Y148_BO5;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_B3 = CLBLM_L_X8Y141_SLICE_X10Y141_BQ;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_B4 = CLBLM_L_X10Y144_SLICE_X12Y144_AO6;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_B5 = CLBLL_L_X4Y143_SLICE_X5Y143_CQ;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_B6 = CLBLM_L_X10Y143_SLICE_X12Y143_DO5;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_D5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_D6 = CLBLM_R_X7Y149_SLICE_X9Y149_C5Q;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_C1 = CLBLM_L_X12Y149_SLICE_X16Y149_CO6;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_C2 = CLBLM_R_X5Y144_SLICE_X7Y144_DQ;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_C3 = CLBLM_L_X8Y142_SLICE_X10Y142_BO5;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_C4 = CLBLM_R_X7Y144_SLICE_X9Y144_BQ;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_C5 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_C6 = CLBLM_R_X7Y148_SLICE_X8Y148_BO5;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_D1 = CLBLM_L_X8Y144_SLICE_X10Y144_AQ;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_D2 = CLBLM_L_X8Y145_SLICE_X10Y145_CO5;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_D3 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_D4 = CLBLM_L_X8Y145_SLICE_X11Y145_AO5;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_D5 = CLBLM_L_X10Y143_SLICE_X12Y143_AO5;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_D6 = CLBLM_L_X8Y143_SLICE_X11Y143_AQ;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_SR = CLBLL_L_X4Y145_SLICE_X5Y145_BO6;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_A1 = CLBLM_R_X5Y154_SLICE_X7Y154_DQ;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_A2 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_A3 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_A5 = CLBLL_L_X4Y142_SLICE_X5Y142_A5Q;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_A6 = 1'b1;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_B1 = CLBLM_R_X5Y146_SLICE_X7Y146_B5Q;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_B2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_B3 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_B4 = CLBLL_L_X4Y152_SLICE_X5Y152_C5Q;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_B5 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_B6 = 1'b1;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_A2 = CLBLM_L_X8Y147_SLICE_X11Y147_A5Q;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_A3 = CLBLM_R_X7Y150_SLICE_X8Y150_AQ;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_C1 = CLBLM_R_X11Y149_SLICE_X14Y149_AQ;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_C2 = CLBLM_L_X10Y144_SLICE_X13Y144_CO6;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_C3 = CLBLM_L_X8Y150_SLICE_X10Y150_A5Q;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_C4 = CLBLM_R_X5Y142_SLICE_X7Y142_CQ;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_C5 = CLBLM_R_X7Y144_SLICE_X9Y144_A5Q;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_C6 = 1'b1;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_A4 = CLBLM_R_X7Y150_SLICE_X8Y150_CQ;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_A5 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_A6 = CLBLM_R_X3Y146_SLICE_X3Y146_CQ;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_D1 = CLBLM_R_X5Y148_SLICE_X6Y148_BQ;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_D2 = CLBLM_L_X12Y149_SLICE_X16Y149_CO6;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_D3 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_D4 = CLBLM_R_X7Y143_SLICE_X8Y143_BQ;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_D5 = CLBLM_L_X10Y143_SLICE_X12Y143_DO6;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_D6 = CLBLM_R_X5Y145_SLICE_X7Y145_BO6;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_SR = CLBLM_R_X7Y148_SLICE_X9Y148_AO5;
  assign LIOB33_X0Y145_IOB_X0Y146_O = CLBLL_L_X2Y148_SLICE_X1Y148_BO6;
  assign LIOB33_X0Y145_IOB_X0Y145_O = CLBLL_L_X2Y146_SLICE_X1Y146_CO6;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_C4 = 1'b1;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_C5 = CLBLM_L_X8Y152_SLICE_X10Y152_DQ;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_B1 = 1'b1;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_C6 = CLBLM_L_X10Y143_SLICE_X12Y143_BO6;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_B2 = CLBLM_L_X10Y152_SLICE_X13Y152_AQ;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_B3 = CLBLM_R_X3Y144_SLICE_X3Y144_CQ;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_B4 = CLBLM_R_X5Y142_SLICE_X7Y142_B5Q;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_A1 = 1'b1;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_A2 = 1'b1;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_A3 = CLBLM_L_X10Y147_SLICE_X13Y147_AQ;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_A5 = 1'b1;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_A6 = 1'b1;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_AX = CLBLM_R_X11Y146_SLICE_X15Y146_BO6;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_B6 = 1'b1;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_B1 = 1'b1;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_B2 = CLBLM_L_X8Y152_SLICE_X11Y152_AQ;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_B3 = 1'b1;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_B4 = 1'b1;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_B6 = 1'b1;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_C2 = 1'b1;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_C3 = CLBLM_L_X8Y152_SLICE_X11Y152_A5Q;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_C4 = 1'b1;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_C5 = 1'b1;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_C6 = 1'b1;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_A2 = CLBLM_R_X7Y149_SLICE_X8Y149_AQ;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_A3 = CLBLM_R_X7Y150_SLICE_X8Y150_AQ;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_A4 = CLBLM_R_X5Y152_SLICE_X6Y152_CQ;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_A5 = CLBLM_R_X7Y150_SLICE_X8Y150_CQ;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_A6 = 1'b1;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_AX = CLBLL_L_X2Y150_SLICE_X1Y150_BO6;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_D1 = 1'b1;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_B1 = CLBLM_R_X3Y152_SLICE_X2Y152_DO6;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_B2 = CLBLM_R_X5Y153_SLICE_X6Y153_AQ;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_B3 = 1'b1;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_B4 = CLBLM_R_X3Y151_SLICE_X3Y151_AQ;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_B5 = CLBLL_L_X4Y153_SLICE_X5Y153_BQ;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_B6 = 1'b1;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_D2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_C1 = 1'b1;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_C2 = CLBLL_L_X4Y152_SLICE_X4Y152_C5Q;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_C1 = 1'b1;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_C2 = 1'b1;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_C3 = CLBLM_R_X3Y148_SLICE_X2Y148_C5Q;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_C4 = 1'b1;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_C5 = 1'b1;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_C6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_C3 = CLBLM_L_X8Y145_SLICE_X11Y145_CO6;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_C4 = CLBLL_L_X2Y149_SLICE_X1Y149_A5Q;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_C6 = CLBLM_L_X10Y152_SLICE_X12Y152_CQ;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_D5 = CLBLM_L_X8Y148_SLICE_X10Y148_A5Q;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_C5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_A6 = CLBLM_L_X8Y152_SLICE_X11Y152_AQ;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_D6 = 1'b1;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_D1 = 1'b1;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_D2 = 1'b1;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_D3 = 1'b1;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_D4 = 1'b1;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_D5 = 1'b1;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_D6 = 1'b1;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_C6 = 1'b1;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_B5 = 1'b1;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_SR = CLBLL_L_X4Y151_SLICE_X4Y151_CO6;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_BX = CLBLL_L_X4Y152_SLICE_X4Y152_BQ;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_C2 = 1'b1;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_C3 = 1'b1;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_C4 = 1'b1;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_C5 = 1'b1;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_C6 = CLBLM_L_X10Y150_SLICE_X13Y150_A5Q;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_CE = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_CX = CLBLM_R_X11Y148_SLICE_X14Y148_BQ;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_D1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_D2 = 1'b1;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_D3 = CLBLM_L_X10Y150_SLICE_X13Y150_AQ;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_D4 = 1'b1;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_D5 = 1'b1;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_D6 = 1'b1;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_DX = CLBLM_R_X7Y151_SLICE_X8Y151_C5Q;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_A1 = CLBLL_L_X2Y148_SLICE_X0Y148_B5Q;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_A2 = CLBLM_R_X5Y149_SLICE_X7Y149_B5Q;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_A3 = CLBLL_L_X4Y151_SLICE_X5Y151_AQ;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_A5 = CLBLL_L_X4Y150_SLICE_X4Y150_AO6;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_A6 = 1'b1;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_AX = CLBLL_L_X4Y151_SLICE_X4Y151_AO6;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_B1 = CLBLL_L_X4Y152_SLICE_X5Y152_AQ;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_B2 = CLBLL_L_X4Y151_SLICE_X5Y151_BQ;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_B4 = 1'b1;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_B5 = CLBLM_L_X10Y143_SLICE_X12Y143_BO5;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_B6 = CLBLM_L_X8Y152_SLICE_X11Y152_A5Q;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_C1 = CLBLM_L_X10Y150_SLICE_X13Y150_AQ;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_C2 = CLBLM_L_X8Y151_SLICE_X10Y151_AQ;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_C3 = CLBLM_R_X3Y145_SLICE_X2Y145_DQ;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_C4 = CLBLM_R_X3Y143_SLICE_X2Y143_AQ;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_C5 = CLBLL_L_X4Y152_SLICE_X5Y152_DQ;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_C6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_D1 = CLBLM_R_X3Y143_SLICE_X2Y143_AQ;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_D2 = CLBLL_L_X4Y151_SLICE_X5Y151_CQ;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_D3 = CLBLM_R_X3Y145_SLICE_X2Y145_DQ;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_D4 = CLBLM_L_X8Y152_SLICE_X11Y152_A5Q;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_D5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_D6 = CLBLM_L_X8Y152_SLICE_X10Y152_AQ;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_B5 = CLBLL_L_X4Y151_SLICE_X5Y151_A5Q;
  assign LIOI3_SING_X0Y150_OLOGIC_X0Y150_D1 = CLBLL_L_X4Y142_SLICE_X4Y142_DO5;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_B6 = 1'b1;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_A1 = CLBLM_L_X8Y148_SLICE_X10Y148_CO6;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_A2 = CLBLM_R_X7Y146_SLICE_X8Y146_BQ;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_A3 = CLBLM_R_X7Y148_SLICE_X8Y148_AQ;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_A4 = CLBLM_L_X8Y148_SLICE_X10Y148_AQ;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_A5 = CLBLM_L_X10Y144_SLICE_X12Y144_AO6;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_A6 = 1'b1;
  assign LIOI3_SING_X0Y150_OLOGIC_X0Y150_T1 = 1'b1;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_AX = CLBLM_L_X10Y145_SLICE_X13Y145_AO6;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_B1 = CLBLM_L_X10Y143_SLICE_X12Y143_AO5;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_B2 = CLBLM_R_X7Y143_SLICE_X8Y143_CQ;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_B3 = CLBLM_R_X5Y146_SLICE_X6Y146_CO6;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_B4 = CLBLM_R_X7Y142_SLICE_X9Y142_CQ;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_B5 = CLBLM_L_X8Y144_SLICE_X11Y144_CO6;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_B6 = CLBLM_L_X10Y143_SLICE_X12Y143_DO6;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_C1 = CLBLM_L_X10Y148_SLICE_X12Y148_BO5;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_C2 = CLBLM_L_X8Y145_SLICE_X10Y145_AO5;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_C3 = CLBLM_L_X10Y145_SLICE_X13Y145_DO6;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_C4 = CLBLL_L_X4Y141_SLICE_X5Y141_A5Q;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_C5 = CLBLM_L_X8Y145_SLICE_X11Y145_DO6;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_C6 = CLBLM_L_X8Y144_SLICE_X11Y144_BO6;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_C1 = CLBLL_L_X4Y152_SLICE_X5Y152_BQ;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_C2 = CLBLM_R_X7Y149_SLICE_X9Y149_C5Q;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_D1 = CLBLL_L_X4Y145_SLICE_X5Y145_AQ;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_D2 = CLBLM_L_X8Y144_SLICE_X10Y144_DO6;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_D3 = 1'b1;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_D4 = CLBLM_L_X10Y143_SLICE_X12Y143_AO5;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_D5 = CLBLM_L_X8Y148_SLICE_X10Y148_CO6;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_D6 = CLBLM_L_X10Y149_SLICE_X12Y149_DQ;
  assign CLBLM_L_X8Y145_SLICE_X11Y145_SR = CLBLM_R_X7Y144_SLICE_X8Y144_DO6;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_A1 = CLBLM_L_X8Y142_SLICE_X10Y142_BO5;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_A2 = CLBLM_L_X8Y144_SLICE_X11Y144_AQ;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_A3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_A4 = CLBLM_R_X7Y145_SLICE_X9Y145_AQ;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_A5 = CLBLM_L_X8Y145_SLICE_X10Y145_CO5;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_A6 = 1'b1;
  assign CLBLM_L_X8Y145_SLICE_X10Y145_AX = CLBLM_R_X7Y146_SLICE_X9Y146_AO6;
endmodule
