module top(
  input LIOB33_SING_X0Y50_IOB_X0Y50_IPAD,
  input LIOB33_X0Y51_IOB_X0Y51_IPAD,
  input LIOB33_X0Y51_IOB_X0Y52_IPAD,
  input LIOB33_X0Y53_IOB_X0Y53_IPAD,
  input LIOB33_X0Y53_IOB_X0Y54_IPAD,
  input LIOB33_X0Y55_IOB_X0Y55_IPAD,
  input LIOB33_X0Y55_IOB_X0Y56_IPAD,
  input LIOB33_X0Y57_IOB_X0Y57_IPAD,
  input LIOB33_X0Y57_IOB_X0Y58_IPAD,
  input LIOB33_X0Y59_IOB_X0Y59_IPAD,
  input LIOB33_X0Y59_IOB_X0Y60_IPAD,
  input LIOB33_X0Y61_IOB_X0Y61_IPAD,
  input LIOB33_X0Y61_IOB_X0Y62_IPAD,
  input LIOB33_X0Y63_IOB_X0Y63_IPAD,
  input LIOB33_X0Y63_IOB_X0Y64_IPAD,
  input LIOB33_X0Y65_IOB_X0Y65_IPAD,
  input LIOB33_X0Y65_IOB_X0Y66_IPAD,
  input LIOB33_X0Y67_IOB_X0Y67_IPAD,
  input LIOB33_X0Y67_IOB_X0Y68_IPAD,
  input LIOB33_X0Y69_IOB_X0Y69_IPAD,
  input LIOB33_X0Y69_IOB_X0Y70_IPAD,
  input LIOB33_X0Y71_IOB_X0Y71_IPAD,
  input LIOB33_X0Y71_IOB_X0Y72_IPAD,
  input LIOB33_X0Y73_IOB_X0Y73_IPAD,
  input LIOB33_X0Y73_IOB_X0Y74_IPAD,
  input LIOB33_X0Y75_IOB_X0Y75_IPAD,
  input LIOB33_X0Y75_IOB_X0Y76_IPAD,
  input LIOB33_X0Y77_IOB_X0Y77_IPAD,
  input LIOB33_X0Y77_IOB_X0Y78_IPAD,
  input LIOB33_X0Y79_IOB_X0Y79_IPAD,
  input RIOB33_SING_X105Y100_IOB_X1Y100_IPAD,
  input RIOB33_SING_X105Y149_IOB_X1Y149_IPAD,
  input RIOB33_X105Y101_IOB_X1Y101_IPAD,
  input RIOB33_X105Y101_IOB_X1Y102_IPAD,
  input RIOB33_X105Y103_IOB_X1Y103_IPAD,
  input RIOB33_X105Y103_IOB_X1Y104_IPAD,
  input RIOB33_X105Y105_IOB_X1Y105_IPAD,
  input RIOB33_X105Y105_IOB_X1Y106_IPAD,
  input RIOB33_X105Y107_IOB_X1Y107_IPAD,
  input RIOB33_X105Y107_IOB_X1Y108_IPAD,
  input RIOB33_X105Y109_IOB_X1Y109_IPAD,
  input RIOB33_X105Y109_IOB_X1Y110_IPAD,
  input RIOB33_X105Y111_IOB_X1Y111_IPAD,
  input RIOB33_X105Y111_IOB_X1Y112_IPAD,
  input RIOB33_X105Y113_IOB_X1Y113_IPAD,
  input RIOB33_X105Y113_IOB_X1Y114_IPAD,
  input RIOB33_X105Y115_IOB_X1Y115_IPAD,
  input RIOB33_X105Y115_IOB_X1Y116_IPAD,
  input RIOB33_X105Y117_IOB_X1Y117_IPAD,
  input RIOB33_X105Y117_IOB_X1Y118_IPAD,
  input RIOB33_X105Y119_IOB_X1Y119_IPAD,
  input RIOB33_X105Y119_IOB_X1Y120_IPAD,
  input RIOB33_X105Y121_IOB_X1Y121_IPAD,
  input RIOB33_X105Y121_IOB_X1Y122_IPAD,
  input RIOB33_X105Y123_IOB_X1Y123_IPAD,
  input RIOB33_X105Y123_IOB_X1Y124_IPAD,
  input RIOB33_X105Y125_IOB_X1Y125_IPAD,
  input RIOB33_X105Y125_IOB_X1Y126_IPAD,
  input RIOB33_X105Y127_IOB_X1Y127_IPAD,
  input RIOB33_X105Y127_IOB_X1Y128_IPAD,
  input RIOB33_X105Y129_IOB_X1Y129_IPAD,
  input RIOB33_X105Y129_IOB_X1Y130_IPAD,
  input RIOB33_X105Y131_IOB_X1Y131_IPAD,
  input RIOB33_X105Y131_IOB_X1Y132_IPAD,
  input RIOB33_X105Y133_IOB_X1Y133_IPAD,
  input RIOB33_X105Y133_IOB_X1Y134_IPAD,
  input RIOB33_X105Y135_IOB_X1Y135_IPAD,
  input RIOB33_X105Y135_IOB_X1Y136_IPAD,
  input RIOB33_X105Y137_IOB_X1Y137_IPAD,
  input RIOB33_X105Y137_IOB_X1Y138_IPAD,
  input RIOB33_X105Y139_IOB_X1Y139_IPAD,
  input RIOB33_X105Y139_IOB_X1Y140_IPAD,
  input RIOB33_X105Y141_IOB_X1Y141_IPAD,
  input RIOB33_X105Y141_IOB_X1Y142_IPAD,
  input RIOB33_X105Y143_IOB_X1Y143_IPAD,
  input RIOB33_X105Y143_IOB_X1Y144_IPAD,
  input RIOB33_X105Y145_IOB_X1Y145_IPAD,
  input RIOB33_X105Y145_IOB_X1Y146_IPAD,
  input RIOB33_X105Y147_IOB_X1Y147_IPAD,
  input RIOB33_X105Y147_IOB_X1Y148_IPAD,
  output LIOB33_SING_X0Y100_IOB_X0Y100_OPAD,
  output LIOB33_SING_X0Y149_IOB_X0Y149_OPAD,
  output LIOB33_SING_X0Y150_IOB_X0Y150_OPAD,
  output LIOB33_SING_X0Y199_IOB_X0Y199_OPAD,
  output LIOB33_X0Y101_IOB_X0Y101_OPAD,
  output LIOB33_X0Y101_IOB_X0Y102_OPAD,
  output LIOB33_X0Y103_IOB_X0Y103_OPAD,
  output LIOB33_X0Y103_IOB_X0Y104_OPAD,
  output LIOB33_X0Y105_IOB_X0Y105_OPAD,
  output LIOB33_X0Y105_IOB_X0Y106_OPAD,
  output LIOB33_X0Y107_IOB_X0Y107_OPAD,
  output LIOB33_X0Y107_IOB_X0Y108_OPAD,
  output LIOB33_X0Y109_IOB_X0Y109_OPAD,
  output LIOB33_X0Y109_IOB_X0Y110_OPAD,
  output LIOB33_X0Y111_IOB_X0Y111_OPAD,
  output LIOB33_X0Y111_IOB_X0Y112_OPAD,
  output LIOB33_X0Y113_IOB_X0Y113_OPAD,
  output LIOB33_X0Y113_IOB_X0Y114_OPAD,
  output LIOB33_X0Y115_IOB_X0Y115_OPAD,
  output LIOB33_X0Y115_IOB_X0Y116_OPAD,
  output LIOB33_X0Y117_IOB_X0Y117_OPAD,
  output LIOB33_X0Y117_IOB_X0Y118_OPAD,
  output LIOB33_X0Y119_IOB_X0Y119_OPAD,
  output LIOB33_X0Y119_IOB_X0Y120_OPAD,
  output LIOB33_X0Y121_IOB_X0Y121_OPAD,
  output LIOB33_X0Y121_IOB_X0Y122_OPAD,
  output LIOB33_X0Y123_IOB_X0Y123_OPAD,
  output LIOB33_X0Y123_IOB_X0Y124_OPAD,
  output LIOB33_X0Y125_IOB_X0Y125_OPAD,
  output LIOB33_X0Y125_IOB_X0Y126_OPAD,
  output LIOB33_X0Y127_IOB_X0Y127_OPAD,
  output LIOB33_X0Y127_IOB_X0Y128_OPAD,
  output LIOB33_X0Y129_IOB_X0Y129_OPAD,
  output LIOB33_X0Y129_IOB_X0Y130_OPAD,
  output LIOB33_X0Y131_IOB_X0Y131_OPAD,
  output LIOB33_X0Y131_IOB_X0Y132_OPAD,
  output LIOB33_X0Y133_IOB_X0Y133_OPAD,
  output LIOB33_X0Y133_IOB_X0Y134_OPAD,
  output LIOB33_X0Y135_IOB_X0Y135_OPAD,
  output LIOB33_X0Y135_IOB_X0Y136_OPAD,
  output LIOB33_X0Y137_IOB_X0Y137_OPAD,
  output LIOB33_X0Y137_IOB_X0Y138_OPAD,
  output LIOB33_X0Y139_IOB_X0Y139_OPAD,
  output LIOB33_X0Y139_IOB_X0Y140_OPAD,
  output LIOB33_X0Y141_IOB_X0Y141_OPAD,
  output LIOB33_X0Y141_IOB_X0Y142_OPAD,
  output LIOB33_X0Y143_IOB_X0Y143_OPAD,
  output LIOB33_X0Y145_IOB_X0Y145_OPAD,
  output LIOB33_X0Y145_IOB_X0Y146_OPAD,
  output LIOB33_X0Y147_IOB_X0Y147_OPAD,
  output LIOB33_X0Y147_IOB_X0Y148_OPAD,
  output LIOB33_X0Y151_IOB_X0Y151_OPAD,
  output LIOB33_X0Y151_IOB_X0Y152_OPAD,
  output LIOB33_X0Y153_IOB_X0Y153_OPAD,
  output LIOB33_X0Y153_IOB_X0Y154_OPAD,
  output LIOB33_X0Y155_IOB_X0Y155_OPAD,
  output LIOB33_X0Y155_IOB_X0Y156_OPAD,
  output LIOB33_X0Y157_IOB_X0Y157_OPAD,
  output LIOB33_X0Y157_IOB_X0Y158_OPAD,
  output LIOB33_X0Y159_IOB_X0Y159_OPAD,
  output LIOB33_X0Y159_IOB_X0Y160_OPAD,
  output LIOB33_X0Y161_IOB_X0Y161_OPAD,
  output LIOB33_X0Y161_IOB_X0Y162_OPAD,
  output LIOB33_X0Y163_IOB_X0Y163_OPAD,
  output LIOB33_X0Y163_IOB_X0Y164_OPAD,
  output LIOB33_X0Y165_IOB_X0Y165_OPAD,
  output LIOB33_X0Y165_IOB_X0Y166_OPAD,
  output LIOB33_X0Y167_IOB_X0Y167_OPAD,
  output LIOB33_X0Y167_IOB_X0Y168_OPAD,
  output LIOB33_X0Y169_IOB_X0Y169_OPAD,
  output LIOB33_X0Y169_IOB_X0Y170_OPAD,
  output LIOB33_X0Y171_IOB_X0Y171_OPAD,
  output LIOB33_X0Y171_IOB_X0Y172_OPAD,
  output LIOB33_X0Y173_IOB_X0Y173_OPAD,
  output LIOB33_X0Y173_IOB_X0Y174_OPAD,
  output LIOB33_X0Y175_IOB_X0Y175_OPAD,
  output LIOB33_X0Y175_IOB_X0Y176_OPAD,
  output LIOB33_X0Y177_IOB_X0Y177_OPAD,
  output LIOB33_X0Y177_IOB_X0Y178_OPAD,
  output LIOB33_X0Y179_IOB_X0Y179_OPAD,
  output LIOB33_X0Y179_IOB_X0Y180_OPAD,
  output LIOB33_X0Y181_IOB_X0Y181_OPAD,
  output LIOB33_X0Y181_IOB_X0Y182_OPAD,
  output LIOB33_X0Y183_IOB_X0Y183_OPAD,
  output LIOB33_X0Y183_IOB_X0Y184_OPAD,
  output LIOB33_X0Y185_IOB_X0Y185_OPAD,
  output LIOB33_X0Y185_IOB_X0Y186_OPAD,
  output LIOB33_X0Y187_IOB_X0Y187_OPAD,
  output LIOB33_X0Y187_IOB_X0Y188_OPAD,
  output LIOB33_X0Y189_IOB_X0Y189_OPAD,
  output LIOB33_X0Y189_IOB_X0Y190_OPAD,
  output LIOB33_X0Y191_IOB_X0Y191_OPAD,
  output LIOB33_X0Y191_IOB_X0Y192_OPAD,
  output LIOB33_X0Y193_IOB_X0Y193_OPAD,
  output LIOB33_X0Y193_IOB_X0Y194_OPAD,
  output LIOB33_X0Y195_IOB_X0Y195_OPAD,
  output LIOB33_X0Y195_IOB_X0Y196_OPAD,
  output LIOB33_X0Y197_IOB_X0Y197_OPAD,
  output LIOB33_X0Y197_IOB_X0Y198_OPAD,
  output LIOB33_X0Y79_IOB_X0Y80_OPAD,
  output RIOB33_SING_X105Y150_IOB_X1Y150_OPAD,
  output RIOB33_SING_X105Y199_IOB_X1Y199_OPAD,
  output RIOB33_X105Y151_IOB_X1Y151_OPAD,
  output RIOB33_X105Y151_IOB_X1Y152_OPAD,
  output RIOB33_X105Y153_IOB_X1Y153_OPAD,
  output RIOB33_X105Y153_IOB_X1Y154_OPAD,
  output RIOB33_X105Y155_IOB_X1Y155_OPAD,
  output RIOB33_X105Y155_IOB_X1Y156_OPAD,
  output RIOB33_X105Y157_IOB_X1Y157_OPAD,
  output RIOB33_X105Y157_IOB_X1Y158_OPAD,
  output RIOB33_X105Y159_IOB_X1Y159_OPAD,
  output RIOB33_X105Y159_IOB_X1Y160_OPAD,
  output RIOB33_X105Y161_IOB_X1Y161_OPAD,
  output RIOB33_X105Y161_IOB_X1Y162_OPAD,
  output RIOB33_X105Y163_IOB_X1Y163_OPAD,
  output RIOB33_X105Y163_IOB_X1Y164_OPAD,
  output RIOB33_X105Y165_IOB_X1Y165_OPAD,
  output RIOB33_X105Y165_IOB_X1Y166_OPAD,
  output RIOB33_X105Y167_IOB_X1Y167_OPAD,
  output RIOB33_X105Y167_IOB_X1Y168_OPAD,
  output RIOB33_X105Y169_IOB_X1Y169_OPAD,
  output RIOB33_X105Y169_IOB_X1Y170_OPAD,
  output RIOB33_X105Y171_IOB_X1Y171_OPAD,
  output RIOB33_X105Y171_IOB_X1Y172_OPAD,
  output RIOB33_X105Y173_IOB_X1Y173_OPAD,
  output RIOB33_X105Y173_IOB_X1Y174_OPAD,
  output RIOB33_X105Y175_IOB_X1Y175_OPAD,
  output RIOB33_X105Y175_IOB_X1Y176_OPAD,
  output RIOB33_X105Y177_IOB_X1Y177_OPAD,
  output RIOB33_X105Y177_IOB_X1Y178_OPAD,
  output RIOB33_X105Y179_IOB_X1Y179_OPAD,
  output RIOB33_X105Y179_IOB_X1Y180_OPAD,
  output RIOB33_X105Y181_IOB_X1Y181_OPAD,
  output RIOB33_X105Y181_IOB_X1Y182_OPAD,
  output RIOB33_X105Y183_IOB_X1Y183_OPAD,
  output RIOB33_X105Y183_IOB_X1Y184_OPAD,
  output RIOB33_X105Y185_IOB_X1Y185_OPAD,
  output RIOB33_X105Y185_IOB_X1Y186_OPAD,
  output RIOB33_X105Y187_IOB_X1Y187_OPAD,
  output RIOB33_X105Y187_IOB_X1Y188_OPAD,
  output RIOB33_X105Y189_IOB_X1Y189_OPAD,
  output RIOB33_X105Y189_IOB_X1Y190_OPAD,
  output RIOB33_X105Y191_IOB_X1Y191_OPAD,
  output RIOB33_X105Y191_IOB_X1Y192_OPAD,
  output RIOB33_X105Y193_IOB_X1Y193_OPAD,
  output RIOB33_X105Y193_IOB_X1Y194_OPAD,
  output RIOB33_X105Y195_IOB_X1Y195_OPAD,
  output RIOB33_X105Y195_IOB_X1Y196_OPAD,
  output RIOB33_X105Y197_IOB_X1Y197_OPAD,
  output RIOB33_X105Y197_IOB_X1Y198_OPAD
  );
  wire [0:0] CLBLL_L_X26Y136_SLICE_X38Y136_A;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X38Y136_A1;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X38Y136_A2;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X38Y136_A3;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X38Y136_A4;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X38Y136_A5;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X38Y136_A6;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X38Y136_AMUX;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X38Y136_AO5;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X38Y136_AO6;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X38Y136_A_CY;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X38Y136_A_XOR;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X38Y136_B;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X38Y136_B1;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X38Y136_B2;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X38Y136_B3;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X38Y136_B4;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X38Y136_B5;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X38Y136_B6;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X38Y136_BO5;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X38Y136_BO6;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X38Y136_B_CY;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X38Y136_B_XOR;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X38Y136_C;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X38Y136_C1;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X38Y136_C2;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X38Y136_C3;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X38Y136_C4;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X38Y136_C5;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X38Y136_C6;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X38Y136_CO5;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X38Y136_CO6;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X38Y136_C_CY;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X38Y136_C_XOR;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X38Y136_D;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X38Y136_D1;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X38Y136_D2;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X38Y136_D3;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X38Y136_D4;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X38Y136_D5;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X38Y136_D6;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X38Y136_DO5;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X38Y136_DO6;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X38Y136_D_CY;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X38Y136_D_XOR;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X39Y136_A;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X39Y136_A1;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X39Y136_A2;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X39Y136_A3;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X39Y136_A4;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X39Y136_A5;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X39Y136_A6;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X39Y136_AO5;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X39Y136_AO6;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X39Y136_A_CY;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X39Y136_A_XOR;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X39Y136_B;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X39Y136_B1;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X39Y136_B2;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X39Y136_B3;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X39Y136_B4;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X39Y136_B5;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X39Y136_B6;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X39Y136_BO5;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X39Y136_BO6;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X39Y136_B_CY;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X39Y136_B_XOR;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X39Y136_C;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X39Y136_C1;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X39Y136_C2;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X39Y136_C3;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X39Y136_C4;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X39Y136_C5;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X39Y136_C6;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X39Y136_CO5;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X39Y136_CO6;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X39Y136_C_CY;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X39Y136_C_XOR;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X39Y136_D;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X39Y136_D1;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X39Y136_D2;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X39Y136_D3;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X39Y136_D4;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X39Y136_D5;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X39Y136_D6;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X39Y136_DO5;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X39Y136_DO6;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X39Y136_D_CY;
  wire [0:0] CLBLL_L_X26Y136_SLICE_X39Y136_D_XOR;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_A;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_A1;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_A2;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_A3;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_A4;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_A5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_A6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_AMUX;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_AO5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_AO6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_A_CY;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_A_XOR;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_B;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_B1;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_B2;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_B3;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_B4;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_B5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_B6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_BMUX;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_BO5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_BO6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_B_CY;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_B_XOR;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_C;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_C1;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_C2;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_C3;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_C4;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_C5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_C6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_CMUX;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_CO5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_CO6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_C_CY;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_C_XOR;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_D;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_D1;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_D2;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_D3;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_D4;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_D5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_D6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_DO5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_DO6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_D_CY;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_D_XOR;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_A;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_A1;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_A2;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_A3;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_A4;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_A5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_A6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_AO5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_AO6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_A_CY;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_A_XOR;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_B;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_B1;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_B2;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_B3;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_B4;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_B5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_B6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_BO5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_BO6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_B_CY;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_B_XOR;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_C;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_C1;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_C2;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_C3;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_C4;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_C5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_C6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_CO5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_CO6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_C_CY;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_C_XOR;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_D;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_D1;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_D2;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_D3;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_D4;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_D5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_D6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_DO5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_DO6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_D_CY;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_D_XOR;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_A;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_A1;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_A2;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_A3;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_A4;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_A5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_A6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_AMUX;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_AO5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_AO6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_A_CY;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_A_XOR;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_B;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_B1;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_B2;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_B3;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_B4;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_B5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_B6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_BO5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_BO6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_B_CY;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_B_XOR;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_C;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_C1;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_C2;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_C3;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_C4;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_C5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_C6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_CO5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_CO6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_C_CY;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_C_XOR;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_D;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_D1;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_D2;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_D3;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_D4;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_D5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_D6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_DO5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_DO6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_D_CY;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_D_XOR;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_A;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_A1;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_A2;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_A3;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_A4;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_A5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_A6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_AMUX;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_AO5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_AO6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_A_CY;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_A_XOR;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_B;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_B1;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_B2;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_B3;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_B4;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_B5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_B6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_BO5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_BO6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_B_CY;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_B_XOR;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_C;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_C1;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_C2;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_C3;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_C4;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_C5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_C6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_CO5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_CO6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_C_CY;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_C_XOR;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_D;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_D1;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_D2;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_D3;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_D4;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_D5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_D6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_DO5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_DO6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_D_CY;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_D_XOR;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_A;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_A1;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_A2;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_A3;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_A4;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_A5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_A6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_AO5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_AO6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_A_CY;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_A_XOR;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_B;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_B1;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_B2;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_B3;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_B4;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_B5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_B6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_BO5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_BO6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_B_CY;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_B_XOR;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_C;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_C1;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_C2;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_C3;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_C4;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_C5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_C6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_CO5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_CO6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_C_CY;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_C_XOR;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_D;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_D1;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_D2;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_D3;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_D4;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_D5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_D6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_DO5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_DO6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_D_CY;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_D_XOR;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_A;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_A1;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_A2;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_A3;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_A4;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_A5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_A6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_AMUX;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_AO5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_AO6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_A_CY;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_A_XOR;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_B;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_B1;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_B2;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_B3;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_B4;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_B5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_B6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_BMUX;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_BO5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_BO6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_B_CY;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_B_XOR;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_C;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_C1;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_C2;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_C3;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_C4;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_C5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_C6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_CMUX;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_CO5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_CO6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_C_CY;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_C_XOR;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_D;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_D1;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_D2;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_D3;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_D4;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_D5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_D6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_DO5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_DO6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_D_CY;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_D_XOR;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A1;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A2;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A3;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A4;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_AMUX;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_AO5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_AO6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A_CY;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A_XOR;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B1;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B2;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B3;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B4;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_BMUX;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_BO5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_BO6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B_CY;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B_XOR;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C1;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C2;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C3;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C4;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_CMUX;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_CO5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_CO6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C_CY;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C_XOR;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D1;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D2;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D3;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D4;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_DO5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_DO6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D_CY;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D_XOR;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A1;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A2;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A3;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A4;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_AO5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_AO6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A_CY;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A_XOR;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B1;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B2;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B3;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B4;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_BMUX;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_BO5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_BO6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B_CY;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B_XOR;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C1;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C2;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C3;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C4;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_CO5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_CO6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C_CY;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C_XOR;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D1;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D2;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D3;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D4;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_DMUX;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_DO5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_DO6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D_CY;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D_XOR;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A1;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A2;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A3;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A4;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_AMUX;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_AO5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_AO6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A_CY;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A_XOR;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B1;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B2;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B3;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B4;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_BMUX;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_BO5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_BO6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B_CY;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B_XOR;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C1;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C2;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C3;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C4;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_CMUX;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_CO5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_CO6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C_CY;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C_XOR;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D1;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D2;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D3;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D4;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_DO5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_DO6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D_CY;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D_XOR;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A1;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A2;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A3;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A4;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_AMUX;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_AO5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_AO6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A_CY;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A_XOR;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B1;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B2;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B3;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B4;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_BO5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_BO6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B_CY;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B_XOR;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C1;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C2;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C3;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C4;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_CMUX;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_CO5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_CO6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C_CY;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C_XOR;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D1;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D2;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D3;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D4;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_DO5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_DO6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D_CY;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D_XOR;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_A;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_A1;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_A2;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_A3;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_A4;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_A5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_A6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_AO5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_AO6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_A_CY;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_A_XOR;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_B;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_B1;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_B2;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_B3;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_B4;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_B5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_B6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_BMUX;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_BO5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_BO6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_B_CY;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_B_XOR;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_C;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_C1;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_C2;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_C3;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_C4;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_C5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_C6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_CO5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_CO6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_C_CY;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_C_XOR;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_D;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_D1;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_D2;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_D3;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_D4;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_D5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_D6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_DO5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_DO6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_D_CY;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_D_XOR;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_A;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_A1;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_A2;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_A3;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_A4;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_A5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_A6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_AMUX;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_AO5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_AO6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_A_CY;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_A_XOR;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_B;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_B1;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_B2;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_B3;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_B4;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_B5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_B6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_BMUX;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_BO5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_BO6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_B_CY;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_B_XOR;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_C;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_C1;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_C2;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_C3;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_C4;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_C5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_C6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_CO5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_CO6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_C_CY;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_C_XOR;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_D;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_D1;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_D2;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_D3;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_D4;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_D5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_D6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_DO5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_DO6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_D_CY;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_D_XOR;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_A;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_A1;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_A2;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_A3;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_A4;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_A5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_A6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_AMUX;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_AO5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_AO6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_A_CY;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_A_XOR;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_B;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_B1;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_B2;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_B3;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_B4;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_B5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_B6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_BO5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_BO6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_B_CY;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_B_XOR;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_C;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_C1;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_C2;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_C3;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_C4;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_C5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_C6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_CO5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_CO6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_C_CY;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_C_XOR;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_D;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_D1;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_D2;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_D3;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_D4;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_D5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_D6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_DO5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_DO6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_D_CY;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_D_XOR;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_A;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_A1;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_A2;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_A3;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_A4;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_A5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_A6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_AO5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_AO6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_A_CY;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_A_XOR;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_B;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_B1;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_B2;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_B3;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_B4;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_B5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_B6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_BO5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_BO6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_B_CY;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_B_XOR;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_C;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_C1;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_C2;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_C3;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_C4;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_C5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_C6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_CO5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_CO6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_C_CY;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_C_XOR;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_D;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_D1;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_D2;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_D3;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_D4;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_D5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_D6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_DO5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_DO6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_D_CY;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_D_XOR;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A1;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A2;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A3;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A4;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_AO5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_AO6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A_CY;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A_XOR;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B1;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B2;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B3;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B4;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_BO5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_BO6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B_CY;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B_XOR;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C1;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C2;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C3;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C4;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_CO5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_CO6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C_CY;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C_XOR;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D1;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D2;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D3;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D4;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_DO5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_DO6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D_CY;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D_XOR;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A1;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A2;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A3;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A4;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_AMUX;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_AO5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_AO6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A_CY;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A_XOR;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B1;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B2;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B3;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B4;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_BO5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_BO6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B_CY;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B_XOR;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C1;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C2;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C3;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C4;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_CMUX;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_CO5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_CO6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C_CY;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C_XOR;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D1;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D2;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D3;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D4;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_DO5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_DO6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D_CY;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D_XOR;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_A;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_A1;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_A2;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_A3;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_A4;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_A5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_A6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_AMUX;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_AO5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_AO6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_A_CY;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_A_XOR;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_B;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_B1;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_B2;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_B3;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_B4;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_B5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_B6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_BO5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_BO6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_B_CY;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_B_XOR;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_C;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_C1;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_C2;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_C3;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_C4;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_C5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_C6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_CO5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_CO6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_C_CY;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_C_XOR;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_D;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_D1;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_D2;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_D3;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_D4;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_D5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_D6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_DO5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_DO6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_D_CY;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X0Y114_D_XOR;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_A;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_A1;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_A2;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_A3;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_A4;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_A5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_A6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_AMUX;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_AO5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_AO6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_A_CY;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_A_XOR;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_B;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_B1;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_B2;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_B3;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_B4;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_B5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_B6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_BO5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_BO6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_B_CY;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_B_XOR;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_C;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_C1;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_C2;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_C3;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_C4;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_C5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_C6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_CO5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_CO6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_C_CY;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_C_XOR;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_D;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_D1;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_D2;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_D3;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_D4;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_D5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_D6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_DO5;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_DO6;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_D_CY;
  wire [0:0] CLBLL_L_X2Y114_SLICE_X1Y114_D_XOR;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_A;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_A1;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_A2;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_A3;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_A4;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_A5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_A6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_AO5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_AO6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_A_CY;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_A_XOR;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_B;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_B1;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_B2;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_B3;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_B4;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_B5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_B6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_BO5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_BO6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_B_CY;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_B_XOR;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_C;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_C1;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_C2;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_C3;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_C4;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_C5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_C6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_CO5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_CO6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_C_CY;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_C_XOR;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_D;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_D1;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_D2;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_D3;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_D4;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_D5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_D6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_DO5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_DO6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_D_CY;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_D_XOR;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_A;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_A1;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_A2;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_A3;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_A4;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_A5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_A6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_AO5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_AO6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_AQ;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_A_CY;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_A_XOR;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_B;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_B1;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_B2;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_B3;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_B4;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_B5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_B6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_BO5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_BO6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_BQ;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_B_CY;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_B_XOR;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_C;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_C1;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_C2;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_C3;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_C4;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_C5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_C6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_CLK;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_CO5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_CO6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_C_CY;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_C_XOR;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_D;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_D1;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_D2;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_D3;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_D4;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_D5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_D6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_DO5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_DO6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_D_CY;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_D_XOR;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A1;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A2;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A3;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A4;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A5Q;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_AMUX;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_AO5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_AO6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_AQ;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_AX;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A_CY;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A_XOR;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B1;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B2;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B3;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B4;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_BMUX;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_BO5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_BO6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B_CY;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B_XOR;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C1;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C2;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C3;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C4;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_CLK;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_CO5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_CO6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_CQ;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C_CY;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C_XOR;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D1;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D2;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D3;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D4;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_DO5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_DO6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_DQ;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D_CY;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D_XOR;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A1;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A2;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A3;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A4;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_AO5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_AO6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_AQ;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A_CY;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A_XOR;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B1;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B2;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B3;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B4;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_BMUX;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_BO5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_BO6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B_CY;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B_XOR;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C1;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C2;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C3;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C4;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_CLK;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_CO5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_CO6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C_CY;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C_XOR;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D1;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D2;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D3;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D4;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_DO5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_DO6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D_CY;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D_XOR;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A1;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A2;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A3;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A4;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_AO5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_AO6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_AQ;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A_CY;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A_XOR;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B1;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B2;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B3;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B4;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_BO5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_BO6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_BQ;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B_CY;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B_XOR;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C1;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C2;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C3;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C4;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_CLK;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_CO5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_CO6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C_CY;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C_XOR;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D1;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D2;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D3;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D4;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_DO5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_DO6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D_CY;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D_XOR;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A1;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A2;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A3;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A4;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_AMUX;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_AO5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_AO6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A_CY;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A_XOR;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B1;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B2;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B3;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B4;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_BO5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_BO6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B_CY;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B_XOR;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C1;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C2;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C3;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C4;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_CO5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_CO6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C_CY;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C_XOR;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D1;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D2;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D3;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D4;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_DO5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_DO6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D_CY;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_AO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_AO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_AQ;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_BO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_BO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_BQ;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_CLK;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_CO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_CO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_DO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_DO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_AO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_AO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_AQ;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_BMUX;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_BO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_BO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_CLK;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_CO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_CO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_DO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_DO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D_XOR;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A1;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A2;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A3;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A4;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_AO5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_AO6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_AQ;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A_CY;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A_XOR;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B1;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B2;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B3;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B4;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B5Q;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_BMUX;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_BO5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_BO6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_BQ;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B_CY;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B_XOR;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C1;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C2;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C3;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C4;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C5Q;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_CLK;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_CMUX;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_CO5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_CO6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_CQ;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C_CY;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C_XOR;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D1;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D2;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D3;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D4;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_DO5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_DO6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D_CY;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D_XOR;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A1;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A2;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A3;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A4;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_AO5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_AO6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_AQ;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_AX;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A_CY;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A_XOR;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B1;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B2;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B3;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B4;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_BO5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_BO6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B_CY;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B_XOR;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C1;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C2;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C3;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C4;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_CLK;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_CMUX;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_CO5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_CO6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C_CY;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C_XOR;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D1;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D2;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D3;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D4;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_DMUX;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_DO5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_DO6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D_CY;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D_XOR;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A1;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A2;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A3;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A4;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_AO5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_AO6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_AQ;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A_CY;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A_XOR;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B1;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B2;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B3;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B4;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_BO5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_BO6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_BQ;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B_CY;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B_XOR;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C1;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C2;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C3;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C4;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_CLK;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_CO5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_CO6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_CQ;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C_CY;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C_XOR;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D1;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D2;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D3;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D4;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_DO5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_DO6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D_CY;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D_XOR;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A1;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A2;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A3;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A4;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_AO5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_AO6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_AQ;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A_CY;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A_XOR;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B1;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B2;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B3;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B4;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_BO5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_BO6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B_CY;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B_XOR;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C1;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C2;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C3;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C4;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_CLK;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_CO5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_CO6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C_CY;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C_XOR;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D1;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D2;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D3;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D4;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_DO5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_DO6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D_CY;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_AO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_AO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_BO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_BO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_BQ;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_CLK;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_CMUX;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_CO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_CO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_DO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_DO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_AO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_AO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_AQ;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_BMUX;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_BO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_BO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_CLK;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_CO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_CO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_DO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_DO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_AO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_AO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_AQ;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_BO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_BO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_BQ;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_CLK;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_CMUX;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_CO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_CO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_DO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_DO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_AO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_AO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_AQ;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B5Q;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_BMUX;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_BO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_BO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_BQ;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_CLK;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_CO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_CO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_DO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_DO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D_XOR;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A1;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A2;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A3;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A4;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_AO5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_AO6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_AQ;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A_CY;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A_XOR;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B1;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B2;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B3;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B4;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_BO5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_BO6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_BQ;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B_CY;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B_XOR;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C1;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C2;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C3;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C4;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_CLK;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_CO5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_CO6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_CQ;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C_CY;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C_XOR;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D1;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D2;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D3;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D4;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_DO5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_DO6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D_CY;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D_XOR;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A1;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A2;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A3;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A4;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_AO5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_AO6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_AQ;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A_CY;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A_XOR;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B1;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B2;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B3;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B4;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_BO5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_BO6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B_CY;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B_XOR;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C1;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C2;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C3;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C4;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_CLK;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_CO5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_CO6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C_CY;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C_XOR;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D1;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D2;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D3;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D4;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_DO5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_DO6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D_CY;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_AO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_AO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_BO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_BO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_CO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_CO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_DO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_DO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A5Q;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_AMUX;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_AO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_AO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_AQ;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_BO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_BO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_BQ;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_CLK;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_CO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_CO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_CQ;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_DO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_DO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D_XOR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A1;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A2;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A3;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A4;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A5Q;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_AMUX;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_AO5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_AO6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_AQ;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_AX;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A_CY;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_A_XOR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B1;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B2;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B3;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B4;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_BMUX;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_BO5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_BO6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B_CY;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_B_XOR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C1;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C2;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C3;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C4;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_CLK;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_CO5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_CO6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C_CY;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_C_XOR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D1;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D2;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D3;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D4;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_DO5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_DO6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D_CY;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X4Y116_D_XOR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A1;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A2;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A3;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A4;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A5Q;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_AMUX;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_AO5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_AO6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_AQ;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_AX;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A_CY;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_A_XOR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B1;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B2;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B3;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B4;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B5Q;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_BMUX;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_BO5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_BO6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_BQ;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B_CY;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_B_XOR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C1;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C2;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C3;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C4;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_CLK;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_CO5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_CO6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C_CY;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_C_XOR;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D1;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D2;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D3;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D4;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_DO5;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_DO6;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D_CY;
  wire [0:0] CLBLL_L_X4Y116_SLICE_X5Y116_D_XOR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A1;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A2;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A3;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A4;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_AO5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_AO6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_AQ;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A_CY;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A_XOR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B1;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B2;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B3;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B4;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_BO5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_BO6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_BQ;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B_CY;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B_XOR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C1;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C2;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C3;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C4;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_CLK;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_CO5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_CO6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_CQ;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C_CY;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C_XOR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D1;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D2;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D3;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D4;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_DO5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_DO6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_DQ;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D_CY;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D_XOR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A1;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A2;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A3;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A4;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_AO5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_AO6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_AQ;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A_CY;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A_XOR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B1;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B2;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B3;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B4;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_BMUX;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_BO5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_BO6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B_CY;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B_XOR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C1;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C2;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C3;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C4;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_CLK;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_CO5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_CO6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C_CY;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C_XOR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D1;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D2;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D3;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D4;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_DO5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_DO6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D_CY;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D_XOR;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_A;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_A1;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_A2;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_A3;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_A4;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_A5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_A5Q;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_A6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_AMUX;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_AO5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_AO6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_AQ;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_AX;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_A_CY;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_A_XOR;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_B;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_B1;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_B2;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_B3;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_B4;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_B5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_B6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_BO5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_BO6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_BQ;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_B_CY;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_B_XOR;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_C;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_C1;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_C2;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_C3;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_C4;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_C5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_C6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_CLK;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_CMUX;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_CO5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_CO6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_C_CY;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_C_XOR;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_D;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_D1;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_D2;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_D3;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_D4;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_D5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_D6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_DMUX;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_DO5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_DO6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_D_CY;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_D_XOR;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_A;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_A1;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_A2;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_A3;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_A4;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_A5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_A6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_AO5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_AO6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_A_CY;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_A_XOR;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_B;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_B1;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_B2;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_B3;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_B4;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_B5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_B6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_BO5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_BO6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_B_CY;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_B_XOR;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_C;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_C1;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_C2;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_C3;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_C4;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_C5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_C6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_CO5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_CO6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_C_CY;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_C_XOR;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_D;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_D1;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_D2;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_D3;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_D4;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_D5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_D6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_DO5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_DO6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_D_CY;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_D_XOR;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A1;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A2;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A3;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A4;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_AO5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_AO6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A_CY;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A_XOR;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B1;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B2;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B3;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B4;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_BO5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_BO6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B_CY;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B_XOR;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C1;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C2;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C3;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C4;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_CO5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_CO6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C_CY;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C_XOR;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D1;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D2;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D3;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D4;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_DO5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_DO6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D_CY;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D_XOR;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A1;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A2;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A3;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A4;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_AO5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_AO6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A_CY;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A_XOR;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B1;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B2;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B3;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B4;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_BO5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_BO6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B_CY;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B_XOR;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C1;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C2;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C3;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C4;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_CO5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_CO6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C_CY;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C_XOR;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D1;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D2;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D3;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D4;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_DO5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_DO6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D_CY;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D_XOR;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_A;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_A1;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_A2;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_A3;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_A4;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_A5;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_A6;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_AO5;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_AO6;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_AQ;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_A_CY;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_A_XOR;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_B;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_B1;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_B2;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_B3;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_B4;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_B5;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_B6;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_BO5;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_BO6;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_B_CY;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_B_XOR;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_C;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_C1;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_C2;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_C3;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_C4;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_C5;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_C6;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_CLK;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_CO5;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_CO6;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_C_CY;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_C_XOR;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_D;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_D1;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_D2;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_D3;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_D4;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_D5;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_D6;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_DO5;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_DO6;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_D_CY;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_D_XOR;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_A;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_A1;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_A2;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_A3;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_A4;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_A5;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_A6;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_AO5;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_AO6;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_A_CY;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_A_XOR;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_B;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_B1;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_B2;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_B3;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_B4;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_B5;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_B6;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_BO5;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_BO6;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_B_CY;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_B_XOR;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_C;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_C1;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_C2;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_C3;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_C4;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_C5;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_C6;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_CO5;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_CO6;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_C_CY;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_C_XOR;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_D;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_D1;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_D2;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_D3;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_D4;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_D5;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_D6;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_DO5;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_DO6;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_D_CY;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_D_XOR;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_A;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_A1;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_A2;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_A3;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_A4;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_A5;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_A6;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_AO5;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_AO6;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_AQ;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_A_CY;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_A_XOR;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_B;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_B1;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_B2;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_B3;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_B4;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_B5;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_B6;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_BO5;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_BO6;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_BQ;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_B_CY;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_B_XOR;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_C;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_C1;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_C2;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_C3;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_C4;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_C5;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_C6;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_CLK;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_CMUX;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_CO5;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_CO6;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_C_CY;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_C_XOR;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_D;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_D1;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_D2;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_D3;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_D4;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_D5;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_D6;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_DO5;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_DO6;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_D_CY;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_D_XOR;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_A;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_A1;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_A2;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_A3;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_A4;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_A5;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_A6;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_AO5;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_AO6;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_A_CY;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_A_XOR;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_B;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_B1;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_B2;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_B3;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_B4;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_B5;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_B6;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_BO5;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_BO6;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_B_CY;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_B_XOR;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_C;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_C1;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_C2;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_C3;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_C4;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_C5;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_C6;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_CO5;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_CO6;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_C_CY;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_C_XOR;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_D;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_D1;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_D2;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_D3;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_D4;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_D5;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_D6;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_DO5;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_DO6;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_D_CY;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_D_XOR;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_A;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_A1;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_A2;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_A3;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_A4;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_A5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_A6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_AO5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_AO6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_AQ;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_A_CY;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_A_XOR;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_B;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_B1;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_B2;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_B3;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_B4;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_B5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_B6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_BMUX;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_BO5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_BO6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_B_CY;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_B_XOR;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_C;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_C1;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_C2;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_C3;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_C4;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_C5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_C6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_CLK;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_CO5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_CO6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_C_CY;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_C_XOR;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_D;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_D1;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_D2;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_D3;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_D4;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_D5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_D6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_DO5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_DO6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_D_CY;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_D_XOR;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_A;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_A1;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_A2;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_A3;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_A4;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_A5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_A6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_AO5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_AO6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_AQ;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_A_CY;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_A_XOR;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_B;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_B1;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_B2;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_B3;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_B4;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_B5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_B6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_BO5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_BO6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_BQ;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_B_CY;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_B_XOR;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_C;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_C1;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_C2;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_C3;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_C4;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_C5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_C6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_CLK;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_CO5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_CO6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_CQ;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_C_CY;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_C_XOR;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_D;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_D1;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_D2;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_D3;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_D4;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_D5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_D6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_DO5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_DO6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_D_CY;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_D_XOR;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_A;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_A1;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_A2;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_A3;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_A4;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_A5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_A6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_AO5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_AO6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_AQ;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_A_CY;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_A_XOR;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_B;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_B1;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_B2;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_B3;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_B4;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_B5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_B6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_BO5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_BO6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_BQ;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_B_CY;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_B_XOR;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_C;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_C1;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_C2;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_C3;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_C4;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_C5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_C6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_CLK;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_CO5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_CO6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_C_CY;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_C_XOR;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_D;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_D1;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_D2;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_D3;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_D4;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_D5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_D6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_DMUX;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_DO5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_DO6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_D_CY;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_D_XOR;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_A;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_A1;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_A2;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_A3;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_A4;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_A5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_A6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_AO5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_AO6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_AQ;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_A_CY;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_A_XOR;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_B;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_B1;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_B2;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_B3;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_B4;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_B5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_B6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_BO5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_BO6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_B_CY;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_B_XOR;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_C;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_C1;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_C2;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_C3;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_C4;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_C5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_C6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_CLK;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_CO5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_CO6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_C_CY;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_C_XOR;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_D;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_D1;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_D2;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_D3;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_D4;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_D5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_D6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_DO5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_DO6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_D_CY;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_D_XOR;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_A;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_A1;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_A2;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_A3;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_A4;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_A5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_A6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_AMUX;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_AO5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_AO6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_A_CY;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_A_XOR;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_B;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_B1;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_B2;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_B3;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_B4;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_B5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_B6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_BO5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_BO6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_BQ;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_B_CY;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_B_XOR;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_C;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_C1;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_C2;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_C3;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_C4;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_C5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_C6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_CLK;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_CO5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_CO6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_CQ;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_C_CY;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_C_XOR;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_D;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_D1;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_D2;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_D3;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_D4;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_D5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_D6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_DO5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_DO6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_D_CY;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_D_XOR;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_A;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_A1;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_A2;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_A3;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_A4;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_A5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_A6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_AO5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_AO6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_AQ;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_A_CY;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_A_XOR;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_B;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_B1;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_B2;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_B3;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_B4;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_B5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_B6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_BO5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_BO6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_B_CY;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_B_XOR;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_C;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_C1;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_C2;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_C3;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_C4;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_C5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_C6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_CLK;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_CO5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_CO6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_C_CY;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_C_XOR;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_D;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_D1;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_D2;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_D3;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_D4;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_D5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_D6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_DO5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_DO6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_D_CY;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_D_XOR;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_A;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_A1;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_A2;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_A3;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_A4;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_A5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_A6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_AO5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_AO6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_AQ;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_A_CY;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_A_XOR;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_B;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_B1;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_B2;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_B3;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_B4;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_B5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_B6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_BO5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_BO6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_BQ;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_B_CY;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_B_XOR;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_C;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_C1;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_C2;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_C3;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_C4;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_C5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_C6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_CLK;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_CMUX;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_CO5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_CO6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_C_CY;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_C_XOR;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_D;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_D1;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_D2;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_D3;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_D4;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_D5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_D6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_DO5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_DO6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_D_CY;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_D_XOR;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_A;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_A1;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_A2;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_A3;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_A4;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_A5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_A6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_AMUX;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_AO5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_AO6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_A_CY;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_A_XOR;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_B;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_B1;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_B2;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_B3;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_B4;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_B5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_B6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_BMUX;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_BO5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_BO6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_B_CY;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_B_XOR;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_C;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_C1;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_C2;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_C3;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_C4;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_C5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_C6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_CO5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_CO6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_C_CY;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_C_XOR;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_D;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_D1;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_D2;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_D3;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_D4;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_D5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_D6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_DMUX;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_DO5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_DO6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_D_CY;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_D_XOR;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_A;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_A1;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_A2;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_A3;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_A4;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_A5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_A6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_AO5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_AO6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_AQ;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_A_CY;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_A_XOR;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_B;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_B1;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_B2;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_B3;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_B4;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_B5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_B5Q;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_B6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_BMUX;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_BO5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_BO6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_BQ;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_B_CY;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_B_XOR;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_C;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_C1;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_C2;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_C3;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_C4;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_C5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_C6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_CLK;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_CMUX;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_CO5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_CO6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_C_CY;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_C_XOR;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_D;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_D1;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_D2;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_D3;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_D4;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_D5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_D6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_DO5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_DO6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_D_CY;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_D_XOR;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_A;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_A1;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_A2;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_A3;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_A4;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_A5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_A6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_AO5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_AO6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_AQ;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_A_CY;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_A_XOR;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_B;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_B1;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_B2;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_B3;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_B4;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_B5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_B6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_BO5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_BO6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_BQ;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_B_CY;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_B_XOR;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_C;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_C1;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_C2;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_C3;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_C4;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_C5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_C6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_CLK;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_CO5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_CO6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_CQ;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_C_CY;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_C_XOR;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_D;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_D1;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_D2;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_D3;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_D4;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_D5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_D6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_DO5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_DO6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_DQ;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_D_CY;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_D_XOR;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_A;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_A1;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_A2;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_A3;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_A4;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_A5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_A5Q;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_A6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_AMUX;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_AO5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_AO6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_AQ;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_AX;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_A_CY;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_A_XOR;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_B;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_B1;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_B2;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_B3;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_B4;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_B5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_B6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_BO5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_BO6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_BQ;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_B_CY;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_B_XOR;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_C;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_C1;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_C2;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_C3;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_C4;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_C5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_C5Q;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_C6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_CLK;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_CMUX;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_CO5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_CO6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_CQ;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_C_CY;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_C_XOR;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_D;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_D1;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_D2;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_D3;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_D4;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_D5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_D6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_DO5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_DO6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_DQ;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_D_CY;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_D_XOR;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_A;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_A1;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_A2;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_A3;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_A4;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_A5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_A6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_AO5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_AO6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_AQ;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_A_CY;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_A_XOR;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_B;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_B1;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_B2;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_B3;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_B4;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_B5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_B6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_BO5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_BO6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_BQ;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_B_CY;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_B_XOR;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_C;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_C1;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_C2;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_C3;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_C4;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_C5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_C5Q;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_C6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_CLK;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_CMUX;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_CO5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_CO6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_CQ;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_C_CY;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_C_XOR;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_D;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_D1;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_D2;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_D3;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_D4;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_D5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_D6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_DO5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_DO6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_D_CY;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_D_XOR;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_A;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_A1;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_A2;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_A3;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_A4;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_A5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_A6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_AO5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_AO6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_AQ;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_A_CY;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_A_XOR;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_B;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_B1;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_B2;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_B3;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_B4;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_B5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_B6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_BO5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_BO6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_BQ;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_B_CY;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_B_XOR;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_C;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_C1;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_C2;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_C3;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_C4;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_C5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_C5Q;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_C6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_CLK;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_CMUX;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_CO5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_CO6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_CQ;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_C_CY;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_C_XOR;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_D;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_D1;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_D2;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_D3;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_D4;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_D5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_D6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_DO5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_DO6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_D_CY;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_D_XOR;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_A;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_A1;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_A2;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_A3;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_A4;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_A5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_A6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_AO5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_AO6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_AQ;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_AX;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_A_CY;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_A_XOR;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_B;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_B1;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_B2;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_B3;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_B4;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_B5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_B6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_BO5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_BO6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_B_CY;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_B_XOR;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_C;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_C1;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_C2;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_C3;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_C4;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_C5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_C6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_CE;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_CLK;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_CO5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_CO6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_C_CY;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_C_XOR;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_D;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_D1;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_D2;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_D3;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_D4;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_D5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_D6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_DO5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_DO6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_D_CY;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_D_XOR;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_SR;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_A;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_A1;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_A2;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_A3;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_A4;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_A5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_A6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_AO5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_AO6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_AQ;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_A_CY;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_A_XOR;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_B;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_B1;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_B2;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_B3;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_B4;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_B5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_B6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_BO5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_BO6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_BQ;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_B_CY;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_B_XOR;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_C;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_C1;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_C2;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_C3;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_C4;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_C5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_C6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_CLK;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_CO5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_CO6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_CQ;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_C_CY;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_C_XOR;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_D;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_D1;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_D2;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_D3;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_D4;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_D5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_D6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_DMUX;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_DO5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_DO6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_D_CY;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_D_XOR;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_A;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_A1;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_A2;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_A3;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_A4;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_A5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_A6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_AO5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_AO6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_AQ;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_A_CY;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_A_XOR;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_B;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_B1;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_B2;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_B3;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_B4;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_B5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_B6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_BO5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_BO6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_BQ;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_B_CY;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_B_XOR;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_C;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_C1;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_C2;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_C3;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_C4;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_C5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_C5Q;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_C6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_CLK;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_CMUX;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_CO5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_CO6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_CQ;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_C_CY;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_C_XOR;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_D;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_D1;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_D2;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_D3;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_D4;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_D5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_D6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_DO5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_DO6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_DQ;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_D_CY;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_D_XOR;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_A;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_A1;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_A2;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_A3;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_A4;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_A5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_A6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_AO5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_AO6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_AQ;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_A_CY;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_A_XOR;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_B;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_B1;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_B2;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_B3;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_B4;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_B5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_B6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_BO5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_BO6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_BQ;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_B_CY;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_B_XOR;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_C;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_C1;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_C2;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_C3;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_C4;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_C5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_C6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_CLK;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_CO5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_CO6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_CQ;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_C_CY;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_C_XOR;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_D;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_D1;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_D2;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_D3;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_D4;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_D5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_D6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_DO5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_DO6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_DQ;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_D_CY;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X12Y114_D_XOR;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_A;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_A1;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_A2;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_A3;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_A4;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_A5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_A6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_AO5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_AO6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_AQ;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_A_CY;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_A_XOR;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_B;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_B1;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_B2;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_B3;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_B4;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_B5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_B6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_BO5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_BO6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_BQ;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_B_CY;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_B_XOR;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_C;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_C1;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_C2;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_C3;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_C4;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_C5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_C6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_CLK;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_CO5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_CO6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_CQ;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_C_CY;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_C_XOR;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_D;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_D1;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_D2;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_D3;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_D4;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_D5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_D6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_DO5;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_DO6;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_D_CY;
  wire [0:0] CLBLM_L_X10Y114_SLICE_X13Y114_D_XOR;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_A;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_A1;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_A2;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_A3;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_A4;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_A5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_A6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_AO5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_AO6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_A_CY;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_A_XOR;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_B;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_B1;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_B2;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_B3;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_B4;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_B5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_B6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_BO5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_BO6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_B_CY;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_B_XOR;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_C;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_C1;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_C2;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_C3;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_C4;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_C5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_C6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_CLK;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_CO5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_CO6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_CQ;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_C_CY;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_C_XOR;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_D;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_D1;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_D2;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_D3;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_D4;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_D5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_D6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_DO5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_DO6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_D_CY;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X12Y115_D_XOR;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_A;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_A1;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_A2;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_A3;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_A4;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_A5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_A6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_AO5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_AO6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_AQ;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_A_CY;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_A_XOR;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_B;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_B1;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_B2;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_B3;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_B4;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_B5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_B6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_BO5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_BO6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_BQ;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_B_CY;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_B_XOR;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_C;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_C1;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_C2;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_C3;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_C4;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_C5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_C6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_CLK;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_CO5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_CO6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_CQ;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_C_CY;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_C_XOR;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_D;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_D1;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_D2;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_D3;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_D4;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_D5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_D6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_DMUX;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_DO5;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_DO6;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_D_CY;
  wire [0:0] CLBLM_L_X10Y115_SLICE_X13Y115_D_XOR;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_A;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_A1;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_A2;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_A3;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_A4;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_A5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_A6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_AO5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_AO6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_A_CY;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_A_XOR;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_B;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_B1;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_B2;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_B3;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_B4;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_B5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_B6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_BO5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_BO6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_BQ;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_B_CY;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_B_XOR;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_C;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_C1;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_C2;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_C3;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_C4;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_C5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_C6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_CLK;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_CO5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_CO6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_CQ;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_C_CY;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_C_XOR;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_D;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_D1;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_D2;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_D3;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_D4;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_D5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_D6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_DMUX;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_DO5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_DO6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_D_CY;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X12Y116_D_XOR;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_A;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_A1;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_A2;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_A3;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_A4;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_A5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_A6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_AO5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_AO6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_AQ;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_A_CY;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_A_XOR;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_B;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_B1;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_B2;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_B3;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_B4;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_B5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_B6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_BO5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_BO6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_BQ;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_B_CY;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_B_XOR;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_C;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_C1;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_C2;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_C3;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_C4;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_C5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_C6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_CLK;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_CO5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_CO6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_CQ;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_C_CY;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_C_XOR;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_D;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_D1;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_D2;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_D3;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_D4;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_D5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_D6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_DO5;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_DO6;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_D_CY;
  wire [0:0] CLBLM_L_X10Y116_SLICE_X13Y116_D_XOR;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_A;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_A1;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_A2;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_A3;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_A4;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_A5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_A5Q;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_A6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_AMUX;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_AO5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_AO6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_AQ;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_A_CY;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_A_XOR;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_B;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_B1;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_B2;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_B3;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_B4;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_B5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_B6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_BO5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_BO6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_BQ;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_B_CY;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_B_XOR;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_C;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_C1;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_C2;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_C3;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_C4;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_C5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_C6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_CLK;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_CO5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_CO6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_C_CY;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_C_XOR;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_D;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_D1;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_D2;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_D3;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_D4;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_D5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_D6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_DO5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_DO6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_D_CY;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_D_XOR;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_A;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_A1;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_A2;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_A3;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_A4;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_A5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_A6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_AMUX;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_AO5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_AO6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_A_CY;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_A_XOR;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_B;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_B1;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_B2;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_B3;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_B4;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_B5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_B6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_BMUX;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_BO5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_BO6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_B_CY;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_B_XOR;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_C;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_C1;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_C2;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_C3;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_C4;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_C5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_C6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_CO5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_CO6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_C_CY;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_C_XOR;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_D;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_D1;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_D2;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_D3;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_D4;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_D5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_D6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_DO5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_DO6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_D_CY;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_D_XOR;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_A;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_A1;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_A2;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_A3;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_A4;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_A5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_A6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_AO5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_AO6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_AQ;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_A_CY;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_A_XOR;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_B;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_B1;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_B2;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_B3;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_B4;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_B5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_B6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_BO5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_BO6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_BQ;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_B_CY;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_B_XOR;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_C;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_C1;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_C2;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_C3;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_C4;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_C5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_C6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_CLK;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_CO5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_CO6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_C_CY;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_C_XOR;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_D;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_D1;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_D2;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_D3;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_D4;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_D5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_D6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_DO5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_DO6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_D_CY;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_D_XOR;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_A;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_A1;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_A2;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_A3;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_A4;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_A5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_A6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_AO5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_AO6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_AQ;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_A_CY;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_A_XOR;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_B;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_B1;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_B2;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_B3;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_B4;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_B5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_B6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_BO5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_BO6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_B_CY;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_B_XOR;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_C;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_C1;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_C2;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_C3;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_C4;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_C5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_C6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_CLK;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_CMUX;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_CO5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_CO6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_C_CY;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_C_XOR;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_D;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_D1;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_D2;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_D3;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_D4;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_D5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_D6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_DO5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_DO6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_D_CY;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_D_XOR;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_A;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_A1;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_A2;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_A3;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_A4;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_A5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_A6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_AO5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_AO6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_AQ;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_A_CY;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_A_XOR;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_B;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_B1;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_B2;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_B3;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_B4;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_B5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_B6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_BO5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_BO6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_B_CY;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_B_XOR;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_C;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_C1;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_C2;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_C3;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_C4;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_C5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_C6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_CLK;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_CMUX;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_CO5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_CO6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_C_CY;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_C_XOR;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_D;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_D1;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_D2;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_D3;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_D4;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_D5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_D6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_DO5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_DO6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_D_CY;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_D_XOR;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_A;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_A1;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_A2;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_A3;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_A4;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_A5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_A6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_AO5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_AO6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_A_CY;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_A_XOR;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_B;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_B1;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_B2;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_B3;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_B4;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_B5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_B6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_BO5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_BO6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_B_CY;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_B_XOR;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_C;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_C1;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_C2;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_C3;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_C4;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_C5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_C6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_CO5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_CO6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_C_CY;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_C_XOR;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_D;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_D1;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_D2;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_D3;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_D4;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_D5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_D6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_DO5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_DO6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_D_CY;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_D_XOR;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_A;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_A1;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_A2;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_A3;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_A4;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_A5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_A6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_AO5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_AO6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_A_CY;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_A_XOR;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_B;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_B1;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_B2;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_B3;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_B4;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_B5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_B6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_BO5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_BO6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_B_CY;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_B_XOR;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_C;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_C1;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_C2;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_C3;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_C4;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_C5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_C6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_CO5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_CO6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_C_CY;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_C_XOR;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_D;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_D1;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_D2;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_D3;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_D4;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_D5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_D6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_DO5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_DO6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_D_CY;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_D_XOR;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_A;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_A1;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_A2;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_A3;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_A4;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_A5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_A6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_AO5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_AO6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_A_CY;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_A_XOR;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_B;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_B1;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_B2;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_B3;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_B4;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_B5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_B6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_BO5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_BO6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_B_CY;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_B_XOR;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_C;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_C1;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_C2;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_C3;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_C4;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_C5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_C6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_CO5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_CO6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_C_CY;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_C_XOR;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_D;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_D1;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_D2;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_D3;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_D4;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_D5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_D6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_DO5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_DO6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_D_CY;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_D_XOR;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_A;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_A1;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_A2;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_A3;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_A4;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_A5;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_A6;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_AO5;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_AO6;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_AQ;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_A_CY;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_A_XOR;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_B;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_B1;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_B2;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_B3;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_B4;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_B5;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_B6;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_BMUX;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_BO5;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_BO6;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_B_CY;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_B_XOR;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_C;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_C1;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_C2;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_C3;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_C4;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_C5;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_C6;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_CLK;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_CMUX;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_CO5;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_CO6;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_C_CY;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_C_XOR;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_D;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_D1;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_D2;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_D3;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_D4;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_D5;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_D6;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_DO5;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_DO6;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_D_CY;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X16Y105_D_XOR;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_A;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_A1;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_A2;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_A3;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_A4;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_A5;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_A6;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_AMUX;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_AO5;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_AO6;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_A_CY;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_A_XOR;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_B;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_B1;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_B2;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_B3;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_B4;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_B5;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_B6;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_BMUX;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_BO5;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_BO6;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_B_CY;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_B_XOR;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_C;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_C1;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_C2;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_C3;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_C4;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_C5;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_C6;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_CO5;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_CO6;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_C_CY;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_C_XOR;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_D;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_D1;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_D2;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_D3;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_D4;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_D5;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_D6;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_DO5;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_DO6;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_D_CY;
  wire [0:0] CLBLM_L_X12Y105_SLICE_X17Y105_D_XOR;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_A;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_A1;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_A2;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_A3;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_A4;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_A5;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_A6;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_AO5;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_AO6;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_AQ;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_A_CY;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_A_XOR;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_B;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_B1;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_B2;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_B3;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_B4;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_B5;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_B6;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_BO5;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_BO6;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_B_CY;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_B_XOR;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_C;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_C1;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_C2;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_C3;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_C4;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_C5;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_C6;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_CLK;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_CO5;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_CO6;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_C_CY;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_C_XOR;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_D;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_D1;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_D2;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_D3;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_D4;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_D5;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_D6;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_DO5;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_DO6;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_D_CY;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X16Y106_D_XOR;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_A;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_A1;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_A2;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_A3;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_A4;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_A5;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_A6;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_AO5;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_AO6;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_AQ;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_A_CY;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_A_XOR;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_B;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_B1;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_B2;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_B3;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_B4;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_B5;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_B6;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_BO5;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_BO6;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_B_CY;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_B_XOR;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_C;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_C1;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_C2;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_C3;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_C4;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_C5;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_C6;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_CLK;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_CO5;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_CO6;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_C_CY;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_C_XOR;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_D;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_D1;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_D2;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_D3;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_D4;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_D5;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_D6;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_DO5;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_DO6;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_D_CY;
  wire [0:0] CLBLM_L_X12Y106_SLICE_X17Y106_D_XOR;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_A;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_A1;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_A2;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_A3;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_A4;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_A5;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_A6;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_AO5;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_AO6;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_AQ;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_A_CY;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_A_XOR;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_B;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_B1;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_B2;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_B3;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_B4;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_B5;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_B6;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_BO5;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_BO6;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_BQ;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_B_CY;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_B_XOR;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_C;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_C1;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_C2;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_C3;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_C4;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_C5;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_C6;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_CLK;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_CO5;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_CO6;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_CQ;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_C_CY;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_C_XOR;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_D;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_D1;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_D2;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_D3;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_D4;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_D5;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_D6;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_DO5;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_DO6;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_DQ;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_D_CY;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_D_XOR;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_A;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_A1;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_A2;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_A3;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_A4;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_A5;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_A6;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_AO5;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_AO6;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_AQ;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_A_CY;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_A_XOR;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_B;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_B1;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_B2;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_B3;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_B4;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_B5;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_B6;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_BO5;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_BO6;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_BQ;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_B_CY;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_B_XOR;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_C;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_C1;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_C2;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_C3;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_C4;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_C5;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_C6;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_CLK;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_CMUX;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_CO5;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_CO6;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_C_CY;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_C_XOR;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_D;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_D1;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_D2;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_D3;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_D4;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_D5;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_D6;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_DMUX;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_DO5;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_DO6;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_D_CY;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_D_XOR;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_A;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_A1;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_A2;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_A3;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_A4;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_A5;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_A6;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_AMUX;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_AO5;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_AO6;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_AQ;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_A_CY;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_A_XOR;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_B;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_B1;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_B2;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_B3;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_B4;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_B5;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_B6;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_BO5;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_BO6;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_BQ;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_B_CY;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_B_XOR;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_C;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_C1;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_C2;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_C3;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_C4;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_C5;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_C6;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_CLK;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_CO5;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_CO6;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_CQ;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_C_CY;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_C_XOR;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_D;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_D1;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_D2;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_D3;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_D4;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_D5;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_D6;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_DO5;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_DO6;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_DQ;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_D_CY;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_D_XOR;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_A;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_A1;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_A2;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_A3;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_A4;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_A5;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_A6;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_AO5;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_AO6;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_AQ;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_A_CY;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_A_XOR;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_B;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_B1;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_B2;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_B3;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_B4;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_B5;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_B6;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_BO5;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_BO6;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_BQ;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_B_CY;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_B_XOR;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_C;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_C1;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_C2;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_C3;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_C4;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_C5;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_C6;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_CLK;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_CMUX;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_CO5;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_CO6;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_C_CY;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_C_XOR;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_D;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_D1;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_D2;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_D3;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_D4;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_D5;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_D6;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_DO5;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_DO6;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_D_CY;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_D_XOR;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_A;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_A1;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_A2;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_A3;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_A4;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_A5;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_A6;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_AO5;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_AO6;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_AQ;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_A_CY;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_A_XOR;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_B;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_B1;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_B2;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_B3;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_B4;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_B5;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_B6;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_BO5;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_BO6;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_BQ;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_B_CY;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_B_XOR;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_C;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_C1;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_C2;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_C3;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_C4;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_C5;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_C6;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_CLK;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_CO5;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_CO6;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_CQ;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_C_CY;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_C_XOR;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_D;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_D1;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_D2;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_D3;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_D4;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_D5;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_D5Q;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_D6;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_DMUX;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_DO5;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_DO6;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_DQ;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_D_CY;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_D_XOR;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_A;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_A1;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_A2;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_A3;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_A4;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_A5;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_A6;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_AO5;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_AO6;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_AQ;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_A_CY;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_A_XOR;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_B;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_B1;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_B2;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_B3;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_B4;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_B5;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_B6;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_BO5;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_BO6;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_BQ;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_B_CY;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_B_XOR;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_C;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_C1;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_C2;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_C3;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_C4;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_C5;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_C6;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_CLK;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_CO5;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_CO6;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_CQ;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_C_CY;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_C_XOR;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_D;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_D1;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_D2;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_D3;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_D4;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_D5;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_D6;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_DO5;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_DO6;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_DQ;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_D_CY;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_D_XOR;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_A;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_A1;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_A2;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_A3;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_A4;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_A5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_A6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_AMUX;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_AO5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_AO6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_AQ;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_AX;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_A_CY;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_A_XOR;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_B;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_B1;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_B2;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_B3;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_B4;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_B5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_B6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_BMUX;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_BO5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_BO6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_B_CY;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_B_XOR;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_C;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_C1;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_C2;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_C3;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_C4;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_C5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_C6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_CE;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_CLK;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_CMUX;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_CO5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_CO6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_C_CY;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_C_XOR;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_D;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_D1;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_D2;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_D3;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_D4;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_D5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_D6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_DMUX;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_DO5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_DO6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_D_CY;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_D_XOR;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_SR;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_A;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_A1;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_A2;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_A3;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_A4;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_A5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_A6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_AO5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_AO6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_AQ;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_A_CY;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_A_XOR;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_B;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_B1;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_B2;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_B3;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_B4;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_B5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_B6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_BO5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_BO6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_BQ;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_B_CY;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_B_XOR;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_C;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_C1;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_C2;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_C3;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_C4;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_C5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_C6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_CLK;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_CO5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_CO6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_CQ;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_C_CY;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_C_XOR;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_D;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_D1;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_D2;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_D3;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_D4;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_D5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_D6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_DO5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_DO6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_DQ;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_D_CY;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_D_XOR;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_A;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_A1;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_A2;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_A3;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_A4;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_A5;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_A6;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_AO5;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_AO6;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_AQ;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_A_CY;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_A_XOR;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_B;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_B1;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_B2;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_B3;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_B4;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_B5;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_B6;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_BO5;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_BO6;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_BQ;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_B_CY;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_B_XOR;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_C;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_C1;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_C2;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_C3;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_C4;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_C5;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_C6;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_CLK;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_CO5;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_CO6;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_CQ;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_C_CY;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_C_XOR;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_D;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_D1;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_D2;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_D3;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_D4;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_D5;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_D6;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_DO5;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_DO6;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_DQ;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_D_CY;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X16Y111_D_XOR;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_A;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_A1;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_A2;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_A3;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_A4;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_A5;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_A6;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_AO5;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_AO6;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_A_CY;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_A_XOR;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_B;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_B1;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_B2;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_B3;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_B4;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_B5;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_B6;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_BO5;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_BO6;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_B_CY;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_B_XOR;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_C;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_C1;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_C2;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_C3;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_C4;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_C5;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_C6;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_CO5;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_CO6;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_C_CY;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_C_XOR;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_D;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_D1;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_D2;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_D3;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_D4;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_D5;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_D6;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_DO5;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_DO6;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_D_CY;
  wire [0:0] CLBLM_L_X12Y111_SLICE_X17Y111_D_XOR;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_A;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_A1;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_A2;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_A3;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_A4;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_A5;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_A5Q;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_A6;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_AMUX;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_AO5;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_AO6;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_AQ;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_AX;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_A_CY;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_A_XOR;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_B;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_B1;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_B2;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_B3;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_B4;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_B5;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_B5Q;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_B6;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_BMUX;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_BO5;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_BO6;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_BQ;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_B_CY;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_B_XOR;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_C;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_C1;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_C2;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_C3;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_C4;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_C5;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_C6;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_CLK;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_CO5;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_CO6;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_CQ;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_C_CY;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_C_XOR;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_D;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_D1;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_D2;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_D3;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_D4;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_D5;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_D6;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_DO5;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_DO6;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_DQ;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_D_CY;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X16Y112_D_XOR;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_A;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_A1;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_A2;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_A3;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_A4;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_A5;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_A5Q;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_A6;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_AMUX;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_AO5;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_AO6;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_AQ;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_AX;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_A_CY;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_A_XOR;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_B;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_B1;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_B2;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_B3;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_B4;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_B5;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_B5Q;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_B6;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_BMUX;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_BO5;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_BO6;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_BQ;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_BX;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_B_CY;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_B_XOR;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_C;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_C1;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_C2;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_C3;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_C4;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_C5;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_C6;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_CLK;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_CMUX;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_CO5;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_CO6;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_C_CY;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_C_XOR;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_D;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_D1;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_D2;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_D3;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_D4;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_D5;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_D6;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_DO5;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_DO6;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_D_CY;
  wire [0:0] CLBLM_L_X12Y112_SLICE_X17Y112_D_XOR;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_A;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_A1;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_A2;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_A3;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_A4;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_A5;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_A6;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_AO5;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_AO6;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_AQ;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_A_CY;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_A_XOR;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_B;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_B1;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_B2;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_B3;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_B4;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_B5;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_B6;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_BO5;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_BO6;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_BQ;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_B_CY;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_B_XOR;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_C;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_C1;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_C2;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_C3;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_C4;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_C5;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_C6;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_CLK;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_CO5;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_CO6;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_CQ;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_C_CY;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_C_XOR;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_D;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_D1;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_D2;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_D3;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_D4;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_D5;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_D6;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_DO5;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_DO6;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_D_CY;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X16Y113_D_XOR;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_A;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_A1;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_A2;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_A3;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_A4;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_A5;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_A6;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_AO5;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_AO6;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_AQ;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_A_CY;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_A_XOR;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_B;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_B1;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_B2;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_B3;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_B4;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_B5;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_B5Q;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_B6;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_BMUX;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_BO5;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_BO6;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_BQ;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_B_CY;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_B_XOR;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_C;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_C1;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_C2;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_C3;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_C4;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_C5;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_C6;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_CLK;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_CO5;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_CO6;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_CQ;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_C_CY;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_C_XOR;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_D;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_D1;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_D2;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_D3;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_D4;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_D5;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_D6;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_DO5;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_DO6;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_D_CY;
  wire [0:0] CLBLM_L_X12Y113_SLICE_X17Y113_D_XOR;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_A;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_A1;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_A2;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_A3;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_A4;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_A5;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_A6;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_AO5;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_AO6;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_AQ;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_A_CY;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_A_XOR;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_B;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_B1;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_B2;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_B3;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_B4;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_B5;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_B6;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_BO5;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_BO6;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_BQ;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_B_CY;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_B_XOR;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_C;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_C1;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_C2;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_C3;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_C4;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_C5;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_C6;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_CLK;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_CO5;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_CO6;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_CQ;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_C_CY;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_C_XOR;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_D;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_D1;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_D2;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_D3;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_D4;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_D5;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_D6;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_DMUX;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_DO5;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_DO6;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_D_CY;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X16Y114_D_XOR;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_A;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_A1;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_A2;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_A3;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_A4;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_A5;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_A6;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_AO5;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_AO6;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_AQ;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_A_CY;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_A_XOR;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_B;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_B1;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_B2;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_B3;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_B4;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_B5;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_B6;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_BO5;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_BO6;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_BQ;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_B_CY;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_B_XOR;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_C;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_C1;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_C2;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_C3;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_C4;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_C5;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_C6;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_CLK;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_CO5;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_CO6;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_C_CY;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_C_XOR;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_D;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_D1;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_D2;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_D3;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_D4;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_D5;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_D6;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_DO5;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_DO6;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_D_CY;
  wire [0:0] CLBLM_L_X12Y114_SLICE_X17Y114_D_XOR;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_A;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_A1;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_A2;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_A3;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_A4;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_A5;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_A6;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_AO5;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_AO6;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_AQ;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_AX;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_A_CY;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_A_XOR;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_B;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_B1;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_B2;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_B3;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_B4;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_B5;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_B6;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_BO5;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_BO6;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_B_CY;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_B_XOR;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_C;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_C1;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_C2;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_C3;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_C4;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_C5;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_C6;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_CLK;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_CO5;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_CO6;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_C_CY;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_C_XOR;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_D;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_D1;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_D2;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_D3;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_D4;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_D5;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_D6;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_DO5;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_DO6;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_D_CY;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X16Y115_D_XOR;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_A;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_A1;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_A2;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_A3;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_A4;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_A5;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_A6;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_AO5;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_AO6;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_A_CY;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_A_XOR;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_B;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_B1;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_B2;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_B3;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_B4;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_B5;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_B6;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_BO5;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_BO6;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_B_CY;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_B_XOR;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_C;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_C1;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_C2;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_C3;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_C4;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_C5;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_C6;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_CO5;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_CO6;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_C_CY;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_C_XOR;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_D;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_D1;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_D2;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_D3;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_D4;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_D5;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_D6;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_DO5;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_DO6;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_D_CY;
  wire [0:0] CLBLM_L_X12Y115_SLICE_X17Y115_D_XOR;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_A;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_A1;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_A2;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_A3;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_A4;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_A5;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_A6;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_AMUX;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_AO5;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_AO6;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_AQ;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_AX;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_A_CY;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_A_XOR;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_B;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_B1;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_B2;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_B3;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_B4;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_B5;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_B6;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_BO5;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_BO6;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_B_CY;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_B_XOR;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_C;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_C1;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_C2;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_C3;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_C4;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_C5;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_C6;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_CE;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_CLK;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_CO5;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_CO6;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_C_CY;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_C_XOR;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_D;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_D1;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_D2;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_D3;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_D4;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_D5;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_D6;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_DO5;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_DO6;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_D_CY;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_D_XOR;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X16Y117_SR;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_A;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_A1;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_A2;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_A3;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_A4;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_A5;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_A6;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_AO5;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_AO6;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_AQ;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_A_CY;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_A_XOR;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_B;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_B1;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_B2;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_B3;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_B4;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_B5;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_B6;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_BO5;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_BO6;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_BQ;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_B_CY;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_B_XOR;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_C;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_C1;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_C2;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_C3;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_C4;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_C5;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_C6;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_CLK;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_CO5;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_CO6;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_C_CY;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_C_XOR;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_D;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_D1;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_D2;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_D3;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_D4;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_D5;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_D6;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_DO5;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_DO6;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_D_CY;
  wire [0:0] CLBLM_L_X12Y117_SLICE_X17Y117_D_XOR;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_A;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_A1;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_A2;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_A3;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_A4;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_A5;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_A6;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_AO5;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_AO6;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_AQ;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_AX;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_A_CY;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_A_XOR;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_B;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_B1;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_B2;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_B3;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_B4;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_B5;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_B6;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_BO5;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_BO6;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_B_CY;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_B_XOR;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_C;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_C1;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_C2;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_C3;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_C4;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_C5;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_C6;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_CE;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_CLK;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_CO5;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_CO6;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_C_CY;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_C_XOR;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_D;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_D1;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_D2;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_D3;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_D4;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_D5;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_D6;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_DO5;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_DO6;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_D_CY;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_D_XOR;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X16Y118_SR;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_A;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_A1;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_A2;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_A3;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_A4;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_A5;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_A6;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_AO5;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_AO6;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_A_CY;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_A_XOR;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_B;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_B1;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_B2;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_B3;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_B4;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_B5;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_B6;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_BO5;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_BO6;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_B_CY;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_B_XOR;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_C;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_C1;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_C2;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_C3;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_C4;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_C5;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_C6;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_CO5;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_CO6;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_C_CY;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_C_XOR;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_D;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_D1;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_D2;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_D3;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_D4;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_D5;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_D6;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_DO5;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_DO6;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_D_CY;
  wire [0:0] CLBLM_L_X12Y118_SLICE_X17Y118_D_XOR;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_A;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_A1;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_A2;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_A3;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_A4;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_A5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_A6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_AO5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_AO6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_A_CY;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_A_XOR;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_B;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_B1;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_B2;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_B3;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_B4;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_B5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_B6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_BO5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_BO6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_B_CY;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_B_XOR;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_C;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_C1;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_C2;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_C3;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_C4;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_C5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_C6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_CO5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_CO6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_C_CY;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_C_XOR;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_D;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_D1;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_D2;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_D3;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_D4;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_D5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_D6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_DO5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_DO6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_D_CY;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_D_XOR;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_A;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_A1;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_A2;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_A3;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_A4;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_A5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_A6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_AMUX;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_AO5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_AO6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_AQ;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_A_CY;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_A_XOR;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_B;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_B1;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_B2;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_B3;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_B4;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_B5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_B6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_BO5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_BO6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_B_CY;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_B_XOR;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_C;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_C1;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_C2;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_C3;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_C4;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_C5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_C6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_CLK;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_CO5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_CO6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_C_CY;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_C_XOR;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_D;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_D1;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_D2;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_D3;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_D4;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_D5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_D6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_DO5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_DO6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_D_CY;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_D_XOR;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_A;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_A1;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_A2;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_A3;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_A4;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_A5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_A6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_AO5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_AO6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_AQ;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_A_CY;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_A_XOR;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_B;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_B1;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_B2;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_B3;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_B4;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_B5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_B6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_BO5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_BO6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_B_CY;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_B_XOR;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_C;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_C1;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_C2;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_C3;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_C4;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_C5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_C6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_CLK;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_CO5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_CO6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_C_CY;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_C_XOR;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_D;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_D1;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_D2;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_D3;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_D4;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_D5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_D6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_DO5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_DO6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_D_CY;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_D_XOR;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_A;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_A1;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_A2;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_A3;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_A4;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_A5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_A6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_AO5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_AO6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_AQ;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_A_CY;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_A_XOR;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_B;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_B1;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_B2;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_B3;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_B4;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_B5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_B6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_BO5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_BO6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_BQ;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_B_CY;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_B_XOR;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_C;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_C1;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_C2;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_C3;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_C4;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_C5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_C6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_CLK;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_CMUX;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_CO5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_CO6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_C_CY;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_C_XOR;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_D;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_D1;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_D2;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_D3;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_D4;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_D5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_D6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_DO5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_DO6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_D_CY;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_D_XOR;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_A;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_A1;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_A2;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_A3;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_A4;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_A5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_A6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_AO5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_AO6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_AQ;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_A_CY;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_A_XOR;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_B;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_B1;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_B2;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_B3;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_B4;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_B5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_B6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_BO5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_BO6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_BQ;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_B_CY;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_B_XOR;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_C;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_C1;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_C2;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_C3;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_C4;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_C5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_C6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_CLK;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_CO5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_CO6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_CQ;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_C_CY;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_C_XOR;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_D;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_D1;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_D2;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_D3;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_D4;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_D5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_D6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_DMUX;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_DO5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_DO6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_D_CY;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_D_XOR;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_A;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_A1;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_A2;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_A3;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_A4;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_A5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_A5Q;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_A6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_AMUX;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_AO5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_AO6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_AQ;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_AX;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_A_CY;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_A_XOR;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_B;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_B1;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_B2;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_B3;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_B4;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_B5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_B6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_BO5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_BO6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_BQ;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_B_CY;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_B_XOR;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_C;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_C1;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_C2;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_C3;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_C4;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_C5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_C6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_CLK;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_CMUX;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_CO5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_CO6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_C_CY;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_C_XOR;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_D;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_D1;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_D2;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_D3;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_D4;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_D5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_D6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_DO5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_DO6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_D_CY;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_D_XOR;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_A;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_A1;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_A2;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_A3;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_A4;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_A5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_A6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_AO5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_AO6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_AQ;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_A_CY;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_A_XOR;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_B;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_B1;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_B2;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_B3;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_B4;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_B5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_B6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_BO5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_BO6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_BQ;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_B_CY;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_B_XOR;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_C;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_C1;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_C2;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_C3;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_C4;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_C5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_C6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_CLK;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_CO5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_CO6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_CQ;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_C_CY;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_C_XOR;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_D;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_D1;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_D2;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_D3;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_D4;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_D5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_D6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_DO5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_DO6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_D_CY;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_D_XOR;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_A;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_A1;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_A2;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_A3;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_A4;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_A5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_A5Q;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_A6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_AMUX;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_AO5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_AO6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_AQ;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_A_CY;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_A_XOR;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_B;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_B1;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_B2;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_B3;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_B4;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_B5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_B5Q;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_B6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_BMUX;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_BO5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_BO6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_BQ;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_B_CY;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_B_XOR;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_C;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_C1;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_C2;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_C3;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_C4;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_C5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_C6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_CLK;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_CO5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_CO6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_CQ;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_C_CY;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_C_XOR;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_D;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_D1;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_D2;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_D3;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_D4;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_D5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_D6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_DMUX;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_DO5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_DO6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_D_CY;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_D_XOR;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_A;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_A1;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_A2;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_A3;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_A4;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_A5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_A6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_AMUX;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_AO5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_AO6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_AQ;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_A_CY;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_A_XOR;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_B;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_B1;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_B2;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_B3;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_B4;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_B5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_B6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_BO5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_BO6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_BQ;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_B_CY;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_B_XOR;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_C;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_C1;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_C2;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_C3;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_C4;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_C5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_C6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_CLK;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_CO5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_CO6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_CQ;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_C_CY;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_C_XOR;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_D;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_D1;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_D2;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_D3;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_D4;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_D5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_D6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_DO5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_DO6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_DQ;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_D_CY;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_D_XOR;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_A;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_A1;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_A2;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_A3;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_A4;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_A5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_A6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_AO5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_AO6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_AQ;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_A_CY;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_A_XOR;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_B;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_B1;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_B2;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_B3;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_B4;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_B5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_B6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_BO5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_BO6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_BQ;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_B_CY;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_B_XOR;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_C;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_C1;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_C2;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_C3;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_C4;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_C5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_C6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_CLK;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_CO5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_CO6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_C_CY;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_C_XOR;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_D;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_D1;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_D2;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_D3;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_D4;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_D5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_D6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_DO5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_DO6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_D_CY;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_D_XOR;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_A;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_A1;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_A2;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_A3;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_A4;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_A5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_A6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_AO5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_AO6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_AQ;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_A_CY;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_A_XOR;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_B;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_B1;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_B2;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_B3;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_B4;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_B5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_B6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_BO5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_BO6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_BQ;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_B_CY;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_B_XOR;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_C;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_C1;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_C2;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_C3;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_C4;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_C5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_C5Q;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_C6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_CLK;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_CMUX;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_CO5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_CO6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_CQ;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_C_CY;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_C_XOR;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_D;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_D1;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_D2;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_D3;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_D4;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_D5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_D6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_DO5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_DO6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_DQ;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_D_CY;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_D_XOR;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_A;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_A1;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_A2;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_A3;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_A4;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_A5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_A5Q;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_A6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_AMUX;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_AO5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_AO6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_AQ;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_AX;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_A_CY;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_A_XOR;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_B;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_B1;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_B2;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_B3;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_B4;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_B5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_B6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_BO5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_BO6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_BQ;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_B_CY;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_B_XOR;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_C;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_C1;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_C2;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_C3;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_C4;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_C5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_C6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_CLK;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_CO5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_CO6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_CQ;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_C_CY;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_C_XOR;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_D;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_D1;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_D2;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_D3;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_D4;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_D5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_D6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_DO5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_DO6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_D_CY;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_D_XOR;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A1;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A2;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A3;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A4;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_AO5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_AO6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_AQ;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A_CY;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A_XOR;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B1;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B2;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B3;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B4;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_BO5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_BO6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_BQ;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B_CY;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B_XOR;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C1;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C2;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C3;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C4;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_CLK;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_CMUX;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_CO5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_CO6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C_CY;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C_XOR;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D1;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D2;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D3;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D4;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_DO5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_DO6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D_CY;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D_XOR;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A1;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A2;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A3;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A4;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A5Q;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_AMUX;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_AO5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_AO6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_AQ;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_AX;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A_CY;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A_XOR;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B1;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B2;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B3;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B4;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_BMUX;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_BO5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_BO6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B_CY;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B_XOR;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C1;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C2;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C3;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C4;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_CLK;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_CO5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_CO6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_CQ;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C_CY;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C_XOR;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D1;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D2;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D3;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D4;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_DO5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_DO6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_DQ;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D_CY;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D_XOR;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A1;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A2;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A3;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A4;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A5Q;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_AMUX;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_AO5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_AO6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_AQ;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A_CY;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A_XOR;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B1;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B2;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B3;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B4;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_BMUX;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_BO5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_BO6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B_CY;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B_XOR;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C1;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C2;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C3;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C4;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_CLK;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_CMUX;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_CO5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_CO6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C_CY;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C_XOR;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D1;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D2;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D3;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D4;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_DMUX;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_DO5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_DO6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D_CY;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D_XOR;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A1;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A2;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A3;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A4;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_AO5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_AO6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_AQ;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A_CY;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A_XOR;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B1;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B2;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B3;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B4;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_BO5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_BO6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_BQ;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B_CY;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B_XOR;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C1;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C2;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C3;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C4;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_CLK;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_CO5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_CO6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_CQ;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C_CY;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C_XOR;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D1;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D2;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D3;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D4;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_DMUX;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_DO5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_DO6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D_CY;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D_XOR;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A1;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A2;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A3;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A4;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A5Q;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_AMUX;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_AO5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_AO6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_AQ;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A_CY;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A_XOR;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B1;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B2;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B3;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B4;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_BO5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_BO6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B_CY;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B_XOR;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C1;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C2;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C3;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C4;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_CLK;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_CO5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_CO6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C_CY;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C_XOR;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D1;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D2;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D3;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D4;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_DO5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_DO6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D_CY;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D_XOR;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A1;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A2;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A3;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A4;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_AMUX;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_AO5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_AO6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A_CY;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A_XOR;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B1;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B2;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B3;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B4;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_BO5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_BO6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B_CY;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B_XOR;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C1;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C2;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C3;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C4;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_CO5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_CO6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C_CY;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C_XOR;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D1;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D2;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D3;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D4;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_DMUX;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_DO5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_DO6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D_CY;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D_XOR;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A1;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A2;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A3;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A4;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_AO5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_AO6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_AQ;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A_CY;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A_XOR;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B1;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B2;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B3;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B4;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_BO5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_BO6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_BQ;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B_CY;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B_XOR;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C1;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C2;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C3;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C4;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_CLK;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_CO5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_CO6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_CQ;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C_CY;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C_XOR;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D1;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D2;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D3;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D4;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D5Q;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_DMUX;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_DO5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_DO6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_DQ;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D_CY;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D_XOR;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A1;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A2;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A3;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A4;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_AO5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_AO6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_AQ;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A_CY;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A_XOR;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B1;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B2;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B3;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B4;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_BO5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_BO6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_BQ;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B_CY;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B_XOR;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C1;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C2;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C3;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C4;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_CLK;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_CO5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_CO6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C_CY;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C_XOR;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D1;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D2;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D3;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D4;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_DO5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_DO6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D_CY;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D_XOR;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_A;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_A1;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_A2;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_A3;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_A4;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_A5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_A6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_AO5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_AO6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_AQ;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_A_CY;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_A_XOR;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_B;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_B1;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_B2;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_B3;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_B4;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_B5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_B6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_BO5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_BO6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_BQ;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_B_CY;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_B_XOR;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_C;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_C1;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_C2;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_C3;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_C4;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_C5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_C6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_CLK;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_CO5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_CO6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_CQ;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_C_CY;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_C_XOR;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_D;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_D1;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_D2;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_D3;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_D4;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_D5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_D6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_DO5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_DO6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_DQ;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_D_CY;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_D_XOR;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_A;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_A1;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_A2;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_A3;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_A4;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_A5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_A6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_AO5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_AO6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_AQ;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_A_CY;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_A_XOR;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_B;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_B1;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_B2;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_B3;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_B4;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_B5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_B5Q;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_B6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_BMUX;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_BO5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_BO6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_BQ;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_B_CY;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_B_XOR;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_C;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_C1;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_C2;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_C3;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_C4;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_C5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_C6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_CLK;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_CO5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_CO6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_CQ;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_C_CY;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_C_XOR;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_D;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_D1;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_D2;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_D3;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_D4;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_D5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_D6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_DO5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_DO6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_D_CY;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_D_XOR;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_A;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_A1;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_A2;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_A3;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_A4;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_A5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_A5Q;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_A6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_AMUX;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_AO5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_AO6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_AQ;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_AX;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_A_CY;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_A_XOR;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_B;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_B1;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_B2;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_B3;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_B4;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_B5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_B6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_BO5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_BO6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_BQ;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_B_CY;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_B_XOR;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_C;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_C1;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_C2;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_C3;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_C4;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_C5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_C6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_CLK;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_CO5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_CO6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_CQ;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_C_CY;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_C_XOR;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_D;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_D1;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_D2;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_D3;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_D4;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_D5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_D6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_DO5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_DO6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_D_CY;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X10Y115_D_XOR;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_A;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_A1;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_A2;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_A3;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_A4;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_A5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_A6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_AO5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_AO6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_AQ;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_A_CY;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_A_XOR;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_B;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_B1;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_B2;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_B3;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_B4;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_B5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_B6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_BO5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_BO6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_BQ;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_B_CY;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_B_XOR;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_C;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_C1;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_C2;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_C3;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_C4;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_C5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_C6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_CLK;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_CO5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_CO6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_C_CY;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_C_XOR;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_D;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_D1;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_D2;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_D3;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_D4;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_D5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_D6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_DO5;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_DO6;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_D_CY;
  wire [0:0] CLBLM_L_X8Y115_SLICE_X11Y115_D_XOR;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_A;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_A1;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_A2;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_A3;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_A4;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_A5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_A6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_AO5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_AO6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_A_CY;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_A_XOR;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_B;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_B1;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_B2;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_B3;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_B4;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_B5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_B6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_BO5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_BO6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_BQ;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_B_CY;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_B_XOR;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_C;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_C1;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_C2;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_C3;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_C4;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_C5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_C6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_CLK;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_CO5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_CO6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_CQ;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_C_CY;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_C_XOR;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_D;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_D1;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_D2;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_D3;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_D4;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_D5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_D6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_DO5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_DO6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_DQ;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_D_CY;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_D_XOR;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_A;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_A1;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_A2;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_A3;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_A4;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_A5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_A6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_AO5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_AO6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_AQ;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_A_CY;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_A_XOR;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_B;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_B1;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_B2;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_B3;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_B4;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_B5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_B6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_BO5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_BO6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_BQ;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_B_CY;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_B_XOR;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_C;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_C1;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_C2;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_C3;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_C4;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_C5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_C6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_CLK;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_CO5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_CO6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_C_CY;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_C_XOR;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_D;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_D1;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_D2;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_D3;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_D4;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_D5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_D6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_DO5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_DO6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_D_CY;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_D_XOR;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_A;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_A1;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_A2;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_A3;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_A4;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_A5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_A6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_AO5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_AO6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_AQ;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_A_CY;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_A_XOR;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_B;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_B1;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_B2;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_B3;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_B4;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_B5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_B6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_BO5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_BO6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_BQ;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_B_CY;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_B_XOR;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_C;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_C1;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_C2;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_C3;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_C4;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_C5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_C6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_CLK;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_CO5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_CO6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_C_CY;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_C_XOR;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_D;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_D1;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_D2;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_D3;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_D4;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_D5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_D6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_DO5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_DO6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_D_CY;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_D_XOR;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_A;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_A1;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_A2;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_A3;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_A4;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_A5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_A6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_AO5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_AO6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_A_CY;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_A_XOR;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_B;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_B1;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_B2;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_B3;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_B4;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_B5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_B6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_BO5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_BO6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_B_CY;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_B_XOR;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_C;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_C1;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_C2;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_C3;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_C4;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_C5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_C6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_CO5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_CO6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_C_CY;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_C_XOR;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_D;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_D1;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_D2;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_D3;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_D4;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_D5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_D6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_DO5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_DO6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_D_CY;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_D_XOR;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_A;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_A1;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_A2;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_A3;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_A4;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_A5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_A6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_AO5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_AO6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_AQ;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_A_CY;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_A_XOR;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_B;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_B1;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_B2;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_B3;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_B4;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_B5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_B6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_BO5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_BO6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_BQ;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_B_CY;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_B_XOR;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_C;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_C1;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_C2;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_C3;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_C4;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_C5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_C6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_CLK;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_CMUX;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_CO5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_CO6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_C_CY;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_C_XOR;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_D;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_D1;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_D2;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_D3;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_D4;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_D5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_D6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_DMUX;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_DO5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_DO6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_D_CY;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_D_XOR;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_A;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_A1;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_A2;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_A3;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_A4;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_A5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_A6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_AO5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_AO6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_A_CY;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_A_XOR;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_B;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_B1;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_B2;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_B3;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_B4;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_B5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_B6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_BO5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_BO6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_B_CY;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_B_XOR;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_C;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_C1;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_C2;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_C3;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_C4;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_C5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_C6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_CO5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_CO6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_C_CY;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_C_XOR;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_D;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_D1;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_D2;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_D3;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_D4;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_D5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_D6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_DO5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_DO6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_D_CY;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_D_XOR;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_A;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_A1;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_A2;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_A3;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_A4;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_A5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_A6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_AMUX;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_AO5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_AO6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_AQ;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_A_CY;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_A_XOR;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_B;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_B1;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_B2;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_B3;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_B4;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_B5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_B6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_BO5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_BO6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_B_CY;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_B_XOR;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_C;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_C1;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_C2;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_C3;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_C4;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_C5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_C6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_CLK;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_CO5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_CO6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_C_CY;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_C_XOR;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_D;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_D1;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_D2;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_D3;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_D4;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_D5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_D6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_DO5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_DO6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_D_CY;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_D_XOR;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_A;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_A1;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_A2;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_A3;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_A4;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_A5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_A6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_AO5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_AO6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_A_CY;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_A_XOR;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_B;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_B1;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_B2;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_B3;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_B4;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_B5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_B6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_BO5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_BO6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_B_CY;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_B_XOR;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_C;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_C1;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_C2;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_C3;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_C4;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_C5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_C6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_CO5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_CO6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_C_CY;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_C_XOR;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_D;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_D1;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_D2;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_D3;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_D4;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_D5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_D6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_DO5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_DO6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_D_CY;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_D_XOR;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_A;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_A1;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_A2;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_A3;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_A4;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_A5;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_A6;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_AO5;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_AO6;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_A_CY;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_A_XOR;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_B;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_B1;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_B2;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_B3;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_B4;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_B5;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_B6;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_BO5;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_BO6;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_B_CY;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_B_XOR;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_C;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_C1;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_C2;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_C3;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_C4;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_C5;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_C6;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_CO5;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_CO6;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_C_CY;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_C_XOR;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_D;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_D1;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_D2;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_D3;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_D4;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_D5;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_D6;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_DO5;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_DO6;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_D_CY;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X162Y138_D_XOR;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_A;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_A1;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_A2;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_A3;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_A4;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_A5;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_A6;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_AO5;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_AO6;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_A_CY;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_A_XOR;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_B;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_B1;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_B2;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_B3;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_B4;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_B5;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_B6;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_BO5;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_BO6;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_B_CY;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_B_XOR;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_C;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_C1;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_C2;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_C3;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_C4;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_C5;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_C6;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_CO5;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_CO6;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_C_CY;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_C_XOR;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_D;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_D1;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_D2;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_D3;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_D4;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_D5;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_D6;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_DO5;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_DO6;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_D_CY;
  wire [0:0] CLBLM_R_X103Y138_SLICE_X163Y138_D_XOR;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A1;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A2;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A3;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A4;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_AO5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_AO6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A_CY;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A_XOR;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B1;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B2;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B3;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B4;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_BO5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_BO6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B_CY;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B_XOR;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C1;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C2;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C3;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C4;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_CO5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_CO6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C_CY;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C_XOR;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D1;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D2;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D3;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D4;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_DO5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_DO6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D_CY;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D_XOR;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A1;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A2;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A3;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A4;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_AO5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_AO6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A_CY;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A_XOR;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B1;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B2;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B3;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B4;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_BO5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_BO6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B_CY;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B_XOR;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C1;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C2;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C3;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C4;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_CO5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_CO6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C_CY;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C_XOR;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D1;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D2;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D3;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D4;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_DO5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_DO6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D_CY;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D_XOR;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_A;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_A1;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_A2;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_A3;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_A4;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_A5;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_A6;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_AO5;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_AO6;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_A_CY;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_A_XOR;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_B;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_B1;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_B2;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_B3;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_B4;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_B5;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_B6;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_BO5;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_BO6;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_B_CY;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_B_XOR;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_C;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_C1;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_C2;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_C3;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_C4;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_C5;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_C6;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_CO5;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_CO6;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_C_CY;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_C_XOR;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_D;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_D1;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_D2;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_D3;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_D4;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_D5;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_D6;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_DO5;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_DO6;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_D_CY;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X162Y170_D_XOR;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_A;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_A1;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_A2;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_A3;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_A4;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_A5;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_A6;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_AMUX;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_AO5;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_AO6;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_A_CY;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_A_XOR;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_B;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_B1;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_B2;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_B3;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_B4;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_B5;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_B6;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_BO5;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_BO6;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_B_CY;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_B_XOR;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_C;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_C1;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_C2;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_C3;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_C4;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_C5;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_C6;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_CO5;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_CO6;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_C_CY;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_C_XOR;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_D;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_D1;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_D2;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_D3;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_D4;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_D5;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_D6;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_DO5;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_DO6;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_D_CY;
  wire [0:0] CLBLM_R_X103Y170_SLICE_X163Y170_D_XOR;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_A;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_A1;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_A2;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_A3;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_A4;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_A5;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_A6;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_AO5;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_AO6;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_A_CY;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_A_XOR;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_B;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_B1;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_B2;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_B3;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_B4;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_B5;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_B6;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_BO5;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_BO6;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_B_CY;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_B_XOR;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_C;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_C1;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_C2;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_C3;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_C4;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_C5;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_C6;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_CO5;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_CO6;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_C_CY;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_C_XOR;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_D;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_D1;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_D2;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_D3;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_D4;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_D5;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_D6;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_DO5;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_DO6;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_D_CY;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_D_XOR;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_A;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_A1;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_A2;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_A3;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_A4;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_A5;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_A6;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_AMUX;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_AO5;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_AO6;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_A_CY;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_A_XOR;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_B;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_B1;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_B2;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_B3;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_B4;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_B5;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_B6;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_BO5;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_BO6;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_B_CY;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_B_XOR;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_C;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_C1;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_C2;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_C3;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_C4;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_C5;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_C6;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_CO5;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_CO6;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_C_CY;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_C_XOR;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_D;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_D1;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_D2;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_D3;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_D4;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_D5;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_D6;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_DO5;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_DO6;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_D_CY;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_D_XOR;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_A;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_A1;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_A2;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_A3;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_A4;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_A5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_A6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_AO5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_AO6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_A_CY;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_A_XOR;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_B;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_B1;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_B2;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_B3;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_B4;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_B5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_B6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_BO5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_BO6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_B_CY;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_B_XOR;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_C;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_C1;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_C2;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_C3;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_C4;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_C5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_C6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_CO5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_CO6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_C_CY;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_C_XOR;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_D;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_D1;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_D2;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_D3;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_D4;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_D5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_D6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_DO5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_DO6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_D_CY;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_D_XOR;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_A;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_A1;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_A2;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_A3;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_A4;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_A5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_A6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_AMUX;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_AO5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_AO6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_A_CY;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_A_XOR;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_B;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_B1;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_B2;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_B3;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_B4;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_B5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_B6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_BO5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_BO6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_B_CY;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_B_XOR;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_C;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_C1;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_C2;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_C3;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_C4;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_C5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_C6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_CO5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_CO6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_C_CY;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_C_XOR;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_D;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_D1;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_D2;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_D3;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_D4;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_D5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_D6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_DO5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_DO6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_D_CY;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_D_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_AO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_AO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_BO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_BO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_CO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_CO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_DO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_DO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_AMUX;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_AO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_AO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_BO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_BO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_CO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_CO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_DO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_DO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D_XOR;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_A;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_A1;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_A2;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_A3;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_A4;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_A5;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_A6;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_AO5;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_AO6;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_AQ;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_A_CY;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_A_XOR;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_B;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_B1;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_B2;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_B3;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_B4;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_B5;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_B6;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_BO5;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_BO6;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_BQ;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_B_CY;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_B_XOR;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_C;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_C1;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_C2;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_C3;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_C4;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_C5;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_C5Q;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_C6;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_CLK;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_CMUX;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_CO5;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_CO6;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_CQ;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_C_CY;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_C_XOR;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_D;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_D1;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_D2;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_D3;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_D4;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_D5;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_D6;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_DO5;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_DO6;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_DQ;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_D_CY;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_D_XOR;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_A;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_A1;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_A2;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_A3;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_A4;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_A5;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_A5Q;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_A6;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_AMUX;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_AO5;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_AO6;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_AQ;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_AX;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_A_CY;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_A_XOR;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_B;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_B1;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_B2;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_B3;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_B4;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_B5;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_B6;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_BO5;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_BO6;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_BQ;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_B_CY;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_B_XOR;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_C;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_C1;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_C2;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_C3;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_C4;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_C5;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_C6;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_CLK;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_CO5;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_CO6;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_CQ;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_C_CY;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_C_XOR;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_D;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_D1;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_D2;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_D3;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_D4;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_D5;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_D6;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_DMUX;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_DO5;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_DO6;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_D_CY;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_D_XOR;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_A;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_A1;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_A2;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_A3;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_A4;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_A5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_A6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_AO5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_AO6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_AQ;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_A_CY;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_A_XOR;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_B;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_B1;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_B2;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_B3;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_B4;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_B5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_B6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_BO5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_BO6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_BQ;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_B_CY;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_B_XOR;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_C;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_C1;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_C2;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_C3;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_C4;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_C5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_C6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_CLK;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_CO5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_CO6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_CQ;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_C_CY;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_C_XOR;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_D;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_D1;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_D2;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_D3;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_D4;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_D5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_D6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_DO5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_DO6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_DQ;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_D_CY;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_D_XOR;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_A;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_A1;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_A2;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_A3;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_A4;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_A5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_A6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_AO5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_AO6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_AQ;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_A_CY;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_A_XOR;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_B;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_B1;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_B2;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_B3;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_B4;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_B5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_B6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_BMUX;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_BO5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_BO6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_B_CY;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_B_XOR;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_C;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_C1;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_C2;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_C3;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_C4;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_C5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_C6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_CLK;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_CMUX;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_CO5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_CO6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_C_CY;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_C_XOR;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_D;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_D1;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_D2;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_D3;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_D4;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_D5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_D6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_DMUX;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_DO5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_DO6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_D_CY;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_D_XOR;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_A;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_A1;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_A2;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_A3;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_A4;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_A5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_A6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_AMUX;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_AO5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_AO6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_A_CY;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_A_XOR;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_B;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_B1;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_B2;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_B3;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_B4;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_B5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_B6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_BO5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_BO6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_B_CY;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_B_XOR;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_C;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_C1;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_C2;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_C3;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_C4;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_C5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_C6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_CO5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_CO6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_C_CY;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_C_XOR;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_D;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_D1;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_D2;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_D3;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_D4;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_D5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_D6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_DO5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_DO6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_D_CY;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_D_XOR;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_A;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_A1;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_A2;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_A3;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_A4;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_A5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_A6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_AO5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_AO6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_AQ;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_A_CY;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_A_XOR;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_B;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_B1;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_B2;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_B3;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_B4;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_B5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_B6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_BO5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_BO6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_BQ;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_B_CY;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_B_XOR;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_C;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_C1;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_C2;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_C3;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_C4;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_C5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_C6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_CLK;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_CO5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_CO6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_CQ;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_C_CY;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_C_XOR;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_D;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_D1;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_D2;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_D3;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_D4;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_D5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_D6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_DO5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_DO6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_D_CY;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_D_XOR;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_A;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_A1;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_A2;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_A3;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_A4;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_A5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_A6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_AO5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_AO6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_AQ;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_A_CY;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_A_XOR;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_B;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_B1;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_B2;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_B3;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_B4;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_B5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_B6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_BMUX;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_BO5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_BO6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_B_CY;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_B_XOR;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_C;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_C1;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_C2;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_C3;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_C4;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_C5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_C6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_CLK;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_CO5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_CO6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_C_CY;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_C_XOR;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_D;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_D1;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_D2;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_D3;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_D4;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_D5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_D6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_DO5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_DO6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_D_CY;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_D_XOR;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_A;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_A1;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_A2;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_A3;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_A4;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_A5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_A6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_AMUX;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_AO5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_AO6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_AQ;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_AX;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_A_CY;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_A_XOR;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_B;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_B1;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_B2;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_B3;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_B4;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_B5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_B6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_BMUX;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_BO5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_BO6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_B_CY;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_B_XOR;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_C;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_C1;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_C2;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_C3;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_C4;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_C5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_C6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_CLK;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_CMUX;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_CO5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_CO6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_C_CY;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_C_XOR;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_D;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_D1;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_D2;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_D3;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_D4;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_D5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_D6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_DO5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_DO6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_D_CY;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_D_XOR;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_A;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_A1;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_A2;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_A3;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_A4;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_A5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_A6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_AO5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_AO6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_AQ;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_A_CY;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_A_XOR;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_B;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_B1;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_B2;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_B3;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_B4;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_B5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_B6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_BO5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_BO6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_BQ;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_B_CY;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_B_XOR;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_C;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_C1;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_C2;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_C3;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_C4;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_C5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_C6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_CLK;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_CO5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_CO6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_C_CY;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_C_XOR;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_D;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_D1;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_D2;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_D3;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_D4;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_D5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_D6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_DO5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_DO6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_D_CY;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_D_XOR;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_A;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_A1;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_A2;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_A3;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_A4;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_A5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_A6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_AMUX;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_AO5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_AO6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_A_CY;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_A_XOR;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_B;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_B1;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_B2;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_B3;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_B4;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_B5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_B6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_BO5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_BO6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_B_CY;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_B_XOR;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_C;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_C1;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_C2;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_C3;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_C4;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_C5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_C6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_CMUX;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_CO5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_CO6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_C_CY;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_C_XOR;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_D;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_D1;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_D2;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_D3;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_D4;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_D5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_D6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_DO5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_DO6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_D_CY;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_D_XOR;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_A;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_A1;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_A2;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_A3;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_A4;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_A5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_A5Q;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_A6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_AMUX;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_AO5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_AO6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_AQ;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_AX;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_A_CY;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_A_XOR;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_B;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_B1;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_B2;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_B3;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_B4;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_B5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_B6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_BMUX;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_BO5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_BO6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_B_CY;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_B_XOR;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_C;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_C1;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_C2;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_C3;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_C4;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_C5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_C6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_CLK;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_CO5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_CO6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_CQ;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_C_CY;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_C_XOR;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_D;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_D1;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_D2;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_D3;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_D4;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_D5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_D5Q;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_D6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_DMUX;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_DO5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_DO6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_DQ;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_D_CY;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_D_XOR;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_A;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_A1;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_A2;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_A3;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_A4;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_A5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_A5Q;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_A6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_AMUX;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_AO5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_AO6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_AQ;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_AX;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_A_CY;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_A_XOR;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_B;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_B1;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_B2;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_B3;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_B4;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_B5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_B6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_BO5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_BO6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_BQ;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_B_CY;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_B_XOR;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_C;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_C1;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_C2;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_C3;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_C4;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_C5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_C6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_CLK;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_CO5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_CO6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_CQ;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_C_CY;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_C_XOR;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_D;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_D1;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_D2;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_D3;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_D4;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_D5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_D6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_DO5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_DO6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_D_CY;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_D_XOR;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_A;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_A1;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_A2;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_A3;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_A4;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_A5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_A6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_AMUX;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_AO5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_AO6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_A_CY;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_A_XOR;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_B;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_B1;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_B2;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_B3;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_B4;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_B5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_B6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_BO5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_BO6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_B_CY;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_B_XOR;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_C;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_C1;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_C2;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_C3;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_C4;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_C5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_C6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_CO5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_CO6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_C_CY;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_C_XOR;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_D;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_D1;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_D2;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_D3;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_D4;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_D5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_D6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_DO5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_DO6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_D_CY;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_D_XOR;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_A;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_A1;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_A2;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_A3;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_A4;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_A5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_A6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_AO5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_AO6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_AQ;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_A_CY;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_A_XOR;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_B;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_B1;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_B2;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_B3;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_B4;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_B5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_B6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_BO5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_BO6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_BQ;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_B_CY;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_B_XOR;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_C;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_C1;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_C2;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_C3;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_C4;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_C5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_C5Q;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_C6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_CLK;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_CMUX;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_CO5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_CO6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_CQ;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_C_CY;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_C_XOR;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_D;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_D1;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_D2;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_D3;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_D4;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_D5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_D6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_DO5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_DO6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_D_CY;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_D_XOR;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_A;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_A1;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_A2;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_A3;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_A4;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_A5;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_A6;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_AMUX;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_AO5;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_AO6;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_A_CY;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_A_XOR;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_B;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_B1;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_B2;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_B3;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_B4;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_B5;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_B5Q;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_B6;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_BMUX;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_BO5;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_BO6;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_BQ;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_B_CY;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_B_XOR;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_C;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_C1;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_C2;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_C3;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_C4;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_C5;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_C5Q;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_C6;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_CLK;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_CMUX;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_CO5;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_CO6;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_CQ;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_C_CY;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_C_XOR;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_D;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_D1;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_D2;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_D3;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_D4;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_D5;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_D6;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_DO5;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_DO6;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_D_CY;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X14Y112_D_XOR;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_A;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_A1;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_A2;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_A3;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_A4;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_A5;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_A6;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_AO5;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_AO6;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_AQ;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_A_CY;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_A_XOR;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_B;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_B1;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_B2;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_B3;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_B4;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_B5;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_B6;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_BO5;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_BO6;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_BQ;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_B_CY;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_B_XOR;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_C;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_C1;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_C2;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_C3;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_C4;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_C5;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_C6;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_CLK;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_CO5;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_CO6;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_C_CY;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_C_XOR;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_D;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_D1;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_D2;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_D3;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_D4;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_D5;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_D6;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_DO5;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_DO6;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_D_CY;
  wire [0:0] CLBLM_R_X11Y112_SLICE_X15Y112_D_XOR;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_A;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_A1;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_A2;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_A3;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_A4;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_A5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_A6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_AO5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_AO6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_AQ;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_A_CY;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_A_XOR;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_B;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_B1;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_B2;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_B3;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_B4;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_B5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_B6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_BO5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_BO6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_BQ;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_B_CY;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_B_XOR;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_C;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_C1;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_C2;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_C3;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_C4;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_C5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_C6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_CLK;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_CO5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_CO6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_CQ;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_C_CY;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_C_XOR;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_D;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_D1;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_D2;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_D3;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_D4;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_D5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_D6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_DO5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_DQ;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_D_CY;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X14Y113_D_XOR;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_A;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_A1;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_A2;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_A3;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_A4;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_A5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_A6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_AO5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_AO6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_AQ;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_A_CY;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_A_XOR;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_B;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_B1;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_B2;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_B3;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_B4;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_B5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_B6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_BO5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_BO6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_BQ;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_B_CY;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_B_XOR;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_C;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_C1;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_C2;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_C3;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_C4;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_C5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_C6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_CLK;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_CO5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_CO6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_CQ;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_C_CY;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_C_XOR;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_D;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_D1;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_D2;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_D3;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_D4;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_D5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_D6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_DO5;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_DO6;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_DQ;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_D_CY;
  wire [0:0] CLBLM_R_X11Y113_SLICE_X15Y113_D_XOR;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_A;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_A1;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_A2;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_A3;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_A4;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_A5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_A6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_AO5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_AO6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_AQ;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_A_CY;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_A_XOR;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_B;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_B1;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_B2;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_B3;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_B4;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_B5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_B6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_BO5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_BO6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_BQ;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_B_CY;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_B_XOR;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_C;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_C1;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_C2;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_C3;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_C4;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_C5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_C6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_CLK;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_CO5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_CO6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_CQ;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_C_CY;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_C_XOR;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_D;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_D1;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_D2;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_D3;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_D4;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_D5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_D6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_DO5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_DO6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_DQ;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_D_CY;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X14Y114_D_XOR;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_A;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_A1;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_A2;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_A3;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_A4;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_A5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_A6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_AO5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_AO6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_A_CY;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_A_XOR;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_B;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_B1;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_B2;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_B3;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_B4;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_B5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_B6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_BO5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_BO6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_B_CY;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_B_XOR;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_C;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_C1;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_C2;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_C3;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_C4;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_C5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_C6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_CO5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_CO6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_C_CY;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_C_XOR;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_D;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_D1;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_D2;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_D3;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_D4;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_D5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_D6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_DO5;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_DO6;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_D_CY;
  wire [0:0] CLBLM_R_X11Y114_SLICE_X15Y114_D_XOR;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_A;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_A1;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_A2;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_A3;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_A4;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_A5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_A6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_AMUX;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_AO5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_AO6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_AQ;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_AX;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_A_CY;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_A_XOR;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_B;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_B1;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_B2;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_B3;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_B4;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_B5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_B6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_BMUX;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_BO5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_BO6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_BQ;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_BX;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_B_CY;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_B_XOR;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_C;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_C1;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_C2;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_C3;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_C4;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_C5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_C6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_CE;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_CLK;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_CO5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_CO6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_C_CY;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_C_XOR;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_D;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_D1;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_D2;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_D3;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_D4;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_D5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_D6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_DO5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_DO6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_D_CY;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_D_XOR;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X14Y115_SR;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_A;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_A1;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_A2;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_A3;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_A4;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_A5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_A6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_AO5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_AO6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_AQ;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_A_CY;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_A_XOR;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_B;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_B1;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_B2;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_B3;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_B4;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_B5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_B5Q;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_B6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_BMUX;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_BO5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_BO6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_BQ;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_B_CY;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_B_XOR;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_C;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_C1;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_C2;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_C3;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_C4;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_C5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_C6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_CLK;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_CO5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_CO6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_CQ;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_C_CY;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_C_XOR;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_D;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_D1;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_D2;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_D3;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_D4;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_D5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_D6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_DMUX;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_DO5;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_DO6;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_D_CY;
  wire [0:0] CLBLM_R_X11Y115_SLICE_X15Y115_D_XOR;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_A;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_A1;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_A2;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_A3;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_A4;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_A5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_A5Q;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_A6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_AMUX;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_AO5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_AO6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_AQ;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_AX;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_A_CY;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_A_XOR;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_B;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_B1;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_B2;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_B3;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_B4;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_B5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_B6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_BO5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_BO6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_BQ;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_B_CY;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_B_XOR;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_C;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_C1;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_C2;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_C3;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_C4;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_C5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_C6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_CLK;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_CO5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_CO6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_C_CY;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_C_XOR;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_D;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_D1;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_D2;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_D3;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_D4;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_D5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_D6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_DO5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_DO6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_D_CY;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X14Y116_D_XOR;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_A;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_A1;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_A2;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_A3;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_A4;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_A5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_A6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_AO5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_AO6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_AQ;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_A_CY;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_A_XOR;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_B;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_B1;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_B2;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_B3;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_B4;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_B5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_B6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_BO5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_BO6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_B_CY;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_B_XOR;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_C;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_C1;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_C2;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_C3;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_C4;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_C5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_C6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_CLK;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_CO5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_CO6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_C_CY;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_C_XOR;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_D;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_D1;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_D2;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_D3;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_D4;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_D5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_D6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_DO5;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_DO6;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_D_CY;
  wire [0:0] CLBLM_R_X11Y116_SLICE_X15Y116_D_XOR;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_A;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_A1;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_A2;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_A3;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_A4;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_A5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_A6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_AO5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_AO6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_A_CY;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_A_XOR;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_B;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_B1;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_B2;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_B3;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_B4;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_B5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_B6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_BO5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_BO6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_B_CY;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_B_XOR;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_C;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_C1;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_C2;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_C3;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_C4;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_C5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_C6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_CO5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_CO6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_C_CY;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_C_XOR;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_D;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_D1;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_D2;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_D3;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_D4;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_D5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_D6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_DO5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_DO6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_D_CY;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X14Y117_D_XOR;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_A;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_A1;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_A2;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_A3;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_A4;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_A5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_A6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_AO5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_AO6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_AQ;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_A_CY;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_A_XOR;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_B;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_B1;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_B2;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_B3;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_B4;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_B5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_B6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_BMUX;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_BO5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_BO6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_B_CY;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_B_XOR;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_C;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_C1;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_C2;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_C3;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_C4;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_C5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_C6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_CLK;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_CO5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_CO6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_CQ;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_C_CY;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_C_XOR;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_D;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_D1;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_D2;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_D3;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_D4;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_D5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_D6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_DO5;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_DO6;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_DQ;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_D_CY;
  wire [0:0] CLBLM_R_X11Y117_SLICE_X15Y117_D_XOR;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_A;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_A1;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_A2;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_A3;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_A4;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_A5;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_A6;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_AO5;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_AO6;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_A_CY;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_A_XOR;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_B;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_B1;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_B2;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_B3;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_B4;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_B5;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_B6;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_BO5;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_BO6;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_B_CY;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_B_XOR;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_C;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_C1;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_C2;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_C3;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_C4;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_C5;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_C6;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_CO5;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_CO6;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_C_CY;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_C_XOR;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_D;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_D1;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_D2;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_D3;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_D4;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_D5;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_D6;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_DO5;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_DO6;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_D_CY;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X14Y118_D_XOR;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_A;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_A1;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_A2;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_A3;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_A4;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_A5;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_A5Q;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_A6;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_AMUX;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_AO5;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_AO6;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_AQ;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_A_CY;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_A_XOR;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_B;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_B1;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_B2;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_B3;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_B4;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_B5;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_B6;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_BO5;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_BO6;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_B_CY;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_B_XOR;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_C;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_C1;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_C2;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_C3;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_C4;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_C5;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_C6;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_CLK;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_CO5;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_CO6;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_C_CY;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_C_XOR;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_D;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_D1;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_D2;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_D3;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_D4;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_D5;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_D6;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_DO5;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_DO6;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_D_CY;
  wire [0:0] CLBLM_R_X11Y118_SLICE_X15Y118_D_XOR;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_A;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_A1;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_A2;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_A3;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_A4;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_A5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_A6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_AO5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_AO6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_AQ;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_A_CY;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_A_XOR;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_B;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_B1;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_B2;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_B3;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_B4;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_B5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_B6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_BO5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_BO6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_B_CY;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_B_XOR;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_C;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_C1;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_C2;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_C3;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_C4;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_C5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_C6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_CLK;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_CO5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_CO6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_C_CY;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_C_XOR;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_D;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_D1;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_D2;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_D3;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_D4;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_D5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_D6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_DO5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_DO6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_D_CY;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_D_XOR;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_A;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_A1;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_A2;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_A3;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_A4;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_A5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_A6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_AO5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_AO6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_A_CY;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_A_XOR;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_B;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_B1;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_B2;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_B3;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_B4;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_B5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_B6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_BO5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_BO6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_B_CY;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_B_XOR;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_C;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_C1;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_C2;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_C3;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_C4;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_C5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_C6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_CO5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_CO6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_C_CY;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_C_XOR;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_D;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_D1;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_D2;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_D3;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_D4;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_D5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_D6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_DO5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_DO6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_D_CY;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_D_XOR;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_A;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_A1;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_A2;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_A3;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_A4;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_A5;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_A6;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_AO5;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_AO6;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_A_CY;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_A_XOR;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_B;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_B1;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_B2;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_B3;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_B4;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_B5;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_B6;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_BO5;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_BO6;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_B_CY;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_B_XOR;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_C;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_C1;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_C2;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_C3;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_C4;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_C5;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_C6;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_CO5;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_CO6;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_C_CY;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_C_XOR;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_D;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_D1;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_D2;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_D3;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_D4;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_D5;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_D6;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_DO5;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_DO6;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_D_CY;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X18Y106_D_XOR;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_A;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_A1;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_A2;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_A3;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_A4;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_A5;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_A6;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_AO5;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_AO6;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_A_CY;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_A_XOR;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_B;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_B1;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_B2;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_B3;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_B4;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_B5;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_B6;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_BO5;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_BO6;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_B_CY;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_B_XOR;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_C;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_C1;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_C2;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_C3;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_C4;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_C5;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_C6;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_CO5;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_CO6;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_C_CY;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_C_XOR;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_D;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_D1;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_D2;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_D3;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_D4;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_D5;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_D6;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_DO5;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_DO6;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_D_CY;
  wire [0:0] CLBLM_R_X13Y106_SLICE_X19Y106_D_XOR;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_A;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_A1;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_A2;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_A3;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_A4;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_A5;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_A6;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_AO5;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_AO6;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_AQ;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_A_CY;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_A_XOR;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_B;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_B1;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_B2;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_B3;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_B4;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_B5;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_B6;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_BMUX;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_BO5;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_BO6;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_B_CY;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_B_XOR;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_C;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_C1;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_C2;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_C3;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_C4;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_C5;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_C6;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_CLK;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_CO5;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_CO6;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_C_CY;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_C_XOR;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_D;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_D1;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_D2;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_D3;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_D4;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_D5;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_D6;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_DO5;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_DO6;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_D_CY;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X18Y107_D_XOR;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_A;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_A1;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_A2;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_A3;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_A4;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_A5;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_A6;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_AO5;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_AO6;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_AQ;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_A_CY;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_A_XOR;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_B;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_B1;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_B2;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_B3;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_B4;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_B5;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_B6;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_BO5;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_BO6;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_BQ;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_B_CY;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_B_XOR;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_C;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_C1;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_C2;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_C3;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_C4;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_C5;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_C6;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_CLK;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_CO5;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_CO6;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_C_CY;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_C_XOR;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_D;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_D1;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_D2;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_D3;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_D4;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_D5;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_D6;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_DO5;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_DO6;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_D_CY;
  wire [0:0] CLBLM_R_X13Y107_SLICE_X19Y107_D_XOR;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_A;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_A1;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_A2;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_A3;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_A4;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_A5;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_A6;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_AO5;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_AO6;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_AQ;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_A_CY;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_A_XOR;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_B;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_B1;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_B2;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_B3;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_B4;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_B5;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_B6;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_BMUX;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_BO5;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_BO6;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_B_CY;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_B_XOR;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_C;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_C1;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_C2;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_C3;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_C4;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_C5;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_C6;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_CLK;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_CMUX;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_CO5;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_CO6;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_C_CY;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_C_XOR;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_D;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_D1;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_D2;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_D3;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_D4;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_D5;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_D6;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_DO5;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_DO6;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_D_CY;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X18Y108_D_XOR;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_A;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_A1;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_A2;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_A3;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_A4;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_A5;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_A6;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_AO5;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_AO6;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_AQ;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_A_CY;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_A_XOR;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_B;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_B1;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_B2;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_B3;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_B4;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_B5;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_B6;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_BO5;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_BO6;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_BQ;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_B_CY;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_B_XOR;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_C;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_C1;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_C2;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_C3;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_C4;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_C5;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_C6;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_CLK;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_CO5;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_CO6;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_C_CY;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_C_XOR;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_D;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_D1;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_D2;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_D3;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_D4;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_D5;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_D6;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_DO5;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_DO6;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_D_CY;
  wire [0:0] CLBLM_R_X13Y108_SLICE_X19Y108_D_XOR;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_A;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_A1;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_A2;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_A3;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_A4;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_A5;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_A6;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_AO5;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_AO6;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_AQ;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_A_CY;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_A_XOR;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_B;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_B1;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_B2;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_B3;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_B4;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_B5;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_B6;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_BMUX;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_BO5;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_BO6;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_B_CY;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_B_XOR;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_C;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_C1;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_C2;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_C3;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_C4;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_C5;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_C6;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_CLK;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_CO5;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_CO6;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_C_CY;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_C_XOR;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_D;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_D1;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_D2;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_D3;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_D4;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_D5;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_D6;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_DO5;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_DO6;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_D_CY;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X18Y109_D_XOR;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_A;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_A1;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_A2;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_A3;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_A4;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_A5;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_A6;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_AO5;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_AO6;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_AQ;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_A_CY;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_A_XOR;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_B;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_B1;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_B2;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_B3;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_B4;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_B5;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_B6;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_BO5;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_BO6;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_BQ;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_B_CY;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_B_XOR;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_C;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_C1;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_C2;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_C3;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_C4;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_C5;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_C6;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_CLK;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_CO5;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_CO6;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_C_CY;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_C_XOR;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_D;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_D1;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_D2;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_D3;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_D4;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_D5;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_D6;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_DO5;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_DO6;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_D_CY;
  wire [0:0] CLBLM_R_X13Y109_SLICE_X19Y109_D_XOR;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_A;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_A1;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_A2;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_A3;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_A4;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_A5;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_A6;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_AO5;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_AO6;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_AQ;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_A_CY;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_A_XOR;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_B;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_B1;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_B2;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_B3;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_B4;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_B5;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_B6;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_BO5;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_BO6;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_BQ;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_B_CY;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_B_XOR;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_C;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_C1;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_C2;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_C3;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_C4;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_C5;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_C6;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_CLK;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_CO5;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_CO6;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_CQ;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_C_CY;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_C_XOR;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_D;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_D1;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_D2;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_D3;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_D4;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_D5;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_D6;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_DMUX;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_DO5;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_DO6;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_D_CY;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X18Y110_D_XOR;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_A;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_A1;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_A2;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_A3;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_A4;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_A5;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_A6;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_AO5;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_AO6;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_AQ;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_A_CY;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_A_XOR;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_B;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_B1;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_B2;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_B3;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_B4;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_B5;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_B6;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_BO5;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_BO6;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_BQ;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_B_CY;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_B_XOR;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_C;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_C1;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_C2;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_C3;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_C4;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_C5;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_C6;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_CLK;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_CO5;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_CO6;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_CQ;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_C_CY;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_C_XOR;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_D;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_D1;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_D2;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_D3;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_D4;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_D5;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_D6;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_DO5;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_DO6;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_D_CY;
  wire [0:0] CLBLM_R_X13Y110_SLICE_X19Y110_D_XOR;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_A;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_A1;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_A2;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_A3;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_A4;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_A5;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_A5Q;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_A6;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_AMUX;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_AO5;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_AO6;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_AQ;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_A_CY;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_A_XOR;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_B;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_B1;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_B2;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_B3;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_B4;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_B5;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_B6;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_BO5;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_BO6;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_BQ;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_B_CY;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_B_XOR;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_C;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_C1;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_C2;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_C3;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_C4;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_C5;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_C6;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_CLK;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_CO5;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_CO6;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_CQ;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_C_CY;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_C_XOR;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_D;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_D1;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_D2;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_D3;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_D4;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_D5;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_D6;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_DO5;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_DO6;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_D_CY;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X18Y112_D_XOR;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_A;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_A1;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_A2;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_A3;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_A4;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_A5;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_A6;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_AO5;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_AO6;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_A_CY;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_A_XOR;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_B;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_B1;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_B2;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_B3;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_B4;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_B5;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_B6;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_BO5;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_BO6;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_B_CY;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_B_XOR;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_C;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_C1;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_C2;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_C3;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_C4;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_C5;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_C6;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_CO5;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_CO6;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_C_CY;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_C_XOR;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_D;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_D1;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_D2;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_D3;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_D4;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_D5;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_D6;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_DO5;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_DO6;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_D_CY;
  wire [0:0] CLBLM_R_X13Y112_SLICE_X19Y112_D_XOR;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_A;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_A1;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_A2;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_A3;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_A4;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_A5;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_A6;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_AO5;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_AO6;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_AQ;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_A_CY;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_A_XOR;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_B;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_B1;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_B2;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_B3;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_B4;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_B5;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_B6;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_BO5;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_BO6;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_BQ;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_B_CY;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_B_XOR;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_C;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_C1;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_C2;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_C3;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_C4;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_C5;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_C6;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_CLK;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_CO5;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_CO6;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_CQ;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_C_CY;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_C_XOR;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_D;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_D1;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_D2;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_D3;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_D4;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_D5;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_D6;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_DO5;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_DO6;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_D_CY;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X18Y113_D_XOR;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_A;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_A1;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_A2;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_A3;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_A4;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_A5;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_A6;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_AO5;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_AO6;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_AQ;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_A_CY;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_A_XOR;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_B;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_B1;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_B2;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_B3;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_B4;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_B5;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_B6;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_BO5;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_BO6;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_B_CY;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_B_XOR;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_C;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_C1;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_C2;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_C3;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_C4;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_C5;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_C6;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_CLK;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_CO5;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_CO6;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_C_CY;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_C_XOR;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_D;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_D1;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_D2;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_D3;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_D4;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_D5;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_D6;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_DO5;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_DO6;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_D_CY;
  wire [0:0] CLBLM_R_X13Y113_SLICE_X19Y113_D_XOR;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_A;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_A1;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_A2;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_A3;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_A4;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_A5;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_A6;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_AMUX;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_AO5;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_AO6;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_AQ;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_AX;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_A_CY;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_A_XOR;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_B;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_B1;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_B2;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_B3;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_B4;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_B5;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_B6;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_BO5;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_BO6;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_BQ;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_BX;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_B_CY;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_B_XOR;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_C;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_C1;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_C2;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_C3;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_C4;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_C5;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_C6;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_CLK;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_CO5;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_CO6;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_C_CY;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_C_XOR;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_D;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_D1;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_D2;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_D3;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_D4;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_D5;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_D6;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_DO5;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_DO6;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_D_CY;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X18Y117_D_XOR;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_A;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_A1;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_A2;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_A3;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_A4;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_A5;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_A6;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_AO5;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_AO6;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_A_CY;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_A_XOR;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_B;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_B1;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_B2;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_B3;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_B4;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_B5;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_B6;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_BO5;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_BO6;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_B_CY;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_B_XOR;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_C;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_C1;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_C2;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_C3;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_C4;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_C5;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_C6;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_CO5;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_CO6;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_C_CY;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_C_XOR;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_D;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_D1;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_D2;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_D3;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_D4;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_D5;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_D6;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_DO5;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_DO6;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_D_CY;
  wire [0:0] CLBLM_R_X13Y117_SLICE_X19Y117_D_XOR;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_A;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_A1;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_A2;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_A3;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_A4;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_A5;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_A6;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_AMUX;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_AO5;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_AO6;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_A_CY;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_A_XOR;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_B;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_B1;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_B2;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_B3;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_B4;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_B5;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_B6;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_BO5;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_BO6;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_B_CY;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_B_XOR;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_C;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_C1;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_C2;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_C3;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_C4;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_C5;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_C6;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_CO5;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_CO6;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_C_CY;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_C_XOR;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_D;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_D1;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_D2;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_D3;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_D4;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_D5;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_D6;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_DO5;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_DO6;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_D_CY;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X18Y118_D_XOR;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_A;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_A1;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_A2;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_A3;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_A4;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_A5;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_A6;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_AO5;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_AO6;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_A_CY;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_A_XOR;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_B;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_B1;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_B2;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_B3;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_B4;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_B5;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_B6;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_BO5;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_BO6;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_B_CY;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_B_XOR;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_C;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_C1;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_C2;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_C3;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_C4;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_C5;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_C6;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_CO5;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_CO6;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_C_CY;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_C_XOR;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_D;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_D1;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_D2;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_D3;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_D4;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_D5;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_D6;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_DO5;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_DO6;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_D_CY;
  wire [0:0] CLBLM_R_X13Y118_SLICE_X19Y118_D_XOR;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X56Y117_A;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X56Y117_A1;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X56Y117_A2;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X56Y117_A3;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X56Y117_A4;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X56Y117_A5;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X56Y117_A6;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X56Y117_AO5;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X56Y117_AO6;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X56Y117_A_CY;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X56Y117_A_XOR;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X56Y117_B;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X56Y117_B1;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X56Y117_B2;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X56Y117_B3;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X56Y117_B4;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X56Y117_B5;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X56Y117_B6;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X56Y117_BO5;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X56Y117_BO6;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X56Y117_B_CY;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X56Y117_B_XOR;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X56Y117_C;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X56Y117_C1;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X56Y117_C2;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X56Y117_C3;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X56Y117_C4;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X56Y117_C5;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X56Y117_C6;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X56Y117_CO5;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X56Y117_CO6;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X56Y117_C_CY;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X56Y117_C_XOR;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X56Y117_D;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X56Y117_D1;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X56Y117_D2;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X56Y117_D3;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X56Y117_D4;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X56Y117_D5;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X56Y117_D6;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X56Y117_DO5;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X56Y117_DO6;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X56Y117_D_CY;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X56Y117_D_XOR;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X57Y117_A;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X57Y117_A1;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X57Y117_A2;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X57Y117_A3;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X57Y117_A4;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X57Y117_A5;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X57Y117_A6;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X57Y117_AO5;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X57Y117_AO6;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X57Y117_A_CY;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X57Y117_A_XOR;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X57Y117_B;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X57Y117_B1;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X57Y117_B2;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X57Y117_B3;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X57Y117_B4;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X57Y117_B5;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X57Y117_B6;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X57Y117_BO5;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X57Y117_BO6;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X57Y117_B_CY;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X57Y117_B_XOR;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X57Y117_C;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X57Y117_C1;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X57Y117_C2;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X57Y117_C3;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X57Y117_C4;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X57Y117_C5;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X57Y117_C6;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X57Y117_CO5;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X57Y117_CO6;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X57Y117_C_CY;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X57Y117_C_XOR;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X57Y117_D;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X57Y117_D1;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X57Y117_D2;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X57Y117_D3;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X57Y117_D4;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X57Y117_D5;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X57Y117_D6;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X57Y117_DO5;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X57Y117_DO6;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X57Y117_D_CY;
  wire [0:0] CLBLM_R_X37Y117_SLICE_X57Y117_D_XOR;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_A;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_A1;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_A2;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_A3;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_A4;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_A5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_A6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_AO5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_AO6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_A_CY;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_A_XOR;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_B;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_B1;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_B2;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_B3;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_B4;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_B5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_B6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_BO5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_BO6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_B_CY;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_B_XOR;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_C;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_C1;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_C2;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_C3;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_C4;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_C5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_C6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_CO5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_CO6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_C_CY;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_C_XOR;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_D;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_D1;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_D2;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_D3;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_D4;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_D5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_D6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_DO5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_DO6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_D_CY;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_D_XOR;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_A;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_A1;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_A2;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_A3;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_A4;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_A5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_A6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_AO5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_AO6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_A_CY;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_A_XOR;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_B;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_B1;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_B2;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_B3;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_B4;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_B5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_B6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_BO5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_BO6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_B_CY;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_B_XOR;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_C;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_C1;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_C2;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_C3;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_C4;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_C5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_C6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_CO5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_CO6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_C_CY;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_C_XOR;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_D;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_D1;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_D2;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_D3;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_D4;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_D5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_D6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_DO5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_DO6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_D_CY;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_D_XOR;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_A;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_A1;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_A2;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_A3;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_A4;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_A5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_A6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_AO5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_AO6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_A_CY;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_A_XOR;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_B;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_B1;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_B2;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_B3;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_B4;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_B5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_B6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_BO5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_BO6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_B_CY;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_B_XOR;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_C;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_C1;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_C2;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_C3;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_C4;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_C5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_C6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_CO5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_CO6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_C_CY;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_C_XOR;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_D;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_D1;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_D2;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_D3;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_D4;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_D5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_D6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_DO5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_DO6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_D_CY;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_D_XOR;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_A;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_A1;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_A2;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_A3;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_A4;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_A5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_A6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_AO5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_AO6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_AQ;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_A_CY;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_A_XOR;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_B;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_B1;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_B2;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_B3;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_B4;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_B5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_B6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_BMUX;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_BO5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_BO6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_B_CY;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_B_XOR;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_C;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_C1;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_C2;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_C3;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_C4;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_C5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_C6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_CLK;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_CO5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_CO6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_C_CY;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_C_XOR;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_D;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_D1;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_D2;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_D3;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_D4;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_D5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_D6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_DO5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_DO6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_D_CY;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_D_XOR;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_A;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_A1;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_A2;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_A3;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_A4;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_A5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_A6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_AO5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_AO6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_A_CY;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_A_XOR;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_B;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_B1;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_B2;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_B3;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_B4;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_B5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_B6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_BO5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_BO6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_B_CY;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_B_XOR;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_C;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_C1;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_C2;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_C3;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_C4;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_C5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_C6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_CMUX;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_CO5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_CO6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_C_CY;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_C_XOR;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_D;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_D1;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_D2;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_D3;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_D4;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_D5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_D6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_DMUX;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_DO5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_DO6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_D_CY;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_D_XOR;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_A;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_A1;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_A2;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_A3;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_A4;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_A5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_A6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_AO5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_AO6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_A_CY;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_A_XOR;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_B;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_B1;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_B2;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_B3;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_B4;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_B5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_B6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_BO5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_BO6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_B_CY;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_B_XOR;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_C;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_C1;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_C2;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_C3;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_C4;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_C5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_C6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_CO5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_CO6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_C_CY;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_C_XOR;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_D;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_D1;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_D2;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_D3;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_D4;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_D5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_D6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_DMUX;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_DO5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_DO6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_D_CY;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_D_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A5Q;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_AMUX;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_AO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_AO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_AQ;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_BO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_BO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_CLK;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_CMUX;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_CO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_CO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_DMUX;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_DO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_DO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_AO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_AO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_BO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_BO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_CO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_CO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_DO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_DO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D_XOR;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A1;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A2;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A3;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A4;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_AMUX;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_AO5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_AO6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A_CY;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A_XOR;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B1;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B2;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B3;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B4;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_BO5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_BO6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B_CY;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B_XOR;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C1;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C2;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C3;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C4;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_CO5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_CO6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C_CY;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C_XOR;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D1;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D2;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D3;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D4;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_DMUX;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_DO5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_DO6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D_CY;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D_XOR;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A1;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A2;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A3;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A4;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_AO5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_AO6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A_CY;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A_XOR;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B1;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B2;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B3;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B4;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_BO5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_BO6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B_CY;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B_XOR;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C1;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C2;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C3;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C4;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_CO5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_CO6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C_CY;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C_XOR;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D1;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D2;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D3;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D4;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_DO5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_DO6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D_CY;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D_XOR;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A1;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A2;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A3;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A4;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_AO5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_AO6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A_CY;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A_XOR;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B1;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B2;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B3;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B4;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_BO5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_BO6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B_CY;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B_XOR;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C1;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C2;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C3;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C4;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_CO5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_CO6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C_CY;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C_XOR;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D1;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D2;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D3;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D4;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_DMUX;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_DO5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_DO6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D_CY;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D_XOR;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A1;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A2;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A3;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A4;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_AO5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_AO6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A_CY;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A_XOR;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B1;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B2;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B3;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B4;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_BO5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_BO6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B_CY;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B_XOR;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C1;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C2;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C3;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C4;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_CO5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_CO6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C_CY;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C_XOR;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D1;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D2;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D3;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D4;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_DO5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_DO6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D_CY;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_AMUX;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_AO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_AO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_BO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_BO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_CO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_CO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_DO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_DO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_AO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_AO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_AQ;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_BMUX;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_BO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_BO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_CLK;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_CO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_CO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_DO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_DO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D_XOR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A1;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A2;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A3;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A4;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_AO5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_AO6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A_CY;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A_XOR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B1;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B2;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B3;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B4;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_BO5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_BO6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B_CY;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B_XOR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C1;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C2;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C3;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C4;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_CO5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_CO6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C_CY;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C_XOR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D1;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D2;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D3;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D4;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_DO5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_DO6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D_CY;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D_XOR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A1;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A2;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A3;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A4;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_AO5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_AO6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_AQ;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A_CY;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A_XOR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B1;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B2;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B3;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B4;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_BO5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_BO6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B_CY;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B_XOR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C1;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C2;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C3;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C4;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_CLK;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_CO5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_CO6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C_CY;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C_XOR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D1;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D2;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D3;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D4;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_DO5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_DO6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D_CY;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D_XOR;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A1;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A2;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A3;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A4;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_AO5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_AO6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_AQ;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A_CY;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_A_XOR;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B1;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B2;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B3;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B4;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_BO5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_BO6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_BQ;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B_CY;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_B_XOR;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C1;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C2;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C3;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C4;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_CLK;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_CMUX;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_CO5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_CO6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C_CY;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_C_XOR;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D1;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D2;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D3;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D4;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_DO5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_DO6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D_CY;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X2Y114_D_XOR;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A1;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A2;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A3;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A4;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_AO5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_AO6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A_CY;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_A_XOR;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B1;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B2;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B3;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B4;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_BO5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_BO6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B_CY;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_B_XOR;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C1;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C2;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C3;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C4;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_CMUX;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_CO5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_CO6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C_CY;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_C_XOR;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D1;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D2;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D3;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D4;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_DO5;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_DO6;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D_CY;
  wire [0:0] CLBLM_R_X3Y114_SLICE_X3Y114_D_XOR;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A1;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A2;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A3;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A4;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_AMUX;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_AO5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_AO6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_AQ;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A_CY;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_A_XOR;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B1;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B2;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B3;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B4;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_BO5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_BO6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B_CY;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_B_XOR;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C1;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C2;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C3;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C4;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_CLK;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_CMUX;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_CO5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_CO6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C_CY;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_C_XOR;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D1;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D2;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D3;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D4;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_DO5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_DO6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D_CY;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X2Y115_D_XOR;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A1;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A2;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A3;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A4;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_AMUX;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_AO5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_AO6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A_CY;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_A_XOR;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B1;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B2;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B3;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B4;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_BMUX;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_BO5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_BO6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B_CY;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_B_XOR;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C1;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C2;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C3;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C4;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_CMUX;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_CO5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_CO6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C_CY;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_C_XOR;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D1;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D2;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D3;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D4;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_DMUX;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_DO5;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_DO6;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D_CY;
  wire [0:0] CLBLM_R_X3Y115_SLICE_X3Y115_D_XOR;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_A;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_A1;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_A2;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_A3;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_A4;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_A5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_A6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_AMUX;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_AO5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_AO6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_A_CY;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_A_XOR;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_B;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_B1;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_B2;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_B3;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_B4;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_B5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_B6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_BO5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_BO6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_B_CY;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_B_XOR;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_C;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_C1;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_C2;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_C3;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_C4;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_C5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_C6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_CO5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_CO6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_C_CY;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_C_XOR;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_D;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_D1;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_D2;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_D3;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_D4;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_D5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_D6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_DO5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_DO6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_D_CY;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X2Y116_D_XOR;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_A;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_A1;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_A2;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_A3;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_A4;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_A5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_A6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_AO5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_AO6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_A_CY;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_A_XOR;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_B;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_B1;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_B2;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_B3;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_B4;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_B5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_B6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_BO5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_BO6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_B_CY;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_B_XOR;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_C;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_C1;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_C2;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_C3;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_C4;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_C5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_C6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_CO5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_CO6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_C_CY;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_C_XOR;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_D;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_D1;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_D2;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_D3;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_D4;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_D5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_D6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_DO5;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_DO6;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_D_CY;
  wire [0:0] CLBLM_R_X3Y116_SLICE_X3Y116_D_XOR;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A1;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A2;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A3;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A4;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_AO5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_AO6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A_CY;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A_XOR;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B1;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B2;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B3;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B4;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_BO5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_BO6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B_CY;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B_XOR;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C1;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C2;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C3;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C4;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_CO5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_CO6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C_CY;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C_XOR;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D1;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D2;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D3;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D4;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_DO5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_DO6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D_CY;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D_XOR;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A1;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A2;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A3;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A4;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_AO5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_AO6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A_CY;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A_XOR;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B1;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B2;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B3;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B4;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_BO5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_BO6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B_CY;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B_XOR;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C1;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C2;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C3;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C4;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_CO5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_CO6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C_CY;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C_XOR;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D1;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D2;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D3;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D4;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_DO5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_DO6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D_CY;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D_XOR;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_A;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_A1;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_A2;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_A3;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_A4;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_A5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_A6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_AO5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_AO6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_AQ;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_A_CY;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_A_XOR;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_B;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_B1;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_B2;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_B3;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_B4;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_B5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_B6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_BO5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_BO6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_BQ;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_B_CY;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_B_XOR;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_C;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_C1;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_C2;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_C3;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_C4;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_C5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_C6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_CLK;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_CO5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_CO6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_C_CY;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_C_XOR;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_D;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_D1;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_D2;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_D3;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_D4;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_D5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_D6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_DO5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_DO6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_D_CY;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_D_XOR;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_A;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_A1;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_A2;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_A3;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_A4;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_A5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_A6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_AO5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_AO6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_AQ;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_A_CY;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_A_XOR;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_B;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_B1;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_B2;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_B3;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_B4;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_B5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_B6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_BO5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_BO6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_BQ;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_B_CY;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_B_XOR;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_C;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_C1;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_C2;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_C3;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_C4;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_C5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_C6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_CLK;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_CO5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_CO6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_C_CY;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_C_XOR;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_D;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_D1;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_D2;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_D3;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_D4;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_D5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_D6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_DO5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_DO6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_D_CY;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_D_XOR;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_A;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_A1;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_A2;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_A3;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_A4;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_A5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_A6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_AO5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_AO6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_AQ;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_A_CY;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_A_XOR;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_B;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_B1;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_B2;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_B3;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_B4;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_B5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_B6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_BO5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_BO6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_BQ;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_B_CY;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_B_XOR;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_C;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_C1;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_C2;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_C3;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_C4;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_C5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_C6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_CLK;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_CO5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_CO6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_CQ;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_C_CY;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_C_XOR;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_D;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_D1;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_D2;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_D3;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_D4;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_D5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_D6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_DO5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_DO6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_DQ;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_D_CY;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_D_XOR;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_A;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_A1;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_A2;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_A3;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_A4;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_A5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_A6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_AO5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_AO6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_AQ;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_A_CY;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_A_XOR;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_B;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_B1;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_B2;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_B3;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_B4;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_B5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_B6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_BMUX;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_BO5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_BO6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_B_CY;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_B_XOR;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_C;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_C1;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_C2;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_C3;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_C4;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_C5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_C6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_CLK;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_CO5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_CO6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_C_CY;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_C_XOR;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_D;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_D1;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_D2;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_D3;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_D4;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_D5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_D6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_DO5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_DO6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_D_CY;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_D_XOR;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_A;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_A1;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_A2;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_A3;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_A4;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_A5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_A6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_AO5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_AO6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_AQ;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_A_CY;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_A_XOR;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_B;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_B1;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_B2;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_B3;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_B4;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_B5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_B6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_BO5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_BO6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_BQ;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_B_CY;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_B_XOR;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_C;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_C1;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_C2;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_C3;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_C4;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_C5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_C6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_CLK;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_CO5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_CO6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_CQ;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_C_CY;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_C_XOR;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_D;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_D1;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_D2;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_D3;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_D4;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_D5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_D6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_DO5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_DO6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_DQ;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_D_CY;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_D_XOR;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_A;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_A1;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_A2;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_A3;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_A4;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_A5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_A6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_AO5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_AO6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_AQ;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_A_CY;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_A_XOR;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_B;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_B1;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_B2;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_B3;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_B4;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_B5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_B5Q;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_B6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_BMUX;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_BO5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_BO6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_BQ;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_B_CY;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_B_XOR;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_C;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_C1;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_C2;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_C3;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_C4;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_C5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_C6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_CLK;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_CMUX;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_CO5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_CO6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_C_CY;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_C_XOR;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_D;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_D1;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_D2;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_D3;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_D4;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_D5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_D6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_DMUX;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_DO5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_DO6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_D_CY;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_D_XOR;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_A;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_A1;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_A2;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_A3;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_A4;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_A5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_A6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_AO5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_AO6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_A_CY;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_A_XOR;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_B;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_B1;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_B2;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_B3;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_B4;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_B5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_B6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_BO5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_BO6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_B_CY;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_B_XOR;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_C;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_C1;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_C2;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_C3;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_C4;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_C5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_C6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_CO5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_CO6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_C_CY;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_C_XOR;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_D;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_D1;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_D2;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_D3;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_D4;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_D5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_D6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_DO5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_DO6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_D_CY;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_D_XOR;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_A;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_A1;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_A2;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_A3;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_A4;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_A5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_A6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_AO5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_AO6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_AQ;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_A_CY;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_A_XOR;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_B;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_B1;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_B2;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_B3;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_B4;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_B5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_B6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_BO5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_BO6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_B_CY;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_B_XOR;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_C;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_C1;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_C2;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_C3;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_C4;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_C5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_C6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_CLK;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_CO5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_CO6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_C_CY;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_C_XOR;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_D;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_D1;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_D2;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_D3;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_D4;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_D5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_D6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_DO5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_DO6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_D_CY;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_D_XOR;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A1;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A2;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A3;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A4;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_AO5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_AO6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_AQ;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A_CY;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A_XOR;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B1;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B2;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B3;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B4;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_BO5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_BO6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_BQ;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B_CY;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B_XOR;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C1;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C2;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C3;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C4;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_CLK;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_CO5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_CO6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_CQ;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C_CY;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C_XOR;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D1;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D2;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D3;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D4;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_DO5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_DO6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_DQ;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D_CY;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D_XOR;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A1;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A2;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A3;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A4;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A5Q;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_AMUX;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_AO5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_AO6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_AQ;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_AX;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A_CY;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A_XOR;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B1;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B2;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B3;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B4;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B5Q;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_BMUX;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_BO5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_BO6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_BQ;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_BX;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B_CY;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B_XOR;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C1;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C2;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C3;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C4;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_CLK;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_CMUX;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_CO5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_CO6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C_CY;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C_XOR;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D1;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D2;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D3;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D4;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_DO5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_DO6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_DQ;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D_CY;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D_XOR;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A1;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A2;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A3;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A4;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_AO5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_AO6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_AQ;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A_CY;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A_XOR;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B1;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B2;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B3;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B4;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B5Q;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_BMUX;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_BO5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_BO6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_BQ;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B_CY;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B_XOR;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C1;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C2;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C3;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C4;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_CLK;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_CO5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_CO6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_CQ;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C_CY;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C_XOR;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D1;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D2;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D3;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D4;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_DO5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_DO6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_DQ;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D_CY;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D_XOR;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A1;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A2;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A3;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A4;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_AO5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_AO6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_AQ;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A_CY;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A_XOR;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B1;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B2;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B3;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B4;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B5Q;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_BMUX;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_BO5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_BO6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_BQ;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B_CY;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B_XOR;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C1;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C2;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C3;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C4;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_CLK;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_CMUX;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_CO5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_CO6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C_CY;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C_XOR;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D1;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D2;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D3;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D4;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_DO5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_DO6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D_CY;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D_XOR;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A1;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A2;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A3;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A4;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_AO5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_AO6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_AQ;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A_CY;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A_XOR;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B1;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B2;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B3;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B4;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_BO5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_BO6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_BQ;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B_CY;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B_XOR;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C1;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C2;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C3;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C4;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_CLK;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_CO5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_CO6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_CQ;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C_CY;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C_XOR;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D1;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D2;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D3;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D4;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_DO5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_DO6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D_CY;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D_XOR;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A1;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A2;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A3;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A4;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_AO5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_AO6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_AQ;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A_CY;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A_XOR;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B1;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B2;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B3;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B4;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_BO5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_BO6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_BQ;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B_CY;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B_XOR;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C1;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C2;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C3;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C4;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_CLK;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_CO5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_CO6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_CQ;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C_CY;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C_XOR;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D1;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D2;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D3;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D4;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_DO5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_DO6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D_CY;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D_XOR;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A1;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A2;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A3;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A4;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_AO5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_AO6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_AQ;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A_CY;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A_XOR;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B1;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B2;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B3;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B4;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_BO5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_BO6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_BQ;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B_CY;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B_XOR;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C1;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C2;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C3;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C4;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_CLK;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_CO5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_CO6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_CQ;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C_CY;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C_XOR;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D1;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D2;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D3;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D4;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_DO5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_DO6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D_CY;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D_XOR;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A1;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A2;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A3;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A4;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_AO5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_AO6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_AQ;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A_CY;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A_XOR;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B1;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B2;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B3;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B4;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_BO5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_BO6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_BQ;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B_CY;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B_XOR;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C1;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C2;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C3;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C4;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_CLK;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_CO5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_CO6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_CQ;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C_CY;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C_XOR;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D1;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D2;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D3;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D4;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_DO5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_DO6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_DQ;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D_CY;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D_XOR;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A1;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A2;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A3;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A4;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_AO5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_AO6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_AQ;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A_CY;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A_XOR;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B1;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B2;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B3;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B4;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_BO5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_BO6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_BQ;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B_CY;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B_XOR;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C1;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C2;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C3;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C4;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_CLK;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_CO5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_CO6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_CQ;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C_CY;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C_XOR;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D1;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D2;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D3;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D4;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_DO5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_DO6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D_CY;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D_XOR;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A1;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A2;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A3;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A4;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_AO5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_AO6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_AQ;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A_CY;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A_XOR;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B1;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B2;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B3;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B4;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_BO5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_BO6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_BQ;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B_CY;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B_XOR;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C1;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C2;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C3;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C4;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_CLK;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_CO5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_CO6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C_CY;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C_XOR;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D1;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D2;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D3;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D4;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_DO5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_DO6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D_CY;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D_XOR;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_A;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_A1;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_A2;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_A3;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_A4;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_A5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_A6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_AO5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_AO6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_AQ;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_A_CY;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_A_XOR;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_B;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_B1;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_B2;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_B3;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_B4;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_B5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_B6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_BO5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_BO6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_B_CY;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_B_XOR;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_C;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_C1;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_C2;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_C3;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_C4;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_C5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_C6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_CLK;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_CO5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_CO6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_C_CY;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_C_XOR;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_D;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_D1;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_D2;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_D3;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_D4;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_D5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_D6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_DO5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_DO6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_D_CY;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_D_XOR;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_A;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_A1;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_A2;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_A3;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_A4;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_A5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_A6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_AO5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_AO6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_AQ;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_A_CY;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_A_XOR;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_B;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_B1;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_B2;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_B3;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_B4;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_B5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_B5Q;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_B6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_BMUX;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_BO5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_BO6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_BQ;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_B_CY;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_B_XOR;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_C;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_C1;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_C2;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_C3;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_C4;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_C5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_C5Q;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_C6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_CLK;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_CMUX;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_CO5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_CO6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_CQ;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_C_CY;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_C_XOR;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_D;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_D1;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_D2;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_D3;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_D4;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_D5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_D6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_DO5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_DO6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_D_CY;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_D_XOR;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A1;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A2;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A3;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A4;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_AO5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_AO6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_AQ;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A_CY;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A_XOR;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B1;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B2;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B3;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B4;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_BO5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_BO6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_BQ;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B_CY;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B_XOR;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C1;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C2;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C3;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C4;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_CLK;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_CO5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_CO6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_CQ;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C_CY;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C_XOR;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D1;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D2;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D3;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D4;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_DMUX;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_DO5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_DO6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D_CY;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D_XOR;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A1;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A2;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A3;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A4;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_AO5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_AO6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_AQ;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A_CY;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A_XOR;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B1;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B2;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B3;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B4;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_BO5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_BO6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_BQ;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B_CY;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B_XOR;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C1;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C2;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C3;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C4;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_CLK;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_CO5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_CO6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C_CY;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C_XOR;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D1;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D2;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D3;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D4;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_DO5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_DO6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D_CY;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D_XOR;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A1;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A2;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A3;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A4;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_AMUX;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_AO5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_AO6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A_CY;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A_XOR;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B1;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B2;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B3;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B4;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_BO5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_BO6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_BQ;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B_CY;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B_XOR;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C1;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C2;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C3;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C4;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_CLK;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_CO5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_CO6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_CQ;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C_CY;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C_XOR;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D1;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D2;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D3;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D4;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D5Q;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_DMUX;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_DO5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_DO6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_DQ;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D_CY;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D_XOR;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A1;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A2;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A3;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A4;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A5Q;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_AMUX;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_AO5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_AO6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_AQ;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_AX;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A_CY;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A_XOR;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B1;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B2;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B3;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B4;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_BO5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_BO6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_BQ;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B_CY;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B_XOR;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C1;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C2;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C3;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C4;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_CLK;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_CMUX;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_CO5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_CO6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C_CY;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C_XOR;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D1;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D2;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D3;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D4;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_DO5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D_CY;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D_XOR;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_A;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_A1;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_A2;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_A3;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_A4;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_A5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_A6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_AO5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_AO6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_A_CY;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_A_XOR;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_B;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_B1;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_B2;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_B3;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_B4;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_B5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_B6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_BO5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_BO6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_B_CY;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_B_XOR;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_C;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_C1;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_C2;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_C3;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_C4;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_C5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_C6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_CO5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_CO6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_C_CY;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_C_XOR;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_D;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_D1;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_D2;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_D3;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_D4;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_D5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_D6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_DO5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_DO6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_D_CY;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_D_XOR;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_A;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_A1;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_A2;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_A3;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_A4;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_A5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_A6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_AO5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_AO6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_AQ;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_A_CY;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_A_XOR;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_B;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_B1;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_B2;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_B3;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_B4;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_B5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_B6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_BO5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_BO6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_B_CY;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_B_XOR;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_C;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_C1;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_C2;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_C3;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_C4;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_C5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_C6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_CLK;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_CO5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_CO6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_C_CY;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_C_XOR;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_D;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_D1;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_D2;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_D3;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_D4;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_D5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_D6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_DO5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_DO6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_D_CY;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_D_XOR;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_A;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_A1;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_A2;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_A3;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_A4;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_A5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_A5Q;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_A6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_AMUX;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_AO5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_AO6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_AQ;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_AX;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_A_CY;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_A_XOR;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_B;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_B1;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_B2;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_B3;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_B4;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_B5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_B6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_BMUX;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_BO5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_BO6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_B_CY;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_B_XOR;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_C;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_C1;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_C2;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_C3;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_C4;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_C5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_C6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_CLK;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_CO5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_CO6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_CQ;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_C_CY;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_C_XOR;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_D;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_D1;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_D2;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_D3;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_D4;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_D5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_D6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_DO5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_DO6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_D_CY;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_D_XOR;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_A;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_A1;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_A2;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_A3;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_A4;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_A5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_A6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_AMUX;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_AO5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_AO6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_AQ;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_A_CY;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_A_XOR;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_B;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_B1;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_B2;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_B3;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_B4;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_B5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_B6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_BO5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_BO6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_BQ;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_B_CY;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_B_XOR;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_C;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_C1;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_C2;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_C3;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_C4;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_C5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_C6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_CLK;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_CO5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_CO6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_CQ;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_C_CY;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_C_XOR;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_D;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_D1;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_D2;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_D3;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_D4;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_D5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_D6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_DO5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_DO6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_D_CY;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_D_XOR;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_A;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_A1;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_A2;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_A3;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_A4;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_A5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_A6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_AO5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_AO6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_AQ;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_A_CY;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_A_XOR;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_B;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_B1;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_B2;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_B3;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_B4;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_B5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_B6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_BO5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_BO6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_BQ;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_B_CY;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_B_XOR;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_C;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_C1;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_C2;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_C3;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_C4;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_C5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_C6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_CLK;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_CO5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_CO6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_CQ;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_C_CY;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_C_XOR;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_D;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_D1;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_D2;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_D3;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_D4;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_D5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_D6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_DO5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_DO6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_D_CY;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_D_XOR;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_A;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_A1;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_A2;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_A3;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_A4;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_A5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_A6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_AO5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_AO6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_AQ;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_A_CY;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_A_XOR;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_B;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_B1;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_B2;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_B3;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_B4;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_B5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_B6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_BO5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_BO6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_BQ;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_B_CY;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_B_XOR;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_C;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_C1;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_C2;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_C3;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_C4;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_C5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_C6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_CLK;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_CO5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_CO6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_CQ;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_C_CY;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_C_XOR;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_D;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_D1;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_D2;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_D3;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_D4;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_D5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_D6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_DMUX;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_DO5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_DO6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_D_CY;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_D_XOR;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_A;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_A1;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_A2;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_A3;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_A4;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_A5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_A6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_AO5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_AO6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_AQ;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_A_CY;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_A_XOR;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_B;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_B1;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_B2;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_B3;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_B4;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_B5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_B6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_BO5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_BO6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_BQ;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_B_CY;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_B_XOR;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_C;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_C1;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_C2;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_C3;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_C4;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_C5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_C6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_CLK;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_CO5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_CO6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_CQ;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_C_CY;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_C_XOR;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_D;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_D1;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_D2;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_D3;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_D4;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_D5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_D6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_DO5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_DO6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_D_CY;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_D_XOR;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_A;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_A1;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_A2;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_A3;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_A4;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_A5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_A6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_AO5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_AO6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_AQ;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_A_CY;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_A_XOR;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_B;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_B1;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_B2;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_B3;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_B4;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_B5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_B6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_BO5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_BO6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_BQ;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_B_CY;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_B_XOR;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_C;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_C1;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_C2;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_C3;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_C4;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_C5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_C5Q;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_C6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_CLK;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_CMUX;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_CO5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_CO6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_CQ;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_C_CY;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_C_XOR;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_D;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_D1;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_D2;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_D3;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_D4;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_D5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_D6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_DO5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_DO6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_D_CY;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_D_XOR;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_A;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_A1;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_A2;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_A3;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_A4;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_A5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_A6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_AO5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_AO6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_AQ;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_A_CY;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_A_XOR;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_B;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_B1;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_B2;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_B3;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_B4;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_B5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_B6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_BO5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_BO6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_BQ;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_B_CY;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_B_XOR;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_C;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_C1;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_C2;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_C3;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_C4;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_C5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_C6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_CLK;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_CO5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_CO6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_CQ;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_C_CY;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_C_XOR;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_D;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_D1;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_D2;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_D3;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_D4;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_D5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_D6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_DMUX;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_DO5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_DO6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_D_CY;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_D_XOR;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_A;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_A1;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_A2;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_A3;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_A4;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_A5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_A6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_AO5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_AO6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_AQ;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_A_CY;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_A_XOR;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_B;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_B1;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_B2;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_B3;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_B4;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_B5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_B6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_BMUX;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_BO5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_BO6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_B_CY;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_B_XOR;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_C;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_C1;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_C2;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_C3;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_C4;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_C5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_C6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_CLK;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_CO5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_CO6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_C_CY;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_C_XOR;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_D;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_D1;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_D2;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_D3;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_D4;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_D5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_D6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_DO5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_DO6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_D_CY;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_D_XOR;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A1;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A2;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A3;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A4;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_AO5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_AO6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_AQ;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A_CY;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A_XOR;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B1;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B2;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B3;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B4;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_BO5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_BO6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_BQ;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B_CY;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B_XOR;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C1;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C2;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C3;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C4;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_CLK;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_CMUX;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_CO5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_CO6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C_CY;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C_XOR;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D1;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D2;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D3;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D4;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_DMUX;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_DO5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_DO6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D_CY;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D_XOR;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A1;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A2;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A3;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A4;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_AO5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_AO6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_AQ;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A_CY;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A_XOR;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B1;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B2;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B3;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B4;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_BO5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_BO6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_BQ;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B_CY;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B_XOR;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C1;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C2;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C3;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C4;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_CLK;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_CO5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_CO6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_CQ;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C_CY;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C_XOR;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D1;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D2;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D3;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D4;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_DO5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_DO6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_DQ;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D_CY;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D_XOR;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A1;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A2;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A3;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A4;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_AO5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_AO6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_AQ;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A_CY;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A_XOR;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B1;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B2;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B3;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B4;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_BO5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_BO6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_BQ;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B_CY;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B_XOR;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C1;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C2;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C3;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C4;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_CLK;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_CO5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_CO6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_CQ;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C_CY;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C_XOR;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D1;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D2;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D3;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D4;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_DMUX;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_DO5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_DO6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D_CY;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D_XOR;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A1;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A2;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A3;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A4;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_AO5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_AO6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_AQ;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A_CY;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A_XOR;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B1;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B2;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B3;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B4;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_BO5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_BO6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_BQ;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B_CY;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B_XOR;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C1;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C2;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C3;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C4;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_CLK;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_CO5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_CO6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C_CY;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C_XOR;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D1;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D2;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D3;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D4;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_DO5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_DO6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D_CY;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D_XOR;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A1;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A2;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A3;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A4;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_AO5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_AO6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_AQ;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A_CY;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A_XOR;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B1;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B2;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B3;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B4;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_BO5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_BO6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_BQ;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B_CY;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B_XOR;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C1;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C2;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C3;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C4;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_CLK;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_CO5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_CO6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_CQ;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C_CY;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C_XOR;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D1;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D2;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D3;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D4;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_DO5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_DO6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_DQ;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D_CY;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D_XOR;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A1;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A2;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A3;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A4;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_AO5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_AO6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_AQ;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A_CY;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A_XOR;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B1;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B2;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B3;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B4;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_BO5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_BO6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_BQ;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B_CY;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B_XOR;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C1;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C2;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C3;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C4;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_CLK;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_CO5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_CO6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_CQ;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C_CY;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C_XOR;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D1;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D2;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D3;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D4;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_DMUX;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_DO5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_DO6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D_CY;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D_XOR;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A1;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A2;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A3;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A4;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_AO5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_AO6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_AQ;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A_CY;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A_XOR;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B1;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B2;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B3;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B4;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_BO5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_BO6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_BQ;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B_CY;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B_XOR;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C1;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C2;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C3;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C4;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C5Q;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_CLK;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_CMUX;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_CO5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_CO6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_CQ;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C_CY;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C_XOR;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D1;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D2;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D3;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D4;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_DO5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_DO6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_DQ;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D_CY;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D_XOR;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A1;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A2;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A3;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A4;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_AO5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_AO6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_AQ;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A_CY;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A_XOR;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B1;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B2;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B3;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B4;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_BO5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_BO6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_BQ;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B_CY;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B_XOR;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C1;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C2;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C3;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C4;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_CLK;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_CO5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_CO6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C_CY;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C_XOR;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D1;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D2;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D3;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D4;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_DO5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_DO6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D_CY;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D_XOR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A1;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A2;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A3;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A4;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_AO5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_AO6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_AQ;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A_CY;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A_XOR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B1;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B2;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B3;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B4;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_BO5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_BO6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_BQ;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B_CY;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B_XOR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C1;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C2;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C3;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C4;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C5Q;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_CLK;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_CMUX;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_CO5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_CO6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_CQ;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C_CY;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C_XOR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D1;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D2;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D3;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D4;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_DO5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_DO6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_DQ;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D_CY;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D_XOR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A1;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A2;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A3;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A4;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A5Q;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_AMUX;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_AO5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_AO6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_AQ;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_AX;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A_CY;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A_XOR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B1;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B2;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B3;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B4;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_BMUX;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_BO5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_BO6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B_CY;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B_XOR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C1;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C2;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C3;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C4;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_CLK;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_CO5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_CO6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C_CY;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C_XOR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D1;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D2;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D3;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D4;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_DO5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_DO6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D_CY;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D_XOR;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A1;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A2;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A3;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A4;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A5Q;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_AMUX;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_AO5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_AO6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_AQ;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A_CY;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A_XOR;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B1;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B2;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B3;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B4;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_BO5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_BO6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_BQ;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B_CY;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B_XOR;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C1;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C2;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C3;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C4;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_CLK;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_CO5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_CO6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_CQ;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C_CY;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C_XOR;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D1;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D2;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D3;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D4;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_DO5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_DO6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D_CY;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D_XOR;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A1;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A2;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A3;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A4;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_AMUX;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_AO5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_AO6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A_CY;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A_XOR;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B1;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B2;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B3;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B4;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_BO5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_BO6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_BQ;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B_CY;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B_XOR;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C1;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C2;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C3;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C4;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_CLK;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_CO5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_CO6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C_CY;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C_XOR;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D1;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D2;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D3;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D4;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_DO5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_DO6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D_CY;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D_XOR;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A1;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A2;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A3;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A4;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_AO5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_AO6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_AQ;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A_CY;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A_XOR;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B1;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B2;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B3;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B4;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B5Q;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_BMUX;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_BO5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_BO6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_BQ;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B_CY;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B_XOR;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C1;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C2;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C3;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C4;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_CLK;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_CO5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_CO6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_CQ;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C_CY;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C_XOR;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D1;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D2;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D3;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D4;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D5Q;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_DMUX;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_DO5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_DO6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_DQ;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D_CY;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D_XOR;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A1;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A2;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A3;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A4;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A5Q;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_AMUX;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_AO5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_AO6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_AQ;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_AX;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A_CY;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A_XOR;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B1;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B2;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B3;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B4;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B5Q;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_BMUX;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_BO5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_BO6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_BQ;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B_CY;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B_XOR;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C1;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C2;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C3;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C4;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_CLK;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_CMUX;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_CO5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_CO6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C_CY;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C_XOR;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D1;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D2;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D3;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D4;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_DO5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_DO6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D_CY;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D_XOR;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_A;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_A1;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_A2;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_A3;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_A4;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_A5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_A6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_AO5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_AO6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_AQ;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_A_CY;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_A_XOR;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_B;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_B1;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_B2;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_B3;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_B4;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_B5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_B6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_BO5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_BO6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_BQ;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_B_CY;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_B_XOR;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_C;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_C1;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_C2;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_C3;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_C4;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_C5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_C6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_CLK;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_CO5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_CO6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_CQ;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_C_CY;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_C_XOR;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_D;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_D1;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_D2;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_D3;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_D4;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_D5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_D6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_DO5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_DO6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_D_CY;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_D_XOR;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_A;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_A1;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_A2;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_A3;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_A4;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_A5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_A6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_AO5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_AO6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_AQ;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_A_CY;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_A_XOR;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_B;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_B1;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_B2;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_B3;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_B4;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_B5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_B6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_BMUX;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_BO5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_BO6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_B_CY;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_B_XOR;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_C;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_C1;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_C2;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_C3;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_C4;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_C5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_C6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_CLK;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_CO5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_CO6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_C_CY;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_C_XOR;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_D;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_D1;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_D2;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_D3;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_D4;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_D5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_D6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_DO5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_DO6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_D_CY;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_D_XOR;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_A;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_A1;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_A2;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_A3;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_A4;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_A5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_A6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_AO5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_AO6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_AQ;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_A_CY;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_A_XOR;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_B;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_B1;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_B2;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_B3;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_B4;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_B5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_B6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_BO5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_BO6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_BQ;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_B_CY;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_B_XOR;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_C;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_C1;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_C2;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_C3;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_C4;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_C5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_C6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_CLK;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_CO5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_CO6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_C_CY;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_C_XOR;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_D;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_D1;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_D2;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_D3;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_D4;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_D5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_D6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_DO5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_DO6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_D_CY;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_D_XOR;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_A;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_A1;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_A2;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_A3;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_A4;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_A5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_A5Q;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_A6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_AMUX;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_AO5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_AO6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_AQ;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_AX;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_A_CY;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_A_XOR;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_B;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_B1;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_B2;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_B3;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_B4;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_B5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_B6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_BO5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_BO6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_BQ;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_B_CY;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_B_XOR;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_C;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_C1;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_C2;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_C3;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_C4;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_C5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_C6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_CLK;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_CMUX;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_CO5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_CO6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_C_CY;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_C_XOR;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_D;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_D1;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_D2;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_D3;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_D4;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_D5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_D6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_DO5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_DO6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_DQ;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_D_CY;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_D_XOR;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_A;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_A1;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_A2;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_A3;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_A4;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_A5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_A6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_AO5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_AO6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_AQ;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_A_CY;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_A_XOR;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_B;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_B1;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_B2;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_B3;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_B4;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_B5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_B6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_BO5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_BO6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_BQ;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_B_CY;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_B_XOR;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_C;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_C1;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_C2;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_C3;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_C4;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_C5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_C6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_CLK;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_CO5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_CO6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_CQ;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_C_CY;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_C_XOR;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_D;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_D1;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_D2;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_D3;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_D4;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_D5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_D6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_DO5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_DO6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_D_CY;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_D_XOR;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_A;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_A1;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_A2;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_A3;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_A4;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_A5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_A6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_AO5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_AO6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_AQ;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_A_CY;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_A_XOR;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_B;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_B1;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_B2;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_B3;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_B4;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_B5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_B6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_BMUX;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_BO5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_BO6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_B_CY;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_B_XOR;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_C;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_C1;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_C2;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_C3;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_C4;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_C5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_C6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_CLK;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_CMUX;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_CO5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_CO6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_C_CY;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_C_XOR;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_D;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_D1;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_D2;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_D3;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_D4;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_D5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_D6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_DO5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_DO6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_D_CY;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_D_XOR;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_A;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_A1;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_A2;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_A3;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_A4;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_A5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_A6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_AO5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_AO6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_A_CY;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_A_XOR;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_B;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_B1;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_B2;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_B3;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_B4;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_B5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_B6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_BO5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_BO6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_B_CY;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_B_XOR;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_C;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_C1;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_C2;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_C3;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_C4;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_C5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_C6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_CO5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_CO6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_C_CY;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_C_XOR;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_D;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_D1;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_D2;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_D3;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_D4;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_D5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_D6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_DO5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_DO6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_D_CY;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_D_XOR;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_A;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_A1;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_A2;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_A3;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_A4;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_A5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_A6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_AMUX;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_AO5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_AO6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_A_CY;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_A_XOR;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_B;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_B1;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_B2;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_B3;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_B4;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_B5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_B6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_BO5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_BO6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_B_CY;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_B_XOR;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_C;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_C1;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_C2;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_C3;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_C4;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_C5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_C6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_CO5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_CO6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_C_CY;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_C_XOR;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_D;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_D1;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_D2;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_D3;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_D4;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_D5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_D6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_DO5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_DO6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_D_CY;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_D_XOR;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE1;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I1;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE1;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S1;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_CE;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_I;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  wire [0:0] LIOB33_SING_X0Y100_IOB_X0Y100_O;
  wire [0:0] LIOB33_SING_X0Y149_IOB_X0Y149_O;
  wire [0:0] LIOB33_SING_X0Y150_IOB_X0Y150_O;
  wire [0:0] LIOB33_SING_X0Y199_IOB_X0Y199_O;
  wire [0:0] LIOB33_SING_X0Y50_IOB_X0Y50_I;
  wire [0:0] LIOB33_X0Y101_IOB_X0Y101_O;
  wire [0:0] LIOB33_X0Y101_IOB_X0Y102_O;
  wire [0:0] LIOB33_X0Y103_IOB_X0Y103_O;
  wire [0:0] LIOB33_X0Y103_IOB_X0Y104_O;
  wire [0:0] LIOB33_X0Y105_IOB_X0Y105_O;
  wire [0:0] LIOB33_X0Y105_IOB_X0Y106_O;
  wire [0:0] LIOB33_X0Y107_IOB_X0Y107_O;
  wire [0:0] LIOB33_X0Y107_IOB_X0Y108_O;
  wire [0:0] LIOB33_X0Y109_IOB_X0Y109_O;
  wire [0:0] LIOB33_X0Y109_IOB_X0Y110_O;
  wire [0:0] LIOB33_X0Y111_IOB_X0Y111_O;
  wire [0:0] LIOB33_X0Y111_IOB_X0Y112_O;
  wire [0:0] LIOB33_X0Y113_IOB_X0Y113_O;
  wire [0:0] LIOB33_X0Y113_IOB_X0Y114_O;
  wire [0:0] LIOB33_X0Y115_IOB_X0Y115_O;
  wire [0:0] LIOB33_X0Y115_IOB_X0Y116_O;
  wire [0:0] LIOB33_X0Y117_IOB_X0Y117_O;
  wire [0:0] LIOB33_X0Y117_IOB_X0Y118_O;
  wire [0:0] LIOB33_X0Y119_IOB_X0Y119_O;
  wire [0:0] LIOB33_X0Y119_IOB_X0Y120_O;
  wire [0:0] LIOB33_X0Y121_IOB_X0Y121_O;
  wire [0:0] LIOB33_X0Y121_IOB_X0Y122_O;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y123_O;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y124_O;
  wire [0:0] LIOB33_X0Y125_IOB_X0Y125_O;
  wire [0:0] LIOB33_X0Y125_IOB_X0Y126_O;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y127_O;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y128_O;
  wire [0:0] LIOB33_X0Y129_IOB_X0Y129_O;
  wire [0:0] LIOB33_X0Y129_IOB_X0Y130_O;
  wire [0:0] LIOB33_X0Y131_IOB_X0Y131_O;
  wire [0:0] LIOB33_X0Y131_IOB_X0Y132_O;
  wire [0:0] LIOB33_X0Y133_IOB_X0Y133_O;
  wire [0:0] LIOB33_X0Y133_IOB_X0Y134_O;
  wire [0:0] LIOB33_X0Y135_IOB_X0Y135_O;
  wire [0:0] LIOB33_X0Y135_IOB_X0Y136_O;
  wire [0:0] LIOB33_X0Y137_IOB_X0Y137_O;
  wire [0:0] LIOB33_X0Y137_IOB_X0Y138_O;
  wire [0:0] LIOB33_X0Y139_IOB_X0Y139_O;
  wire [0:0] LIOB33_X0Y139_IOB_X0Y140_O;
  wire [0:0] LIOB33_X0Y141_IOB_X0Y141_O;
  wire [0:0] LIOB33_X0Y141_IOB_X0Y142_O;
  wire [0:0] LIOB33_X0Y143_IOB_X0Y143_O;
  wire [0:0] LIOB33_X0Y145_IOB_X0Y145_O;
  wire [0:0] LIOB33_X0Y145_IOB_X0Y146_O;
  wire [0:0] LIOB33_X0Y147_IOB_X0Y147_O;
  wire [0:0] LIOB33_X0Y147_IOB_X0Y148_O;
  wire [0:0] LIOB33_X0Y151_IOB_X0Y151_O;
  wire [0:0] LIOB33_X0Y151_IOB_X0Y152_O;
  wire [0:0] LIOB33_X0Y153_IOB_X0Y153_O;
  wire [0:0] LIOB33_X0Y153_IOB_X0Y154_O;
  wire [0:0] LIOB33_X0Y155_IOB_X0Y155_O;
  wire [0:0] LIOB33_X0Y155_IOB_X0Y156_O;
  wire [0:0] LIOB33_X0Y157_IOB_X0Y157_O;
  wire [0:0] LIOB33_X0Y157_IOB_X0Y158_O;
  wire [0:0] LIOB33_X0Y159_IOB_X0Y159_O;
  wire [0:0] LIOB33_X0Y159_IOB_X0Y160_O;
  wire [0:0] LIOB33_X0Y161_IOB_X0Y161_O;
  wire [0:0] LIOB33_X0Y161_IOB_X0Y162_O;
  wire [0:0] LIOB33_X0Y163_IOB_X0Y163_O;
  wire [0:0] LIOB33_X0Y163_IOB_X0Y164_O;
  wire [0:0] LIOB33_X0Y165_IOB_X0Y165_O;
  wire [0:0] LIOB33_X0Y165_IOB_X0Y166_O;
  wire [0:0] LIOB33_X0Y167_IOB_X0Y167_O;
  wire [0:0] LIOB33_X0Y167_IOB_X0Y168_O;
  wire [0:0] LIOB33_X0Y169_IOB_X0Y169_O;
  wire [0:0] LIOB33_X0Y169_IOB_X0Y170_O;
  wire [0:0] LIOB33_X0Y171_IOB_X0Y171_O;
  wire [0:0] LIOB33_X0Y171_IOB_X0Y172_O;
  wire [0:0] LIOB33_X0Y173_IOB_X0Y173_O;
  wire [0:0] LIOB33_X0Y173_IOB_X0Y174_O;
  wire [0:0] LIOB33_X0Y175_IOB_X0Y175_O;
  wire [0:0] LIOB33_X0Y175_IOB_X0Y176_O;
  wire [0:0] LIOB33_X0Y177_IOB_X0Y177_O;
  wire [0:0] LIOB33_X0Y177_IOB_X0Y178_O;
  wire [0:0] LIOB33_X0Y179_IOB_X0Y179_O;
  wire [0:0] LIOB33_X0Y179_IOB_X0Y180_O;
  wire [0:0] LIOB33_X0Y181_IOB_X0Y181_O;
  wire [0:0] LIOB33_X0Y181_IOB_X0Y182_O;
  wire [0:0] LIOB33_X0Y183_IOB_X0Y183_O;
  wire [0:0] LIOB33_X0Y183_IOB_X0Y184_O;
  wire [0:0] LIOB33_X0Y185_IOB_X0Y185_O;
  wire [0:0] LIOB33_X0Y185_IOB_X0Y186_O;
  wire [0:0] LIOB33_X0Y187_IOB_X0Y187_O;
  wire [0:0] LIOB33_X0Y187_IOB_X0Y188_O;
  wire [0:0] LIOB33_X0Y189_IOB_X0Y189_O;
  wire [0:0] LIOB33_X0Y189_IOB_X0Y190_O;
  wire [0:0] LIOB33_X0Y191_IOB_X0Y191_O;
  wire [0:0] LIOB33_X0Y191_IOB_X0Y192_O;
  wire [0:0] LIOB33_X0Y193_IOB_X0Y193_O;
  wire [0:0] LIOB33_X0Y193_IOB_X0Y194_O;
  wire [0:0] LIOB33_X0Y195_IOB_X0Y195_O;
  wire [0:0] LIOB33_X0Y195_IOB_X0Y196_O;
  wire [0:0] LIOB33_X0Y197_IOB_X0Y197_O;
  wire [0:0] LIOB33_X0Y197_IOB_X0Y198_O;
  wire [0:0] LIOB33_X0Y51_IOB_X0Y51_I;
  wire [0:0] LIOB33_X0Y51_IOB_X0Y52_I;
  wire [0:0] LIOB33_X0Y53_IOB_X0Y53_I;
  wire [0:0] LIOB33_X0Y53_IOB_X0Y54_I;
  wire [0:0] LIOB33_X0Y55_IOB_X0Y55_I;
  wire [0:0] LIOB33_X0Y55_IOB_X0Y56_I;
  wire [0:0] LIOB33_X0Y57_IOB_X0Y57_I;
  wire [0:0] LIOB33_X0Y57_IOB_X0Y58_I;
  wire [0:0] LIOB33_X0Y59_IOB_X0Y59_I;
  wire [0:0] LIOB33_X0Y59_IOB_X0Y60_I;
  wire [0:0] LIOB33_X0Y61_IOB_X0Y61_I;
  wire [0:0] LIOB33_X0Y61_IOB_X0Y62_I;
  wire [0:0] LIOB33_X0Y63_IOB_X0Y63_I;
  wire [0:0] LIOB33_X0Y63_IOB_X0Y64_I;
  wire [0:0] LIOB33_X0Y65_IOB_X0Y65_I;
  wire [0:0] LIOB33_X0Y65_IOB_X0Y66_I;
  wire [0:0] LIOB33_X0Y67_IOB_X0Y67_I;
  wire [0:0] LIOB33_X0Y67_IOB_X0Y68_I;
  wire [0:0] LIOB33_X0Y69_IOB_X0Y69_I;
  wire [0:0] LIOB33_X0Y69_IOB_X0Y70_I;
  wire [0:0] LIOB33_X0Y71_IOB_X0Y71_I;
  wire [0:0] LIOB33_X0Y71_IOB_X0Y72_I;
  wire [0:0] LIOB33_X0Y73_IOB_X0Y73_I;
  wire [0:0] LIOB33_X0Y73_IOB_X0Y74_I;
  wire [0:0] LIOB33_X0Y75_IOB_X0Y75_I;
  wire [0:0] LIOB33_X0Y75_IOB_X0Y76_I;
  wire [0:0] LIOB33_X0Y77_IOB_X0Y77_I;
  wire [0:0] LIOB33_X0Y77_IOB_X0Y78_I;
  wire [0:0] LIOB33_X0Y79_IOB_X0Y79_I;
  wire [0:0] LIOB33_X0Y79_IOB_X0Y80_O;
  wire [0:0] LIOI3_SING_X0Y100_OLOGIC_X0Y100_D1;
  wire [0:0] LIOI3_SING_X0Y100_OLOGIC_X0Y100_OQ;
  wire [0:0] LIOI3_SING_X0Y100_OLOGIC_X0Y100_T1;
  wire [0:0] LIOI3_SING_X0Y100_OLOGIC_X0Y100_TQ;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_D1;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_OQ;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_T1;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_TQ;
  wire [0:0] LIOI3_SING_X0Y150_OLOGIC_X0Y150_D1;
  wire [0:0] LIOI3_SING_X0Y150_OLOGIC_X0Y150_OQ;
  wire [0:0] LIOI3_SING_X0Y150_OLOGIC_X0Y150_T1;
  wire [0:0] LIOI3_SING_X0Y150_OLOGIC_X0Y150_TQ;
  wire [0:0] LIOI3_SING_X0Y199_OLOGIC_X0Y199_D1;
  wire [0:0] LIOI3_SING_X0Y199_OLOGIC_X0Y199_OQ;
  wire [0:0] LIOI3_SING_X0Y199_OLOGIC_X0Y199_T1;
  wire [0:0] LIOI3_SING_X0Y199_OLOGIC_X0Y199_TQ;
  wire [0:0] LIOI3_SING_X0Y50_ILOGIC_X0Y50_D;
  wire [0:0] LIOI3_SING_X0Y50_ILOGIC_X0Y50_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y57_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y57_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y58_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y58_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y69_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y69_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y70_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y70_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y63_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y63_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y64_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y64_O;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y101_D1;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y101_OQ;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y101_T1;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y101_TQ;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y102_D1;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y102_OQ;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y102_T1;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y102_TQ;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y103_D1;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y103_OQ;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y103_T1;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y103_TQ;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y104_D1;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y104_OQ;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y104_T1;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y104_TQ;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y105_D1;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y105_OQ;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y105_T1;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y105_TQ;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y106_D1;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y106_OQ;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y106_T1;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y106_TQ;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y109_D1;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y109_OQ;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y109_T1;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y109_TQ;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y110_D1;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y110_OQ;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y110_T1;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y110_TQ;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_D1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_OQ;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_T1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_TQ;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y112_D1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y112_OQ;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y112_T1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y112_TQ;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y115_D1;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y115_OQ;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y115_T1;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y115_TQ;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y116_D1;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y116_OQ;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y116_T1;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y116_TQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y117_D1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y117_OQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y117_T1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y117_TQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_D1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_OQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_T1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_TQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_D1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_OQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_T1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_TQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_D1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_OQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_T1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_TQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_D1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_OQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_T1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_TQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_D1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_OQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_T1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_TQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_D1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_OQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_T1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_TQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_D1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_OQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_T1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_TQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_D1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_OQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_T1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_TQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_D1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_OQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_T1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_TQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_D1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_OQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_T1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_TQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_D1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_OQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_T1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_TQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_D1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_OQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_T1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_TQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_D1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_OQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_T1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_TQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_D1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_OQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_T1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_TQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_D1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_OQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_T1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_TQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_D1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_OQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_T1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_TQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_D1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_OQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_T1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_TQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_D1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_OQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_T1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_TQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_D1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_OQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_T1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_TQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_D1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_OQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_T1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_TQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_D1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_OQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_T1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_TQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_D1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_OQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_T1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_TQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_D1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_OQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_T1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_TQ;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y151_D1;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y151_OQ;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y151_T1;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y151_TQ;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y152_D1;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y152_OQ;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y152_T1;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y152_TQ;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y153_D1;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y153_OQ;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y153_T1;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y153_TQ;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y154_D1;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y154_OQ;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y154_T1;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y154_TQ;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y155_D1;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y155_OQ;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y155_T1;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y155_TQ;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y156_D1;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y156_OQ;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y156_T1;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y156_TQ;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y159_D1;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y159_OQ;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y159_T1;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y159_TQ;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y160_D1;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y160_OQ;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y160_T1;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y160_TQ;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y161_D1;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y161_OQ;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y161_T1;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y161_TQ;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y162_D1;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y162_OQ;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y162_T1;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y162_TQ;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y165_D1;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y165_OQ;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y165_T1;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y165_TQ;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y166_D1;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y166_OQ;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y166_T1;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y166_TQ;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y167_D1;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y167_OQ;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y167_T1;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y167_TQ;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y168_D1;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y168_OQ;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y168_T1;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y168_TQ;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y171_D1;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y171_OQ;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y171_T1;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y171_TQ;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y172_D1;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y172_OQ;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y172_T1;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y172_TQ;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y173_D1;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y173_OQ;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y173_T1;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y173_TQ;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y174_D1;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y174_OQ;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y174_T1;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y174_TQ;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y175_D1;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y175_OQ;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y175_T1;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y175_TQ;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y176_D1;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y176_OQ;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y176_T1;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y176_TQ;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y177_D1;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y177_OQ;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y177_T1;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y177_TQ;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y178_D1;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y178_OQ;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y178_T1;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y178_TQ;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y179_D1;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y179_OQ;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y179_T1;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y179_TQ;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y180_D1;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y180_OQ;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y180_T1;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y180_TQ;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y183_D1;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y183_OQ;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y183_T1;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y183_TQ;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y184_D1;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y184_OQ;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y184_T1;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y184_TQ;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y185_D1;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y185_OQ;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y185_T1;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y185_TQ;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y186_D1;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y186_OQ;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y186_T1;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y186_TQ;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y189_D1;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y189_OQ;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y189_T1;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y189_TQ;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y190_D1;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y190_OQ;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y190_T1;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y190_TQ;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y191_D1;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y191_OQ;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y191_T1;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y191_TQ;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y192_D1;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y192_OQ;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y192_T1;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y192_TQ;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y195_D1;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y195_OQ;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y195_T1;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y195_TQ;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y196_D1;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y196_OQ;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y196_T1;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y196_TQ;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y197_D1;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y197_OQ;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y197_T1;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y197_TQ;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y198_D1;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y198_OQ;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y198_T1;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y198_TQ;
  wire [0:0] LIOI3_X0Y51_ILOGIC_X0Y51_D;
  wire [0:0] LIOI3_X0Y51_ILOGIC_X0Y51_O;
  wire [0:0] LIOI3_X0Y51_ILOGIC_X0Y52_D;
  wire [0:0] LIOI3_X0Y51_ILOGIC_X0Y52_O;
  wire [0:0] LIOI3_X0Y53_ILOGIC_X0Y53_D;
  wire [0:0] LIOI3_X0Y53_ILOGIC_X0Y53_O;
  wire [0:0] LIOI3_X0Y53_ILOGIC_X0Y54_D;
  wire [0:0] LIOI3_X0Y53_ILOGIC_X0Y54_O;
  wire [0:0] LIOI3_X0Y55_ILOGIC_X0Y55_D;
  wire [0:0] LIOI3_X0Y55_ILOGIC_X0Y55_O;
  wire [0:0] LIOI3_X0Y55_ILOGIC_X0Y56_D;
  wire [0:0] LIOI3_X0Y55_ILOGIC_X0Y56_O;
  wire [0:0] LIOI3_X0Y59_ILOGIC_X0Y59_D;
  wire [0:0] LIOI3_X0Y59_ILOGIC_X0Y59_O;
  wire [0:0] LIOI3_X0Y59_ILOGIC_X0Y60_D;
  wire [0:0] LIOI3_X0Y59_ILOGIC_X0Y60_O;
  wire [0:0] LIOI3_X0Y61_ILOGIC_X0Y61_D;
  wire [0:0] LIOI3_X0Y61_ILOGIC_X0Y61_O;
  wire [0:0] LIOI3_X0Y61_ILOGIC_X0Y62_D;
  wire [0:0] LIOI3_X0Y61_ILOGIC_X0Y62_O;
  wire [0:0] LIOI3_X0Y65_ILOGIC_X0Y65_D;
  wire [0:0] LIOI3_X0Y65_ILOGIC_X0Y65_O;
  wire [0:0] LIOI3_X0Y65_ILOGIC_X0Y66_D;
  wire [0:0] LIOI3_X0Y65_ILOGIC_X0Y66_O;
  wire [0:0] LIOI3_X0Y67_ILOGIC_X0Y67_D;
  wire [0:0] LIOI3_X0Y67_ILOGIC_X0Y67_O;
  wire [0:0] LIOI3_X0Y67_ILOGIC_X0Y68_D;
  wire [0:0] LIOI3_X0Y67_ILOGIC_X0Y68_O;
  wire [0:0] LIOI3_X0Y71_ILOGIC_X0Y71_D;
  wire [0:0] LIOI3_X0Y71_ILOGIC_X0Y71_O;
  wire [0:0] LIOI3_X0Y71_ILOGIC_X0Y72_D;
  wire [0:0] LIOI3_X0Y71_ILOGIC_X0Y72_O;
  wire [0:0] LIOI3_X0Y73_ILOGIC_X0Y73_D;
  wire [0:0] LIOI3_X0Y73_ILOGIC_X0Y73_O;
  wire [0:0] LIOI3_X0Y73_ILOGIC_X0Y74_D;
  wire [0:0] LIOI3_X0Y73_ILOGIC_X0Y74_O;
  wire [0:0] LIOI3_X0Y75_ILOGIC_X0Y75_D;
  wire [0:0] LIOI3_X0Y75_ILOGIC_X0Y75_O;
  wire [0:0] LIOI3_X0Y75_ILOGIC_X0Y76_D;
  wire [0:0] LIOI3_X0Y75_ILOGIC_X0Y76_O;
  wire [0:0] LIOI3_X0Y77_ILOGIC_X0Y77_D;
  wire [0:0] LIOI3_X0Y77_ILOGIC_X0Y77_O;
  wire [0:0] LIOI3_X0Y77_ILOGIC_X0Y78_D;
  wire [0:0] LIOI3_X0Y77_ILOGIC_X0Y78_O;
  wire [0:0] LIOI3_X0Y79_ILOGIC_X0Y79_D;
  wire [0:0] LIOI3_X0Y79_ILOGIC_X0Y79_O;
  wire [0:0] LIOI3_X0Y79_OLOGIC_X0Y80_D1;
  wire [0:0] LIOI3_X0Y79_OLOGIC_X0Y80_OQ;
  wire [0:0] LIOI3_X0Y79_OLOGIC_X0Y80_T1;
  wire [0:0] LIOI3_X0Y79_OLOGIC_X0Y80_TQ;
  wire [0:0] RIOB33_SING_X105Y100_IOB_X1Y100_I;
  wire [0:0] RIOB33_SING_X105Y149_IOB_X1Y149_I;
  wire [0:0] RIOB33_SING_X105Y150_IOB_X1Y150_O;
  wire [0:0] RIOB33_SING_X105Y199_IOB_X1Y199_O;
  wire [0:0] RIOB33_X105Y101_IOB_X1Y101_I;
  wire [0:0] RIOB33_X105Y101_IOB_X1Y102_I;
  wire [0:0] RIOB33_X105Y103_IOB_X1Y103_I;
  wire [0:0] RIOB33_X105Y103_IOB_X1Y104_I;
  wire [0:0] RIOB33_X105Y105_IOB_X1Y105_I;
  wire [0:0] RIOB33_X105Y105_IOB_X1Y106_I;
  wire [0:0] RIOB33_X105Y107_IOB_X1Y107_I;
  wire [0:0] RIOB33_X105Y107_IOB_X1Y108_I;
  wire [0:0] RIOB33_X105Y109_IOB_X1Y109_I;
  wire [0:0] RIOB33_X105Y109_IOB_X1Y110_I;
  wire [0:0] RIOB33_X105Y111_IOB_X1Y111_I;
  wire [0:0] RIOB33_X105Y111_IOB_X1Y112_I;
  wire [0:0] RIOB33_X105Y113_IOB_X1Y113_I;
  wire [0:0] RIOB33_X105Y113_IOB_X1Y114_I;
  wire [0:0] RIOB33_X105Y115_IOB_X1Y115_I;
  wire [0:0] RIOB33_X105Y115_IOB_X1Y116_I;
  wire [0:0] RIOB33_X105Y117_IOB_X1Y117_I;
  wire [0:0] RIOB33_X105Y117_IOB_X1Y118_I;
  wire [0:0] RIOB33_X105Y119_IOB_X1Y119_I;
  wire [0:0] RIOB33_X105Y119_IOB_X1Y120_I;
  wire [0:0] RIOB33_X105Y121_IOB_X1Y121_I;
  wire [0:0] RIOB33_X105Y121_IOB_X1Y122_I;
  wire [0:0] RIOB33_X105Y123_IOB_X1Y123_I;
  wire [0:0] RIOB33_X105Y123_IOB_X1Y124_I;
  wire [0:0] RIOB33_X105Y125_IOB_X1Y125_I;
  wire [0:0] RIOB33_X105Y125_IOB_X1Y126_I;
  wire [0:0] RIOB33_X105Y127_IOB_X1Y127_I;
  wire [0:0] RIOB33_X105Y127_IOB_X1Y128_I;
  wire [0:0] RIOB33_X105Y129_IOB_X1Y129_I;
  wire [0:0] RIOB33_X105Y129_IOB_X1Y130_I;
  wire [0:0] RIOB33_X105Y131_IOB_X1Y131_I;
  wire [0:0] RIOB33_X105Y131_IOB_X1Y132_I;
  wire [0:0] RIOB33_X105Y133_IOB_X1Y133_I;
  wire [0:0] RIOB33_X105Y133_IOB_X1Y134_I;
  wire [0:0] RIOB33_X105Y135_IOB_X1Y135_I;
  wire [0:0] RIOB33_X105Y135_IOB_X1Y136_I;
  wire [0:0] RIOB33_X105Y137_IOB_X1Y137_I;
  wire [0:0] RIOB33_X105Y137_IOB_X1Y138_I;
  wire [0:0] RIOB33_X105Y139_IOB_X1Y139_I;
  wire [0:0] RIOB33_X105Y139_IOB_X1Y140_I;
  wire [0:0] RIOB33_X105Y141_IOB_X1Y141_I;
  wire [0:0] RIOB33_X105Y141_IOB_X1Y142_I;
  wire [0:0] RIOB33_X105Y143_IOB_X1Y143_I;
  wire [0:0] RIOB33_X105Y143_IOB_X1Y144_I;
  wire [0:0] RIOB33_X105Y145_IOB_X1Y145_I;
  wire [0:0] RIOB33_X105Y145_IOB_X1Y146_I;
  wire [0:0] RIOB33_X105Y147_IOB_X1Y147_I;
  wire [0:0] RIOB33_X105Y147_IOB_X1Y148_I;
  wire [0:0] RIOB33_X105Y151_IOB_X1Y151_O;
  wire [0:0] RIOB33_X105Y151_IOB_X1Y152_O;
  wire [0:0] RIOB33_X105Y153_IOB_X1Y153_O;
  wire [0:0] RIOB33_X105Y153_IOB_X1Y154_O;
  wire [0:0] RIOB33_X105Y155_IOB_X1Y155_O;
  wire [0:0] RIOB33_X105Y155_IOB_X1Y156_O;
  wire [0:0] RIOB33_X105Y157_IOB_X1Y157_O;
  wire [0:0] RIOB33_X105Y157_IOB_X1Y158_O;
  wire [0:0] RIOB33_X105Y159_IOB_X1Y159_O;
  wire [0:0] RIOB33_X105Y159_IOB_X1Y160_O;
  wire [0:0] RIOB33_X105Y161_IOB_X1Y161_O;
  wire [0:0] RIOB33_X105Y161_IOB_X1Y162_O;
  wire [0:0] RIOB33_X105Y163_IOB_X1Y163_O;
  wire [0:0] RIOB33_X105Y163_IOB_X1Y164_O;
  wire [0:0] RIOB33_X105Y165_IOB_X1Y165_O;
  wire [0:0] RIOB33_X105Y165_IOB_X1Y166_O;
  wire [0:0] RIOB33_X105Y167_IOB_X1Y167_O;
  wire [0:0] RIOB33_X105Y167_IOB_X1Y168_O;
  wire [0:0] RIOB33_X105Y169_IOB_X1Y169_O;
  wire [0:0] RIOB33_X105Y169_IOB_X1Y170_O;
  wire [0:0] RIOB33_X105Y171_IOB_X1Y171_O;
  wire [0:0] RIOB33_X105Y171_IOB_X1Y172_O;
  wire [0:0] RIOB33_X105Y173_IOB_X1Y173_O;
  wire [0:0] RIOB33_X105Y173_IOB_X1Y174_O;
  wire [0:0] RIOB33_X105Y175_IOB_X1Y175_O;
  wire [0:0] RIOB33_X105Y175_IOB_X1Y176_O;
  wire [0:0] RIOB33_X105Y177_IOB_X1Y177_O;
  wire [0:0] RIOB33_X105Y177_IOB_X1Y178_O;
  wire [0:0] RIOB33_X105Y179_IOB_X1Y179_O;
  wire [0:0] RIOB33_X105Y179_IOB_X1Y180_O;
  wire [0:0] RIOB33_X105Y181_IOB_X1Y181_O;
  wire [0:0] RIOB33_X105Y181_IOB_X1Y182_O;
  wire [0:0] RIOB33_X105Y183_IOB_X1Y183_O;
  wire [0:0] RIOB33_X105Y183_IOB_X1Y184_O;
  wire [0:0] RIOB33_X105Y185_IOB_X1Y185_O;
  wire [0:0] RIOB33_X105Y185_IOB_X1Y186_O;
  wire [0:0] RIOB33_X105Y187_IOB_X1Y187_O;
  wire [0:0] RIOB33_X105Y187_IOB_X1Y188_O;
  wire [0:0] RIOB33_X105Y189_IOB_X1Y189_O;
  wire [0:0] RIOB33_X105Y189_IOB_X1Y190_O;
  wire [0:0] RIOB33_X105Y191_IOB_X1Y191_O;
  wire [0:0] RIOB33_X105Y191_IOB_X1Y192_O;
  wire [0:0] RIOB33_X105Y193_IOB_X1Y193_O;
  wire [0:0] RIOB33_X105Y193_IOB_X1Y194_O;
  wire [0:0] RIOB33_X105Y195_IOB_X1Y195_O;
  wire [0:0] RIOB33_X105Y195_IOB_X1Y196_O;
  wire [0:0] RIOB33_X105Y197_IOB_X1Y197_O;
  wire [0:0] RIOB33_X105Y197_IOB_X1Y198_O;
  wire [0:0] RIOI3_SING_X105Y100_ILOGIC_X1Y100_D;
  wire [0:0] RIOI3_SING_X105Y100_ILOGIC_X1Y100_O;
  wire [0:0] RIOI3_SING_X105Y149_ILOGIC_X1Y149_D;
  wire [0:0] RIOI3_SING_X105Y149_ILOGIC_X1Y149_O;
  wire [0:0] RIOI3_SING_X105Y150_OLOGIC_X1Y150_D1;
  wire [0:0] RIOI3_SING_X105Y150_OLOGIC_X1Y150_OQ;
  wire [0:0] RIOI3_SING_X105Y150_OLOGIC_X1Y150_T1;
  wire [0:0] RIOI3_SING_X105Y150_OLOGIC_X1Y150_TQ;
  wire [0:0] RIOI3_SING_X105Y199_OLOGIC_X1Y199_D1;
  wire [0:0] RIOI3_SING_X105Y199_OLOGIC_X1Y199_OQ;
  wire [0:0] RIOI3_SING_X105Y199_OLOGIC_X1Y199_T1;
  wire [0:0] RIOI3_SING_X105Y199_OLOGIC_X1Y199_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y131_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y131_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y132_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y132_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y143_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y143_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y144_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y144_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y114_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y114_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y137_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y137_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y138_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y138_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_TQ;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y101_D;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y101_O;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y102_D;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y102_O;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y103_D;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y103_O;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y104_D;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y104_O;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y105_D;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y105_O;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y106_D;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y106_O;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y109_D;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y109_O;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y110_D;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y110_O;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y111_D;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y111_O;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y112_D;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y112_O;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y115_D;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y115_O;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y116_D;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y116_O;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y117_D;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y117_O;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y118_D;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y118_O;
  wire [0:0] RIOI3_X105Y121_ILOGIC_X1Y121_D;
  wire [0:0] RIOI3_X105Y121_ILOGIC_X1Y121_O;
  wire [0:0] RIOI3_X105Y121_ILOGIC_X1Y122_D;
  wire [0:0] RIOI3_X105Y121_ILOGIC_X1Y122_O;
  wire [0:0] RIOI3_X105Y123_ILOGIC_X1Y123_D;
  wire [0:0] RIOI3_X105Y123_ILOGIC_X1Y123_O;
  wire [0:0] RIOI3_X105Y123_ILOGIC_X1Y124_D;
  wire [0:0] RIOI3_X105Y123_ILOGIC_X1Y124_O;
  wire [0:0] RIOI3_X105Y125_ILOGIC_X1Y125_D;
  wire [0:0] RIOI3_X105Y125_ILOGIC_X1Y125_O;
  wire [0:0] RIOI3_X105Y125_ILOGIC_X1Y126_D;
  wire [0:0] RIOI3_X105Y125_ILOGIC_X1Y126_O;
  wire [0:0] RIOI3_X105Y127_ILOGIC_X1Y127_D;
  wire [0:0] RIOI3_X105Y127_ILOGIC_X1Y127_O;
  wire [0:0] RIOI3_X105Y127_ILOGIC_X1Y128_D;
  wire [0:0] RIOI3_X105Y127_ILOGIC_X1Y128_O;
  wire [0:0] RIOI3_X105Y129_ILOGIC_X1Y129_D;
  wire [0:0] RIOI3_X105Y129_ILOGIC_X1Y129_O;
  wire [0:0] RIOI3_X105Y129_ILOGIC_X1Y130_D;
  wire [0:0] RIOI3_X105Y129_ILOGIC_X1Y130_O;
  wire [0:0] RIOI3_X105Y133_ILOGIC_X1Y133_D;
  wire [0:0] RIOI3_X105Y133_ILOGIC_X1Y133_O;
  wire [0:0] RIOI3_X105Y133_ILOGIC_X1Y134_D;
  wire [0:0] RIOI3_X105Y133_ILOGIC_X1Y134_O;
  wire [0:0] RIOI3_X105Y135_ILOGIC_X1Y135_D;
  wire [0:0] RIOI3_X105Y135_ILOGIC_X1Y135_O;
  wire [0:0] RIOI3_X105Y135_ILOGIC_X1Y136_D;
  wire [0:0] RIOI3_X105Y135_ILOGIC_X1Y136_O;
  wire [0:0] RIOI3_X105Y139_ILOGIC_X1Y139_D;
  wire [0:0] RIOI3_X105Y139_ILOGIC_X1Y139_O;
  wire [0:0] RIOI3_X105Y139_ILOGIC_X1Y140_D;
  wire [0:0] RIOI3_X105Y139_ILOGIC_X1Y140_O;
  wire [0:0] RIOI3_X105Y141_ILOGIC_X1Y141_D;
  wire [0:0] RIOI3_X105Y141_ILOGIC_X1Y141_O;
  wire [0:0] RIOI3_X105Y141_ILOGIC_X1Y142_D;
  wire [0:0] RIOI3_X105Y141_ILOGIC_X1Y142_O;
  wire [0:0] RIOI3_X105Y145_ILOGIC_X1Y145_D;
  wire [0:0] RIOI3_X105Y145_ILOGIC_X1Y145_O;
  wire [0:0] RIOI3_X105Y145_ILOGIC_X1Y146_D;
  wire [0:0] RIOI3_X105Y145_ILOGIC_X1Y146_O;
  wire [0:0] RIOI3_X105Y147_ILOGIC_X1Y147_D;
  wire [0:0] RIOI3_X105Y147_ILOGIC_X1Y147_O;
  wire [0:0] RIOI3_X105Y147_ILOGIC_X1Y148_D;
  wire [0:0] RIOI3_X105Y147_ILOGIC_X1Y148_O;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y151_D1;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y151_OQ;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y151_T1;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y151_TQ;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y152_D1;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y152_OQ;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y152_T1;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y152_TQ;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y153_D1;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y153_OQ;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y153_T1;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y153_TQ;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y154_D1;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y154_OQ;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y154_T1;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y154_TQ;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y155_D1;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y155_OQ;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y155_T1;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y155_TQ;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y156_D1;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y156_OQ;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y156_T1;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y156_TQ;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y159_D1;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y159_OQ;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y159_T1;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y159_TQ;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y160_D1;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y160_OQ;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y160_T1;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y160_TQ;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y161_D1;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y161_OQ;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y161_T1;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y161_TQ;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y162_D1;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y162_OQ;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y162_T1;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y162_TQ;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y165_D1;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y165_OQ;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y165_T1;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y165_TQ;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y166_D1;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y166_OQ;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y166_T1;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y166_TQ;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y167_D1;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y167_OQ;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y167_T1;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y167_TQ;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y168_D1;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y168_OQ;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y168_T1;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y168_TQ;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y171_D1;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y171_OQ;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y171_T1;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y171_TQ;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y172_D1;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y172_OQ;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y172_T1;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y172_TQ;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y173_D1;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y173_OQ;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y173_T1;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y173_TQ;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y174_D1;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y174_OQ;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y174_T1;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y174_TQ;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y175_D1;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y175_OQ;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y175_T1;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y175_TQ;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y176_D1;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y176_OQ;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y176_T1;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y176_TQ;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y177_D1;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y177_OQ;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y177_T1;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y177_TQ;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y178_D1;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y178_OQ;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y178_T1;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y178_TQ;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y179_D1;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y179_OQ;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y179_T1;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y179_TQ;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y180_D1;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y180_OQ;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y180_T1;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y180_TQ;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y183_D1;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y183_OQ;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y183_T1;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y183_TQ;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y184_D1;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y184_OQ;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y184_T1;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y184_TQ;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y185_D1;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y185_OQ;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y185_T1;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y185_TQ;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y186_D1;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y186_OQ;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y186_T1;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y186_TQ;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y189_D1;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y189_OQ;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y189_T1;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y189_TQ;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y190_D1;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y190_OQ;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y190_T1;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y190_TQ;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y191_D1;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y191_OQ;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y191_T1;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y191_TQ;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y192_D1;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y192_OQ;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y192_T1;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y192_TQ;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y195_D1;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y195_OQ;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y195_T1;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y195_TQ;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y196_D1;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y196_OQ;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y196_T1;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y196_TQ;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y197_D1;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y197_OQ;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y197_T1;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y197_TQ;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y198_D1;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y198_OQ;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y198_T1;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y198_TQ;


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y106_SLICE_X0Y106_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y106_SLICE_X0Y106_DO5),
.O6(CLBLL_L_X2Y106_SLICE_X0Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffeefffefffeff)
  ) CLBLL_L_X2Y106_SLICE_X0Y106_CLUT (
.I0(RIOB33_X105Y129_IOB_X1Y129_I),
.I1(RIOB33_X105Y127_IOB_X1Y128_I),
.I2(CLBLM_R_X3Y109_SLICE_X2Y109_CO6),
.I3(RIOB33_X105Y137_IOB_X1Y137_I),
.I4(CLBLM_R_X3Y110_SLICE_X2Y110_DO6),
.I5(1'b1),
.O5(CLBLL_L_X2Y106_SLICE_X0Y106_CO5),
.O6(CLBLL_L_X2Y106_SLICE_X0Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffdfdfffdfffd)
  ) CLBLL_L_X2Y106_SLICE_X0Y106_BLUT (
.I0(RIOB33_X105Y137_IOB_X1Y137_I),
.I1(RIOB33_X105Y129_IOB_X1Y129_I),
.I2(RIOB33_X105Y127_IOB_X1Y128_I),
.I3(CLBLM_R_X3Y111_SLICE_X2Y111_CO6),
.I4(CLBLL_L_X2Y111_SLICE_X1Y111_DO6),
.I5(1'b1),
.O5(CLBLL_L_X2Y106_SLICE_X0Y106_BO5),
.O6(CLBLL_L_X2Y106_SLICE_X0Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffdfffdfffffff5)
  ) CLBLL_L_X2Y106_SLICE_X0Y106_ALUT (
.I0(RIOB33_X105Y137_IOB_X1Y137_I),
.I1(CLBLM_R_X3Y108_SLICE_X2Y108_DO6),
.I2(RIOB33_X105Y129_IOB_X1Y129_I),
.I3(RIOB33_X105Y127_IOB_X1Y128_I),
.I4(CLBLM_R_X3Y110_SLICE_X3Y110_DO6),
.I5(1'b1),
.O5(CLBLL_L_X2Y106_SLICE_X0Y106_AO5),
.O6(CLBLL_L_X2Y106_SLICE_X0Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y106_SLICE_X1Y106_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y106_SLICE_X1Y106_DO5),
.O6(CLBLL_L_X2Y106_SLICE_X1Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y106_SLICE_X1Y106_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y106_SLICE_X1Y106_CO5),
.O6(CLBLL_L_X2Y106_SLICE_X1Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y106_SLICE_X1Y106_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y106_SLICE_X1Y106_BO5),
.O6(CLBLL_L_X2Y106_SLICE_X1Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y106_SLICE_X1Y106_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y106_SLICE_X1Y106_AO5),
.O6(CLBLL_L_X2Y106_SLICE_X1Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y107_SLICE_X0Y107_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y107_SLICE_X0Y107_DO5),
.O6(CLBLL_L_X2Y107_SLICE_X0Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y107_SLICE_X0Y107_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y107_SLICE_X0Y107_CO5),
.O6(CLBLL_L_X2Y107_SLICE_X0Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y107_SLICE_X0Y107_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y107_SLICE_X0Y107_BO5),
.O6(CLBLL_L_X2Y107_SLICE_X0Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcfffffffeeffff)
  ) CLBLL_L_X2Y107_SLICE_X0Y107_ALUT (
.I0(CLBLL_L_X4Y107_SLICE_X5Y107_DO6),
.I1(RIOB33_X105Y129_IOB_X1Y129_I),
.I2(CLBLL_L_X2Y110_SLICE_X1Y110_DO6),
.I3(RIOB33_X105Y127_IOB_X1Y128_I),
.I4(RIOB33_X105Y137_IOB_X1Y137_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y107_SLICE_X0Y107_AO5),
.O6(CLBLL_L_X2Y107_SLICE_X0Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y107_SLICE_X1Y107_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y107_SLICE_X1Y107_DO5),
.O6(CLBLL_L_X2Y107_SLICE_X1Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y107_SLICE_X1Y107_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y107_SLICE_X1Y107_CO5),
.O6(CLBLL_L_X2Y107_SLICE_X1Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y107_SLICE_X1Y107_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y107_SLICE_X1Y107_BO5),
.O6(CLBLL_L_X2Y107_SLICE_X1Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hafafafaf23dcdc23)
  ) CLBLL_L_X2Y107_SLICE_X1Y107_ALUT (
.I0(RIOB33_X105Y129_IOB_X1Y129_I),
.I1(CLBLM_R_X3Y107_SLICE_X3Y107_AQ),
.I2(RIOB33_X105Y137_IOB_X1Y137_I),
.I3(CLBLL_L_X4Y107_SLICE_X5Y107_DO6),
.I4(CLBLM_R_X5Y106_SLICE_X7Y106_CO6),
.I5(1'b1),
.O5(CLBLL_L_X2Y107_SLICE_X1Y107_AO5),
.O6(CLBLL_L_X2Y107_SLICE_X1Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y108_SLICE_X0Y108_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y108_SLICE_X0Y108_DO5),
.O6(CLBLL_L_X2Y108_SLICE_X0Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y108_SLICE_X0Y108_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y108_SLICE_X0Y108_CO5),
.O6(CLBLL_L_X2Y108_SLICE_X0Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y108_SLICE_X0Y108_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y108_SLICE_X0Y108_BO5),
.O6(CLBLL_L_X2Y108_SLICE_X0Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y108_SLICE_X0Y108_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y108_SLICE_X0Y108_AO5),
.O6(CLBLL_L_X2Y108_SLICE_X0Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000010000000000)
  ) CLBLL_L_X2Y108_SLICE_X1Y108_DLUT (
.I0(RIOB33_X105Y133_IOB_X1Y133_I),
.I1(RIOB33_X105Y131_IOB_X1Y132_I),
.I2(CLBLL_L_X2Y114_SLICE_X0Y114_AO5),
.I3(CLBLL_L_X4Y115_SLICE_X5Y115_BQ),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(RIOB33_X105Y133_IOB_X1Y134_I),
.O5(CLBLL_L_X2Y108_SLICE_X1Y108_DO5),
.O6(CLBLL_L_X2Y108_SLICE_X1Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffbaffffffbaba)
  ) CLBLL_L_X2Y108_SLICE_X1Y108_CLUT (
.I0(CLBLM_R_X3Y111_SLICE_X3Y111_AO6),
.I1(CLBLL_L_X2Y109_SLICE_X0Y109_AO6),
.I2(LIOB33_X0Y67_IOB_X0Y67_I),
.I3(CLBLL_L_X2Y108_SLICE_X1Y108_AO6),
.I4(CLBLL_L_X2Y108_SLICE_X1Y108_DO6),
.I5(CLBLM_R_X7Y106_SLICE_X8Y106_AQ),
.O5(CLBLL_L_X2Y108_SLICE_X1Y108_CO5),
.O6(CLBLL_L_X2Y108_SLICE_X1Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffafffffeeffff)
  ) CLBLL_L_X2Y108_SLICE_X1Y108_BLUT (
.I0(RIOB33_X105Y131_IOB_X1Y132_I),
.I1(CLBLM_R_X3Y116_SLICE_X3Y116_AO6),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(RIOB33_X105Y133_IOB_X1Y134_I),
.I4(RIOB33_X105Y133_IOB_X1Y133_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y108_SLICE_X1Y108_BO5),
.O6(CLBLL_L_X2Y108_SLICE_X1Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff7ffffffffffbf)
  ) CLBLL_L_X2Y108_SLICE_X1Y108_ALUT (
.I0(RIOB33_X105Y131_IOB_X1Y132_I),
.I1(RIOB33_X105Y133_IOB_X1Y134_I),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(CLBLL_L_X2Y114_SLICE_X0Y114_AO6),
.I4(RIOB33_X105Y133_IOB_X1Y133_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y108_SLICE_X1Y108_AO5),
.O6(CLBLL_L_X2Y108_SLICE_X1Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h005000ff00500050)
  ) CLBLL_L_X2Y109_SLICE_X0Y109_DLUT (
.I0(CLBLL_L_X2Y112_SLICE_X0Y112_AO6),
.I1(1'b1),
.I2(LIOB33_X0Y67_IOB_X0Y67_I),
.I3(CLBLL_L_X2Y114_SLICE_X0Y114_AO5),
.I4(CLBLL_L_X2Y112_SLICE_X0Y112_AO5),
.I5(CLBLL_L_X4Y115_SLICE_X5Y115_BQ),
.O5(CLBLL_L_X2Y109_SLICE_X0Y109_DO5),
.O6(CLBLL_L_X2Y109_SLICE_X0Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'habaeabaaaeaeaaae)
  ) CLBLL_L_X2Y109_SLICE_X0Y109_CLUT (
.I0(CLBLL_L_X2Y107_SLICE_X1Y107_AO6),
.I1(RIOB33_X105Y133_IOB_X1Y134_I),
.I2(CLBLL_L_X2Y114_SLICE_X0Y114_AO5),
.I3(RIOB33_X105Y133_IOB_X1Y133_I),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(RIOB33_X105Y131_IOB_X1Y132_I),
.O5(CLBLL_L_X2Y109_SLICE_X0Y109_CO5),
.O6(CLBLL_L_X2Y109_SLICE_X0Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff1104ffefffef)
  ) CLBLL_L_X2Y109_SLICE_X0Y109_BLUT (
.I0(CLBLM_R_X3Y116_SLICE_X3Y116_AO6),
.I1(RIOB33_X105Y133_IOB_X1Y134_I),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(RIOB33_X105Y133_IOB_X1Y133_I),
.I4(CLBLL_L_X2Y109_SLICE_X0Y109_CO6),
.I5(1'b1),
.O5(CLBLL_L_X2Y109_SLICE_X0Y109_BO5),
.O6(CLBLL_L_X2Y109_SLICE_X0Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdffffffeeffffff)
  ) CLBLL_L_X2Y109_SLICE_X0Y109_ALUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(RIOB33_X105Y133_IOB_X1Y134_I),
.I2(CLBLL_L_X2Y114_SLICE_X0Y114_AO5),
.I3(RIOB33_X105Y133_IOB_X1Y133_I),
.I4(RIOB33_X105Y131_IOB_X1Y132_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y109_SLICE_X0Y109_AO5),
.O6(CLBLL_L_X2Y109_SLICE_X0Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff4444f4f4)
  ) CLBLL_L_X2Y109_SLICE_X1Y109_DLUT (
.I0(CLBLL_L_X2Y114_SLICE_X1Y114_AO6),
.I1(CLBLL_L_X4Y115_SLICE_X5Y115_BQ),
.I2(LIOB33_X0Y67_IOB_X0Y67_I),
.I3(1'b1),
.I4(CLBLL_L_X2Y109_SLICE_X0Y109_AO6),
.I5(CLBLM_R_X3Y111_SLICE_X3Y111_AO6),
.O5(CLBLL_L_X2Y109_SLICE_X1Y109_DO5),
.O6(CLBLL_L_X2Y109_SLICE_X1Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffefffffff)
  ) CLBLL_L_X2Y109_SLICE_X1Y109_CLUT (
.I0(CLBLL_L_X2Y112_SLICE_X1Y112_AO6),
.I1(CLBLL_L_X2Y109_SLICE_X0Y109_CO6),
.I2(CLBLL_L_X2Y110_SLICE_X0Y110_BO5),
.I3(CLBLL_L_X2Y110_SLICE_X1Y110_AO5),
.I4(CLBLL_L_X2Y108_SLICE_X1Y108_BO5),
.I5(CLBLL_L_X2Y111_SLICE_X1Y111_BO6),
.O5(CLBLL_L_X2Y109_SLICE_X1Y109_CO5),
.O6(CLBLL_L_X2Y109_SLICE_X1Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0200000000000000)
  ) CLBLL_L_X2Y109_SLICE_X1Y109_BLUT (
.I0(CLBLL_L_X2Y108_SLICE_X1Y108_BO5),
.I1(CLBLL_L_X2Y111_SLICE_X1Y111_BO6),
.I2(CLBLL_L_X2Y109_SLICE_X0Y109_CO6),
.I3(CLBLL_L_X2Y110_SLICE_X0Y110_BO5),
.I4(CLBLL_L_X2Y111_SLICE_X1Y111_AO5),
.I5(CLBLL_L_X2Y110_SLICE_X1Y110_AO5),
.O5(CLBLL_L_X2Y109_SLICE_X1Y109_BO5),
.O6(CLBLL_L_X2Y109_SLICE_X1Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0200000000000000)
  ) CLBLL_L_X2Y109_SLICE_X1Y109_ALUT (
.I0(CLBLL_L_X2Y108_SLICE_X1Y108_BO5),
.I1(CLBLL_L_X2Y111_SLICE_X1Y111_BO6),
.I2(CLBLL_L_X2Y109_SLICE_X0Y109_CO6),
.I3(CLBLL_L_X2Y108_SLICE_X1Y108_AO5),
.I4(CLBLL_L_X2Y110_SLICE_X0Y110_BO5),
.I5(CLBLL_L_X2Y110_SLICE_X1Y110_AO5),
.O5(CLBLL_L_X2Y109_SLICE_X1Y109_AO5),
.O6(CLBLL_L_X2Y109_SLICE_X1Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y110_SLICE_X0Y110_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y110_SLICE_X0Y110_DO5),
.O6(CLBLL_L_X2Y110_SLICE_X0Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00001022fffffffd)
  ) CLBLL_L_X2Y110_SLICE_X0Y110_CLUT (
.I0(RIOB33_X105Y133_IOB_X1Y133_I),
.I1(RIOB33_X105Y131_IOB_X1Y132_I),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(RIOB33_X105Y133_IOB_X1Y134_I),
.I4(CLBLM_R_X3Y116_SLICE_X3Y116_AO6),
.I5(1'b1),
.O5(CLBLL_L_X2Y110_SLICE_X0Y110_CO5),
.O6(CLBLL_L_X2Y110_SLICE_X0Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffbffffffeffffff)
  ) CLBLL_L_X2Y110_SLICE_X0Y110_BLUT (
.I0(CLBLM_R_X3Y116_SLICE_X3Y116_AO6),
.I1(RIOB33_X105Y131_IOB_X1Y132_I),
.I2(RIOB33_X105Y133_IOB_X1Y133_I),
.I3(RIOB33_X105Y133_IOB_X1Y134_I),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y110_SLICE_X0Y110_BO5),
.O6(CLBLL_L_X2Y110_SLICE_X0Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00a00000dfdfdfdf)
  ) CLBLL_L_X2Y110_SLICE_X0Y110_ALUT (
.I0(RIOB33_X105Y133_IOB_X1Y133_I),
.I1(RIOB33_X105Y133_IOB_X1Y134_I),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(CLBLL_L_X2Y114_SLICE_X0Y114_AO6),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y110_SLICE_X0Y110_AO5),
.O6(CLBLL_L_X2Y110_SLICE_X0Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000ff00ff00)
  ) CLBLL_L_X2Y110_SLICE_X1Y110_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X3Y110_SLICE_X2Y110_CO6),
.I4(1'b1),
.I5(CLBLL_L_X2Y112_SLICE_X1Y112_BO6),
.O5(CLBLL_L_X2Y110_SLICE_X1Y110_DO5),
.O6(CLBLL_L_X2Y110_SLICE_X1Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffdfffff)
  ) CLBLL_L_X2Y110_SLICE_X1Y110_CLUT (
.I0(CLBLL_L_X2Y111_SLICE_X1Y111_AO6),
.I1(CLBLL_L_X2Y110_SLICE_X0Y110_CO6),
.I2(CLBLL_L_X2Y110_SLICE_X0Y110_BO6),
.I3(CLBLL_L_X2Y109_SLICE_X0Y109_CO6),
.I4(CLBLL_L_X2Y110_SLICE_X1Y110_AO6),
.I5(CLBLL_L_X2Y111_SLICE_X1Y111_BO6),
.O5(CLBLL_L_X2Y110_SLICE_X1Y110_CO5),
.O6(CLBLL_L_X2Y110_SLICE_X1Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000400000000)
  ) CLBLL_L_X2Y110_SLICE_X1Y110_BLUT (
.I0(CLBLL_L_X2Y112_SLICE_X0Y112_CO6),
.I1(CLBLL_L_X2Y108_SLICE_X1Y108_AO5),
.I2(CLBLL_L_X2Y110_SLICE_X0Y110_AO6),
.I3(CLBLL_L_X2Y110_SLICE_X0Y110_CO6),
.I4(CLBLL_L_X2Y109_SLICE_X0Y109_CO6),
.I5(CLBLL_L_X2Y110_SLICE_X1Y110_AO5),
.O5(CLBLL_L_X2Y110_SLICE_X1Y110_BO5),
.O6(CLBLL_L_X2Y110_SLICE_X1Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffeffffffecfff)
  ) CLBLL_L_X2Y110_SLICE_X1Y110_ALUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(CLBLM_R_X3Y116_SLICE_X3Y116_AO6),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(RIOB33_X105Y133_IOB_X1Y133_I),
.I4(RIOB33_X105Y133_IOB_X1Y134_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y110_SLICE_X1Y110_AO5),
.O6(CLBLL_L_X2Y110_SLICE_X1Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y111_SLICE_X0Y111_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y111_SLICE_X0Y111_DO5),
.O6(CLBLL_L_X2Y111_SLICE_X0Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000a000000044)
  ) CLBLL_L_X2Y111_SLICE_X0Y111_CLUT (
.I0(RIOB33_X105Y131_IOB_X1Y132_I),
.I1(CLBLM_R_X5Y110_SLICE_X7Y110_AQ),
.I2(LIOB33_X0Y57_IOB_X0Y58_I),
.I3(CLBLL_L_X2Y114_SLICE_X0Y114_AO5),
.I4(CLBLL_L_X2Y112_SLICE_X1Y112_DO6),
.I5(RIOB33_X105Y131_IOB_X1Y131_I),
.O5(CLBLL_L_X2Y111_SLICE_X0Y111_CO5),
.O6(CLBLL_L_X2Y111_SLICE_X0Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haafaaaaeaaaaaaaa)
  ) CLBLL_L_X2Y111_SLICE_X0Y111_BLUT (
.I0(CLBLL_L_X2Y112_SLICE_X0Y112_CO6),
.I1(RIOB33_X105Y133_IOB_X1Y134_I),
.I2(RIOB33_X105Y133_IOB_X1Y133_I),
.I3(CLBLL_L_X2Y114_SLICE_X0Y114_AO6),
.I4(RIOB33_X105Y131_IOB_X1Y132_I),
.I5(RIOB33_X105Y131_IOB_X1Y131_I),
.O5(CLBLL_L_X2Y111_SLICE_X0Y111_BO5),
.O6(CLBLL_L_X2Y111_SLICE_X0Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0200000000000000)
  ) CLBLL_L_X2Y111_SLICE_X0Y111_ALUT (
.I0(RIOB33_X105Y131_IOB_X1Y132_I),
.I1(CLBLL_L_X2Y114_SLICE_X0Y114_AO5),
.I2(RIOB33_X105Y133_IOB_X1Y134_I),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(RIOB33_X105Y133_IOB_X1Y133_I),
.I5(LIOB33_X0Y67_IOB_X0Y68_I),
.O5(CLBLL_L_X2Y111_SLICE_X0Y111_AO5),
.O6(CLBLL_L_X2Y111_SLICE_X0Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffcdffcdcd)
  ) CLBLL_L_X2Y111_SLICE_X1Y111_DLUT (
.I0(CLBLL_L_X2Y109_SLICE_X0Y109_BO6),
.I1(CLBLM_R_X3Y111_SLICE_X2Y111_BO6),
.I2(CLBLL_L_X2Y111_SLICE_X0Y111_BO6),
.I3(CLBLM_R_X3Y112_SLICE_X3Y112_BO6),
.I4(CLBLM_R_X7Y115_SLICE_X9Y115_AQ),
.I5(CLBLM_R_X3Y111_SLICE_X2Y111_AO6),
.O5(CLBLL_L_X2Y111_SLICE_X1Y111_DO5),
.O6(CLBLL_L_X2Y111_SLICE_X1Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLL_L_X2Y111_SLICE_X1Y111_CLUT (
.I0(CLBLL_L_X2Y113_SLICE_X0Y113_AO6),
.I1(CLBLM_R_X3Y111_SLICE_X2Y111_BO6),
.I2(CLBLM_R_X3Y113_SLICE_X3Y113_DO6),
.I3(CLBLM_R_X3Y112_SLICE_X2Y112_CO6),
.I4(CLBLL_L_X4Y109_SLICE_X4Y109_CO6),
.I5(CLBLL_L_X2Y110_SLICE_X1Y110_BO6),
.O5(CLBLL_L_X2Y111_SLICE_X1Y111_CO5),
.O6(CLBLL_L_X2Y111_SLICE_X1Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h20212000ffffdfff)
  ) CLBLL_L_X2Y111_SLICE_X1Y111_BLUT (
.I0(RIOB33_X105Y131_IOB_X1Y132_I),
.I1(CLBLL_L_X2Y114_SLICE_X0Y114_AO6),
.I2(RIOB33_X105Y133_IOB_X1Y133_I),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(RIOB33_X105Y133_IOB_X1Y134_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y111_SLICE_X1Y111_BO5),
.O6(CLBLL_L_X2Y111_SLICE_X1Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffefffffffffd)
  ) CLBLL_L_X2Y111_SLICE_X1Y111_ALUT (
.I0(RIOB33_X105Y131_IOB_X1Y132_I),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(CLBLM_R_X3Y116_SLICE_X3Y116_AO6),
.I3(RIOB33_X105Y133_IOB_X1Y134_I),
.I4(RIOB33_X105Y133_IOB_X1Y133_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y111_SLICE_X1Y111_AO5),
.O6(CLBLL_L_X2Y111_SLICE_X1Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y112_SLICE_X0Y112_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y112_SLICE_X0Y112_DO5),
.O6(CLBLL_L_X2Y112_SLICE_X0Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000200)
  ) CLBLL_L_X2Y112_SLICE_X0Y112_CLUT (
.I0(RIOB33_X105Y135_IOB_X1Y136_I),
.I1(RIOB33_X105Y129_IOB_X1Y130_I),
.I2(CLBLL_L_X2Y107_SLICE_X1Y107_AO6),
.I3(RIOB33_X105Y135_IOB_X1Y135_I),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(CLBLL_L_X2Y110_SLICE_X0Y110_AO5),
.O5(CLBLL_L_X2Y112_SLICE_X0Y112_CO5),
.O6(CLBLL_L_X2Y112_SLICE_X0Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000080000000)
  ) CLBLL_L_X2Y112_SLICE_X0Y112_BLUT (
.I0(RIOB33_X105Y131_IOB_X1Y132_I),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(CLBLL_L_X4Y109_SLICE_X4Y109_BQ),
.I3(RIOB33_X105Y133_IOB_X1Y134_I),
.I4(RIOB33_X105Y133_IOB_X1Y133_I),
.I5(CLBLL_L_X2Y114_SLICE_X0Y114_AO6),
.O5(CLBLL_L_X2Y112_SLICE_X0Y112_BO5),
.O6(CLBLL_L_X2Y112_SLICE_X0Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff7fff7ffefffeff)
  ) CLBLL_L_X2Y112_SLICE_X0Y112_ALUT (
.I0(RIOB33_X105Y133_IOB_X1Y133_I),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(RIOB33_X105Y133_IOB_X1Y134_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y112_SLICE_X0Y112_AO5),
.O6(CLBLL_L_X2Y112_SLICE_X0Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0fffff0f0ffff)
  ) CLBLL_L_X2Y112_SLICE_X1Y112_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(RIOB33_X105Y133_IOB_X1Y133_I),
.I3(1'b1),
.I4(RIOB33_X105Y133_IOB_X1Y134_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y112_SLICE_X1Y112_DO5),
.O6(CLBLL_L_X2Y112_SLICE_X1Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00f0aafa00f0aafa)
  ) CLBLL_L_X2Y112_SLICE_X1Y112_CLUT (
.I0(CLBLL_L_X4Y109_SLICE_X4Y109_BQ),
.I1(1'b1),
.I2(CLBLM_L_X10Y114_SLICE_X13Y114_AQ),
.I3(CLBLM_R_X3Y112_SLICE_X3Y112_BO5),
.I4(CLBLM_R_X3Y112_SLICE_X2Y112_AO5),
.I5(1'b1),
.O5(CLBLL_L_X2Y112_SLICE_X1Y112_CO5),
.O6(CLBLL_L_X2Y112_SLICE_X1Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffefe)
  ) CLBLL_L_X2Y112_SLICE_X1Y112_BLUT (
.I0(CLBLL_L_X2Y113_SLICE_X1Y113_DO6),
.I1(CLBLL_L_X2Y114_SLICE_X1Y114_BO6),
.I2(CLBLM_R_X3Y113_SLICE_X3Y113_DO6),
.I3(1'b1),
.I4(CLBLL_L_X4Y109_SLICE_X4Y109_CO6),
.I5(CLBLL_L_X2Y112_SLICE_X1Y112_CO6),
.O5(CLBLL_L_X2Y112_SLICE_X1Y112_BO5),
.O6(CLBLL_L_X2Y112_SLICE_X1Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000004000000)
  ) CLBLL_L_X2Y112_SLICE_X1Y112_ALUT (
.I0(CLBLL_L_X2Y109_SLICE_X0Y109_AO5),
.I1(RIOB33_X105Y135_IOB_X1Y135_I),
.I2(RIOB33_X105Y129_IOB_X1Y129_I),
.I3(RIOB33_X105Y137_IOB_X1Y137_I),
.I4(RIOB33_X105Y135_IOB_X1Y136_I),
.I5(RIOB33_X105Y129_IOB_X1Y130_I),
.O5(CLBLL_L_X2Y112_SLICE_X1Y112_AO5),
.O6(CLBLL_L_X2Y112_SLICE_X1Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0010000000000000)
  ) CLBLL_L_X2Y113_SLICE_X0Y113_DLUT (
.I0(RIOB33_X105Y133_IOB_X1Y134_I),
.I1(RIOB33_X105Y133_IOB_X1Y133_I),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(CLBLM_R_X3Y116_SLICE_X3Y116_AO6),
.I4(CLBLM_L_X10Y114_SLICE_X13Y114_AQ),
.I5(RIOB33_X105Y131_IOB_X1Y132_I),
.O5(CLBLL_L_X2Y113_SLICE_X0Y113_DO5),
.O6(CLBLL_L_X2Y113_SLICE_X0Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0400040001010000)
  ) CLBLL_L_X2Y113_SLICE_X0Y113_CLUT (
.I0(CLBLL_L_X2Y114_SLICE_X0Y114_AO5),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(CLBLL_L_X2Y112_SLICE_X1Y112_DO6),
.I3(LIOB33_X0Y53_IOB_X0Y54_I),
.I4(CLBLM_R_X5Y115_SLICE_X6Y115_CQ),
.I5(RIOB33_X105Y131_IOB_X1Y132_I),
.O5(CLBLL_L_X2Y113_SLICE_X0Y113_CO5),
.O6(CLBLL_L_X2Y113_SLICE_X0Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0100000000000000)
  ) CLBLL_L_X2Y113_SLICE_X0Y113_BLUT (
.I0(RIOB33_X105Y133_IOB_X1Y134_I),
.I1(CLBLL_L_X2Y114_SLICE_X0Y114_AO5),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(RIOB33_X105Y133_IOB_X1Y133_I),
.I4(LIOB33_X0Y69_IOB_X0Y70_I),
.I5(RIOB33_X105Y131_IOB_X1Y132_I),
.O5(CLBLL_L_X2Y113_SLICE_X0Y113_BO5),
.O6(CLBLL_L_X2Y113_SLICE_X0Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLL_L_X2Y113_SLICE_X0Y113_ALUT (
.I0(CLBLL_L_X2Y113_SLICE_X0Y113_DO6),
.I1(CLBLM_R_X3Y113_SLICE_X2Y113_BO6),
.I2(CLBLL_L_X2Y113_SLICE_X1Y113_CO6),
.I3(CLBLL_L_X2Y113_SLICE_X0Y113_BO6),
.I4(CLBLL_L_X2Y112_SLICE_X0Y112_BO6),
.I5(CLBLL_L_X2Y113_SLICE_X0Y113_CO6),
.O5(CLBLL_L_X2Y113_SLICE_X0Y113_AO5),
.O6(CLBLL_L_X2Y113_SLICE_X0Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffdfffcfff5fff0)
  ) CLBLL_L_X2Y113_SLICE_X1Y113_DLUT (
.I0(CLBLL_L_X2Y113_SLICE_X1Y113_AO6),
.I1(CLBLL_L_X2Y107_SLICE_X1Y107_AO6),
.I2(CLBLL_L_X2Y112_SLICE_X0Y112_CO6),
.I3(CLBLL_L_X2Y113_SLICE_X1Y113_CO6),
.I4(CLBLL_L_X4Y114_SLICE_X4Y114_AQ),
.I5(CLBLL_L_X4Y110_SLICE_X5Y110_AQ),
.O5(CLBLL_L_X2Y113_SLICE_X1Y113_DO5),
.O6(CLBLL_L_X2Y113_SLICE_X1Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0133010100330000)
  ) CLBLL_L_X2Y113_SLICE_X1Y113_CLUT (
.I0(CLBLM_R_X3Y115_SLICE_X3Y115_AO6),
.I1(CLBLL_L_X2Y114_SLICE_X0Y114_AO5),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(CLBLL_L_X2Y112_SLICE_X0Y112_AO6),
.I4(LIOB33_X0Y59_IOB_X0Y59_I),
.I5(CLBLM_R_X3Y114_SLICE_X2Y114_BQ),
.O5(CLBLL_L_X2Y113_SLICE_X1Y113_CO5),
.O6(CLBLL_L_X2Y113_SLICE_X1Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000080000)
  ) CLBLL_L_X2Y113_SLICE_X1Y113_BLUT (
.I0(RIOB33_X105Y135_IOB_X1Y135_I),
.I1(RIOB33_X105Y137_IOB_X1Y137_I),
.I2(RIOB33_X105Y129_IOB_X1Y129_I),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(RIOB33_X105Y135_IOB_X1Y136_I),
.I5(RIOB33_X105Y129_IOB_X1Y130_I),
.O5(CLBLL_L_X2Y113_SLICE_X1Y113_BO5),
.O6(CLBLL_L_X2Y113_SLICE_X1Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdfffffffbffffff)
  ) CLBLL_L_X2Y113_SLICE_X1Y113_ALUT (
.I0(RIOB33_X105Y133_IOB_X1Y133_I),
.I1(RIOB33_X105Y131_IOB_X1Y132_I),
.I2(CLBLL_L_X2Y114_SLICE_X0Y114_AO5),
.I3(RIOB33_X105Y133_IOB_X1Y134_I),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y113_SLICE_X1Y113_AO5),
.O6(CLBLL_L_X2Y113_SLICE_X1Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y114_SLICE_X0Y114_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y114_SLICE_X0Y114_DO5),
.O6(CLBLL_L_X2Y114_SLICE_X0Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y114_SLICE_X0Y114_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y114_SLICE_X0Y114_CO5),
.O6(CLBLL_L_X2Y114_SLICE_X0Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0202000033023300)
  ) CLBLL_L_X2Y114_SLICE_X0Y114_BLUT (
.I0(RIOB33_X105Y131_IOB_X1Y132_I),
.I1(CLBLL_L_X2Y114_SLICE_X0Y114_AO5),
.I2(CLBLM_R_X3Y115_SLICE_X3Y115_AO6),
.I3(LIOB33_X0Y71_IOB_X0Y71_I),
.I4(LIOB33_X0Y55_IOB_X0Y55_I),
.I5(CLBLL_L_X2Y109_SLICE_X0Y109_AO5),
.O5(CLBLL_L_X2Y114_SLICE_X0Y114_BO5),
.O6(CLBLL_L_X2Y114_SLICE_X0Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffbfffffffffff7)
  ) CLBLL_L_X2Y114_SLICE_X0Y114_ALUT (
.I0(RIOB33_X105Y135_IOB_X1Y135_I),
.I1(RIOB33_X105Y137_IOB_X1Y137_I),
.I2(RIOB33_X105Y129_IOB_X1Y129_I),
.I3(RIOB33_X105Y129_IOB_X1Y130_I),
.I4(RIOB33_X105Y135_IOB_X1Y136_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y114_SLICE_X0Y114_AO5),
.O6(CLBLL_L_X2Y114_SLICE_X0Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y114_SLICE_X1Y114_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y114_SLICE_X1Y114_DO5),
.O6(CLBLL_L_X2Y114_SLICE_X1Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y114_SLICE_X1Y114_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y114_SLICE_X1Y114_CO5),
.O6(CLBLL_L_X2Y114_SLICE_X1Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3300f3f0bbaafbfa)
  ) CLBLL_L_X2Y114_SLICE_X1Y114_BLUT (
.I0(LIOB33_X0Y53_IOB_X0Y54_I),
.I1(CLBLL_L_X2Y114_SLICE_X1Y114_AO5),
.I2(CLBLM_R_X5Y115_SLICE_X6Y115_CQ),
.I3(LIOB33_X0Y69_IOB_X0Y70_I),
.I4(CLBLL_L_X2Y114_SLICE_X1Y114_AO6),
.I5(CLBLL_L_X2Y113_SLICE_X1Y113_AO5),
.O5(CLBLL_L_X2Y114_SLICE_X1Y114_BO5),
.O6(CLBLL_L_X2Y114_SLICE_X1Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffeffffdffff)
  ) CLBLL_L_X2Y114_SLICE_X1Y114_ALUT (
.I0(RIOB33_X105Y131_IOB_X1Y132_I),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(RIOB33_X105Y133_IOB_X1Y134_I),
.I3(CLBLL_L_X2Y114_SLICE_X0Y114_AO5),
.I4(RIOB33_X105Y133_IOB_X1Y133_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y114_SLICE_X1Y114_AO5),
.O6(CLBLL_L_X2Y114_SLICE_X1Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y106_SLICE_X4Y106_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y106_SLICE_X4Y106_DO5),
.O6(CLBLL_L_X4Y106_SLICE_X4Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y106_SLICE_X4Y106_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y106_SLICE_X4Y106_CO5),
.O6(CLBLL_L_X4Y106_SLICE_X4Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y106_SLICE_X4Y106_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y106_SLICE_X4Y106_BO5),
.O6(CLBLL_L_X4Y106_SLICE_X4Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y106_SLICE_X4Y106_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y106_SLICE_X4Y106_AO5),
.O6(CLBLL_L_X4Y106_SLICE_X4Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y106_SLICE_X5Y106_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y106_SLICE_X5Y106_AO6),
.Q(CLBLL_L_X4Y106_SLICE_X5Y106_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y106_SLICE_X5Y106_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y106_SLICE_X5Y106_BO6),
.Q(CLBLL_L_X4Y106_SLICE_X5Y106_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000040000)
  ) CLBLL_L_X4Y106_SLICE_X5Y106_DLUT (
.I0(RIOB33_X105Y133_IOB_X1Y133_I),
.I1(RIOB33_X105Y131_IOB_X1Y132_I),
.I2(RIOB33_X105Y133_IOB_X1Y134_I),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(CLBLM_L_X12Y106_SLICE_X16Y106_AQ),
.I5(CLBLM_R_X3Y116_SLICE_X3Y116_AO6),
.O5(CLBLL_L_X4Y106_SLICE_X5Y106_DO5),
.O6(CLBLL_L_X4Y106_SLICE_X5Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0200000000000000)
  ) CLBLL_L_X4Y106_SLICE_X5Y106_CLUT (
.I0(RIOB33_X105Y133_IOB_X1Y133_I),
.I1(CLBLM_R_X3Y116_SLICE_X3Y116_AO6),
.I2(RIOB33_X105Y133_IOB_X1Y134_I),
.I3(RIOB33_X105Y131_IOB_X1Y132_I),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(CLBLM_R_X5Y106_SLICE_X6Y106_AQ),
.O5(CLBLL_L_X4Y106_SLICE_X5Y106_CO5),
.O6(CLBLL_L_X4Y106_SLICE_X5Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0f5f5a0a0a0a0)
  ) CLBLL_L_X4Y106_SLICE_X5Y106_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(1'b1),
.I2(CLBLL_L_X4Y106_SLICE_X5Y106_AQ),
.I3(1'b1),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X7Y108_SLICE_X8Y108_CQ),
.O5(CLBLL_L_X4Y106_SLICE_X5Y106_BO5),
.O6(CLBLL_L_X4Y106_SLICE_X5Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aaccaaf0aaf0)
  ) CLBLL_L_X4Y106_SLICE_X5Y106_ALUT (
.I0(CLBLM_R_X5Y107_SLICE_X6Y107_CQ),
.I1(CLBLM_R_X3Y110_SLICE_X2Y110_DO6),
.I2(CLBLL_L_X4Y106_SLICE_X5Y106_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X7Y105_SLICE_X8Y105_BO5),
.O5(CLBLL_L_X4Y106_SLICE_X5Y106_AO5),
.O6(CLBLL_L_X4Y106_SLICE_X5Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y107_SLICE_X4Y107_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y107_SLICE_X4Y107_BO6),
.Q(CLBLL_L_X4Y107_SLICE_X4Y107_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y107_SLICE_X4Y107_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y107_SLICE_X4Y107_AO6),
.Q(CLBLL_L_X4Y107_SLICE_X4Y107_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y107_SLICE_X4Y107_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y107_SLICE_X4Y107_CO6),
.Q(CLBLL_L_X4Y107_SLICE_X4Y107_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y107_SLICE_X4Y107_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y107_SLICE_X4Y107_DO6),
.Q(CLBLL_L_X4Y107_SLICE_X4Y107_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hddccdccc11001000)
  ) CLBLL_L_X4Y107_SLICE_X4Y107_DLUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLL_L_X4Y107_SLICE_X4Y107_DQ),
.I3(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.I4(CLBLM_L_X10Y108_SLICE_X13Y108_AQ),
.I5(CLBLM_R_X3Y109_SLICE_X2Y109_A5Q),
.O5(CLBLL_L_X4Y107_SLICE_X4Y107_DO5),
.O6(CLBLL_L_X4Y107_SLICE_X4Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcf40c04fcf40c04)
  ) CLBLL_L_X4Y107_SLICE_X4Y107_CLUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLL_L_X4Y107_SLICE_X4Y107_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.I4(CLBLL_L_X4Y110_SLICE_X4Y110_CQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y107_SLICE_X4Y107_CO5),
.O6(CLBLL_L_X4Y107_SLICE_X4Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0e4a033ff33ff)
  ) CLBLL_L_X4Y107_SLICE_X4Y107_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y105_SLICE_X8Y105_CQ),
.I2(CLBLL_L_X4Y109_SLICE_X4Y109_AQ),
.I3(CLBLL_L_X4Y110_SLICE_X4Y110_AQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y107_SLICE_X4Y107_BO5),
.O6(CLBLL_L_X4Y107_SLICE_X4Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbbb8b8b88bb8b8b)
  ) CLBLL_L_X4Y107_SLICE_X4Y107_ALUT (
.I0(CLBLM_L_X10Y108_SLICE_X13Y108_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(LIOB33_X0Y53_IOB_X0Y53_I),
.I3(CLBLL_L_X4Y113_SLICE_X4Y113_BQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X3Y109_SLICE_X2Y109_AQ),
.O5(CLBLL_L_X4Y107_SLICE_X4Y107_AO5),
.O6(CLBLL_L_X4Y107_SLICE_X4Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y107_SLICE_X5Y107_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y107_SLICE_X5Y107_AO6),
.Q(CLBLL_L_X4Y107_SLICE_X5Y107_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hc33c3cc33cc3c33c)
  ) CLBLL_L_X4Y107_SLICE_X5Y107_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y108_SLICE_X2Y108_DO6),
.I2(CLBLL_L_X2Y111_SLICE_X1Y111_DO6),
.I3(CLBLM_R_X3Y110_SLICE_X3Y110_DO6),
.I4(CLBLL_L_X4Y107_SLICE_X5Y107_BO5),
.I5(CLBLL_L_X2Y110_SLICE_X1Y110_DO6),
.O5(CLBLL_L_X4Y107_SLICE_X5Y107_DO5),
.O6(CLBLL_L_X4Y107_SLICE_X5Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000080000)
  ) CLBLL_L_X4Y107_SLICE_X5Y107_CLUT (
.I0(RIOB33_X105Y133_IOB_X1Y133_I),
.I1(CLBLM_R_X7Y109_SLICE_X8Y109_AQ),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(RIOB33_X105Y133_IOB_X1Y134_I),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(CLBLM_R_X3Y116_SLICE_X3Y116_AO6),
.O5(CLBLL_L_X4Y107_SLICE_X5Y107_CO5),
.O6(CLBLL_L_X4Y107_SLICE_X5Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffff005aa5a55a)
  ) CLBLL_L_X4Y107_SLICE_X5Y107_BLUT (
.I0(CLBLM_R_X3Y109_SLICE_X2Y109_CO6),
.I1(1'b1),
.I2(CLBLM_R_X3Y110_SLICE_X2Y110_DO6),
.I3(CLBLM_R_X3Y110_SLICE_X3Y110_AO6),
.I4(CLBLM_R_X3Y111_SLICE_X2Y111_CO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y107_SLICE_X5Y107_BO5),
.O6(CLBLL_L_X4Y107_SLICE_X5Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff0ffaa00f000aa)
  ) CLBLL_L_X4Y107_SLICE_X5Y107_ALUT (
.I0(CLBLM_R_X5Y107_SLICE_X6Y107_CQ),
.I1(1'b1),
.I2(CLBLL_L_X4Y107_SLICE_X5Y107_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLL_L_X4Y112_SLICE_X4Y112_CO5),
.I5(CLBLM_R_X5Y107_SLICE_X6Y107_DQ),
.O5(CLBLL_L_X4Y107_SLICE_X5Y107_AO5),
.O6(CLBLL_L_X4Y107_SLICE_X5Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y108_SLICE_X4Y108_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y108_SLICE_X4Y108_AO6),
.Q(CLBLL_L_X4Y108_SLICE_X4Y108_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y108_SLICE_X4Y108_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y108_SLICE_X4Y108_BO6),
.Q(CLBLL_L_X4Y108_SLICE_X4Y108_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000045404540)
  ) CLBLL_L_X4Y108_SLICE_X4Y108_DLUT (
.I0(CLBLL_L_X2Y110_SLICE_X0Y110_AO5),
.I1(CLBLL_L_X4Y107_SLICE_X5Y107_AQ),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(CLBLL_L_X4Y108_SLICE_X4Y108_BQ),
.I4(1'b1),
.I5(CLBLM_R_X3Y116_SLICE_X3Y116_AO6),
.O5(CLBLL_L_X4Y108_SLICE_X4Y108_DO5),
.O6(CLBLL_L_X4Y108_SLICE_X4Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0405ffffffff)
  ) CLBLL_L_X4Y108_SLICE_X4Y108_CLUT (
.I0(LIOB33_X0Y53_IOB_X0Y53_I),
.I1(CLBLM_R_X3Y109_SLICE_X2Y109_AQ),
.I2(CLBLM_R_X5Y110_SLICE_X6Y110_B5Q),
.I3(CLBLL_L_X4Y113_SLICE_X4Y113_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLL_L_X4Y108_SLICE_X4Y108_CO5),
.O6(CLBLL_L_X4Y108_SLICE_X4Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'heeaaeeaaeca0eca0)
  ) CLBLL_L_X4Y108_SLICE_X4Y108_BLUT (
.I0(CLBLL_L_X4Y112_SLICE_X4Y112_CO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X7Y107_SLICE_X9Y107_CQ),
.I3(CLBLM_R_X5Y114_SLICE_X7Y114_CQ),
.I4(1'b1),
.I5(CLBLL_L_X4Y108_SLICE_X4Y108_BQ),
.O5(CLBLL_L_X4Y108_SLICE_X4Y108_BO5),
.O6(CLBLL_L_X4Y108_SLICE_X4Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbeaffaa51405500)
  ) CLBLL_L_X4Y108_SLICE_X4Y108_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLL_L_X4Y110_SLICE_X4Y110_AQ),
.I2(CLBLL_L_X4Y108_SLICE_X4Y108_AQ),
.I3(CLBLM_R_X7Y106_SLICE_X9Y106_AQ),
.I4(CLBLM_R_X7Y105_SLICE_X8Y105_CQ),
.I5(CLBLL_L_X4Y108_SLICE_X4Y108_BQ),
.O5(CLBLL_L_X4Y108_SLICE_X4Y108_AO5),
.O6(CLBLL_L_X4Y108_SLICE_X4Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000aa303030ba)
  ) CLBLL_L_X4Y108_SLICE_X5Y108_DLUT (
.I0(CLBLM_R_X7Y108_SLICE_X8Y108_BQ),
.I1(CLBLL_L_X2Y114_SLICE_X0Y114_AO6),
.I2(CLBLM_R_X5Y107_SLICE_X7Y107_B5Q),
.I3(CLBLM_R_X3Y116_SLICE_X3Y116_AO6),
.I4(CLBLL_L_X2Y109_SLICE_X0Y109_AO5),
.I5(CLBLL_L_X2Y108_SLICE_X1Y108_BO6),
.O5(CLBLL_L_X4Y108_SLICE_X5Y108_DO5),
.O6(CLBLL_L_X4Y108_SLICE_X5Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h1111000011f100f0)
  ) CLBLL_L_X4Y108_SLICE_X5Y108_CLUT (
.I0(CLBLL_L_X2Y112_SLICE_X0Y112_AO6),
.I1(CLBLM_R_X3Y116_SLICE_X3Y116_AO6),
.I2(CLBLM_R_X5Y109_SLICE_X7Y109_BQ),
.I3(CLBLL_L_X2Y114_SLICE_X0Y114_AO6),
.I4(CLBLM_R_X5Y105_SLICE_X7Y105_AQ),
.I5(CLBLL_L_X2Y108_SLICE_X1Y108_BO6),
.O5(CLBLL_L_X4Y108_SLICE_X5Y108_CO5),
.O6(CLBLL_L_X4Y108_SLICE_X5Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffbbaafffffbfa)
  ) CLBLL_L_X4Y108_SLICE_X5Y108_BLUT (
.I0(CLBLL_L_X4Y112_SLICE_X5Y112_CO6),
.I1(CLBLL_L_X2Y110_SLICE_X0Y110_BO6),
.I2(CLBLM_R_X7Y106_SLICE_X8Y106_CQ),
.I3(CLBLM_R_X5Y111_SLICE_X6Y111_BQ),
.I4(CLBLL_L_X4Y107_SLICE_X5Y107_CO6),
.I5(CLBLL_L_X2Y108_SLICE_X1Y108_AO5),
.O5(CLBLL_L_X4Y108_SLICE_X5Y108_BO5),
.O6(CLBLL_L_X4Y108_SLICE_X5Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00cc00cc05550fff)
  ) CLBLL_L_X4Y108_SLICE_X5Y108_ALUT (
.I0(CLBLL_L_X2Y111_SLICE_X1Y111_DO6),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X3Y110_SLICE_X3Y110_DO6),
.I3(CLBLM_R_X3Y109_SLICE_X2Y109_CO6),
.I4(CLBLM_R_X3Y108_SLICE_X2Y108_DO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y108_SLICE_X5Y108_AO5),
.O6(CLBLL_L_X4Y108_SLICE_X5Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y109_SLICE_X4Y109_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y109_SLICE_X4Y109_AO6),
.Q(CLBLL_L_X4Y109_SLICE_X4Y109_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y109_SLICE_X4Y109_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y109_SLICE_X4Y109_BO6),
.Q(CLBLL_L_X4Y109_SLICE_X4Y109_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff75ff75ff30ff30)
  ) CLBLL_L_X4Y109_SLICE_X4Y109_DLUT (
.I0(CLBLL_L_X2Y108_SLICE_X1Y108_AO6),
.I1(CLBLM_R_X3Y112_SLICE_X3Y112_BO6),
.I2(CLBLM_R_X11Y114_SLICE_X14Y114_AQ),
.I3(CLBLL_L_X4Y108_SLICE_X4Y108_DO6),
.I4(1'b1),
.I5(CLBLM_R_X7Y108_SLICE_X8Y108_AQ),
.O5(CLBLL_L_X4Y109_SLICE_X4Y109_DO5),
.O6(CLBLL_L_X4Y109_SLICE_X4Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5dff5d5d0cff0c0c)
  ) CLBLL_L_X4Y109_SLICE_X4Y109_CLUT (
.I0(CLBLL_L_X2Y108_SLICE_X1Y108_AO6),
.I1(CLBLM_R_X7Y109_SLICE_X9Y109_BQ),
.I2(CLBLL_L_X2Y110_SLICE_X0Y110_BO5),
.I3(CLBLL_L_X2Y111_SLICE_X1Y111_AO5),
.I4(CLBLM_L_X12Y112_SLICE_X16Y112_AQ),
.I5(CLBLM_R_X7Y107_SLICE_X8Y107_AQ),
.O5(CLBLL_L_X4Y109_SLICE_X4Y109_CO5),
.O6(CLBLL_L_X4Y109_SLICE_X4Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf044f044f044f0ee)
  ) CLBLL_L_X4Y109_SLICE_X4Y109_BLUT (
.I0(CLBLM_R_X7Y105_SLICE_X8Y105_BO5),
.I1(CLBLL_L_X4Y109_SLICE_X4Y109_BQ),
.I2(CLBLM_L_X12Y110_SLICE_X17Y110_BQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLL_L_X2Y110_SLICE_X1Y110_DO6),
.O5(CLBLL_L_X4Y109_SLICE_X4Y109_BO5),
.O6(CLBLL_L_X4Y109_SLICE_X4Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffa8a8a8a8a8a8)
  ) CLBLL_L_X4Y109_SLICE_X4Y109_ALUT (
.I0(CLBLL_L_X4Y112_SLICE_X4Y112_CO6),
.I1(CLBLL_L_X4Y110_SLICE_X4Y110_BQ),
.I2(CLBLL_L_X4Y109_SLICE_X4Y109_AQ),
.I3(1'b1),
.I4(CLBLM_R_X5Y111_SLICE_X7Y111_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLL_L_X4Y109_SLICE_X4Y109_AO5),
.O6(CLBLL_L_X4Y109_SLICE_X4Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y109_SLICE_X5Y109_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y109_SLICE_X5Y109_AO6),
.Q(CLBLL_L_X4Y109_SLICE_X5Y109_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0fafcfef00aaccee)
  ) CLBLL_L_X4Y109_SLICE_X5Y109_DLUT (
.I0(CLBLL_L_X4Y109_SLICE_X4Y109_AQ),
.I1(CLBLM_R_X7Y115_SLICE_X8Y115_AQ),
.I2(CLBLM_R_X3Y112_SLICE_X2Y112_AO5),
.I3(CLBLL_L_X2Y110_SLICE_X0Y110_BO5),
.I4(CLBLL_L_X2Y111_SLICE_X1Y111_AO5),
.I5(CLBLM_R_X5Y107_SLICE_X6Y107_AQ),
.O5(CLBLL_L_X4Y109_SLICE_X5Y109_DO5),
.O6(CLBLL_L_X4Y109_SLICE_X5Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000080)
  ) CLBLL_L_X4Y109_SLICE_X5Y109_CLUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(CLBLM_L_X12Y109_SLICE_X16Y109_D5Q),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(RIOB33_X105Y133_IOB_X1Y134_I),
.I4(RIOB33_X105Y133_IOB_X1Y133_I),
.I5(CLBLM_R_X3Y116_SLICE_X3Y116_AO6),
.O5(CLBLL_L_X4Y109_SLICE_X5Y109_CO5),
.O6(CLBLL_L_X4Y109_SLICE_X5Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffdcffdcdc)
  ) CLBLL_L_X4Y109_SLICE_X5Y109_BLUT (
.I0(CLBLM_R_X3Y112_SLICE_X2Y112_AO5),
.I1(CLBLL_L_X4Y106_SLICE_X5Y106_DO6),
.I2(CLBLL_L_X4Y106_SLICE_X5Y106_AQ),
.I3(CLBLL_L_X2Y110_SLICE_X0Y110_BO5),
.I4(CLBLL_L_X4Y113_SLICE_X5Y113_AQ),
.I5(CLBLL_L_X4Y109_SLICE_X5Y109_CO6),
.O5(CLBLL_L_X4Y109_SLICE_X5Y109_BO5),
.O6(CLBLL_L_X4Y109_SLICE_X5Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbbbb8b8bb88b888)
  ) CLBLL_L_X4Y109_SLICE_X5Y109_ALUT (
.I0(CLBLM_R_X5Y109_SLICE_X7Y109_DQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLL_L_X4Y109_SLICE_X5Y109_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_R_X7Y113_SLICE_X9Y113_DO6),
.I5(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.O5(CLBLL_L_X4Y109_SLICE_X5Y109_AO5),
.O6(CLBLL_L_X4Y109_SLICE_X5Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y110_SLICE_X4Y110_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y110_SLICE_X4Y110_BO5),
.Q(CLBLL_L_X4Y110_SLICE_X4Y110_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y110_SLICE_X4Y110_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y110_SLICE_X4Y110_CO5),
.Q(CLBLL_L_X4Y110_SLICE_X4Y110_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y110_SLICE_X4Y110_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y110_SLICE_X4Y110_AO6),
.Q(CLBLL_L_X4Y110_SLICE_X4Y110_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y110_SLICE_X4Y110_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y110_SLICE_X4Y110_BO6),
.Q(CLBLL_L_X4Y110_SLICE_X4Y110_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y110_SLICE_X4Y110_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y110_SLICE_X4Y110_CO6),
.Q(CLBLL_L_X4Y110_SLICE_X4Y110_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7733773355005500)
  ) CLBLL_L_X4Y110_SLICE_X4Y110_DLUT (
.I0(CLBLL_L_X2Y110_SLICE_X0Y110_CO5),
.I1(CLBLM_R_X3Y112_SLICE_X3Y112_BO6),
.I2(1'b1),
.I3(CLBLM_L_X10Y111_SLICE_X13Y111_AQ),
.I4(1'b1),
.I5(CLBLM_L_X10Y114_SLICE_X13Y114_BQ),
.O5(CLBLL_L_X4Y110_SLICE_X4Y110_DO5),
.O6(CLBLL_L_X4Y110_SLICE_X4Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f3c0c0bb88bb88)
  ) CLBLL_L_X4Y110_SLICE_X4Y110_CLUT (
.I0(CLBLM_R_X5Y110_SLICE_X6Y110_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLL_L_X4Y107_SLICE_X4Y107_A5Q),
.I3(CLBLL_L_X2Y111_SLICE_X1Y111_DO6),
.I4(CLBLM_R_X3Y108_SLICE_X2Y108_DO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y110_SLICE_X4Y110_CO5),
.O6(CLBLL_L_X4Y110_SLICE_X4Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hddcc1100fc30fc30)
  ) CLBLL_L_X4Y110_SLICE_X4Y110_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLL_L_X4Y107_SLICE_X4Y107_A5Q),
.I3(CLBLM_R_X5Y109_SLICE_X7Y109_A5Q),
.I4(CLBLL_L_X4Y110_SLICE_X5Y110_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y110_SLICE_X4Y110_BO5),
.O6(CLBLL_L_X4Y110_SLICE_X4Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff050005ff050005)
  ) CLBLL_L_X4Y110_SLICE_X4Y110_ALUT (
.I0(CLBLL_L_X4Y110_SLICE_X4Y110_B5Q),
.I1(1'b1),
.I2(CLBLM_R_X7Y105_SLICE_X8Y105_CQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLL_L_X4Y110_SLICE_X4Y110_C5Q),
.I5(1'b1),
.O5(CLBLL_L_X4Y110_SLICE_X4Y110_AO5),
.O6(CLBLL_L_X4Y110_SLICE_X4Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y110_SLICE_X5Y110_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y110_SLICE_X8Y110_DO6),
.Q(CLBLL_L_X4Y110_SLICE_X5Y110_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffff7f3fffff5f0)
  ) CLBLL_L_X4Y110_SLICE_X5Y110_DLUT (
.I0(CLBLL_L_X2Y110_SLICE_X0Y110_CO5),
.I1(CLBLM_R_X3Y112_SLICE_X3Y112_BO6),
.I2(CLBLM_R_X5Y114_SLICE_X6Y114_CO6),
.I3(CLBLM_L_X8Y111_SLICE_X11Y111_AQ),
.I4(CLBLL_L_X4Y108_SLICE_X5Y108_DO6),
.I5(CLBLL_L_X4Y111_SLICE_X4Y111_AQ),
.O5(CLBLL_L_X4Y110_SLICE_X5Y110_DO5),
.O6(CLBLL_L_X4Y110_SLICE_X5Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff4fff4fffffff4)
  ) CLBLL_L_X4Y110_SLICE_X5Y110_CLUT (
.I0(CLBLL_L_X2Y108_SLICE_X1Y108_AO5),
.I1(CLBLM_R_X5Y109_SLICE_X7Y109_DQ),
.I2(CLBLM_R_X5Y112_SLICE_X6Y112_DO6),
.I3(CLBLL_L_X4Y106_SLICE_X5Y106_CO6),
.I4(CLBLM_L_X8Y113_SLICE_X10Y113_AQ),
.I5(CLBLL_L_X2Y110_SLICE_X0Y110_BO5),
.O5(CLBLL_L_X4Y110_SLICE_X5Y110_CO5),
.O6(CLBLL_L_X4Y110_SLICE_X5Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h4f4f4444ff4fff44)
  ) CLBLL_L_X4Y110_SLICE_X5Y110_BLUT (
.I0(CLBLM_R_X3Y112_SLICE_X2Y112_AO5),
.I1(CLBLM_R_X5Y112_SLICE_X7Y112_AQ),
.I2(CLBLL_L_X2Y111_SLICE_X1Y111_AO5),
.I3(CLBLM_R_X7Y112_SLICE_X8Y112_AQ),
.I4(CLBLM_L_X8Y116_SLICE_X10Y116_DQ),
.I5(CLBLM_R_X3Y112_SLICE_X3Y112_BO5),
.O5(CLBLL_L_X4Y110_SLICE_X5Y110_BO5),
.O6(CLBLL_L_X4Y110_SLICE_X5Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3233030033330000)
  ) CLBLL_L_X4Y110_SLICE_X5Y110_ALUT (
.I0(CLBLM_R_X5Y110_SLICE_X7Y110_B5Q),
.I1(CLBLM_L_X8Y110_SLICE_X11Y110_BO5),
.I2(CLBLM_R_X5Y115_SLICE_X7Y115_CO6),
.I3(CLBLM_R_X5Y111_SLICE_X7Y111_AQ),
.I4(CLBLM_R_X5Y110_SLICE_X7Y110_BQ),
.I5(CLBLL_L_X4Y113_SLICE_X5Y113_BQ),
.O5(CLBLL_L_X4Y110_SLICE_X5Y110_AO5),
.O6(CLBLL_L_X4Y110_SLICE_X5Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y111_SLICE_X4Y111_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y111_SLICE_X4Y111_AO6),
.Q(CLBLL_L_X4Y111_SLICE_X4Y111_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y111_SLICE_X4Y111_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y111_SLICE_X4Y111_BO6),
.Q(CLBLL_L_X4Y111_SLICE_X4Y111_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y111_SLICE_X4Y111_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y111_SLICE_X4Y111_CO6),
.Q(CLBLL_L_X4Y111_SLICE_X4Y111_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h50dc50dcffff50dc)
  ) CLBLL_L_X4Y111_SLICE_X4Y111_DLUT (
.I0(CLBLL_L_X2Y108_SLICE_X1Y108_AO6),
.I1(CLBLL_L_X4Y114_SLICE_X4Y114_BQ),
.I2(CLBLM_R_X5Y111_SLICE_X6Y111_AQ),
.I3(CLBLL_L_X2Y111_SLICE_X1Y111_AO5),
.I4(CLBLM_R_X7Y114_SLICE_X8Y114_BQ),
.I5(CLBLL_L_X2Y110_SLICE_X0Y110_BO5),
.O5(CLBLL_L_X4Y111_SLICE_X4Y111_DO5),
.O6(CLBLL_L_X4Y111_SLICE_X4Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff5cff0c005c000c)
  ) CLBLL_L_X4Y111_SLICE_X4Y111_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLL_L_X4Y111_SLICE_X4Y111_CQ),
.I2(CLBLM_R_X7Y105_SLICE_X8Y105_BO5),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X3Y111_SLICE_X2Y111_CO6),
.I5(CLBLM_R_X7Y110_SLICE_X8Y110_CQ),
.O5(CLBLL_L_X4Y111_SLICE_X4Y111_CO5),
.O6(CLBLL_L_X4Y111_SLICE_X4Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccff0ff000)
  ) CLBLL_L_X4Y111_SLICE_X4Y111_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y109_SLICE_X6Y109_BQ),
.I2(CLBLL_L_X4Y112_SLICE_X4Y112_CO5),
.I3(CLBLM_R_X5Y111_SLICE_X6Y111_CQ),
.I4(CLBLL_L_X4Y111_SLICE_X4Y111_BQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLL_L_X4Y111_SLICE_X4Y111_BO5),
.O6(CLBLL_L_X4Y111_SLICE_X4Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfceefcee30223022)
  ) CLBLL_L_X4Y111_SLICE_X4Y111_ALUT (
.I0(CLBLM_R_X5Y112_SLICE_X7Y112_CQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLL_L_X4Y111_SLICE_X4Y111_AQ),
.I3(CLBLL_L_X4Y116_SLICE_X4Y116_BO6),
.I4(1'b1),
.I5(CLBLM_R_X5Y109_SLICE_X7Y109_B5Q),
.O5(CLBLL_L_X4Y111_SLICE_X4Y111_AO5),
.O6(CLBLL_L_X4Y111_SLICE_X4Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y111_SLICE_X5Y111_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y111_SLICE_X5Y111_AO6),
.Q(CLBLL_L_X4Y111_SLICE_X5Y111_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffbfffa)
  ) CLBLL_L_X4Y111_SLICE_X5Y111_DLUT (
.I0(CLBLL_L_X4Y108_SLICE_X5Y108_CO6),
.I1(CLBLL_L_X2Y111_SLICE_X1Y111_AO6),
.I2(CLBLL_L_X4Y114_SLICE_X5Y114_DO6),
.I3(CLBLM_R_X5Y113_SLICE_X7Y113_CO6),
.I4(CLBLM_R_X7Y111_SLICE_X9Y111_BQ),
.I5(CLBLL_L_X4Y113_SLICE_X5Y113_CO6),
.O5(CLBLL_L_X4Y111_SLICE_X5Y111_DO5),
.O6(CLBLL_L_X4Y111_SLICE_X5Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h4444444451114444)
  ) CLBLL_L_X4Y111_SLICE_X5Y111_CLUT (
.I0(CLBLM_L_X8Y110_SLICE_X11Y110_BO5),
.I1(CLBLL_L_X4Y113_SLICE_X5Y113_BQ),
.I2(CLBLM_R_X5Y110_SLICE_X7Y110_B5Q),
.I3(CLBLM_R_X5Y110_SLICE_X7Y110_BQ),
.I4(CLBLM_R_X5Y111_SLICE_X7Y111_AQ),
.I5(CLBLM_R_X5Y115_SLICE_X7Y115_CO6),
.O5(CLBLL_L_X4Y111_SLICE_X5Y111_CO5),
.O6(CLBLL_L_X4Y111_SLICE_X5Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h2000000000000000)
  ) CLBLL_L_X4Y111_SLICE_X5Y111_BLUT (
.I0(CLBLM_R_X5Y110_SLICE_X7Y110_B5Q),
.I1(CLBLM_R_X11Y112_SLICE_X15Y112_CO6),
.I2(CLBLM_R_X5Y111_SLICE_X7Y111_AQ),
.I3(CLBLL_L_X4Y113_SLICE_X5Y113_BQ),
.I4(CLBLM_R_X5Y115_SLICE_X7Y115_CO6),
.I5(CLBLM_R_X5Y110_SLICE_X7Y110_BQ),
.O5(CLBLL_L_X4Y111_SLICE_X5Y111_BO5),
.O6(CLBLL_L_X4Y111_SLICE_X5Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff54fffc005400fc)
  ) CLBLL_L_X4Y111_SLICE_X5Y111_ALUT (
.I0(CLBLL_L_X4Y110_SLICE_X4Y110_AQ),
.I1(CLBLM_R_X5Y105_SLICE_X7Y105_BQ),
.I2(CLBLL_L_X4Y111_SLICE_X5Y111_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y105_SLICE_X8Y105_CQ),
.I5(CLBLM_R_X5Y110_SLICE_X7Y110_BQ),
.O5(CLBLL_L_X4Y111_SLICE_X5Y111_AO5),
.O6(CLBLL_L_X4Y111_SLICE_X5Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y112_SLICE_X4Y112_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y112_SLICE_X4Y112_AO6),
.Q(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y112_SLICE_X4Y112_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y112_SLICE_X4Y112_BO6),
.Q(CLBLL_L_X4Y112_SLICE_X4Y112_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdfdfcfcfffdfffc)
  ) CLBLL_L_X4Y112_SLICE_X4Y112_DLUT (
.I0(CLBLL_L_X2Y108_SLICE_X1Y108_AO6),
.I1(CLBLM_R_X3Y114_SLICE_X2Y114_DO6),
.I2(CLBLL_L_X4Y112_SLICE_X5Y112_BO6),
.I3(CLBLM_L_X10Y111_SLICE_X12Y111_C5Q),
.I4(CLBLL_L_X4Y111_SLICE_X5Y111_AQ),
.I5(CLBLM_R_X3Y112_SLICE_X3Y112_BO5),
.O5(CLBLL_L_X4Y112_SLICE_X4Y112_DO5),
.O6(CLBLL_L_X4Y112_SLICE_X4Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h44444044ccccc0cc)
  ) CLBLL_L_X4Y112_SLICE_X4Y112_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLM_R_X11Y113_SLICE_X14Y113_CQ),
.I4(CLBLL_L_X4Y114_SLICE_X4Y114_BQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y112_SLICE_X4Y112_CO5),
.O6(CLBLL_L_X4Y112_SLICE_X4Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffeeffccaaaa0000)
  ) CLBLL_L_X4Y112_SLICE_X4Y112_BLUT (
.I0(CLBLL_L_X4Y117_SLICE_X4Y117_DQ),
.I1(CLBLL_L_X4Y112_SLICE_X4Y112_BQ),
.I2(1'b1),
.I3(CLBLM_R_X5Y109_SLICE_X7Y109_A5Q),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLL_L_X4Y112_SLICE_X4Y112_CO6),
.O5(CLBLL_L_X4Y112_SLICE_X4Y112_BO5),
.O6(CLBLL_L_X4Y112_SLICE_X4Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00a8a8ff00a8a8)
  ) CLBLL_L_X4Y112_SLICE_X4Y112_ALUT (
.I0(CLBLL_L_X4Y116_SLICE_X4Y116_BO6),
.I1(CLBLM_L_X8Y108_SLICE_X10Y108_BQ),
.I2(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.I3(CLBLL_L_X4Y111_SLICE_X4Y111_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y112_SLICE_X4Y112_AO5),
.O6(CLBLL_L_X4Y112_SLICE_X4Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y112_SLICE_X5Y112_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y112_SLICE_X5Y112_AO6),
.Q(CLBLL_L_X4Y112_SLICE_X5Y112_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffbbffbb)
  ) CLBLL_L_X4Y112_SLICE_X5Y112_DLUT (
.I0(CLBLM_R_X7Y108_SLICE_X8Y108_CQ),
.I1(CLBLM_R_X11Y113_SLICE_X14Y113_CQ),
.I2(1'b1),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(1'b1),
.I5(CLBLL_L_X4Y114_SLICE_X4Y114_BQ),
.O5(CLBLL_L_X4Y112_SLICE_X5Y112_DO5),
.O6(CLBLL_L_X4Y112_SLICE_X5Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0705030007050300)
  ) CLBLL_L_X4Y112_SLICE_X5Y112_CLUT (
.I0(CLBLL_L_X2Y112_SLICE_X0Y112_AO6),
.I1(CLBLL_L_X2Y112_SLICE_X0Y112_AO5),
.I2(CLBLL_L_X2Y114_SLICE_X0Y114_AO6),
.I3(CLBLM_R_X7Y112_SLICE_X8Y112_DQ),
.I4(RIOB33_X105Y111_IOB_X1Y112_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y112_SLICE_X5Y112_CO5),
.O6(CLBLL_L_X4Y112_SLICE_X5Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000011100010)
  ) CLBLL_L_X4Y112_SLICE_X5Y112_BLUT (
.I0(CLBLL_L_X26Y136_SLICE_X38Y136_AO6),
.I1(RIOB33_X105Y135_IOB_X1Y135_I),
.I2(CLBLL_L_X4Y112_SLICE_X5Y112_AQ),
.I3(RIOB33_X105Y135_IOB_X1Y136_I),
.I4(CLBLM_R_X7Y106_SLICE_X8Y106_BQ),
.I5(CLBLL_L_X2Y112_SLICE_X0Y112_AO5),
.O5(CLBLL_L_X4Y112_SLICE_X5Y112_BO5),
.O6(CLBLL_L_X4Y112_SLICE_X5Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffa8a8a8ffa8a8a8)
  ) CLBLL_L_X4Y112_SLICE_X5Y112_ALUT (
.I0(CLBLL_L_X4Y112_SLICE_X4Y112_CO6),
.I1(CLBLM_R_X7Y112_SLICE_X9Y112_AQ),
.I2(CLBLL_L_X4Y112_SLICE_X5Y112_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X11Y110_SLICE_X14Y110_D5Q),
.I5(1'b1),
.O5(CLBLL_L_X4Y112_SLICE_X5Y112_AO5),
.O6(CLBLL_L_X4Y112_SLICE_X5Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y113_SLICE_X4Y113_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y113_SLICE_X4Y113_AO6),
.Q(CLBLL_L_X4Y113_SLICE_X4Y113_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y113_SLICE_X4Y113_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y113_SLICE_X4Y113_BO6),
.Q(CLBLL_L_X4Y113_SLICE_X4Y113_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0050005000550000)
  ) CLBLL_L_X4Y113_SLICE_X4Y113_DLUT (
.I0(CLBLM_R_X3Y116_SLICE_X3Y116_AO6),
.I1(1'b1),
.I2(CLBLL_L_X4Y113_SLICE_X4Y113_AQ),
.I3(CLBLL_L_X2Y110_SLICE_X0Y110_AO5),
.I4(CLBLM_R_X5Y113_SLICE_X6Y113_AQ),
.I5(RIOB33_X105Y131_IOB_X1Y131_I),
.O5(CLBLL_L_X4Y113_SLICE_X4Y113_DO5),
.O6(CLBLL_L_X4Y113_SLICE_X4Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf2ff00000d0d0d0d)
  ) CLBLL_L_X4Y113_SLICE_X4Y113_CLUT (
.I0(CLBLM_R_X3Y115_SLICE_X2Y115_AQ),
.I1(CLBLM_R_X3Y109_SLICE_X2Y109_A5Q),
.I2(CLBLL_L_X4Y113_SLICE_X5Y113_B5Q),
.I3(CLBLM_L_X12Y113_SLICE_X17Y113_BQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y113_SLICE_X4Y113_CO5),
.O6(CLBLL_L_X4Y113_SLICE_X4Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'heccccccc20000000)
  ) CLBLL_L_X4Y113_SLICE_X4Y113_BLUT (
.I0(CLBLL_L_X4Y116_SLICE_X5Y116_A5Q),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X5Y112_SLICE_X6Y112_AQ),
.I3(CLBLL_L_X4Y114_SLICE_X4Y114_AQ),
.I4(CLBLM_R_X3Y112_SLICE_X3Y112_AQ),
.I5(CLBLM_R_X11Y113_SLICE_X14Y113_AQ),
.O5(CLBLL_L_X4Y113_SLICE_X4Y113_BO5),
.O6(CLBLL_L_X4Y113_SLICE_X4Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haafcaa30aafcaa30)
  ) CLBLL_L_X4Y113_SLICE_X4Y113_ALUT (
.I0(CLBLM_R_X5Y114_SLICE_X7Y114_AQ),
.I1(CLBLL_L_X4Y112_SLICE_X4Y112_CO5),
.I2(CLBLL_L_X4Y113_SLICE_X4Y113_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X5Y105_SLICE_X6Y105_BQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y113_SLICE_X4Y113_AO5),
.O6(CLBLL_L_X4Y113_SLICE_X4Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y113_SLICE_X5Y113_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y113_SLICE_X5Y113_BO5),
.Q(CLBLL_L_X4Y113_SLICE_X5Y113_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y113_SLICE_X5Y113_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y113_SLICE_X5Y113_AO6),
.Q(CLBLL_L_X4Y113_SLICE_X5Y113_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y113_SLICE_X5Y113_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y113_SLICE_X5Y113_BO6),
.Q(CLBLL_L_X4Y113_SLICE_X5Y113_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0030003000100010)
  ) CLBLL_L_X4Y113_SLICE_X5Y113_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X5Y111_SLICE_X6Y111_DO6),
.I2(CLBLM_R_X5Y115_SLICE_X7Y115_CO6),
.I3(CLBLM_R_X11Y112_SLICE_X15Y112_CO6),
.I4(1'b1),
.I5(CLBLL_L_X4Y113_SLICE_X4Y113_CO5),
.O5(CLBLL_L_X4Y113_SLICE_X5Y113_DO5),
.O6(CLBLL_L_X4Y113_SLICE_X5Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h000011d1000000c0)
  ) CLBLL_L_X4Y113_SLICE_X5Y113_CLUT (
.I0(CLBLM_R_X3Y116_SLICE_X3Y116_AO6),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(RIOB33_X105Y107_IOB_X1Y107_I),
.I3(CLBLL_L_X2Y114_SLICE_X0Y114_AO6),
.I4(CLBLL_L_X2Y110_SLICE_X0Y110_AO5),
.I5(CLBLM_R_X7Y113_SLICE_X8Y113_BQ),
.O5(CLBLL_L_X4Y113_SLICE_X5Y113_CO5),
.O6(CLBLL_L_X4Y113_SLICE_X5Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafaaaaafc0cfc0c)
  ) CLBLL_L_X4Y113_SLICE_X5Y113_BLUT (
.I0(CLBLL_L_X4Y111_SLICE_X5Y111_CO6),
.I1(CLBLL_L_X4Y111_SLICE_X5Y111_BO6),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y112_SLICE_X9Y112_AQ),
.I4(CLBLM_L_X12Y113_SLICE_X16Y113_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y113_SLICE_X5Y113_BO5),
.O6(CLBLL_L_X4Y113_SLICE_X5Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffa00faff500050)
  ) CLBLL_L_X4Y113_SLICE_X5Y113_ALUT (
.I0(CLBLL_L_X4Y112_SLICE_X4Y112_CO5),
.I1(1'b1),
.I2(CLBLL_L_X4Y113_SLICE_X5Y113_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLL_L_X4Y113_SLICE_X4Y113_AQ),
.I5(CLBLM_R_X7Y115_SLICE_X9Y115_A5Q),
.O5(CLBLL_L_X4Y113_SLICE_X5Y113_AO5),
.O6(CLBLL_L_X4Y113_SLICE_X5Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y114_SLICE_X4Y114_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y114_SLICE_X4Y114_AO6),
.Q(CLBLL_L_X4Y114_SLICE_X4Y114_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y114_SLICE_X4Y114_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y114_SLICE_X4Y114_BO6),
.Q(CLBLL_L_X4Y114_SLICE_X4Y114_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y114_SLICE_X4Y114_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y114_SLICE_X4Y114_CO6),
.Q(CLBLL_L_X4Y114_SLICE_X4Y114_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000800000)
  ) CLBLL_L_X4Y114_SLICE_X4Y114_DLUT (
.I0(RIOB33_X105Y133_IOB_X1Y133_I),
.I1(RIOB33_X105Y133_IOB_X1Y134_I),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(CLBLL_L_X2Y114_SLICE_X0Y114_AO6),
.I4(CLBLM_R_X7Y110_SLICE_X8Y110_AQ),
.I5(RIOB33_X105Y131_IOB_X1Y131_I),
.O5(CLBLL_L_X4Y114_SLICE_X4Y114_DO5),
.O6(CLBLL_L_X4Y114_SLICE_X4Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f0eef000f0ee)
  ) CLBLL_L_X4Y114_SLICE_X4Y114_CLUT (
.I0(CLBLM_R_X7Y113_SLICE_X9Y113_A5Q),
.I1(CLBLL_L_X4Y114_SLICE_X4Y114_CQ),
.I2(CLBLM_R_X5Y112_SLICE_X7Y112_CQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLL_L_X4Y113_SLICE_X5Y113_DO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y114_SLICE_X4Y114_CO5),
.O6(CLBLL_L_X4Y114_SLICE_X4Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hef45aa00ee44aa00)
  ) CLBLL_L_X4Y114_SLICE_X4Y114_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLL_L_X4Y114_SLICE_X4Y114_BQ),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLL_L_X4Y111_SLICE_X4Y111_CQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X11Y113_SLICE_X14Y113_CQ),
.O5(CLBLL_L_X4Y114_SLICE_X4Y114_BO5),
.O6(CLBLL_L_X4Y114_SLICE_X4Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccfcccfc00f000f0)
  ) CLBLL_L_X4Y114_SLICE_X4Y114_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y114_SLICE_X8Y114_AQ),
.I2(CLBLL_L_X4Y114_SLICE_X4Y114_AQ),
.I3(CLBLL_L_X4Y108_SLICE_X4Y108_CO6),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLL_L_X4Y114_SLICE_X4Y114_AO5),
.O6(CLBLL_L_X4Y114_SLICE_X4Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y114_SLICE_X5Y114_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y114_SLICE_X5Y114_AO6),
.Q(CLBLL_L_X4Y114_SLICE_X5Y114_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h1131113100300030)
  ) CLBLL_L_X4Y114_SLICE_X5Y114_DLUT (
.I0(CLBLL_L_X2Y112_SLICE_X0Y112_AO5),
.I1(CLBLL_L_X2Y114_SLICE_X0Y114_AO6),
.I2(RIOB33_X105Y115_IOB_X1Y115_I),
.I3(CLBLL_L_X2Y109_SLICE_X0Y109_AO5),
.I4(1'b1),
.I5(CLBLM_L_X10Y113_SLICE_X13Y113_DQ),
.O5(CLBLL_L_X4Y114_SLICE_X5Y114_DO5),
.O6(CLBLL_L_X4Y114_SLICE_X5Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffbfffbfff)
  ) CLBLL_L_X4Y114_SLICE_X5Y114_CLUT (
.I0(CLBLM_R_X5Y111_SLICE_X6Y111_DO6),
.I1(CLBLM_R_X3Y114_SLICE_X2Y114_BQ),
.I2(CLBLM_R_X3Y113_SLICE_X3Y113_AQ),
.I3(CLBLM_R_X5Y115_SLICE_X7Y115_CO6),
.I4(1'b1),
.I5(CLBLM_R_X11Y112_SLICE_X15Y112_CO6),
.O5(CLBLL_L_X4Y114_SLICE_X5Y114_CO5),
.O6(CLBLL_L_X4Y114_SLICE_X5Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000008000000000)
  ) CLBLL_L_X4Y114_SLICE_X5Y114_BLUT (
.I0(CLBLM_R_X3Y113_SLICE_X3Y113_AQ),
.I1(CLBLM_R_X5Y115_SLICE_X7Y115_CO6),
.I2(CLBLL_L_X4Y114_SLICE_X5Y114_AQ),
.I3(CLBLM_R_X5Y111_SLICE_X6Y111_DO6),
.I4(CLBLM_R_X11Y112_SLICE_X15Y112_CO6),
.I5(CLBLM_R_X3Y114_SLICE_X2Y114_BQ),
.O5(CLBLL_L_X4Y114_SLICE_X5Y114_BO5),
.O6(CLBLL_L_X4Y114_SLICE_X5Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hb888b8888b888b88)
  ) CLBLL_L_X4Y114_SLICE_X5Y114_ALUT (
.I0(CLBLM_R_X11Y110_SLICE_X14Y110_CQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLL_L_X4Y114_SLICE_X5Y114_AQ),
.I3(CLBLL_L_X4Y113_SLICE_X4Y113_CO6),
.I4(1'b1),
.I5(CLBLL_L_X4Y114_SLICE_X5Y114_CO6),
.O5(CLBLL_L_X4Y114_SLICE_X5Y114_AO5),
.O6(CLBLL_L_X4Y114_SLICE_X5Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y115_SLICE_X4Y115_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y115_SLICE_X4Y115_DO5),
.O6(CLBLL_L_X4Y115_SLICE_X4Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y115_SLICE_X4Y115_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y115_SLICE_X4Y115_CO5),
.O6(CLBLL_L_X4Y115_SLICE_X4Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y115_SLICE_X4Y115_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y115_SLICE_X4Y115_BO5),
.O6(CLBLL_L_X4Y115_SLICE_X4Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000004000000000)
  ) CLBLL_L_X4Y115_SLICE_X4Y115_ALUT (
.I0(RIOB33_X105Y133_IOB_X1Y133_I),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(CLBLM_R_X5Y111_SLICE_X7Y111_BQ),
.I3(RIOB33_X105Y133_IOB_X1Y134_I),
.I4(CLBLM_R_X3Y116_SLICE_X3Y116_AO6),
.I5(RIOB33_X105Y131_IOB_X1Y132_I),
.O5(CLBLL_L_X4Y115_SLICE_X4Y115_AO5),
.O6(CLBLL_L_X4Y115_SLICE_X4Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y115_SLICE_X5Y115_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y115_SLICE_X5Y115_AO5),
.Q(CLBLL_L_X4Y115_SLICE_X5Y115_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y115_SLICE_X5Y115_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y115_SLICE_X5Y115_AO6),
.Q(CLBLL_L_X4Y115_SLICE_X5Y115_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y115_SLICE_X5Y115_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y115_SLICE_X5Y115_BO6),
.Q(CLBLL_L_X4Y115_SLICE_X5Y115_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y115_SLICE_X5Y115_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y115_SLICE_X5Y115_CO6),
.Q(CLBLL_L_X4Y115_SLICE_X5Y115_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y115_SLICE_X5Y115_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y115_SLICE_X5Y115_DO5),
.O6(CLBLL_L_X4Y115_SLICE_X5Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaacfcfaaaac0c0)
  ) CLBLL_L_X4Y115_SLICE_X5Y115_CLUT (
.I0(CLBLL_L_X4Y116_SLICE_X5Y116_AQ),
.I1(CLBLL_L_X4Y115_SLICE_X5Y115_CQ),
.I2(CLBLL_L_X4Y113_SLICE_X5Y113_DO6),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X5Y110_SLICE_X6Y110_BQ),
.O5(CLBLL_L_X4Y115_SLICE_X5Y115_CO5),
.O6(CLBLL_L_X4Y115_SLICE_X5Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff54ff5400540054)
  ) CLBLL_L_X4Y115_SLICE_X5Y115_BLUT (
.I0(CLBLL_L_X4Y113_SLICE_X5Y113_DO6),
.I1(CLBLL_L_X4Y115_SLICE_X5Y115_BQ),
.I2(CLBLL_L_X4Y116_SLICE_X4Y116_A5Q),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLL_L_X4Y115_SLICE_X5Y115_A5Q),
.O5(CLBLL_L_X4Y115_SLICE_X5Y115_BO5),
.O6(CLBLL_L_X4Y115_SLICE_X5Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaa00aaf0ccf0cc)
  ) CLBLL_L_X4Y115_SLICE_X5Y115_ALUT (
.I0(CLBLM_R_X3Y110_SLICE_X2Y110_DO6),
.I1(CLBLM_R_X3Y109_SLICE_X2Y109_CO6),
.I2(CLBLM_L_X8Y117_SLICE_X10Y117_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y117_SLICE_X9Y117_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y115_SLICE_X5Y115_AO5),
.O6(CLBLL_L_X4Y115_SLICE_X5Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y116_SLICE_X4Y116_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y117_SLICE_X5Y117_BO6),
.Q(CLBLL_L_X4Y116_SLICE_X4Y116_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y116_SLICE_X4Y116_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y116_SLICE_X4Y116_AO6),
.Q(CLBLL_L_X4Y116_SLICE_X4Y116_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y116_SLICE_X4Y116_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y116_SLICE_X4Y116_DO5),
.O6(CLBLL_L_X4Y116_SLICE_X4Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y116_SLICE_X4Y116_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y116_SLICE_X4Y116_CO5),
.O6(CLBLL_L_X4Y116_SLICE_X4Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccc0cc44444444)
  ) CLBLL_L_X4Y116_SLICE_X4Y116_BLUT (
.I0(CLBLM_R_X5Y116_SLICE_X6Y116_DQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLM_R_X11Y113_SLICE_X14Y113_CQ),
.I4(CLBLM_L_X12Y112_SLICE_X16Y112_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y116_SLICE_X4Y116_BO5),
.O6(CLBLL_L_X4Y116_SLICE_X4Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff04ff4000040040)
  ) CLBLL_L_X4Y116_SLICE_X4Y116_ALUT (
.I0(CLBLM_R_X5Y116_SLICE_X6Y116_DQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLL_L_X4Y116_SLICE_X4Y116_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLL_L_X4Y117_SLICE_X5Y117_BO5),
.I5(CLBLL_L_X4Y113_SLICE_X5Y113_B5Q),
.O5(CLBLL_L_X4Y116_SLICE_X4Y116_AO5),
.O6(CLBLL_L_X4Y116_SLICE_X4Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y116_SLICE_X5Y116_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y116_SLICE_X6Y116_AO6),
.Q(CLBLL_L_X4Y116_SLICE_X5Y116_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y116_SLICE_X5Y116_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y116_SLICE_X5Y116_BO5),
.Q(CLBLL_L_X4Y116_SLICE_X5Y116_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y116_SLICE_X5Y116_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y116_SLICE_X5Y116_AO6),
.Q(CLBLL_L_X4Y116_SLICE_X5Y116_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y116_SLICE_X5Y116_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y116_SLICE_X5Y116_BO6),
.Q(CLBLL_L_X4Y116_SLICE_X5Y116_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y116_SLICE_X5Y116_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y116_SLICE_X5Y116_DO5),
.O6(CLBLL_L_X4Y116_SLICE_X5Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y116_SLICE_X5Y116_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y116_SLICE_X5Y116_CO5),
.O6(CLBLL_L_X4Y116_SLICE_X5Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafa5050dd88dd88)
  ) CLBLL_L_X4Y116_SLICE_X5Y116_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLL_L_X4Y116_SLICE_X5Y116_BQ),
.I2(RIOB33_X105Y127_IOB_X1Y127_I),
.I3(CLBLM_R_X7Y117_SLICE_X9Y117_BQ),
.I4(CLBLL_L_X4Y111_SLICE_X5Y111_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y116_SLICE_X5Y116_BO5),
.O6(CLBLL_L_X4Y116_SLICE_X5Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc05cc00cc50cc00)
  ) CLBLL_L_X4Y116_SLICE_X5Y116_ALUT (
.I0(CLBLM_R_X5Y116_SLICE_X6Y116_DQ),
.I1(CLBLM_L_X8Y114_SLICE_X10Y114_BQ),
.I2(CLBLL_L_X4Y116_SLICE_X5Y116_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLL_L_X4Y118_SLICE_X4Y118_A5Q),
.O5(CLBLL_L_X4Y116_SLICE_X5Y116_AO5),
.O6(CLBLL_L_X4Y116_SLICE_X5Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y117_SLICE_X4Y117_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y117_SLICE_X4Y117_AO6),
.Q(CLBLL_L_X4Y117_SLICE_X4Y117_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y117_SLICE_X4Y117_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y117_SLICE_X4Y117_BO6),
.Q(CLBLL_L_X4Y117_SLICE_X4Y117_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y117_SLICE_X4Y117_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y117_SLICE_X4Y117_CO6),
.Q(CLBLL_L_X4Y117_SLICE_X4Y117_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y117_SLICE_X4Y117_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y117_SLICE_X4Y117_DO6),
.Q(CLBLL_L_X4Y117_SLICE_X4Y117_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h888d888888d88888)
  ) CLBLL_L_X4Y117_SLICE_X4Y117_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y116_SLICE_X8Y116_BQ),
.I2(CLBLL_L_X4Y117_SLICE_X4Y117_DQ),
.I3(CLBLM_R_X5Y116_SLICE_X6Y116_DQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLL_L_X4Y118_SLICE_X4Y118_DO5),
.O5(CLBLL_L_X4Y117_SLICE_X4Y117_DO5),
.O6(CLBLL_L_X4Y117_SLICE_X4Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hbf15ff55ea40aa00)
  ) CLBLL_L_X4Y117_SLICE_X4Y117_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLL_L_X4Y116_SLICE_X4Y116_AQ),
.I2(CLBLL_L_X4Y117_SLICE_X5Y117_BO5),
.I3(CLBLM_R_X7Y106_SLICE_X9Y106_AQ),
.I4(CLBLL_L_X4Y117_SLICE_X4Y117_BQ),
.I5(CLBLM_R_X5Y116_SLICE_X6Y116_DQ),
.O5(CLBLL_L_X4Y117_SLICE_X4Y117_CO5),
.O6(CLBLL_L_X4Y117_SLICE_X4Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff002828ff008888)
  ) CLBLL_L_X4Y117_SLICE_X4Y117_BLUT (
.I0(CLBLL_L_X4Y116_SLICE_X4Y116_BO5),
.I1(CLBLL_L_X4Y117_SLICE_X4Y117_BQ),
.I2(CLBLL_L_X4Y116_SLICE_X4Y116_AQ),
.I3(CLBLM_R_X5Y110_SLICE_X6Y110_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLL_L_X4Y117_SLICE_X5Y117_BO5),
.O5(CLBLL_L_X4Y117_SLICE_X4Y117_BO5),
.O6(CLBLL_L_X4Y117_SLICE_X4Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000028a028a0)
  ) CLBLL_L_X4Y117_SLICE_X4Y117_ALUT (
.I0(CLBLL_L_X4Y116_SLICE_X4Y116_BO5),
.I1(CLBLL_L_X4Y117_SLICE_X4Y117_DQ),
.I2(CLBLL_L_X4Y117_SLICE_X4Y117_AQ),
.I3(CLBLL_L_X4Y118_SLICE_X4Y118_DO5),
.I4(CLBLM_R_X5Y111_SLICE_X7Y111_BQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLL_L_X4Y117_SLICE_X4Y117_AO5),
.O6(CLBLL_L_X4Y117_SLICE_X4Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y117_SLICE_X5Y117_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y117_SLICE_X5Y117_AO6),
.Q(CLBLL_L_X4Y117_SLICE_X5Y117_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y117_SLICE_X5Y117_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y117_SLICE_X5Y117_DO5),
.O6(CLBLL_L_X4Y117_SLICE_X5Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y117_SLICE_X5Y117_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y117_SLICE_X5Y117_CO5),
.O6(CLBLL_L_X4Y117_SLICE_X5Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f3c0c0a000a000)
  ) CLBLL_L_X4Y117_SLICE_X5Y117_BLUT (
.I0(CLBLL_L_X4Y118_SLICE_X4Y118_DO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLL_L_X4Y117_SLICE_X5Y117_AQ),
.I3(CLBLL_L_X4Y118_SLICE_X4Y118_BQ),
.I4(CLBLM_R_X5Y116_SLICE_X7Y116_BQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y117_SLICE_X5Y117_BO5),
.O6(CLBLL_L_X4Y117_SLICE_X5Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff4800000048)
  ) CLBLL_L_X4Y117_SLICE_X5Y117_ALUT (
.I0(CLBLL_L_X4Y118_SLICE_X4Y118_DO6),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLL_L_X4Y117_SLICE_X5Y117_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X5Y116_SLICE_X6Y116_DQ),
.I5(CLBLM_L_X8Y115_SLICE_X10Y115_A5Q),
.O5(CLBLL_L_X4Y117_SLICE_X5Y117_AO5),
.O6(CLBLL_L_X4Y117_SLICE_X5Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y118_SLICE_X4Y118_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y118_SLICE_X4Y118_CO6),
.Q(CLBLL_L_X4Y118_SLICE_X4Y118_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y118_SLICE_X4Y118_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y118_SLICE_X4Y118_AO6),
.Q(CLBLL_L_X4Y118_SLICE_X4Y118_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y118_SLICE_X4Y118_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y118_SLICE_X4Y118_BO6),
.Q(CLBLL_L_X4Y118_SLICE_X4Y118_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000088008800)
  ) CLBLL_L_X4Y118_SLICE_X4Y118_DLUT (
.I0(CLBLL_L_X4Y116_SLICE_X5Y116_AQ),
.I1(CLBLL_L_X4Y118_SLICE_X4Y118_AQ),
.I2(CLBLL_L_X4Y117_SLICE_X4Y117_DQ),
.I3(CLBLL_L_X4Y118_SLICE_X4Y118_A5Q),
.I4(CLBLL_L_X4Y117_SLICE_X4Y117_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y118_SLICE_X4Y118_DO5),
.O6(CLBLL_L_X4Y118_SLICE_X4Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaba001010101010)
  ) CLBLL_L_X4Y118_SLICE_X4Y118_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y116_SLICE_X6Y116_DQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLL_L_X4Y118_SLICE_X4Y118_A5Q),
.I4(CLBLM_R_X7Y118_SLICE_X9Y118_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y118_SLICE_X4Y118_CO5),
.O6(CLBLL_L_X4Y118_SLICE_X4Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00000f2f80208)
  ) CLBLL_L_X4Y118_SLICE_X4Y118_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLL_L_X4Y118_SLICE_X4Y118_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X3Y118_SLICE_X3Y118_AO6),
.I4(CLBLM_L_X10Y117_SLICE_X12Y117_BQ),
.I5(CLBLM_R_X5Y116_SLICE_X6Y116_DQ),
.O5(CLBLL_L_X4Y118_SLICE_X4Y118_BO5),
.O6(CLBLL_L_X4Y118_SLICE_X4Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbe3caa00eeccaa00)
  ) CLBLL_L_X4Y118_SLICE_X4Y118_ALUT (
.I0(CLBLL_L_X4Y114_SLICE_X4Y114_CQ),
.I1(CLBLL_L_X4Y118_SLICE_X4Y118_AQ),
.I2(CLBLL_L_X4Y116_SLICE_X5Y116_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLL_L_X4Y118_SLICE_X4Y118_CO5),
.I5(CLBLL_L_X4Y118_SLICE_X4Y118_A5Q),
.O5(CLBLL_L_X4Y118_SLICE_X4Y118_AO5),
.O6(CLBLL_L_X4Y118_SLICE_X4Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y118_SLICE_X5Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y118_SLICE_X5Y118_DO5),
.O6(CLBLL_L_X4Y118_SLICE_X5Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y118_SLICE_X5Y118_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y118_SLICE_X5Y118_CO5),
.O6(CLBLL_L_X4Y118_SLICE_X5Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y118_SLICE_X5Y118_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y118_SLICE_X5Y118_BO5),
.O6(CLBLL_L_X4Y118_SLICE_X5Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y118_SLICE_X5Y118_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y118_SLICE_X5Y118_AO5),
.O6(CLBLL_L_X4Y118_SLICE_X5Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X26Y136_SLICE_X38Y136_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X26Y136_SLICE_X38Y136_DO5),
.O6(CLBLL_L_X26Y136_SLICE_X38Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X26Y136_SLICE_X38Y136_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X26Y136_SLICE_X38Y136_CO5),
.O6(CLBLL_L_X26Y136_SLICE_X38Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X26Y136_SLICE_X38Y136_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X26Y136_SLICE_X38Y136_BO5),
.O6(CLBLL_L_X26Y136_SLICE_X38Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcfffcfffffffcc)
  ) CLBLL_L_X26Y136_SLICE_X38Y136_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y129_IOB_X1Y130_I),
.I2(RIOB33_X105Y137_IOB_X1Y137_I),
.I3(RIOB33_X105Y129_IOB_X1Y129_I),
.I4(RIOB33_X105Y127_IOB_X1Y128_I),
.I5(1'b1),
.O5(CLBLL_L_X26Y136_SLICE_X38Y136_AO5),
.O6(CLBLL_L_X26Y136_SLICE_X38Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X26Y136_SLICE_X39Y136_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X26Y136_SLICE_X39Y136_DO5),
.O6(CLBLL_L_X26Y136_SLICE_X39Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X26Y136_SLICE_X39Y136_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X26Y136_SLICE_X39Y136_CO5),
.O6(CLBLL_L_X26Y136_SLICE_X39Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X26Y136_SLICE_X39Y136_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X26Y136_SLICE_X39Y136_BO5),
.O6(CLBLL_L_X26Y136_SLICE_X39Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X26Y136_SLICE_X39Y136_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X26Y136_SLICE_X39Y136_AO5),
.O6(CLBLL_L_X26Y136_SLICE_X39Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y126_SLICE_X78Y126_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y126_SLICE_X78Y126_DO5),
.O6(CLBLL_L_X52Y126_SLICE_X78Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y126_SLICE_X78Y126_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y126_SLICE_X78Y126_CO5),
.O6(CLBLL_L_X52Y126_SLICE_X78Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y126_SLICE_X78Y126_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y126_SLICE_X78Y126_BO5),
.O6(CLBLL_L_X52Y126_SLICE_X78Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00ff00ff00ff)
  ) CLBLL_L_X52Y126_SLICE_X78Y126_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(RIOB33_X105Y123_IOB_X1Y124_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y126_SLICE_X78Y126_AO5),
.O6(CLBLL_L_X52Y126_SLICE_X78Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y126_SLICE_X79Y126_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y126_SLICE_X79Y126_DO5),
.O6(CLBLL_L_X52Y126_SLICE_X79Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y126_SLICE_X79Y126_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y126_SLICE_X79Y126_CO5),
.O6(CLBLL_L_X52Y126_SLICE_X79Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y126_SLICE_X79Y126_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y126_SLICE_X79Y126_BO5),
.O6(CLBLL_L_X52Y126_SLICE_X79Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y126_SLICE_X79Y126_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y126_SLICE_X79Y126_AO5),
.O6(CLBLL_L_X52Y126_SLICE_X79Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y104_SLICE_X10Y104_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y104_SLICE_X10Y104_DO5),
.O6(CLBLM_L_X8Y104_SLICE_X10Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y104_SLICE_X10Y104_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y104_SLICE_X10Y104_CO5),
.O6(CLBLM_L_X8Y104_SLICE_X10Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y104_SLICE_X10Y104_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y104_SLICE_X10Y104_BO5),
.O6(CLBLM_L_X8Y104_SLICE_X10Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h77ff77ffffffffff)
  ) CLBLM_L_X8Y104_SLICE_X10Y104_ALUT (
.I0(CLBLM_L_X8Y114_SLICE_X11Y114_B5Q),
.I1(CLBLM_L_X10Y104_SLICE_X12Y104_CO6),
.I2(1'b1),
.I3(CLBLM_L_X10Y106_SLICE_X12Y106_BO6),
.I4(1'b1),
.I5(CLBLM_L_X12Y110_SLICE_X16Y110_DO5),
.O5(CLBLM_L_X8Y104_SLICE_X10Y104_AO5),
.O6(CLBLM_L_X8Y104_SLICE_X10Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y104_SLICE_X11Y104_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y104_SLICE_X11Y104_AO6),
.Q(CLBLM_L_X8Y104_SLICE_X11Y104_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y104_SLICE_X11Y104_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y104_SLICE_X11Y104_DO5),
.O6(CLBLM_L_X8Y104_SLICE_X11Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y104_SLICE_X11Y104_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y104_SLICE_X11Y104_CO5),
.O6(CLBLM_L_X8Y104_SLICE_X11Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffaffaaffa)
  ) CLBLM_L_X8Y104_SLICE_X11Y104_BLUT (
.I0(CLBLM_L_X8Y105_SLICE_X11Y105_DO6),
.I1(1'b1),
.I2(CLBLM_R_X5Y105_SLICE_X6Y105_AQ),
.I3(CLBLM_L_X8Y105_SLICE_X11Y105_BQ),
.I4(1'b1),
.I5(CLBLM_L_X8Y105_SLICE_X10Y105_CO6),
.O5(CLBLM_L_X8Y104_SLICE_X11Y104_BO5),
.O6(CLBLM_L_X8Y104_SLICE_X11Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0f0c0000ffcc)
  ) CLBLM_L_X8Y104_SLICE_X11Y104_ALUT (
.I0(CLBLM_L_X10Y110_SLICE_X13Y110_CQ),
.I1(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.I2(CLBLM_L_X8Y105_SLICE_X11Y105_CO6),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y104_SLICE_X11Y104_AO5),
.O6(CLBLM_L_X8Y104_SLICE_X11Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y105_SLICE_X10Y105_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y105_SLICE_X10Y105_AO6),
.Q(CLBLM_L_X8Y105_SLICE_X10Y105_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffeeffeeffeeffee)
  ) CLBLM_L_X8Y105_SLICE_X10Y105_DLUT (
.I0(CLBLM_R_X7Y105_SLICE_X9Y105_BQ),
.I1(CLBLM_L_X8Y105_SLICE_X10Y105_AQ),
.I2(1'b1),
.I3(CLBLM_L_X8Y105_SLICE_X11Y105_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y105_SLICE_X10Y105_DO5),
.O6(CLBLM_L_X8Y105_SLICE_X10Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5faf5faff5faf5fa)
  ) CLBLM_L_X8Y105_SLICE_X10Y105_CLUT (
.I0(CLBLM_R_X7Y105_SLICE_X9Y105_BQ),
.I1(1'b1),
.I2(CLBLM_R_X7Y107_SLICE_X8Y107_BQ),
.I3(CLBLM_L_X8Y106_SLICE_X10Y106_AQ),
.I4(1'b1),
.I5(CLBLM_L_X10Y110_SLICE_X13Y110_BQ),
.O5(CLBLM_L_X8Y105_SLICE_X10Y105_CO5),
.O6(CLBLM_L_X8Y105_SLICE_X10Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3c3cc3c3c3c33c3c)
  ) CLBLM_L_X8Y105_SLICE_X10Y105_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y107_SLICE_X10Y107_AQ),
.I2(CLBLM_R_X7Y107_SLICE_X8Y107_BQ),
.I3(1'b1),
.I4(CLBLM_L_X8Y106_SLICE_X11Y106_AQ),
.I5(CLBLM_R_X5Y105_SLICE_X6Y105_AQ),
.O5(CLBLM_L_X8Y105_SLICE_X10Y105_BO5),
.O6(CLBLM_L_X8Y105_SLICE_X10Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaf333c000)
  ) CLBLM_L_X8Y105_SLICE_X10Y105_ALUT (
.I0(CLBLM_R_X7Y117_SLICE_X9Y117_DQ),
.I1(CLBLM_L_X10Y106_SLICE_X12Y106_BO6),
.I2(CLBLM_L_X8Y105_SLICE_X10Y105_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X7Y105_SLICE_X9Y105_BQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y105_SLICE_X10Y105_AO5),
.O6(CLBLM_L_X8Y105_SLICE_X10Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y105_SLICE_X11Y105_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y105_SLICE_X11Y105_AO6),
.Q(CLBLM_L_X8Y105_SLICE_X11Y105_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y105_SLICE_X11Y105_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y105_SLICE_X11Y105_BO6),
.Q(CLBLM_L_X8Y105_SLICE_X11Y105_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h77dd77ddbbeebbee)
  ) CLBLM_L_X8Y105_SLICE_X11Y105_DLUT (
.I0(CLBLM_L_X8Y106_SLICE_X11Y106_AQ),
.I1(CLBLM_L_X8Y105_SLICE_X11Y105_AQ),
.I2(1'b1),
.I3(CLBLM_L_X8Y107_SLICE_X10Y107_AQ),
.I4(1'b1),
.I5(CLBLM_L_X10Y107_SLICE_X12Y107_AQ),
.O5(CLBLM_L_X8Y105_SLICE_X11Y105_DO5),
.O6(CLBLM_L_X8Y105_SLICE_X11Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0504504050400504)
  ) CLBLM_L_X8Y105_SLICE_X11Y105_CLUT (
.I0(CLBLM_L_X8Y104_SLICE_X11Y104_AQ),
.I1(CLBLM_R_X3Y108_SLICE_X2Y108_DO6),
.I2(CLBLM_R_X11Y106_SLICE_X14Y106_AQ),
.I3(CLBLM_L_X10Y112_SLICE_X12Y112_DO6),
.I4(CLBLM_L_X10Y108_SLICE_X12Y108_BQ),
.I5(CLBLM_L_X8Y106_SLICE_X10Y106_DO6),
.O5(CLBLM_L_X8Y105_SLICE_X11Y105_CO5),
.O6(CLBLM_L_X8Y105_SLICE_X11Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf088f0fff088f000)
  ) CLBLM_L_X8Y105_SLICE_X11Y105_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X8Y105_SLICE_X11Y105_BQ),
.I2(CLBLM_R_X5Y105_SLICE_X6Y105_BQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y106_SLICE_X12Y106_BO6),
.I5(CLBLM_L_X8Y106_SLICE_X11Y106_BQ),
.O5(CLBLM_L_X8Y105_SLICE_X11Y105_BO5),
.O6(CLBLM_L_X8Y105_SLICE_X11Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffa0ffcc00a000cc)
  ) CLBLM_L_X8Y105_SLICE_X11Y105_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X8Y107_SLICE_X10Y107_BQ),
.I2(CLBLM_L_X8Y105_SLICE_X11Y105_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y106_SLICE_X12Y106_BO6),
.I5(CLBLM_L_X12Y107_SLICE_X16Y107_AQ),
.O5(CLBLM_L_X8Y105_SLICE_X11Y105_AO5),
.O6(CLBLM_L_X8Y105_SLICE_X11Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y106_SLICE_X10Y106_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y106_SLICE_X10Y106_AO6),
.Q(CLBLM_L_X8Y106_SLICE_X10Y106_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y106_SLICE_X10Y106_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y106_SLICE_X10Y106_BO6),
.Q(CLBLM_L_X8Y106_SLICE_X10Y106_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y106_SLICE_X10Y106_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y106_SLICE_X10Y106_CO6),
.Q(CLBLM_L_X8Y106_SLICE_X10Y106_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h9696696969699696)
  ) CLBLM_L_X8Y106_SLICE_X10Y106_DLUT (
.I0(CLBLM_L_X8Y105_SLICE_X10Y105_BO6),
.I1(CLBLM_L_X8Y106_SLICE_X10Y106_AQ),
.I2(CLBLM_L_X8Y110_SLICE_X11Y110_DQ),
.I3(1'b1),
.I4(CLBLM_R_X5Y107_SLICE_X7Y107_AQ),
.I5(CLBLM_L_X8Y113_SLICE_X10Y113_BQ),
.O5(CLBLM_L_X8Y106_SLICE_X10Y106_DO5),
.O6(CLBLM_L_X8Y106_SLICE_X10Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0cccc00cc)
  ) CLBLM_L_X8Y106_SLICE_X10Y106_CLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y106_SLICE_X10Y106_CQ),
.I2(CLBLM_R_X5Y107_SLICE_X7Y107_B5Q),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y106_SLICE_X10Y106_CO5),
.O6(CLBLM_L_X8Y106_SLICE_X10Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0000066cc)
  ) CLBLM_L_X8Y106_SLICE_X10Y106_BLUT (
.I0(CLBLM_R_X7Y107_SLICE_X8Y107_DO6),
.I1(CLBLM_L_X8Y106_SLICE_X10Y106_BQ),
.I2(CLBLM_L_X8Y110_SLICE_X11Y110_CQ),
.I3(CLBLM_R_X7Y105_SLICE_X9Y105_CQ),
.I4(CLBLM_L_X10Y113_SLICE_X13Y113_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y106_SLICE_X10Y106_BO5),
.O6(CLBLM_L_X8Y106_SLICE_X10Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffcc00ccfacc50)
  ) CLBLM_L_X8Y106_SLICE_X10Y106_ALUT (
.I0(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.I1(CLBLM_L_X12Y112_SLICE_X16Y112_CQ),
.I2(CLBLM_L_X8Y106_SLICE_X10Y106_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y106_SLICE_X9Y106_BQ),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_L_X8Y106_SLICE_X10Y106_AO5),
.O6(CLBLM_L_X8Y106_SLICE_X10Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y106_SLICE_X11Y106_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y106_SLICE_X11Y106_CO6),
.Q(CLBLM_L_X8Y106_SLICE_X11Y106_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y106_SLICE_X11Y106_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y106_SLICE_X11Y106_AO6),
.Q(CLBLM_L_X8Y106_SLICE_X11Y106_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y106_SLICE_X11Y106_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y106_SLICE_X11Y106_BO6),
.Q(CLBLM_L_X8Y106_SLICE_X11Y106_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5a5affffffff5a5a)
  ) CLBLM_L_X8Y106_SLICE_X11Y106_DLUT (
.I0(CLBLM_L_X8Y110_SLICE_X11Y110_DQ),
.I1(1'b1),
.I2(CLBLM_L_X10Y107_SLICE_X12Y107_BQ),
.I3(1'b1),
.I4(CLBLM_L_X10Y106_SLICE_X13Y106_CQ),
.I5(CLBLM_L_X8Y113_SLICE_X10Y113_BQ),
.O5(CLBLM_L_X8Y106_SLICE_X11Y106_DO5),
.O6(CLBLM_L_X8Y106_SLICE_X11Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccff003355f555f5)
  ) CLBLM_L_X8Y106_SLICE_X11Y106_CLUT (
.I0(CLBLM_R_X7Y106_SLICE_X8Y106_CQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X8Y114_SLICE_X11Y114_B5Q),
.I3(CLBLM_L_X10Y104_SLICE_X12Y104_BO6),
.I4(CLBLM_L_X10Y107_SLICE_X12Y107_BQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y106_SLICE_X11Y106_CO5),
.O6(CLBLM_L_X8Y106_SLICE_X11Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hef45af05ea40aa00)
  ) CLBLM_L_X8Y106_SLICE_X11Y106_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y106_SLICE_X11Y106_BQ),
.I2(CLBLM_L_X10Y106_SLICE_X12Y106_BO6),
.I3(CLBLM_L_X8Y109_SLICE_X11Y109_AQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_L_X10Y106_SLICE_X13Y106_CQ),
.O5(CLBLM_L_X8Y106_SLICE_X11Y106_BO5),
.O6(CLBLM_L_X8Y106_SLICE_X11Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcc3300fedc3210)
  ) CLBLM_L_X8Y106_SLICE_X11Y106_ALUT (
.I0(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X8Y106_SLICE_X11Y106_AQ),
.I3(CLBLM_L_X10Y106_SLICE_X13Y106_AQ),
.I4(CLBLM_L_X8Y109_SLICE_X10Y109_DQ),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_L_X8Y106_SLICE_X11Y106_AO5),
.O6(CLBLM_L_X8Y106_SLICE_X11Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y107_SLICE_X10Y107_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y107_SLICE_X10Y107_AO6),
.Q(CLBLM_L_X8Y107_SLICE_X10Y107_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y107_SLICE_X10Y107_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y107_SLICE_X10Y107_BO6),
.Q(CLBLM_L_X8Y107_SLICE_X10Y107_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y107_SLICE_X10Y107_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y107_SLICE_X10Y107_CO6),
.Q(CLBLM_L_X8Y107_SLICE_X10Y107_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h33333333f3f3f3f3)
  ) CLBLM_L_X8Y107_SLICE_X10Y107_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y107_SLICE_X10Y107_CQ),
.I2(RIOB33_X105Y141_IOB_X1Y142_I),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X8Y119_SLICE_X10Y119_AQ),
.O5(CLBLM_L_X8Y107_SLICE_X10Y107_DO5),
.O6(CLBLM_L_X8Y107_SLICE_X10Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf7f70707f7f50705)
  ) CLBLM_L_X8Y107_SLICE_X10Y107_CLUT (
.I0(CLBLM_L_X8Y107_SLICE_X10Y107_DO6),
.I1(CLBLM_L_X10Y107_SLICE_X12Y107_CO6),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X11Y108_SLICE_X14Y108_BO6),
.I4(CLBLM_L_X12Y106_SLICE_X16Y106_AQ),
.I5(CLBLM_R_X3Y108_SLICE_X2Y108_BO6),
.O5(CLBLM_L_X8Y107_SLICE_X10Y107_CO5),
.O6(CLBLM_L_X8Y107_SLICE_X10Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haacfaac0aa0faa00)
  ) CLBLM_L_X8Y107_SLICE_X10Y107_BLUT (
.I0(CLBLM_L_X10Y111_SLICE_X12Y111_CQ),
.I1(CLBLM_L_X8Y107_SLICE_X10Y107_BQ),
.I2(CLBLM_L_X10Y106_SLICE_X12Y106_BO6),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y110_SLICE_X13Y110_BQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X8Y107_SLICE_X10Y107_BO5),
.O6(CLBLM_L_X8Y107_SLICE_X10Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffcc00ccfacc50)
  ) CLBLM_L_X8Y107_SLICE_X10Y107_ALUT (
.I0(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.I1(CLBLM_L_X10Y109_SLICE_X12Y109_AQ),
.I2(CLBLM_L_X8Y107_SLICE_X10Y107_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y108_SLICE_X10Y108_DQ),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_L_X8Y107_SLICE_X10Y107_AO5),
.O6(CLBLM_L_X8Y107_SLICE_X10Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y107_SLICE_X11Y107_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y107_SLICE_X11Y107_AO5),
.Q(CLBLM_L_X8Y107_SLICE_X11Y107_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y107_SLICE_X11Y107_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y107_SLICE_X11Y107_BO5),
.Q(CLBLM_L_X8Y107_SLICE_X11Y107_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y107_SLICE_X11Y107_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y107_SLICE_X11Y107_AO6),
.Q(CLBLM_L_X8Y107_SLICE_X11Y107_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y107_SLICE_X11Y107_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y107_SLICE_X11Y107_BO6),
.Q(CLBLM_L_X8Y107_SLICE_X11Y107_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y107_SLICE_X11Y107_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y107_SLICE_X11Y107_CO6),
.Q(CLBLM_L_X8Y107_SLICE_X11Y107_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ffffff00fffd)
  ) CLBLM_L_X8Y107_SLICE_X11Y107_DLUT (
.I0(CLBLM_L_X8Y106_SLICE_X11Y106_CO5),
.I1(CLBLM_R_X5Y110_SLICE_X7Y110_DO6),
.I2(CLBLL_L_X4Y107_SLICE_X5Y107_DO6),
.I3(CLBLM_L_X8Y107_SLICE_X11Y107_A5Q),
.I4(CLBLM_L_X10Y107_SLICE_X13Y107_CO6),
.I5(CLBLM_R_X11Y111_SLICE_X14Y111_BO6),
.O5(CLBLM_L_X8Y107_SLICE_X11Y107_DO5),
.O6(CLBLM_L_X8Y107_SLICE_X11Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffaeeea55504440)
  ) CLBLM_L_X8Y107_SLICE_X11Y107_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y107_SLICE_X11Y107_CQ),
.I2(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_L_X10Y107_SLICE_X12Y107_DO6),
.I5(CLBLM_L_X8Y110_SLICE_X10Y110_BQ),
.O5(CLBLM_L_X8Y107_SLICE_X11Y107_CO5),
.O6(CLBLM_L_X8Y107_SLICE_X11Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hddccddcc11aa00aa)
  ) CLBLM_L_X8Y107_SLICE_X11Y107_BLUT (
.I0(CLBLM_L_X8Y107_SLICE_X11Y107_B5Q),
.I1(CLBLM_L_X8Y107_SLICE_X11Y107_BQ),
.I2(1'b1),
.I3(CLBLM_L_X8Y107_SLICE_X11Y107_DO6),
.I4(CLBLM_L_X8Y107_SLICE_X11Y107_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X8Y107_SLICE_X11Y107_BO5),
.O6(CLBLM_L_X8Y107_SLICE_X11Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h22f000f011ff5500)
  ) CLBLM_L_X8Y107_SLICE_X11Y107_ALUT (
.I0(CLBLM_L_X8Y107_SLICE_X11Y107_B5Q),
.I1(CLBLM_L_X8Y107_SLICE_X11Y107_BQ),
.I2(CLBLM_L_X8Y107_SLICE_X11Y107_AQ),
.I3(CLBLM_L_X8Y107_SLICE_X11Y107_DO6),
.I4(CLBLM_L_X8Y107_SLICE_X11Y107_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X8Y107_SLICE_X11Y107_AO5),
.O6(CLBLM_L_X8Y107_SLICE_X11Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y108_SLICE_X10Y108_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y108_SLICE_X10Y108_AO6),
.Q(CLBLM_L_X8Y108_SLICE_X10Y108_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y108_SLICE_X10Y108_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y108_SLICE_X10Y108_BO6),
.Q(CLBLM_L_X8Y108_SLICE_X10Y108_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y108_SLICE_X10Y108_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y108_SLICE_X10Y108_CO6),
.Q(CLBLM_L_X8Y108_SLICE_X10Y108_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y108_SLICE_X10Y108_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y108_SLICE_X10Y108_DO6),
.Q(CLBLM_L_X8Y108_SLICE_X10Y108_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff00a8000000a8)
  ) CLBLM_L_X8Y108_SLICE_X10Y108_DLUT (
.I0(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.I1(CLBLM_L_X8Y108_SLICE_X10Y108_CQ),
.I2(CLBLM_L_X8Y108_SLICE_X10Y108_DQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLL_L_X4Y110_SLICE_X4Y110_BQ),
.O5(CLBLM_L_X8Y108_SLICE_X10Y108_DO5),
.O6(CLBLM_L_X8Y108_SLICE_X10Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa0000f0ff)
  ) CLBLM_L_X8Y108_SLICE_X10Y108_CLUT (
.I0(CLBLM_R_X5Y115_SLICE_X6Y115_AQ),
.I1(1'b1),
.I2(CLBLM_L_X8Y119_SLICE_X10Y119_AQ),
.I3(RIOB33_X105Y141_IOB_X1Y142_I),
.I4(CLBLM_L_X10Y108_SLICE_X12Y108_DO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y108_SLICE_X10Y108_CO5),
.O6(CLBLM_L_X8Y108_SLICE_X10Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000505ff005050)
  ) CLBLM_L_X8Y108_SLICE_X10Y108_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(1'b1),
.I2(CLBLM_R_X11Y110_SLICE_X15Y110_BQ),
.I3(CLBLM_L_X8Y106_SLICE_X10Y106_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y108_SLICE_X10Y108_AO5),
.O5(CLBLM_L_X8Y108_SLICE_X10Y108_BO5),
.O6(CLBLM_L_X8Y108_SLICE_X10Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0aa88aa88aa88)
  ) CLBLM_L_X8Y108_SLICE_X10Y108_ALUT (
.I0(RIOB33_X105Y121_IOB_X1Y121_I),
.I1(CLBLM_L_X8Y107_SLICE_X11Y107_CQ),
.I2(CLBLL_L_X4Y114_SLICE_X4Y114_AQ),
.I3(CLBLM_L_X10Y112_SLICE_X12Y112_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y108_SLICE_X10Y108_AO5),
.O6(CLBLM_L_X8Y108_SLICE_X10Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y108_SLICE_X11Y108_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y108_SLICE_X11Y108_AO6),
.Q(CLBLM_L_X8Y108_SLICE_X11Y108_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y108_SLICE_X11Y108_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y108_SLICE_X11Y108_BO6),
.Q(CLBLM_L_X8Y108_SLICE_X11Y108_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000110011)
  ) CLBLM_L_X8Y108_SLICE_X11Y108_DLUT (
.I0(CLBLL_L_X4Y107_SLICE_X4Y107_CQ),
.I1(CLBLM_L_X8Y106_SLICE_X10Y106_CQ),
.I2(1'b1),
.I3(CLBLM_L_X8Y108_SLICE_X11Y108_AQ),
.I4(1'b1),
.I5(CLBLM_L_X10Y113_SLICE_X13Y113_BQ),
.O5(CLBLM_L_X8Y108_SLICE_X11Y108_DO5),
.O6(CLBLM_L_X8Y108_SLICE_X11Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f05050f0c0)
  ) CLBLM_L_X8Y108_SLICE_X11Y108_CLUT (
.I0(CLBLM_L_X8Y108_SLICE_X11Y108_BQ),
.I1(CLBLM_L_X10Y112_SLICE_X12Y112_DO6),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLM_R_X3Y110_SLICE_X3Y110_DO6),
.I4(CLBLM_L_X8Y108_SLICE_X11Y108_DO6),
.I5(CLBLM_R_X13Y112_SLICE_X18Y112_BQ),
.O5(CLBLM_L_X8Y108_SLICE_X11Y108_CO5),
.O6(CLBLM_L_X8Y108_SLICE_X11Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfe0ef404ff0ff000)
  ) CLBLM_L_X8Y108_SLICE_X11Y108_BLUT (
.I0(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.I1(CLBLM_R_X7Y108_SLICE_X9Y108_CO6),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X11Y110_SLICE_X15Y110_CQ),
.I4(CLBLM_L_X8Y108_SLICE_X11Y108_BQ),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_L_X8Y108_SLICE_X11Y108_BO5),
.O6(CLBLM_L_X8Y108_SLICE_X11Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcca0cca0ccaaccaa)
  ) CLBLM_L_X8Y108_SLICE_X11Y108_ALUT (
.I0(CLBLM_L_X8Y108_SLICE_X11Y108_AQ),
.I1(CLBLM_L_X8Y108_SLICE_X11Y108_BQ),
.I2(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_L_X8Y108_SLICE_X11Y108_AO5),
.O6(CLBLM_L_X8Y108_SLICE_X11Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y109_SLICE_X10Y109_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y109_SLICE_X10Y109_CO5),
.Q(CLBLM_L_X8Y109_SLICE_X10Y109_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y109_SLICE_X10Y109_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y109_SLICE_X10Y109_AO6),
.Q(CLBLM_L_X8Y109_SLICE_X10Y109_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y109_SLICE_X10Y109_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y109_SLICE_X10Y109_BO6),
.Q(CLBLM_L_X8Y109_SLICE_X10Y109_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y109_SLICE_X10Y109_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y109_SLICE_X10Y109_CO6),
.Q(CLBLM_L_X8Y109_SLICE_X10Y109_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y109_SLICE_X10Y109_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y109_SLICE_X10Y109_DO6),
.Q(CLBLM_L_X8Y109_SLICE_X10Y109_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hdddddd88d8d8d888)
  ) CLBLM_L_X8Y109_SLICE_X10Y109_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y106_SLICE_X6Y106_DQ),
.I2(CLBLM_L_X8Y109_SLICE_X10Y109_DQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.I5(CLBLM_R_X7Y109_SLICE_X8Y109_DO6),
.O5(CLBLM_L_X8Y109_SLICE_X10Y109_DO5),
.O6(CLBLM_L_X8Y109_SLICE_X10Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hdddd8888e4e4e4e4)
  ) CLBLM_L_X8Y109_SLICE_X10Y109_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y109_SLICE_X11Y109_A5Q),
.I2(CLBLM_R_X7Y109_SLICE_X9Y109_AQ),
.I3(1'b1),
.I4(CLBLM_R_X5Y109_SLICE_X6Y109_CQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y109_SLICE_X10Y109_CO5),
.O6(CLBLM_L_X8Y109_SLICE_X10Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0c000cff0c000c)
  ) CLBLM_L_X8Y109_SLICE_X10Y109_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y109_SLICE_X10Y109_BQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y109_SLICE_X10Y109_C5Q),
.I5(1'b1),
.O5(CLBLM_L_X8Y109_SLICE_X10Y109_BO5),
.O6(CLBLM_L_X8Y109_SLICE_X10Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccaaccf0ccaaccf0)
  ) CLBLM_L_X8Y109_SLICE_X10Y109_ALUT (
.I0(CLBLM_L_X10Y108_SLICE_X12Y108_CQ),
.I1(CLBLM_R_X11Y111_SLICE_X15Y111_C5Q),
.I2(CLBLM_L_X8Y109_SLICE_X10Y109_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLL_L_X4Y112_SLICE_X4Y112_CO5),
.I5(1'b1),
.O5(CLBLM_L_X8Y109_SLICE_X10Y109_AO5),
.O6(CLBLM_L_X8Y109_SLICE_X10Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y109_SLICE_X11Y109_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y111_SLICE_X10Y111_BO6),
.Q(CLBLM_L_X8Y109_SLICE_X11Y109_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y109_SLICE_X11Y109_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y109_SLICE_X11Y109_AO6),
.Q(CLBLM_L_X8Y109_SLICE_X11Y109_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y109_SLICE_X11Y109_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y109_SLICE_X11Y109_BO6),
.Q(CLBLM_L_X8Y109_SLICE_X11Y109_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y109_SLICE_X11Y109_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y109_SLICE_X11Y109_CO6),
.Q(CLBLM_L_X8Y109_SLICE_X11Y109_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h201f201f201f201f)
  ) CLBLM_L_X8Y109_SLICE_X11Y109_DLUT (
.I0(CLBLM_R_X5Y117_SLICE_X7Y117_AQ),
.I1(CLBLM_R_X11Y112_SLICE_X14Y112_BQ),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLM_L_X8Y107_SLICE_X11Y107_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y109_SLICE_X11Y109_DO5),
.O6(CLBLM_L_X8Y109_SLICE_X11Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0f5a0e4a0f5a0e4)
  ) CLBLM_L_X8Y109_SLICE_X11Y109_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y109_SLICE_X11Y109_CQ),
.I2(CLBLM_R_X7Y106_SLICE_X9Y106_CQ),
.I3(CLBLM_R_X5Y115_SLICE_X7Y115_CO6),
.I4(CLBLM_L_X12Y110_SLICE_X17Y110_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y109_SLICE_X11Y109_CO5),
.O6(CLBLM_L_X8Y109_SLICE_X11Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcfc5c5c0cfc5c5)
  ) CLBLM_L_X8Y109_SLICE_X11Y109_BLUT (
.I0(CLBLM_L_X8Y106_SLICE_X11Y106_A5Q),
.I1(CLBLM_R_X13Y117_SLICE_X18Y117_AQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X5Y109_SLICE_X6Y109_CQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_L_X8Y109_SLICE_X10Y109_CQ),
.O5(CLBLM_L_X8Y109_SLICE_X11Y109_BO5),
.O6(CLBLM_L_X8Y109_SLICE_X11Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heca0eeaaeeaaeca0)
  ) CLBLM_L_X8Y109_SLICE_X11Y109_ALUT (
.I0(CLBLM_L_X8Y104_SLICE_X11Y104_AO5),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X8Y109_SLICE_X11Y109_AQ),
.I3(CLBLM_L_X8Y108_SLICE_X10Y108_BQ),
.I4(CLBLM_L_X8Y111_SLICE_X10Y111_CO6),
.I5(CLBLM_L_X8Y108_SLICE_X11Y108_CO6),
.O5(CLBLM_L_X8Y109_SLICE_X11Y109_AO5),
.O6(CLBLM_L_X8Y109_SLICE_X11Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y110_SLICE_X10Y110_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y110_SLICE_X10Y110_AO6),
.Q(CLBLM_L_X8Y110_SLICE_X10Y110_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y110_SLICE_X10Y110_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y110_SLICE_X10Y110_BO6),
.Q(CLBLM_L_X8Y110_SLICE_X10Y110_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaaffaacc88cc88)
  ) CLBLM_L_X8Y110_SLICE_X10Y110_DLUT (
.I0(CLBLM_L_X10Y104_SLICE_X12Y104_AQ),
.I1(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.I2(1'b1),
.I3(CLBLM_R_X7Y116_SLICE_X8Y116_CQ),
.I4(1'b1),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_L_X8Y110_SLICE_X10Y110_DO5),
.O6(CLBLM_L_X8Y110_SLICE_X10Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000fcfc0000ffaa)
  ) CLBLM_L_X8Y110_SLICE_X10Y110_CLUT (
.I0(CLBLM_R_X7Y110_SLICE_X9Y110_BQ),
.I1(CLBLM_R_X7Y105_SLICE_X9Y105_AQ),
.I2(CLBLM_L_X8Y110_SLICE_X10Y110_AQ),
.I3(CLBLM_R_X7Y105_SLICE_X8Y105_A5Q),
.I4(CLBLM_L_X10Y113_SLICE_X13Y113_CQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y110_SLICE_X10Y110_CO5),
.O6(CLBLM_L_X8Y110_SLICE_X10Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa00003c3c)
  ) CLBLM_L_X8Y110_SLICE_X10Y110_BLUT (
.I0(CLBLM_L_X12Y111_SLICE_X16Y111_BQ),
.I1(CLBLM_L_X8Y110_SLICE_X10Y110_BQ),
.I2(CLBLM_R_X7Y108_SLICE_X9Y108_BO6),
.I3(1'b1),
.I4(CLBLM_L_X10Y113_SLICE_X13Y113_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y110_SLICE_X10Y110_BO5),
.O6(CLBLM_L_X8Y110_SLICE_X10Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff3333fcec3020)
  ) CLBLM_L_X8Y110_SLICE_X10Y110_ALUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X8Y110_SLICE_X10Y110_AQ),
.I3(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.I4(CLBLM_R_X11Y105_SLICE_X14Y105_DQ),
.I5(CLBLM_R_X7Y110_SLICE_X9Y110_DO6),
.O5(CLBLM_L_X8Y110_SLICE_X10Y110_AO5),
.O6(CLBLM_L_X8Y110_SLICE_X10Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y110_SLICE_X11Y110_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y110_SLICE_X11Y110_BO6),
.Q(CLBLM_L_X8Y110_SLICE_X11Y110_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y110_SLICE_X11Y110_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y110_SLICE_X11Y110_AO6),
.Q(CLBLM_L_X8Y110_SLICE_X11Y110_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y110_SLICE_X11Y110_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y110_SLICE_X11Y110_CO6),
.Q(CLBLM_L_X8Y110_SLICE_X11Y110_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y110_SLICE_X11Y110_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y110_SLICE_X11Y110_DO6),
.Q(CLBLM_L_X8Y110_SLICE_X11Y110_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccaaaaaaf0)
  ) CLBLM_L_X8Y110_SLICE_X11Y110_DLUT (
.I0(CLBLM_R_X11Y113_SLICE_X14Y113_AQ),
.I1(CLBLM_L_X12Y108_SLICE_X17Y108_AQ),
.I2(CLBLM_L_X8Y110_SLICE_X11Y110_DQ),
.I3(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y110_SLICE_X11Y110_DO5),
.O6(CLBLM_L_X8Y110_SLICE_X11Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000555c555c)
  ) CLBLM_L_X8Y110_SLICE_X11Y110_CLUT (
.I0(CLBLM_L_X8Y112_SLICE_X11Y112_AO6),
.I1(CLBLM_L_X8Y110_SLICE_X11Y110_CQ),
.I2(RIOB33_X105Y117_IOB_X1Y118_I),
.I3(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.I4(CLBLM_L_X8Y110_SLICE_X10Y110_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y110_SLICE_X11Y110_CO5),
.O6(CLBLM_L_X8Y110_SLICE_X11Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0ccf000ffbbffbb)
  ) CLBLM_L_X8Y110_SLICE_X11Y110_BLUT (
.I0(CLBLM_L_X12Y113_SLICE_X17Y113_BQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_L_X8Y107_SLICE_X11Y107_CQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y110_SLICE_X11Y110_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X8Y110_SLICE_X11Y110_BO5),
.O6(CLBLM_L_X8Y110_SLICE_X11Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfd31fd31ec20ec20)
  ) CLBLM_L_X8Y110_SLICE_X11Y110_ALUT (
.I0(CLBLL_L_X4Y116_SLICE_X4Y116_BO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X8Y110_SLICE_X11Y110_AQ),
.I3(CLBLM_L_X8Y106_SLICE_X11Y106_BQ),
.I4(1'b1),
.I5(CLBLM_L_X8Y115_SLICE_X10Y115_CQ),
.O5(CLBLM_L_X8Y110_SLICE_X11Y110_AO5),
.O6(CLBLM_L_X8Y110_SLICE_X11Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y111_SLICE_X10Y111_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y111_SLICE_X10Y111_AO5),
.Q(CLBLM_L_X8Y111_SLICE_X10Y111_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y111_SLICE_X10Y111_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y111_SLICE_X10Y111_AO6),
.Q(CLBLM_L_X8Y111_SLICE_X10Y111_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffef0000ff001010)
  ) CLBLM_L_X8Y111_SLICE_X10Y111_DLUT (
.I0(CLBLM_L_X8Y111_SLICE_X11Y111_DO5),
.I1(CLBLM_L_X8Y114_SLICE_X10Y114_CQ),
.I2(CLBLM_L_X10Y112_SLICE_X12Y112_BQ),
.I3(CLBLM_R_X11Y111_SLICE_X15Y111_BQ),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(CLBLM_R_X7Y112_SLICE_X8Y112_BQ),
.O5(CLBLM_L_X8Y111_SLICE_X10Y111_DO5),
.O6(CLBLM_L_X8Y111_SLICE_X10Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h1ed2ee22e12d11dd)
  ) CLBLM_L_X8Y111_SLICE_X10Y111_CLUT (
.I0(CLBLM_L_X8Y112_SLICE_X10Y112_DO6),
.I1(CLBLM_L_X8Y111_SLICE_X10Y111_AQ),
.I2(CLBLM_L_X8Y111_SLICE_X11Y111_DO6),
.I3(CLBLM_L_X12Y106_SLICE_X17Y106_AQ),
.I4(CLBLM_L_X8Y112_SLICE_X11Y112_AO5),
.I5(CLBLM_R_X7Y105_SLICE_X8Y105_CQ),
.O5(CLBLM_L_X8Y111_SLICE_X10Y111_CO5),
.O6(CLBLM_L_X8Y111_SLICE_X10Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'he2e2e2c0aaaaaa00)
  ) CLBLM_L_X8Y111_SLICE_X10Y111_BLUT (
.I0(RIOB33_X105Y121_IOB_X1Y121_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X8Y106_SLICE_X10Y106_AQ),
.I3(CLBLM_R_X7Y111_SLICE_X9Y111_AQ),
.I4(CLBLM_R_X5Y109_SLICE_X6Y109_DQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y111_SLICE_X10Y111_BO5),
.O6(CLBLM_L_X8Y111_SLICE_X10Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa30aa30f0fff000)
  ) CLBLM_L_X8Y111_SLICE_X10Y111_ALUT (
.I0(CLBLM_L_X12Y110_SLICE_X17Y110_CQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_L_X8Y111_SLICE_X10Y111_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X3Y111_SLICE_X2Y111_CO6),
.I5(1'b1),
.O5(CLBLM_L_X8Y111_SLICE_X10Y111_AO5),
.O6(CLBLM_L_X8Y111_SLICE_X10Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y111_SLICE_X11Y111_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y111_SLICE_X11Y111_AO6),
.Q(CLBLM_L_X8Y111_SLICE_X11Y111_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y111_SLICE_X11Y111_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y111_SLICE_X11Y111_BO6),
.Q(CLBLM_L_X8Y111_SLICE_X11Y111_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y111_SLICE_X11Y111_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y111_SLICE_X11Y111_CO6),
.Q(CLBLM_L_X8Y111_SLICE_X11Y111_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h11111111bbbbbbbb)
  ) CLBLM_L_X8Y111_SLICE_X11Y111_DLUT (
.I0(CLBLM_R_X7Y111_SLICE_X8Y111_CQ),
.I1(CLBLM_R_X7Y117_SLICE_X9Y117_DQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y111_SLICE_X11Y111_DO5),
.O6(CLBLM_L_X8Y111_SLICE_X11Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f055550000)
  ) CLBLM_L_X8Y111_SLICE_X11Y111_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(1'b1),
.I2(CLBLM_R_X5Y110_SLICE_X7Y110_B5Q),
.I3(1'b1),
.I4(CLBLM_R_X13Y112_SLICE_X18Y112_BQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y111_SLICE_X11Y111_CO5),
.O6(CLBLM_L_X8Y111_SLICE_X11Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0ffccaa88)
  ) CLBLM_L_X8Y111_SLICE_X11Y111_BLUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_L_X8Y111_SLICE_X11Y111_BQ),
.I2(CLBLM_R_X11Y106_SLICE_X15Y106_AQ),
.I3(CLBLM_L_X8Y112_SLICE_X11Y112_DO6),
.I4(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y111_SLICE_X11Y111_BO5),
.O6(CLBLM_L_X8Y111_SLICE_X11Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccff00f000)
  ) CLBLM_L_X8Y111_SLICE_X11Y111_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y111_SLICE_X8Y111_CQ),
.I2(CLBLM_L_X8Y111_SLICE_X11Y111_AQ),
.I3(CLBLL_L_X4Y116_SLICE_X4Y116_BO6),
.I4(CLBLM_L_X12Y110_SLICE_X17Y110_CQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y111_SLICE_X11Y111_AO5),
.O6(CLBLM_L_X8Y111_SLICE_X11Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y112_SLICE_X10Y112_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y112_SLICE_X10Y112_AO5),
.Q(CLBLM_L_X8Y112_SLICE_X10Y112_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y112_SLICE_X10Y112_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y112_SLICE_X10Y112_AO6),
.Q(CLBLM_L_X8Y112_SLICE_X10Y112_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555555555555554)
  ) CLBLM_L_X8Y112_SLICE_X10Y112_DLUT (
.I0(CLBLM_L_X12Y106_SLICE_X17Y106_AQ),
.I1(CLBLM_L_X10Y110_SLICE_X12Y110_DO6),
.I2(CLBLM_R_X7Y113_SLICE_X8Y113_DQ),
.I3(CLBLM_L_X8Y112_SLICE_X11Y112_BO6),
.I4(CLBLM_L_X8Y118_SLICE_X10Y118_BQ),
.I5(CLBLM_R_X7Y115_SLICE_X8Y115_BQ),
.O5(CLBLM_L_X8Y112_SLICE_X10Y112_DO5),
.O6(CLBLM_L_X8Y112_SLICE_X10Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hbfff1555eaaa4000)
  ) CLBLM_L_X8Y112_SLICE_X10Y112_CLUT (
.I0(RIOB33_X105Y121_IOB_X1Y121_I),
.I1(CLBLM_L_X8Y114_SLICE_X10Y114_CQ),
.I2(CLBLM_L_X8Y111_SLICE_X11Y111_DO6),
.I3(CLBLM_L_X10Y112_SLICE_X12Y112_BQ),
.I4(CLBLM_R_X7Y115_SLICE_X8Y115_CQ),
.I5(CLBLM_R_X7Y115_SLICE_X8Y115_BQ),
.O5(CLBLM_L_X8Y112_SLICE_X10Y112_CO5),
.O6(CLBLM_L_X8Y112_SLICE_X10Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h1f1f1f5c1f1f1f1f)
  ) CLBLM_L_X8Y112_SLICE_X10Y112_BLUT (
.I0(CLBLM_R_X11Y112_SLICE_X14Y112_CQ),
.I1(CLBLM_R_X7Y113_SLICE_X8Y113_DQ),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLM_L_X10Y112_SLICE_X12Y112_BQ),
.I4(CLBLM_L_X8Y111_SLICE_X11Y111_DO5),
.I5(CLBLM_L_X8Y114_SLICE_X10Y114_CQ),
.O5(CLBLM_L_X8Y112_SLICE_X10Y112_BO5),
.O6(CLBLM_L_X8Y112_SLICE_X10Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'he2e2e2e2fccc3000)
  ) CLBLM_L_X8Y112_SLICE_X10Y112_ALUT (
.I0(CLBLM_L_X8Y115_SLICE_X10Y115_A5Q),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X7Y112_SLICE_X9Y112_BQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_L_X8Y105_SLICE_X10Y105_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y112_SLICE_X10Y112_AO5),
.O6(CLBLM_L_X8Y112_SLICE_X10Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbff0b0ff4f00400)
  ) CLBLM_L_X8Y112_SLICE_X11Y112_DLUT (
.I0(CLBLM_R_X7Y117_SLICE_X9Y117_DQ),
.I1(CLBLM_R_X7Y111_SLICE_X8Y111_CQ),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLM_L_X8Y112_SLICE_X11Y112_AO5),
.I4(CLBLM_L_X10Y112_SLICE_X12Y112_CQ),
.I5(CLBLM_L_X8Y115_SLICE_X10Y115_BQ),
.O5(CLBLM_L_X8Y112_SLICE_X11Y112_DO5),
.O6(CLBLM_L_X8Y112_SLICE_X11Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafa0000bafa0c00)
  ) CLBLM_L_X8Y112_SLICE_X11Y112_CLUT (
.I0(CLBLM_R_X5Y109_SLICE_X6Y109_DQ),
.I1(CLBLM_L_X10Y112_SLICE_X12Y112_BQ),
.I2(CLBLM_L_X8Y118_SLICE_X10Y118_BQ),
.I3(CLBLM_L_X8Y114_SLICE_X10Y114_CQ),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(CLBLM_L_X8Y111_SLICE_X11Y111_DO5),
.O5(CLBLM_L_X8Y112_SLICE_X11Y112_CO5),
.O6(CLBLM_L_X8Y112_SLICE_X11Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_L_X8Y112_SLICE_X11Y112_BLUT (
.I0(CLBLM_R_X7Y112_SLICE_X8Y112_BQ),
.I1(CLBLM_L_X8Y114_SLICE_X11Y114_BQ),
.I2(CLBLM_L_X12Y113_SLICE_X17Y113_B5Q),
.I3(CLBLM_L_X8Y115_SLICE_X10Y115_BQ),
.I4(CLBLM_L_X10Y111_SLICE_X12Y111_BQ),
.I5(CLBLM_L_X8Y109_SLICE_X10Y109_BQ),
.O5(CLBLM_L_X8Y112_SLICE_X11Y112_BO5),
.O6(CLBLM_L_X8Y112_SLICE_X11Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3336333355005500)
  ) CLBLM_L_X8Y112_SLICE_X11Y112_ALUT (
.I0(CLBLM_L_X8Y114_SLICE_X10Y114_CQ),
.I1(CLBLM_L_X8Y114_SLICE_X11Y114_BQ),
.I2(CLBLM_R_X7Y111_SLICE_X8Y111_CQ),
.I3(CLBLM_L_X10Y112_SLICE_X12Y112_BQ),
.I4(CLBLM_R_X7Y117_SLICE_X9Y117_DQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y112_SLICE_X11Y112_AO5),
.O6(CLBLM_L_X8Y112_SLICE_X11Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y113_SLICE_X10Y113_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y113_SLICE_X10Y113_DO5),
.Q(CLBLM_L_X8Y113_SLICE_X10Y113_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y113_SLICE_X10Y113_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y113_SLICE_X10Y113_AO6),
.Q(CLBLM_L_X8Y113_SLICE_X10Y113_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y113_SLICE_X10Y113_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y113_SLICE_X10Y113_BO6),
.Q(CLBLM_L_X8Y113_SLICE_X10Y113_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y113_SLICE_X10Y113_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y113_SLICE_X10Y113_CO6),
.Q(CLBLM_L_X8Y113_SLICE_X10Y113_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y113_SLICE_X10Y113_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y113_SLICE_X10Y113_DO6),
.Q(CLBLM_L_X8Y113_SLICE_X10Y113_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcf03cf038888b8b8)
  ) CLBLM_L_X8Y113_SLICE_X10Y113_DLUT (
.I0(CLBLM_L_X10Y111_SLICE_X13Y111_C5Q),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(RIOB33_X105Y119_IOB_X1Y119_I),
.I3(CLBLM_R_X5Y111_SLICE_X6Y111_CQ),
.I4(CLBLM_L_X8Y113_SLICE_X10Y113_D5Q),
.I5(1'b1),
.O5(CLBLM_L_X8Y113_SLICE_X10Y113_DO5),
.O6(CLBLM_L_X8Y113_SLICE_X10Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa000f0f00)
  ) CLBLM_L_X8Y113_SLICE_X10Y113_CLUT (
.I0(CLBLM_R_X11Y114_SLICE_X14Y114_AQ),
.I1(1'b1),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_L_X8Y112_SLICE_X11Y112_CO6),
.I4(CLBLM_R_X5Y113_SLICE_X6Y113_BQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y113_SLICE_X10Y113_CO5),
.O6(CLBLM_L_X8Y113_SLICE_X10Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00aaaaacac)
  ) CLBLM_L_X8Y113_SLICE_X10Y113_BLUT (
.I0(CLBLM_L_X10Y113_SLICE_X12Y113_CQ),
.I1(CLBLM_L_X8Y113_SLICE_X10Y113_BQ),
.I2(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.I3(CLBLM_R_X7Y114_SLICE_X9Y114_BQ),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y113_SLICE_X10Y113_BO5),
.O6(CLBLM_L_X8Y113_SLICE_X10Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00d8d8ff00d8d8)
  ) CLBLM_L_X8Y113_SLICE_X10Y113_ALUT (
.I0(CLBLL_L_X4Y112_SLICE_X4Y112_CO5),
.I1(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I2(CLBLM_L_X8Y113_SLICE_X10Y113_AQ),
.I3(CLBLM_L_X10Y106_SLICE_X13Y106_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y113_SLICE_X10Y113_AO5),
.O6(CLBLM_L_X8Y113_SLICE_X10Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y113_SLICE_X11Y113_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y113_SLICE_X11Y113_AO6),
.Q(CLBLM_L_X8Y113_SLICE_X11Y113_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y113_SLICE_X11Y113_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y113_SLICE_X11Y113_BO6),
.Q(CLBLM_L_X8Y113_SLICE_X11Y113_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6699669999669966)
  ) CLBLM_L_X8Y113_SLICE_X11Y113_DLUT (
.I0(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I1(CLBLM_L_X12Y108_SLICE_X16Y108_AQ),
.I2(1'b1),
.I3(CLBLM_L_X8Y113_SLICE_X11Y113_AQ),
.I4(1'b1),
.I5(CLBLM_R_X7Y115_SLICE_X9Y115_A5Q),
.O5(CLBLM_L_X8Y113_SLICE_X11Y113_DO5),
.O6(CLBLM_L_X8Y113_SLICE_X11Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hc8c8c8c88cc8c8c8)
  ) CLBLM_L_X8Y113_SLICE_X11Y113_CLUT (
.I0(CLBLM_R_X13Y112_SLICE_X18Y112_CQ),
.I1(RIOB33_X105Y121_IOB_X1Y121_I),
.I2(CLBLM_L_X12Y113_SLICE_X17Y113_B5Q),
.I3(CLBLM_L_X8Y114_SLICE_X10Y114_CQ),
.I4(CLBLM_L_X8Y111_SLICE_X11Y111_DO6),
.I5(CLBLM_L_X10Y112_SLICE_X12Y112_BQ),
.O5(CLBLM_L_X8Y113_SLICE_X11Y113_CO5),
.O6(CLBLM_L_X8Y113_SLICE_X11Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55fa50ee44ea40)
  ) CLBLM_L_X8Y113_SLICE_X11Y113_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y113_SLICE_X11Y113_BQ),
.I2(RIOB33_X105Y117_IOB_X1Y118_I),
.I3(CLBLM_L_X8Y113_SLICE_X10Y113_BQ),
.I4(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.I5(CLBLM_L_X8Y113_SLICE_X11Y113_CO6),
.O5(CLBLM_L_X8Y113_SLICE_X11Y113_BO5),
.O6(CLBLM_L_X8Y113_SLICE_X11Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf505f000fa0af000)
  ) CLBLM_L_X8Y113_SLICE_X11Y113_ALUT (
.I0(CLBLM_L_X8Y113_SLICE_X11Y113_DO6),
.I1(1'b1),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y114_SLICE_X10Y114_DQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_L_X8Y108_SLICE_X11Y108_CO6),
.O5(CLBLM_L_X8Y113_SLICE_X11Y113_AO5),
.O6(CLBLM_L_X8Y113_SLICE_X11Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y114_SLICE_X10Y114_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y114_SLICE_X10Y114_AO6),
.Q(CLBLM_L_X8Y114_SLICE_X10Y114_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y114_SLICE_X10Y114_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y114_SLICE_X10Y114_BO6),
.Q(CLBLM_L_X8Y114_SLICE_X10Y114_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y114_SLICE_X10Y114_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y114_SLICE_X10Y114_CO6),
.Q(CLBLM_L_X8Y114_SLICE_X10Y114_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y114_SLICE_X10Y114_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y114_SLICE_X10Y114_DO6),
.Q(CLBLM_L_X8Y114_SLICE_X10Y114_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00aaf0aaf0)
  ) CLBLM_L_X8Y114_SLICE_X10Y114_DLUT (
.I0(CLBLM_R_X7Y118_SLICE_X8Y118_BQ),
.I1(1'b1),
.I2(CLBLM_L_X10Y112_SLICE_X12Y112_CQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X8Y114_SLICE_X10Y114_DO5),
.O6(CLBLM_L_X8Y114_SLICE_X10Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaeeaaaa00440000)
  ) CLBLM_L_X8Y114_SLICE_X10Y114_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y114_SLICE_X10Y114_CQ),
.I2(1'b1),
.I3(CLBLM_R_X7Y112_SLICE_X8Y112_CQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_L_X8Y115_SLICE_X10Y115_BQ),
.O5(CLBLM_L_X8Y114_SLICE_X10Y114_CO5),
.O6(CLBLM_L_X8Y114_SLICE_X10Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000ff0ffc0c)
  ) CLBLM_L_X8Y114_SLICE_X10Y114_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y114_SLICE_X10Y114_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y113_SLICE_X9Y113_A5Q),
.I4(CLBLM_L_X12Y113_SLICE_X16Y113_BQ),
.I5(CLBLM_R_X5Y115_SLICE_X7Y115_CO6),
.O5(CLBLM_L_X8Y114_SLICE_X10Y114_BO5),
.O6(CLBLM_L_X8Y114_SLICE_X10Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaccccf0f0)
  ) CLBLM_L_X8Y114_SLICE_X10Y114_ALUT (
.I0(CLBLM_R_X11Y113_SLICE_X15Y113_DQ),
.I1(CLBLM_R_X5Y113_SLICE_X6Y113_BQ),
.I2(CLBLM_L_X8Y114_SLICE_X10Y114_AQ),
.I3(1'b1),
.I4(CLBLL_L_X4Y112_SLICE_X4Y112_CO5),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y114_SLICE_X10Y114_AO5),
.O6(CLBLM_L_X8Y114_SLICE_X10Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y114_SLICE_X11Y114_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y114_SLICE_X11Y114_BO5),
.Q(CLBLM_L_X8Y114_SLICE_X11Y114_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y114_SLICE_X11Y114_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y114_SLICE_X11Y114_AO6),
.Q(CLBLM_L_X8Y114_SLICE_X11Y114_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y114_SLICE_X11Y114_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y114_SLICE_X11Y114_BO6),
.Q(CLBLM_L_X8Y114_SLICE_X11Y114_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y114_SLICE_X11Y114_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y114_SLICE_X11Y114_CO6),
.Q(CLBLM_L_X8Y114_SLICE_X11Y114_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000555500005595)
  ) CLBLM_L_X8Y114_SLICE_X11Y114_DLUT (
.I0(CLBLM_L_X10Y111_SLICE_X12Y111_BQ),
.I1(CLBLM_R_X7Y111_SLICE_X8Y111_CQ),
.I2(CLBLM_R_X7Y117_SLICE_X9Y117_DQ),
.I3(CLBLM_L_X8Y114_SLICE_X10Y114_CQ),
.I4(CLBLM_R_X5Y117_SLICE_X7Y117_AQ),
.I5(CLBLM_L_X10Y112_SLICE_X12Y112_BQ),
.O5(CLBLM_L_X8Y114_SLICE_X11Y114_DO5),
.O6(CLBLM_L_X8Y114_SLICE_X11Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00aa3caa3c)
  ) CLBLM_L_X8Y114_SLICE_X11Y114_CLUT (
.I0(CLBLM_L_X8Y115_SLICE_X11Y115_AQ),
.I1(CLBLM_L_X10Y114_SLICE_X12Y114_BQ),
.I2(CLBLM_L_X8Y111_SLICE_X10Y111_BO5),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X8Y114_SLICE_X11Y114_CO5),
.O6(CLBLM_L_X8Y114_SLICE_X11Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fc000ccacacaca)
  ) CLBLM_L_X8Y114_SLICE_X11Y114_BLUT (
.I0(CLBLM_L_X8Y109_SLICE_X11Y109_BQ),
.I1(CLBLM_L_X8Y114_SLICE_X11Y114_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_L_X12Y117_SLICE_X17Y117_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y114_SLICE_X11Y114_BO5),
.O6(CLBLM_L_X8Y114_SLICE_X11Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccaaa0aaa0)
  ) CLBLM_L_X8Y114_SLICE_X11Y114_ALUT (
.I0(CLBLL_L_X4Y116_SLICE_X4Y116_BO6),
.I1(CLBLM_L_X8Y111_SLICE_X11Y111_CQ),
.I2(CLBLM_L_X8Y114_SLICE_X11Y114_AQ),
.I3(CLBLM_R_X7Y115_SLICE_X9Y115_BQ),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y114_SLICE_X11Y114_AO5),
.O6(CLBLM_L_X8Y114_SLICE_X11Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y115_SLICE_X10Y115_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y115_SLICE_X14Y115_AO6),
.Q(CLBLM_L_X8Y115_SLICE_X10Y115_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y115_SLICE_X10Y115_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y115_SLICE_X10Y115_AO6),
.Q(CLBLM_L_X8Y115_SLICE_X10Y115_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y115_SLICE_X10Y115_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y115_SLICE_X10Y115_BO6),
.Q(CLBLM_L_X8Y115_SLICE_X10Y115_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y115_SLICE_X10Y115_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y115_SLICE_X10Y115_CO6),
.Q(CLBLM_L_X8Y115_SLICE_X10Y115_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffbfff)
  ) CLBLM_L_X8Y115_SLICE_X10Y115_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I2(CLBLM_L_X10Y115_SLICE_X12Y115_CQ),
.I3(CLBLM_L_X10Y115_SLICE_X13Y115_DO5),
.I4(CLBLL_L_X4Y114_SLICE_X4Y114_BQ),
.I5(CLBLM_R_X7Y111_SLICE_X9Y111_CQ),
.O5(CLBLM_L_X8Y115_SLICE_X10Y115_DO5),
.O6(CLBLM_L_X8Y115_SLICE_X10Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa0caa0caa0caa0c)
  ) CLBLM_L_X8Y115_SLICE_X10Y115_CLUT (
.I0(CLBLM_L_X8Y114_SLICE_X10Y114_AQ),
.I1(CLBLM_L_X8Y116_SLICE_X11Y116_BQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y115_SLICE_X10Y115_CO5),
.O6(CLBLM_L_X8Y115_SLICE_X10Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000c0cff000c0c)
  ) CLBLM_L_X8Y115_SLICE_X10Y115_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y115_SLICE_X10Y115_BQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X7Y111_SLICE_X9Y111_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y115_SLICE_X10Y115_BO5),
.O6(CLBLM_L_X8Y115_SLICE_X10Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccfafacccc0000)
  ) CLBLM_L_X8Y115_SLICE_X10Y115_ALUT (
.I0(CLBLM_L_X10Y115_SLICE_X13Y115_BQ),
.I1(CLBLM_R_X11Y118_SLICE_X15Y118_AQ),
.I2(CLBLM_L_X8Y115_SLICE_X10Y115_AQ),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y115_SLICE_X9Y115_DO6),
.O5(CLBLM_L_X8Y115_SLICE_X10Y115_AO5),
.O6(CLBLM_L_X8Y115_SLICE_X10Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y115_SLICE_X11Y115_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y115_SLICE_X11Y115_AO6),
.Q(CLBLM_L_X8Y115_SLICE_X11Y115_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y115_SLICE_X11Y115_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y115_SLICE_X11Y115_BO6),
.Q(CLBLM_L_X8Y115_SLICE_X11Y115_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000300000000)
  ) CLBLM_L_X8Y115_SLICE_X11Y115_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X12Y112_SLICE_X17Y112_BQ),
.I2(CLBLM_L_X12Y112_SLICE_X16Y112_AQ),
.I3(CLBLM_L_X8Y116_SLICE_X11Y116_BQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X7Y115_SLICE_X9Y115_BQ),
.O5(CLBLM_L_X8Y115_SLICE_X11Y115_DO5),
.O6(CLBLM_L_X8Y115_SLICE_X11Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8800000000000000)
  ) CLBLM_L_X8Y115_SLICE_X11Y115_CLUT (
.I0(CLBLM_L_X10Y114_SLICE_X12Y114_BQ),
.I1(CLBLM_L_X8Y114_SLICE_X11Y114_CQ),
.I2(1'b1),
.I3(CLBLM_L_X8Y115_SLICE_X10Y115_CQ),
.I4(CLBLM_L_X8Y115_SLICE_X11Y115_DO6),
.I5(CLBLM_R_X13Y117_SLICE_X18Y117_BQ),
.O5(CLBLM_L_X8Y115_SLICE_X11Y115_CO5),
.O6(CLBLM_L_X8Y115_SLICE_X11Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hafafacaca0a0a0a0)
  ) CLBLM_L_X8Y115_SLICE_X11Y115_BLUT (
.I0(CLBLM_R_X5Y109_SLICE_X6Y109_CQ),
.I1(CLBLM_L_X8Y115_SLICE_X11Y115_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(CLBLM_L_X8Y115_SLICE_X10Y115_AQ),
.I5(CLBLM_R_X7Y115_SLICE_X9Y115_DO6),
.O5(CLBLM_L_X8Y115_SLICE_X11Y115_BO5),
.O6(CLBLM_L_X8Y115_SLICE_X11Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffaffeaaafaaaea)
  ) CLBLM_L_X8Y115_SLICE_X11Y115_ALUT (
.I0(CLBLM_R_X7Y112_SLICE_X9Y112_DO6),
.I1(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.I2(CLBLM_L_X8Y115_SLICE_X11Y115_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLM_R_X5Y116_SLICE_X7Y116_A5Q),
.O5(CLBLM_L_X8Y115_SLICE_X11Y115_AO5),
.O6(CLBLM_L_X8Y115_SLICE_X11Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y116_SLICE_X10Y116_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y116_SLICE_X10Y116_AO6),
.Q(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y116_SLICE_X10Y116_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y116_SLICE_X10Y116_BO6),
.Q(CLBLM_L_X8Y116_SLICE_X10Y116_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y116_SLICE_X10Y116_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y116_SLICE_X10Y116_CO6),
.Q(CLBLM_L_X8Y116_SLICE_X10Y116_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y116_SLICE_X10Y116_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y116_SLICE_X10Y116_DO6),
.Q(CLBLM_L_X8Y116_SLICE_X10Y116_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdfccccc31300000)
  ) CLBLM_L_X8Y116_SLICE_X10Y116_DLUT (
.I0(RIOB33_X105Y121_IOB_X1Y121_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X8Y116_SLICE_X10Y116_DQ),
.I3(CLBLM_R_X11Y113_SLICE_X14Y113_CQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_L_X10Y115_SLICE_X13Y115_CQ),
.O5(CLBLM_L_X8Y116_SLICE_X10Y116_DO5),
.O6(CLBLM_L_X8Y116_SLICE_X10Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa0caaffaa0caa00)
  ) CLBLM_L_X8Y116_SLICE_X10Y116_CLUT (
.I0(CLBLM_R_X7Y115_SLICE_X9Y115_B5Q),
.I1(CLBLM_L_X8Y116_SLICE_X10Y116_CQ),
.I2(CLBLM_L_X10Y117_SLICE_X13Y117_AO5),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y118_SLICE_X8Y118_DO6),
.I5(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.O5(CLBLM_L_X8Y116_SLICE_X10Y116_CO5),
.O6(CLBLM_L_X8Y116_SLICE_X10Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff005050d8d8)
  ) CLBLM_L_X8Y116_SLICE_X10Y116_BLUT (
.I0(CLBLM_R_X7Y118_SLICE_X8Y118_DO6),
.I1(CLBLM_L_X8Y116_SLICE_X10Y116_BQ),
.I2(CLBLM_L_X8Y117_SLICE_X10Y117_AQ),
.I3(CLBLM_R_X5Y112_SLICE_X6Y112_AQ),
.I4(CLBLM_L_X10Y117_SLICE_X13Y117_AO5),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y116_SLICE_X10Y116_BO5),
.O6(CLBLM_L_X8Y116_SLICE_X10Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff010001ff000000)
  ) CLBLM_L_X8Y116_SLICE_X10Y116_ALUT (
.I0(CLBLM_L_X8Y113_SLICE_X10Y113_DQ),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X5Y112_SLICE_X7Y112_BQ),
.I5(RIOB33_X105Y119_IOB_X1Y119_I),
.O5(CLBLM_L_X8Y116_SLICE_X10Y116_AO5),
.O6(CLBLM_L_X8Y116_SLICE_X10Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y116_SLICE_X11Y116_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y116_SLICE_X11Y116_AO6),
.Q(CLBLM_L_X8Y116_SLICE_X11Y116_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y116_SLICE_X11Y116_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y116_SLICE_X11Y116_BO6),
.Q(CLBLM_L_X8Y116_SLICE_X11Y116_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0ff00ff00ff00ff0)
  ) CLBLM_L_X8Y116_SLICE_X11Y116_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X13Y117_SLICE_X18Y117_BQ),
.I3(CLBLM_R_X5Y112_SLICE_X7Y112_CQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y116_SLICE_X11Y116_DO5),
.O6(CLBLM_L_X8Y116_SLICE_X11Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h333311333f3f153f)
  ) CLBLM_L_X8Y116_SLICE_X11Y116_CLUT (
.I0(CLBLM_R_X7Y114_SLICE_X8Y114_A5Q),
.I1(CLBLM_L_X10Y115_SLICE_X13Y115_CQ),
.I2(CLBLM_R_X7Y118_SLICE_X8Y118_CQ),
.I3(CLBLM_L_X8Y118_SLICE_X10Y118_AQ),
.I4(CLBLM_R_X11Y117_SLICE_X15Y117_AQ),
.I5(CLBLM_L_X10Y119_SLICE_X12Y119_AQ),
.O5(CLBLM_L_X8Y116_SLICE_X11Y116_CO5),
.O6(CLBLM_L_X8Y116_SLICE_X11Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f022f099f044)
  ) CLBLM_L_X8Y116_SLICE_X11Y116_BLUT (
.I0(CLBLM_L_X8Y116_SLICE_X11Y116_DO6),
.I1(CLBLM_L_X8Y116_SLICE_X11Y116_BQ),
.I2(CLBLM_L_X10Y117_SLICE_X12Y117_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X12Y112_SLICE_X17Y112_BQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X8Y116_SLICE_X11Y116_BO5),
.O6(CLBLM_L_X8Y116_SLICE_X11Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0cacacaca)
  ) CLBLM_L_X8Y116_SLICE_X11Y116_ALUT (
.I0(CLBLM_R_X7Y116_SLICE_X8Y116_BQ),
.I1(CLBLM_L_X12Y108_SLICE_X17Y108_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X10Y116_SLICE_X12Y116_DO6),
.O5(CLBLM_L_X8Y116_SLICE_X11Y116_AO5),
.O6(CLBLM_L_X8Y116_SLICE_X11Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y117_SLICE_X10Y117_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y117_SLICE_X10Y117_AO6),
.Q(CLBLM_L_X8Y117_SLICE_X10Y117_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y117_SLICE_X10Y117_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y117_SLICE_X10Y117_BO6),
.Q(CLBLM_L_X8Y117_SLICE_X10Y117_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffcccc)
  ) CLBLM_L_X8Y117_SLICE_X10Y117_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y119_SLICE_X12Y119_AQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X7Y118_SLICE_X8Y118_CQ),
.I5(CLBLM_R_X7Y114_SLICE_X8Y114_A5Q),
.O5(CLBLM_L_X8Y117_SLICE_X10Y117_DO5),
.O6(CLBLM_L_X8Y117_SLICE_X10Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0f5f0f1f0f)
  ) CLBLM_L_X8Y117_SLICE_X10Y117_CLUT (
.I0(CLBLM_L_X10Y116_SLICE_X12Y116_DO6),
.I1(CLBLM_R_X11Y117_SLICE_X15Y117_AQ),
.I2(CLBLM_L_X8Y117_SLICE_X10Y117_BQ),
.I3(CLBLM_R_X7Y116_SLICE_X8Y116_BQ),
.I4(CLBLM_L_X8Y117_SLICE_X10Y117_DO6),
.I5(CLBLM_R_X7Y116_SLICE_X9Y116_CO6),
.O5(CLBLM_L_X8Y117_SLICE_X10Y117_CO5),
.O6(CLBLM_L_X8Y117_SLICE_X10Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaf3c0aaaaf3f3)
  ) CLBLM_L_X8Y117_SLICE_X10Y117_BLUT (
.I0(CLBLM_R_X13Y113_SLICE_X18Y113_BQ),
.I1(CLBLM_L_X10Y117_SLICE_X13Y117_AO5),
.I2(CLBLM_R_X7Y110_SLICE_X8Y110_DO5),
.I3(CLBLM_L_X8Y118_SLICE_X10Y118_DO5),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y117_SLICE_X10Y117_CO6),
.O5(CLBLM_L_X8Y117_SLICE_X10Y117_BO5),
.O6(CLBLM_L_X8Y117_SLICE_X10Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0075752020)
  ) CLBLM_L_X8Y117_SLICE_X10Y117_ALUT (
.I0(CLBLM_R_X7Y118_SLICE_X8Y118_DO6),
.I1(CLBLM_L_X10Y117_SLICE_X13Y117_AO5),
.I2(CLBLM_L_X8Y117_SLICE_X10Y117_AQ),
.I3(CLBLM_R_X5Y116_SLICE_X7Y116_BQ),
.I4(CLBLM_L_X10Y116_SLICE_X13Y116_BQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y117_SLICE_X10Y117_AO5),
.O6(CLBLM_L_X8Y117_SLICE_X10Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y117_SLICE_X11Y117_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y117_SLICE_X11Y117_DO5),
.O6(CLBLM_L_X8Y117_SLICE_X11Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y117_SLICE_X11Y117_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y117_SLICE_X11Y117_CO5),
.O6(CLBLM_L_X8Y117_SLICE_X11Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y117_SLICE_X11Y117_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y117_SLICE_X11Y117_BO5),
.O6(CLBLM_L_X8Y117_SLICE_X11Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y117_SLICE_X11Y117_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y117_SLICE_X11Y117_AO5),
.O6(CLBLM_L_X8Y117_SLICE_X11Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y118_SLICE_X10Y118_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y118_SLICE_X10Y118_AO6),
.Q(CLBLM_L_X8Y118_SLICE_X10Y118_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y118_SLICE_X10Y118_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y118_SLICE_X10Y118_BO6),
.Q(CLBLM_L_X8Y118_SLICE_X10Y118_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7ddd7ddd03000300)
  ) CLBLM_L_X8Y118_SLICE_X10Y118_DLUT (
.I0(CLBLM_L_X10Y117_SLICE_X13Y117_CO6),
.I1(CLBLM_L_X8Y118_SLICE_X10Y118_AQ),
.I2(CLBLM_R_X7Y118_SLICE_X8Y118_CQ),
.I3(CLBLM_L_X10Y119_SLICE_X12Y119_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y118_SLICE_X10Y118_DO5),
.O6(CLBLM_L_X8Y118_SLICE_X10Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0503f1ffcfc0000)
  ) CLBLM_L_X8Y118_SLICE_X10Y118_CLUT (
.I0(CLBLM_R_X7Y114_SLICE_X8Y114_A5Q),
.I1(CLBLM_L_X10Y119_SLICE_X12Y119_AQ),
.I2(CLBLM_L_X8Y118_SLICE_X10Y118_AQ),
.I3(CLBLM_R_X11Y117_SLICE_X15Y117_AQ),
.I4(CLBLM_R_X7Y118_SLICE_X8Y118_CQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y118_SLICE_X10Y118_CO5),
.O6(CLBLM_L_X8Y118_SLICE_X10Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fcf0fc000c000c)
  ) CLBLM_L_X8Y118_SLICE_X10Y118_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y118_SLICE_X10Y118_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(1'b1),
.I5(CLBLM_R_X7Y117_SLICE_X8Y117_BQ),
.O5(CLBLM_L_X8Y118_SLICE_X10Y118_BO5),
.O6(CLBLM_L_X8Y118_SLICE_X10Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00fa50aa00be14)
  ) CLBLM_L_X8Y118_SLICE_X10Y118_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y117_SLICE_X13Y117_CO6),
.I2(CLBLM_L_X8Y118_SLICE_X10Y118_AQ),
.I3(CLBLM_L_X8Y116_SLICE_X11Y116_BQ),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(CLBLM_L_X8Y118_SLICE_X10Y118_CO6),
.O5(CLBLM_L_X8Y118_SLICE_X10Y118_AO5),
.O6(CLBLM_L_X8Y118_SLICE_X10Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y118_SLICE_X11Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y118_SLICE_X11Y118_DO5),
.O6(CLBLM_L_X8Y118_SLICE_X11Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y118_SLICE_X11Y118_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y118_SLICE_X11Y118_CO5),
.O6(CLBLM_L_X8Y118_SLICE_X11Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y118_SLICE_X11Y118_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y118_SLICE_X11Y118_BO5),
.O6(CLBLM_L_X8Y118_SLICE_X11Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y118_SLICE_X11Y118_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y118_SLICE_X11Y118_AO5),
.O6(CLBLM_L_X8Y118_SLICE_X11Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y119_SLICE_X10Y119_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y119_SLICE_X10Y119_AO6),
.Q(CLBLM_L_X8Y119_SLICE_X10Y119_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y119_SLICE_X10Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y119_SLICE_X10Y119_DO5),
.O6(CLBLM_L_X8Y119_SLICE_X10Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y119_SLICE_X10Y119_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y119_SLICE_X10Y119_CO5),
.O6(CLBLM_L_X8Y119_SLICE_X10Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y119_SLICE_X10Y119_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y119_SLICE_X10Y119_BO5),
.O6(CLBLM_L_X8Y119_SLICE_X10Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hb8bb888800ff0000)
  ) CLBLM_L_X8Y119_SLICE_X10Y119_ALUT (
.I0(CLBLM_L_X10Y115_SLICE_X13Y115_BQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X8Y119_SLICE_X10Y119_AQ),
.I3(RIOB33_X105Y141_IOB_X1Y142_I),
.I4(CLBLM_L_X12Y112_SLICE_X16Y112_B5Q),
.I5(1'b1),
.O5(CLBLM_L_X8Y119_SLICE_X10Y119_AO5),
.O6(CLBLM_L_X8Y119_SLICE_X10Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y119_SLICE_X11Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y119_SLICE_X11Y119_DO5),
.O6(CLBLM_L_X8Y119_SLICE_X11Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y119_SLICE_X11Y119_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y119_SLICE_X11Y119_CO5),
.O6(CLBLM_L_X8Y119_SLICE_X11Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y119_SLICE_X11Y119_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y119_SLICE_X11Y119_BO5),
.O6(CLBLM_L_X8Y119_SLICE_X11Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y119_SLICE_X11Y119_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y119_SLICE_X11Y119_AO5),
.O6(CLBLM_L_X8Y119_SLICE_X11Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y104_SLICE_X12Y104_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y104_SLICE_X12Y104_AO6),
.Q(CLBLM_L_X10Y104_SLICE_X12Y104_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y104_SLICE_X12Y104_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y104_SLICE_X12Y104_DO5),
.O6(CLBLM_L_X10Y104_SLICE_X12Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffff5f0faf0)
  ) CLBLM_L_X10Y104_SLICE_X12Y104_CLUT (
.I0(CLBLM_R_X3Y108_SLICE_X3Y108_CO6),
.I1(1'b1),
.I2(CLBLM_L_X10Y105_SLICE_X12Y105_DO6),
.I3(CLBLM_L_X12Y110_SLICE_X16Y110_DO5),
.I4(CLBLM_L_X10Y105_SLICE_X13Y105_CO6),
.I5(CLBLM_L_X8Y104_SLICE_X11Y104_BO6),
.O5(CLBLM_L_X10Y104_SLICE_X12Y104_CO5),
.O6(CLBLM_L_X10Y104_SLICE_X12Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h02ff01ffffffffff)
  ) CLBLM_L_X10Y104_SLICE_X12Y104_BLUT (
.I0(CLBLM_L_X10Y105_SLICE_X13Y105_CO6),
.I1(CLBLM_L_X8Y104_SLICE_X11Y104_BO6),
.I2(CLBLM_L_X10Y105_SLICE_X12Y105_DO6),
.I3(CLBLM_L_X12Y110_SLICE_X16Y110_DO5),
.I4(CLBLM_R_X3Y108_SLICE_X3Y108_CO6),
.I5(CLBLM_L_X10Y106_SLICE_X12Y106_BO6),
.O5(CLBLM_L_X10Y104_SLICE_X12Y104_BO5),
.O6(CLBLM_L_X10Y104_SLICE_X12Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8888888888d888d8)
  ) CLBLM_L_X10Y104_SLICE_X12Y104_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y106_SLICE_X13Y106_BQ),
.I2(CLBLM_L_X10Y104_SLICE_X12Y104_AQ),
.I3(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.I4(1'b1),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_L_X10Y104_SLICE_X12Y104_AO5),
.O6(CLBLM_L_X10Y104_SLICE_X12Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y104_SLICE_X13Y104_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y104_SLICE_X13Y104_DO5),
.O6(CLBLM_L_X10Y104_SLICE_X13Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y104_SLICE_X13Y104_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y104_SLICE_X13Y104_CO5),
.O6(CLBLM_L_X10Y104_SLICE_X13Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y104_SLICE_X13Y104_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y104_SLICE_X13Y104_BO5),
.O6(CLBLM_L_X10Y104_SLICE_X13Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y104_SLICE_X13Y104_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y104_SLICE_X13Y104_AO5),
.O6(CLBLM_L_X10Y104_SLICE_X13Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y105_SLICE_X12Y105_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y105_SLICE_X12Y105_AO6),
.Q(CLBLM_L_X10Y105_SLICE_X12Y105_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y105_SLICE_X12Y105_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y105_SLICE_X12Y105_BO6),
.Q(CLBLM_L_X10Y105_SLICE_X12Y105_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff7dffbeff7dffbe)
  ) CLBLM_L_X10Y105_SLICE_X12Y105_DLUT (
.I0(CLBLM_L_X8Y106_SLICE_X11Y106_BQ),
.I1(CLBLM_L_X10Y108_SLICE_X12Y108_BQ),
.I2(CLBLM_L_X8Y107_SLICE_X10Y107_BQ),
.I3(CLBLM_L_X8Y106_SLICE_X11Y106_DO6),
.I4(CLBLM_R_X11Y106_SLICE_X14Y106_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y105_SLICE_X12Y105_DO5),
.O6(CLBLM_L_X10Y105_SLICE_X12Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0040000080800000)
  ) CLBLM_L_X10Y105_SLICE_X12Y105_CLUT (
.I0(CLBLM_L_X10Y106_SLICE_X12Y106_AQ),
.I1(CLBLM_L_X10Y105_SLICE_X12Y105_AQ),
.I2(CLBLM_R_X11Y105_SLICE_X14Y105_CQ),
.I3(CLBLM_R_X5Y115_SLICE_X7Y115_CO6),
.I4(CLBLM_R_X11Y105_SLICE_X14Y105_C5Q),
.I5(1'b1),
.O5(CLBLM_L_X10Y105_SLICE_X12Y105_CO5),
.O6(CLBLM_L_X10Y105_SLICE_X12Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffd800d8ff500050)
  ) CLBLM_L_X10Y105_SLICE_X12Y105_BLUT (
.I0(CLBLM_L_X10Y106_SLICE_X12Y106_BO6),
.I1(CLBLM_L_X10Y105_SLICE_X12Y105_BQ),
.I2(CLBLM_L_X8Y105_SLICE_X10Y105_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X11Y106_SLICE_X14Y106_AQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X10Y105_SLICE_X12Y105_BO5),
.O6(CLBLM_L_X10Y105_SLICE_X12Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffa0ff82a0a08282)
  ) CLBLM_L_X10Y105_SLICE_X12Y105_ALUT (
.I0(CLBLM_R_X7Y106_SLICE_X9Y106_DO6),
.I1(CLBLM_R_X5Y115_SLICE_X7Y115_CO6),
.I2(CLBLM_L_X10Y105_SLICE_X12Y105_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y105_SLICE_X12Y105_CO5),
.I5(CLBLM_L_X8Y107_SLICE_X10Y107_CQ),
.O5(CLBLM_L_X10Y105_SLICE_X12Y105_AO5),
.O6(CLBLM_L_X10Y105_SLICE_X12Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffeeffee)
  ) CLBLM_L_X10Y105_SLICE_X13Y105_DLUT (
.I0(CLBLM_L_X10Y107_SLICE_X12Y107_AQ),
.I1(CLBLM_R_X11Y105_SLICE_X14Y105_AQ),
.I2(1'b1),
.I3(CLBLM_L_X8Y105_SLICE_X11Y105_BQ),
.I4(1'b1),
.I5(CLBLM_L_X10Y105_SLICE_X12Y105_BQ),
.O5(CLBLM_L_X10Y105_SLICE_X13Y105_DO5),
.O6(CLBLM_L_X10Y105_SLICE_X13Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h9999999999998989)
  ) CLBLM_L_X10Y105_SLICE_X13Y105_CLUT (
.I0(CLBLM_R_X11Y105_SLICE_X14Y105_BQ),
.I1(CLBLM_L_X10Y111_SLICE_X13Y111_BQ),
.I2(CLBLM_L_X10Y106_SLICE_X12Y106_DO6),
.I3(1'b1),
.I4(CLBLM_L_X10Y105_SLICE_X13Y105_DO6),
.I5(CLBLM_L_X8Y105_SLICE_X10Y105_DO6),
.O5(CLBLM_L_X10Y105_SLICE_X13Y105_CO5),
.O6(CLBLM_L_X10Y105_SLICE_X13Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888a2228888)
  ) CLBLM_L_X10Y105_SLICE_X13Y105_BLUT (
.I0(CLBLM_R_X7Y106_SLICE_X9Y106_DO6),
.I1(CLBLM_R_X11Y105_SLICE_X14Y105_CQ),
.I2(CLBLM_L_X10Y106_SLICE_X12Y106_AQ),
.I3(CLBLM_R_X11Y105_SLICE_X14Y105_C5Q),
.I4(CLBLM_L_X10Y105_SLICE_X12Y105_AQ),
.I5(CLBLM_R_X5Y115_SLICE_X7Y115_CO6),
.O5(CLBLM_L_X10Y105_SLICE_X13Y105_BO5),
.O6(CLBLM_L_X10Y105_SLICE_X13Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00a288aa00)
  ) CLBLM_L_X10Y105_SLICE_X13Y105_ALUT (
.I0(CLBLM_R_X7Y106_SLICE_X9Y106_DO6),
.I1(CLBLM_R_X11Y105_SLICE_X14Y105_CQ),
.I2(CLBLM_L_X10Y106_SLICE_X12Y106_AQ),
.I3(CLBLM_R_X11Y105_SLICE_X14Y105_C5Q),
.I4(CLBLM_L_X10Y105_SLICE_X12Y105_AQ),
.I5(CLBLM_R_X5Y115_SLICE_X7Y115_CO6),
.O5(CLBLM_L_X10Y105_SLICE_X13Y105_AO5),
.O6(CLBLM_L_X10Y105_SLICE_X13Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y106_SLICE_X12Y106_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y106_SLICE_X12Y106_AO6),
.Q(CLBLM_L_X10Y106_SLICE_X12Y106_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000001)
  ) CLBLM_L_X10Y106_SLICE_X12Y106_DLUT (
.I0(CLBLM_L_X10Y110_SLICE_X13Y110_AQ),
.I1(CLBLM_L_X10Y110_SLICE_X13Y110_BQ),
.I2(CLBLM_L_X8Y106_SLICE_X11Y106_BQ),
.I3(CLBLM_L_X10Y106_SLICE_X13Y106_CQ),
.I4(CLBLM_L_X10Y107_SLICE_X12Y107_BQ),
.I5(CLBLM_L_X8Y107_SLICE_X10Y107_BQ),
.O5(CLBLM_L_X10Y106_SLICE_X12Y106_DO5),
.O6(CLBLM_L_X10Y106_SLICE_X12Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00a5a58787)
  ) CLBLM_L_X10Y106_SLICE_X12Y106_CLUT (
.I0(CLBLM_R_X11Y110_SLICE_X14Y110_AQ),
.I1(CLBLM_R_X3Y108_SLICE_X2Y108_DO6),
.I2(CLBLM_R_X5Y107_SLICE_X7Y107_AQ),
.I3(CLBLM_L_X10Y105_SLICE_X13Y105_CO6),
.I4(CLBLM_L_X10Y112_SLICE_X12Y112_DO6),
.I5(CLBLM_L_X12Y110_SLICE_X16Y110_DO5),
.O5(CLBLM_L_X10Y106_SLICE_X12Y106_CO5),
.O6(CLBLM_L_X10Y106_SLICE_X12Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00030000aaa8aaaa)
  ) CLBLM_L_X10Y106_SLICE_X12Y106_BLUT (
.I0(CLBLM_L_X10Y107_SLICE_X12Y107_BQ),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_L_X10Y113_SLICE_X13Y113_AQ),
.I3(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.I4(CLBLM_R_X7Y105_SLICE_X8Y105_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y106_SLICE_X12Y106_BO5),
.O6(CLBLM_L_X10Y106_SLICE_X12Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000feaa5400)
  ) CLBLM_L_X10Y106_SLICE_X12Y106_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y105_SLICE_X12Y105_CO6),
.I2(CLBLM_L_X10Y106_SLICE_X12Y106_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_L_X8Y115_SLICE_X10Y115_AQ),
.I5(CLBLM_L_X10Y111_SLICE_X12Y111_CQ),
.O5(CLBLM_L_X10Y106_SLICE_X12Y106_AO5),
.O6(CLBLM_L_X10Y106_SLICE_X12Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y106_SLICE_X13Y106_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y106_SLICE_X13Y106_AO6),
.Q(CLBLM_L_X10Y106_SLICE_X13Y106_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y106_SLICE_X13Y106_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y106_SLICE_X13Y106_BO6),
.Q(CLBLM_L_X10Y106_SLICE_X13Y106_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y106_SLICE_X13Y106_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y106_SLICE_X13Y106_CO6),
.Q(CLBLM_L_X10Y106_SLICE_X13Y106_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff7f33dfcc5f00)
  ) CLBLM_L_X10Y106_SLICE_X13Y106_DLUT (
.I0(CLBLM_L_X12Y105_SLICE_X17Y105_AO6),
.I1(CLBLL_L_X4Y107_SLICE_X4Y107_BO5),
.I2(CLBLM_R_X11Y105_SLICE_X15Y105_BQ),
.I3(CLBLM_L_X12Y107_SLICE_X17Y107_BQ),
.I4(CLBLM_L_X8Y106_SLICE_X10Y106_BQ),
.I5(CLBLM_R_X5Y107_SLICE_X6Y107_BQ),
.O5(CLBLM_L_X10Y106_SLICE_X13Y106_DO5),
.O6(CLBLM_L_X10Y106_SLICE_X13Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0bbf011f011f011)
  ) CLBLM_L_X10Y106_SLICE_X13Y106_CLUT (
.I0(CLBLM_L_X10Y106_SLICE_X12Y106_BO6),
.I1(CLBLM_L_X10Y106_SLICE_X12Y106_CO6),
.I2(CLBLM_R_X13Y109_SLICE_X19Y109_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y106_SLICE_X13Y106_CQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X10Y106_SLICE_X13Y106_CO5),
.O6(CLBLM_L_X10Y106_SLICE_X13Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa00cc00cc)
  ) CLBLM_L_X10Y106_SLICE_X13Y106_BLUT (
.I0(CLBLM_R_X7Y107_SLICE_X9Y107_C5Q),
.I1(CLBLM_L_X10Y106_SLICE_X13Y106_BQ),
.I2(1'b1),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y106_SLICE_X13Y106_BO5),
.O6(CLBLM_L_X10Y106_SLICE_X13Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00aaccaac0)
  ) CLBLM_L_X10Y106_SLICE_X13Y106_ALUT (
.I0(CLBLM_R_X11Y106_SLICE_X14Y106_CQ),
.I1(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.I2(CLBLM_L_X10Y106_SLICE_X13Y106_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y107_SLICE_X13Y107_AQ),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_L_X10Y106_SLICE_X13Y106_AO5),
.O6(CLBLM_L_X10Y106_SLICE_X13Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y107_SLICE_X12Y107_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y107_SLICE_X12Y107_AO6),
.Q(CLBLM_L_X10Y107_SLICE_X12Y107_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y107_SLICE_X12Y107_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y107_SLICE_X12Y107_BO6),
.Q(CLBLM_L_X10Y107_SLICE_X12Y107_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0aaa2aaa2)
  ) CLBLM_L_X10Y107_SLICE_X12Y107_DLUT (
.I0(CLBLM_L_X10Y104_SLICE_X12Y104_AQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_L_X10Y110_SLICE_X12Y110_CO6),
.I3(CLBLM_R_X3Y108_SLICE_X2Y108_DO6),
.I4(1'b1),
.I5(CLBLM_R_X7Y116_SLICE_X8Y116_CQ),
.O5(CLBLM_L_X10Y107_SLICE_X12Y107_DO5),
.O6(CLBLM_L_X10Y107_SLICE_X12Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000003aaaaaaab)
  ) CLBLM_L_X10Y107_SLICE_X12Y107_CLUT (
.I0(RIOB33_X105Y141_IOB_X1Y142_I),
.I1(CLBLM_R_X5Y115_SLICE_X7Y115_CO6),
.I2(CLBLM_L_X10Y112_SLICE_X12Y112_DO6),
.I3(CLBLM_R_X3Y108_SLICE_X2Y108_DO6),
.I4(CLBLM_R_X11Y108_SLICE_X15Y108_DO6),
.I5(CLBLM_L_X8Y119_SLICE_X10Y119_AQ),
.O5(CLBLM_L_X10Y107_SLICE_X12Y107_CO5),
.O6(CLBLM_L_X10Y107_SLICE_X12Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffa0cc0000a0cc)
  ) CLBLM_L_X10Y107_SLICE_X12Y107_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X8Y105_SLICE_X11Y105_BQ),
.I2(CLBLM_L_X10Y107_SLICE_X12Y107_BQ),
.I3(CLBLM_L_X10Y106_SLICE_X12Y106_BO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X11Y116_SLICE_X14Y116_BQ),
.O5(CLBLM_L_X10Y107_SLICE_X12Y107_BO5),
.O6(CLBLM_L_X10Y107_SLICE_X12Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaf000aaaacccc)
  ) CLBLM_L_X10Y107_SLICE_X12Y107_ALUT (
.I0(CLBLM_L_X8Y108_SLICE_X10Y108_CQ),
.I1(CLBLM_L_X10Y107_SLICE_X12Y107_BQ),
.I2(CLBLM_L_X10Y107_SLICE_X12Y107_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X10Y106_SLICE_X12Y106_BO6),
.O5(CLBLM_L_X10Y107_SLICE_X12Y107_AO5),
.O6(CLBLM_L_X10Y107_SLICE_X12Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y107_SLICE_X13Y107_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y107_SLICE_X13Y107_AO6),
.Q(CLBLM_L_X10Y107_SLICE_X13Y107_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_L_X10Y107_SLICE_X13Y107_DLUT (
.I0(CLBLL_L_X2Y108_SLICE_X1Y108_AO6),
.I1(CLBLM_R_X11Y106_SLICE_X14Y106_CQ),
.I2(CLBLM_L_X12Y105_SLICE_X17Y105_CO6),
.I3(CLBLM_R_X7Y114_SLICE_X9Y114_CO6),
.I4(CLBLM_R_X11Y106_SLICE_X15Y106_CO5),
.I5(CLBLM_L_X10Y107_SLICE_X13Y107_BO6),
.O5(CLBLM_L_X10Y107_SLICE_X13Y107_DO5),
.O6(CLBLM_L_X10Y107_SLICE_X13Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000010)
  ) CLBLM_L_X10Y107_SLICE_X13Y107_CLUT (
.I0(CLBLM_L_X10Y105_SLICE_X12Y105_CO5),
.I1(CLBLM_L_X8Y115_SLICE_X11Y115_BQ),
.I2(CLBLM_L_X10Y105_SLICE_X12Y105_AQ),
.I3(CLBLM_R_X5Y115_SLICE_X7Y115_DO6),
.I4(CLBLM_L_X10Y107_SLICE_X13Y107_DO6),
.I5(CLBLM_R_X3Y107_SLICE_X3Y107_CO6),
.O5(CLBLM_L_X10Y107_SLICE_X13Y107_CO5),
.O6(CLBLM_L_X10Y107_SLICE_X13Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffd)
  ) CLBLM_L_X10Y107_SLICE_X13Y107_BLUT (
.I0(CLBLM_L_X10Y106_SLICE_X12Y106_BO5),
.I1(CLBLM_L_X8Y107_SLICE_X11Y107_BQ),
.I2(CLBLM_R_X11Y105_SLICE_X15Y105_BQ),
.I3(CLBLM_L_X12Y110_SLICE_X17Y110_BQ),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(CLBLM_R_X11Y107_SLICE_X14Y107_BO6),
.O5(CLBLM_L_X10Y107_SLICE_X13Y107_BO5),
.O6(CLBLM_L_X10Y107_SLICE_X13Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000f0ccf0ff)
  ) CLBLM_L_X10Y107_SLICE_X13Y107_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y119_SLICE_X10Y119_AQ),
.I2(CLBLM_R_X7Y106_SLICE_X8Y106_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y141_IOB_X1Y142_I),
.I5(CLBLM_L_X10Y108_SLICE_X13Y108_BO6),
.O5(CLBLM_L_X10Y107_SLICE_X13Y107_AO5),
.O6(CLBLM_L_X10Y107_SLICE_X13Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y108_SLICE_X12Y108_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y108_SLICE_X12Y108_BO6),
.Q(CLBLM_L_X10Y108_SLICE_X12Y108_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y108_SLICE_X12Y108_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y108_SLICE_X12Y108_CO6),
.Q(CLBLM_L_X10Y108_SLICE_X12Y108_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000033335a55)
  ) CLBLM_L_X10Y108_SLICE_X12Y108_DLUT (
.I0(CLBLM_L_X10Y110_SLICE_X12Y110_AQ),
.I1(CLBLM_L_X8Y112_SLICE_X10Y112_AQ),
.I2(CLBLM_R_X11Y108_SLICE_X15Y108_AO5),
.I3(CLBLM_L_X10Y108_SLICE_X12Y108_AO5),
.I4(CLBLM_R_X5Y115_SLICE_X7Y115_CO6),
.I5(CLBLM_L_X8Y108_SLICE_X10Y108_CQ),
.O5(CLBLM_L_X10Y108_SLICE_X12Y108_DO5),
.O6(CLBLM_L_X10Y108_SLICE_X12Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000ff005a5a)
  ) CLBLM_L_X10Y108_SLICE_X12Y108_CLUT (
.I0(CLBLM_L_X10Y110_SLICE_X12Y110_CO5),
.I1(1'b1),
.I2(CLBLM_R_X5Y108_SLICE_X7Y108_AQ),
.I3(CLBLM_R_X11Y105_SLICE_X15Y105_A5Q),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X10Y108_SLICE_X12Y108_CO5),
.O6(CLBLM_L_X10Y108_SLICE_X12Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00aaaaff00acac)
  ) CLBLM_L_X10Y108_SLICE_X12Y108_BLUT (
.I0(CLBLM_R_X5Y112_SLICE_X6Y112_CQ),
.I1(CLBLM_L_X10Y108_SLICE_X12Y108_BQ),
.I2(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.I3(CLBLM_R_X11Y108_SLICE_X14Y108_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_L_X10Y108_SLICE_X12Y108_BO5),
.O6(CLBLM_L_X10Y108_SLICE_X12Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdff020030303030)
  ) CLBLM_L_X10Y108_SLICE_X12Y108_ALUT (
.I0(CLBLM_L_X10Y105_SLICE_X12Y105_AQ),
.I1(CLBLM_R_X11Y105_SLICE_X14Y105_C5Q),
.I2(CLBLM_L_X10Y106_SLICE_X12Y106_AQ),
.I3(CLBLM_R_X11Y105_SLICE_X14Y105_CQ),
.I4(CLBLM_L_X8Y115_SLICE_X10Y115_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y108_SLICE_X12Y108_AO5),
.O6(CLBLM_L_X10Y108_SLICE_X12Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y108_SLICE_X13Y108_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y108_SLICE_X13Y108_AO6),
.Q(CLBLM_L_X10Y108_SLICE_X13Y108_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0eff00f100f10eff)
  ) CLBLM_L_X10Y108_SLICE_X13Y108_DLUT (
.I0(CLBLM_R_X3Y110_SLICE_X2Y110_BO6),
.I1(CLBLL_L_X4Y107_SLICE_X5Y107_BO6),
.I2(CLBLM_R_X5Y115_SLICE_X7Y115_DO6),
.I3(CLBLM_R_X7Y107_SLICE_X9Y107_C5Q),
.I4(CLBLM_L_X10Y109_SLICE_X13Y109_BO5),
.I5(CLBLM_L_X8Y109_SLICE_X11Y109_CQ),
.O5(CLBLM_L_X10Y108_SLICE_X13Y108_DO5),
.O6(CLBLM_L_X10Y108_SLICE_X13Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h000011140000bbbe)
  ) CLBLM_L_X10Y108_SLICE_X13Y108_CLUT (
.I0(CLBLM_R_X5Y115_SLICE_X7Y115_CO6),
.I1(CLBLM_L_X8Y115_SLICE_X11Y115_BQ),
.I2(CLBLM_L_X10Y109_SLICE_X13Y109_AO5),
.I3(CLBLM_R_X11Y105_SLICE_X14Y105_CQ),
.I4(CLBLM_L_X10Y108_SLICE_X13Y108_AQ),
.I5(CLBLM_R_X13Y112_SLICE_X18Y112_A5Q),
.O5(CLBLM_L_X10Y108_SLICE_X13Y108_CO5),
.O6(CLBLM_L_X10Y108_SLICE_X13Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0207070202020707)
  ) CLBLM_L_X10Y108_SLICE_X13Y108_BLUT (
.I0(CLBLM_R_X5Y115_SLICE_X7Y115_CO6),
.I1(CLBLM_R_X11Y108_SLICE_X15Y108_AQ),
.I2(CLBLM_L_X10Y107_SLICE_X13Y107_AQ),
.I3(CLBLM_L_X10Y109_SLICE_X13Y109_AO5),
.I4(CLBLM_L_X12Y110_SLICE_X17Y110_AQ),
.I5(CLBLM_R_X11Y105_SLICE_X14Y105_CQ),
.O5(CLBLM_L_X10Y108_SLICE_X13Y108_BO5),
.O6(CLBLM_L_X10Y108_SLICE_X13Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0cfc0cfcf)
  ) CLBLM_L_X10Y108_SLICE_X13Y108_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X13Y110_SLICE_X19Y110_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y119_SLICE_X10Y119_AQ),
.I4(RIOB33_X105Y141_IOB_X1Y142_I),
.I5(CLBLM_L_X10Y108_SLICE_X13Y108_CO6),
.O5(CLBLM_L_X10Y108_SLICE_X13Y108_AO5),
.O6(CLBLM_L_X10Y108_SLICE_X13Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y109_SLICE_X12Y109_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y109_SLICE_X12Y109_AO6),
.Q(CLBLM_L_X10Y109_SLICE_X12Y109_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y109_SLICE_X12Y109_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y109_SLICE_X12Y109_BO6),
.Q(CLBLM_L_X10Y109_SLICE_X12Y109_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00dd005d00)
  ) CLBLM_L_X10Y109_SLICE_X12Y109_DLUT (
.I0(CLBLM_L_X10Y104_SLICE_X12Y104_AQ),
.I1(CLBLM_L_X10Y110_SLICE_X12Y110_CO5),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_L_X8Y104_SLICE_X11Y104_AO5),
.I4(CLBLM_R_X3Y111_SLICE_X2Y111_CO6),
.I5(CLBLM_R_X7Y116_SLICE_X8Y116_CQ),
.O5(CLBLM_L_X10Y109_SLICE_X12Y109_DO5),
.O6(CLBLM_L_X10Y109_SLICE_X12Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcedfcece33003300)
  ) CLBLM_L_X10Y109_SLICE_X12Y109_CLUT (
.I0(CLBLM_L_X10Y104_SLICE_X12Y104_AQ),
.I1(CLBLM_R_X7Y116_SLICE_X8Y116_CQ),
.I2(CLBLM_L_X8Y109_SLICE_X11Y109_DO6),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X3Y111_SLICE_X2Y111_CO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y109_SLICE_X12Y109_CO5),
.O6(CLBLM_L_X10Y109_SLICE_X12Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf808f808f808f808)
  ) CLBLM_L_X10Y109_SLICE_X12Y109_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X10Y109_SLICE_X12Y109_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X5Y108_SLICE_X7Y108_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y109_SLICE_X12Y109_BO5),
.O6(CLBLM_L_X10Y109_SLICE_X12Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc00ffcccc00f0)
  ) CLBLM_L_X10Y109_SLICE_X12Y109_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y116_SLICE_X8Y116_CQ),
.I2(CLBLM_L_X10Y109_SLICE_X12Y109_AQ),
.I3(CLBLM_R_X5Y115_SLICE_X7Y115_CO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X10Y114_SLICE_X12Y114_CQ),
.O5(CLBLM_L_X10Y109_SLICE_X12Y109_AO5),
.O6(CLBLM_L_X10Y109_SLICE_X12Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hab57a854a854ab57)
  ) CLBLM_L_X10Y109_SLICE_X13Y109_DLUT (
.I0(CLBLM_R_X11Y111_SLICE_X15Y111_C5Q),
.I1(CLBLM_R_X3Y107_SLICE_X3Y107_CO6),
.I2(CLBLM_R_X5Y115_SLICE_X7Y115_DO6),
.I3(CLBLM_R_X11Y115_SLICE_X15Y115_BQ),
.I4(CLBLM_L_X10Y109_SLICE_X13Y109_AO6),
.I5(CLBLM_L_X10Y109_SLICE_X13Y109_BO6),
.O5(CLBLM_L_X10Y109_SLICE_X13Y109_DO5),
.O6(CLBLM_L_X10Y109_SLICE_X13Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000a8ff0000a8a8)
  ) CLBLM_L_X10Y109_SLICE_X13Y109_CLUT (
.I0(RIOB33_X105Y121_IOB_X1Y121_I),
.I1(CLBLM_R_X11Y111_SLICE_X15Y111_BQ),
.I2(CLBLM_L_X8Y109_SLICE_X11Y109_AQ),
.I3(CLBLL_L_X2Y110_SLICE_X1Y110_DO6),
.I4(CLBLM_R_X7Y109_SLICE_X8Y109_DO5),
.I5(CLBLM_L_X10Y109_SLICE_X12Y109_CO5),
.O5(CLBLM_L_X10Y109_SLICE_X13Y109_CO5),
.O6(CLBLM_L_X10Y109_SLICE_X13Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ef1008080000)
  ) CLBLM_L_X10Y109_SLICE_X13Y109_BLUT (
.I0(CLBLM_L_X10Y105_SLICE_X12Y105_AQ),
.I1(CLBLM_R_X11Y105_SLICE_X14Y105_C5Q),
.I2(CLBLM_L_X10Y106_SLICE_X12Y106_AQ),
.I3(CLBLM_R_X7Y110_SLICE_X8Y110_CQ),
.I4(CLBLM_R_X11Y105_SLICE_X14Y105_CQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y109_SLICE_X13Y109_BO5),
.O6(CLBLM_L_X10Y109_SLICE_X13Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfeff0100fbfbfbfb)
  ) CLBLM_L_X10Y109_SLICE_X13Y109_ALUT (
.I0(CLBLM_L_X10Y105_SLICE_X12Y105_AQ),
.I1(CLBLM_R_X11Y105_SLICE_X14Y105_C5Q),
.I2(CLBLM_L_X10Y106_SLICE_X12Y106_AQ),
.I3(CLBLM_R_X11Y105_SLICE_X14Y105_CQ),
.I4(CLBLM_L_X10Y115_SLICE_X13Y115_BQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y109_SLICE_X13Y109_AO5),
.O6(CLBLM_L_X10Y109_SLICE_X13Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y110_SLICE_X12Y110_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y110_SLICE_X12Y110_BO5),
.Q(CLBLM_L_X10Y110_SLICE_X12Y110_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y110_SLICE_X12Y110_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y110_SLICE_X12Y110_AO6),
.Q(CLBLM_L_X10Y110_SLICE_X12Y110_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y110_SLICE_X12Y110_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y110_SLICE_X12Y110_BO6),
.Q(CLBLM_L_X10Y110_SLICE_X12Y110_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffcfffc)
  ) CLBLM_L_X10Y110_SLICE_X12Y110_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y106_SLICE_X13Y106_BQ),
.I2(CLBLM_L_X10Y110_SLICE_X12Y110_BQ),
.I3(CLBLM_L_X8Y110_SLICE_X11Y110_A5Q),
.I4(1'b1),
.I5(CLBLM_L_X10Y109_SLICE_X12Y109_BQ),
.O5(CLBLM_L_X10Y110_SLICE_X12Y110_DO5),
.O6(CLBLM_L_X10Y110_SLICE_X12Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafa0000ccccff00)
  ) CLBLM_L_X10Y110_SLICE_X12Y110_CLUT (
.I0(CLBLM_L_X10Y113_SLICE_X12Y113_BQ),
.I1(CLBLM_R_X13Y112_SLICE_X18Y112_CQ),
.I2(CLBLM_L_X10Y112_SLICE_X12Y112_CQ),
.I3(CLBLM_L_X8Y110_SLICE_X11Y110_CQ),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y110_SLICE_X12Y110_CO5),
.O6(CLBLM_L_X10Y110_SLICE_X12Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf8f80808cfc0cfc0)
  ) CLBLM_L_X10Y110_SLICE_X12Y110_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X10Y110_SLICE_X12Y110_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X5Y110_SLICE_X6Y110_AQ),
.I4(CLBLM_L_X10Y107_SLICE_X12Y107_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y110_SLICE_X12Y110_BO5),
.O6(CLBLM_L_X10Y110_SLICE_X12Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000aaa0aaa0)
  ) CLBLM_L_X10Y110_SLICE_X12Y110_ALUT (
.I0(CLBLM_R_X7Y115_SLICE_X9Y115_DO6),
.I1(1'b1),
.I2(CLBLM_L_X10Y110_SLICE_X12Y110_AQ),
.I3(CLBLM_R_X7Y110_SLICE_X8Y110_CQ),
.I4(CLBLM_L_X8Y108_SLICE_X10Y108_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y110_SLICE_X12Y110_AO5),
.O6(CLBLM_L_X10Y110_SLICE_X12Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y110_SLICE_X13Y110_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y110_SLICE_X13Y110_AO6),
.Q(CLBLM_L_X10Y110_SLICE_X13Y110_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y110_SLICE_X13Y110_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y110_SLICE_X13Y110_BO6),
.Q(CLBLM_L_X10Y110_SLICE_X13Y110_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y110_SLICE_X13Y110_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y110_SLICE_X13Y110_CO6),
.Q(CLBLM_L_X10Y110_SLICE_X13Y110_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y110_SLICE_X13Y110_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y110_SLICE_X13Y110_DO6),
.Q(CLBLM_L_X10Y110_SLICE_X13Y110_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbbaaaaa11100000)
  ) CLBLM_L_X10Y110_SLICE_X13Y110_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_L_X10Y110_SLICE_X13Y110_DQ),
.I3(CLBLM_L_X10Y109_SLICE_X12Y109_CO6),
.I4(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.I5(CLBLM_L_X8Y111_SLICE_X11Y111_AQ),
.O5(CLBLM_L_X10Y110_SLICE_X13Y110_DO5),
.O6(CLBLM_L_X10Y110_SLICE_X13Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffeefaea55445040)
  ) CLBLM_L_X10Y110_SLICE_X13Y110_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y110_SLICE_X13Y110_CQ),
.I2(RIOB33_X105Y117_IOB_X1Y118_I),
.I3(CLBLM_L_X10Y109_SLICE_X12Y109_CO6),
.I4(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.I5(CLBLM_L_X10Y112_SLICE_X12Y112_BQ),
.O5(CLBLM_L_X10Y110_SLICE_X13Y110_CO5),
.O6(CLBLM_L_X10Y110_SLICE_X13Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaccf0aaaa00f0)
  ) CLBLM_L_X10Y110_SLICE_X13Y110_BLUT (
.I0(CLBLM_L_X10Y118_SLICE_X12Y118_BQ),
.I1(CLBLM_L_X10Y110_SLICE_X13Y110_BQ),
.I2(CLBLM_L_X10Y107_SLICE_X12Y107_AQ),
.I3(CLBLM_L_X10Y106_SLICE_X12Y106_BO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X10Y110_SLICE_X13Y110_BO5),
.O6(CLBLM_L_X10Y110_SLICE_X13Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hacafaca0a0afa0a0)
  ) CLBLM_L_X10Y110_SLICE_X13Y110_ALUT (
.I0(CLBLM_R_X7Y111_SLICE_X8Y111_AQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y106_SLICE_X12Y106_BO6),
.I4(CLBLM_R_X11Y105_SLICE_X14Y105_AQ),
.I5(CLBLM_L_X10Y110_SLICE_X13Y110_AQ),
.O5(CLBLM_L_X10Y110_SLICE_X13Y110_AO5),
.O6(CLBLM_L_X10Y110_SLICE_X13Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y111_SLICE_X12Y111_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y113_SLICE_X12Y113_DO6),
.Q(CLBLM_L_X10Y111_SLICE_X12Y111_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y111_SLICE_X12Y111_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y111_SLICE_X12Y111_CO5),
.Q(CLBLM_L_X10Y111_SLICE_X12Y111_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y111_SLICE_X12Y111_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y111_SLICE_X12Y111_AO6),
.Q(CLBLM_L_X10Y111_SLICE_X12Y111_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y111_SLICE_X12Y111_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y111_SLICE_X12Y111_BO6),
.Q(CLBLM_L_X10Y111_SLICE_X12Y111_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y111_SLICE_X12Y111_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y111_SLICE_X12Y111_CO6),
.Q(CLBLM_L_X10Y111_SLICE_X12Y111_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y111_SLICE_X12Y111_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y111_SLICE_X12Y111_DO6),
.Q(CLBLM_L_X10Y111_SLICE_X12Y111_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0f5a0f5a0)
  ) CLBLM_L_X10Y111_SLICE_X12Y111_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(1'b1),
.I2(CLBLM_L_X10Y108_SLICE_X12Y108_BQ),
.I3(CLBLM_L_X8Y112_SLICE_X10Y112_A5Q),
.I4(1'b1),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X10Y111_SLICE_X12Y111_DO5),
.O6(CLBLM_L_X10Y111_SLICE_X12Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd88dd88f5f5a0a0)
  ) CLBLM_L_X10Y111_SLICE_X12Y111_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X11Y109_SLICE_X14Y109_BQ),
.I2(CLBLM_R_X11Y110_SLICE_X15Y110_BQ),
.I3(CLBLM_R_X13Y113_SLICE_X18Y113_AQ),
.I4(CLBLM_L_X8Y117_SLICE_X10Y117_BQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y111_SLICE_X12Y111_CO5),
.O6(CLBLM_L_X10Y111_SLICE_X12Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc0cfc0cf000f000)
  ) CLBLM_L_X10Y111_SLICE_X12Y111_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y111_SLICE_X12Y111_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y113_SLICE_X11Y113_BQ),
.I4(1'b1),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X10Y111_SLICE_X12Y111_BO5),
.O6(CLBLM_L_X10Y111_SLICE_X12Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a3a0a3a0aca0ac)
  ) CLBLM_L_X10Y111_SLICE_X12Y111_ALUT (
.I0(CLBLM_L_X10Y114_SLICE_X12Y114_DQ),
.I1(CLBLM_L_X10Y110_SLICE_X12Y110_CO6),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(1'b1),
.I5(CLBLM_R_X5Y109_SLICE_X7Y109_AQ),
.O5(CLBLM_L_X10Y111_SLICE_X12Y111_AO5),
.O6(CLBLM_L_X10Y111_SLICE_X12Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y111_SLICE_X13Y111_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y111_SLICE_X13Y111_CO5),
.Q(CLBLM_L_X10Y111_SLICE_X13Y111_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y111_SLICE_X13Y111_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y111_SLICE_X13Y111_AO6),
.Q(CLBLM_L_X10Y111_SLICE_X13Y111_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y111_SLICE_X13Y111_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y111_SLICE_X13Y111_BO6),
.Q(CLBLM_L_X10Y111_SLICE_X13Y111_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y111_SLICE_X13Y111_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y111_SLICE_X13Y111_CO6),
.Q(CLBLM_L_X10Y111_SLICE_X13Y111_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00f300ff00b300ff)
  ) CLBLM_L_X10Y111_SLICE_X13Y111_DLUT (
.I0(CLBLM_L_X10Y111_SLICE_X13Y111_C5Q),
.I1(CLBLL_L_X2Y110_SLICE_X1Y110_DO6),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLM_R_X7Y109_SLICE_X8Y109_DO5),
.I4(CLBLM_L_X10Y109_SLICE_X12Y109_CO5),
.I5(CLBLM_L_X8Y111_SLICE_X11Y111_BQ),
.O5(CLBLM_L_X10Y111_SLICE_X13Y111_DO5),
.O6(CLBLM_L_X10Y111_SLICE_X13Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5a0f5a08888d8d8)
  ) CLBLM_L_X10Y111_SLICE_X13Y111_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y106_SLICE_X10Y106_BQ),
.I2(CLBLM_R_X11Y111_SLICE_X15Y111_AQ),
.I3(RIOB33_X105Y103_IOB_X1Y103_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y111_SLICE_X13Y111_CO5),
.O6(CLBLM_L_X10Y111_SLICE_X13Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffca0a0000ca0a)
  ) CLBLM_L_X10Y111_SLICE_X13Y111_BLUT (
.I0(CLBLM_L_X10Y110_SLICE_X13Y110_AQ),
.I1(CLBLM_L_X10Y111_SLICE_X13Y111_BQ),
.I2(CLBLM_L_X10Y106_SLICE_X12Y106_BO6),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y114_SLICE_X11Y114_AQ),
.O5(CLBLM_L_X10Y111_SLICE_X13Y111_BO5),
.O6(CLBLM_L_X10Y111_SLICE_X13Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfe54aa00fe54aa00)
  ) CLBLM_L_X10Y111_SLICE_X13Y111_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X11Y115_SLICE_X15Y115_AQ),
.I2(CLBLM_L_X10Y111_SLICE_X13Y111_AQ),
.I3(CLBLM_R_X11Y106_SLICE_X14Y106_BQ),
.I4(CLBLL_L_X4Y116_SLICE_X4Y116_BO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y111_SLICE_X13Y111_AO5),
.O6(CLBLM_L_X10Y111_SLICE_X13Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y112_SLICE_X12Y112_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y112_SLICE_X12Y112_CO5),
.Q(CLBLM_L_X10Y112_SLICE_X12Y112_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y112_SLICE_X12Y112_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y112_SLICE_X12Y112_AO6),
.Q(CLBLM_L_X10Y112_SLICE_X12Y112_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y112_SLICE_X12Y112_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y112_SLICE_X12Y112_BO6),
.Q(CLBLM_L_X10Y112_SLICE_X12Y112_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y112_SLICE_X12Y112_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y112_SLICE_X12Y112_CO6),
.Q(CLBLM_L_X10Y112_SLICE_X12Y112_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000000c000c)
  ) CLBLM_L_X10Y112_SLICE_X12Y112_DLUT (
.I0(1'b1),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(CLBLM_R_X13Y113_SLICE_X18Y113_DO6),
.I3(RIOB33_X105Y135_IOB_X1Y135_I),
.I4(1'b1),
.I5(RIOB33_X105Y135_IOB_X1Y136_I),
.O5(CLBLM_L_X10Y112_SLICE_X12Y112_DO5),
.O6(CLBLM_L_X10Y112_SLICE_X12Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hb1a0b1a0ff55aa00)
  ) CLBLM_L_X10Y112_SLICE_X12Y112_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X7Y118_SLICE_X8Y118_CQ),
.I3(CLBLM_L_X10Y111_SLICE_X12Y111_DQ),
.I4(CLBLM_L_X12Y112_SLICE_X16Y112_B5Q),
.I5(1'b1),
.O5(CLBLM_L_X10Y112_SLICE_X12Y112_CO5),
.O6(CLBLM_L_X10Y112_SLICE_X12Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fc000cf0f00000)
  ) CLBLM_L_X10Y112_SLICE_X12Y112_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y112_SLICE_X12Y112_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y112_SLICE_X8Y112_CQ),
.I4(CLBLM_L_X12Y112_SLICE_X16Y112_BQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X10Y112_SLICE_X12Y112_BO5),
.O6(CLBLM_L_X10Y112_SLICE_X12Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0fffff0f0eeff)
  ) CLBLM_L_X10Y112_SLICE_X12Y112_ALUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(CLBLM_R_X13Y113_SLICE_X18Y113_DO6),
.I2(CLBLM_L_X8Y110_SLICE_X11Y110_A5Q),
.I3(RIOB33_X105Y135_IOB_X1Y136_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y135_IOB_X1Y135_I),
.O5(CLBLM_L_X10Y112_SLICE_X12Y112_AO5),
.O6(CLBLM_L_X10Y112_SLICE_X12Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y112_SLICE_X13Y112_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y77_IOB_X0Y77_I),
.D(CLBLM_R_X7Y115_SLICE_X9Y115_A5Q),
.Q(CLBLM_L_X10Y112_SLICE_X13Y112_AQ),
.R(CLBLM_L_X12Y117_SLICE_X16Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffefefefe)
  ) CLBLM_L_X10Y112_SLICE_X13Y112_DLUT (
.I0(CLBLM_R_X11Y112_SLICE_X14Y112_BQ),
.I1(CLBLM_R_X7Y112_SLICE_X9Y112_BQ),
.I2(CLBLM_L_X10Y111_SLICE_X13Y111_C5Q),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X12Y111_SLICE_X16Y111_DQ),
.O5(CLBLM_L_X10Y112_SLICE_X13Y112_DO5),
.O6(CLBLM_L_X10Y112_SLICE_X13Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffcfffffffc)
  ) CLBLM_L_X10Y112_SLICE_X13Y112_CLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y111_SLICE_X12Y111_DQ),
.I2(CLBLM_L_X10Y112_SLICE_X12Y112_CQ),
.I3(CLBLM_L_X8Y112_SLICE_X10Y112_A5Q),
.I4(CLBLM_R_X11Y111_SLICE_X15Y111_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y112_SLICE_X13Y112_CO5),
.O6(CLBLM_L_X10Y112_SLICE_X13Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_L_X10Y112_SLICE_X13Y112_BLUT (
.I0(CLBLM_L_X10Y112_SLICE_X13Y112_DO6),
.I1(CLBLM_R_X7Y110_SLICE_X8Y110_BQ),
.I2(CLBLM_L_X12Y112_SLICE_X17Y112_DO6),
.I3(CLBLM_R_X11Y112_SLICE_X14Y112_DO6),
.I4(CLBLM_R_X5Y114_SLICE_X7Y114_BQ),
.I5(CLBLM_R_X11Y112_SLICE_X15Y112_BQ),
.O5(CLBLM_L_X10Y112_SLICE_X13Y112_BO5),
.O6(CLBLM_L_X10Y112_SLICE_X13Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_L_X10Y112_SLICE_X13Y112_ALUT (
.I0(CLBLM_R_X11Y112_SLICE_X14Y112_CQ),
.I1(CLBLM_R_X13Y112_SLICE_X18Y112_CQ),
.I2(CLBLM_R_X5Y109_SLICE_X6Y109_DQ),
.I3(CLBLM_L_X10Y112_SLICE_X13Y112_BO6),
.I4(CLBLM_R_X7Y112_SLICE_X8Y112_C5Q),
.I5(CLBLM_L_X10Y112_SLICE_X13Y112_CO6),
.O5(CLBLM_L_X10Y112_SLICE_X13Y112_AO5),
.O6(CLBLM_L_X10Y112_SLICE_X13Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y113_SLICE_X12Y113_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y113_SLICE_X12Y113_AO6),
.Q(CLBLM_L_X10Y113_SLICE_X12Y113_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y113_SLICE_X12Y113_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y113_SLICE_X12Y113_BO6),
.Q(CLBLM_L_X10Y113_SLICE_X12Y113_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y113_SLICE_X12Y113_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y113_SLICE_X12Y113_CO6),
.Q(CLBLM_L_X10Y113_SLICE_X12Y113_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa50ea400f0f3f3f)
  ) CLBLM_L_X10Y113_SLICE_X12Y113_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X12Y113_SLICE_X17Y113_CQ),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLM_L_X8Y107_SLICE_X10Y107_BQ),
.I4(CLBLM_R_X5Y114_SLICE_X7Y114_BQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y113_SLICE_X12Y113_DO5),
.O6(CLBLM_L_X10Y113_SLICE_X12Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa00fc0000)
  ) CLBLM_L_X10Y113_SLICE_X12Y113_CLUT (
.I0(CLBLM_L_X10Y111_SLICE_X12Y111_AQ),
.I1(CLBLM_L_X10Y113_SLICE_X12Y113_CQ),
.I2(CLBLM_R_X11Y109_SLICE_X14Y109_BQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y113_SLICE_X12Y113_CO5),
.O6(CLBLM_L_X10Y113_SLICE_X12Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffa5550eeea4440)
  ) CLBLM_L_X10Y113_SLICE_X12Y113_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y113_SLICE_X12Y113_BQ),
.I2(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I5(CLBLM_L_X8Y112_SLICE_X11Y112_CO6),
.O5(CLBLM_L_X10Y113_SLICE_X12Y113_BO5),
.O6(CLBLM_L_X10Y113_SLICE_X12Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbb88888bbb88888)
  ) CLBLM_L_X10Y113_SLICE_X12Y113_ALUT (
.I0(CLBLM_L_X10Y110_SLICE_X13Y110_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y113_SLICE_X12Y113_AQ),
.I3(CLBLM_R_X11Y110_SLICE_X15Y110_BQ),
.I4(CLBLL_L_X4Y116_SLICE_X4Y116_BO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y113_SLICE_X12Y113_AO5),
.O6(CLBLM_L_X10Y113_SLICE_X12Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y113_SLICE_X13Y113_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y113_SLICE_X13Y113_CO5),
.Q(CLBLM_L_X10Y113_SLICE_X13Y113_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y113_SLICE_X13Y113_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y113_SLICE_X13Y113_AO6),
.Q(CLBLM_L_X10Y113_SLICE_X13Y113_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y113_SLICE_X13Y113_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y113_SLICE_X13Y113_BO6),
.Q(CLBLM_L_X10Y113_SLICE_X13Y113_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y113_SLICE_X13Y113_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y113_SLICE_X13Y113_CO6),
.Q(CLBLM_L_X10Y113_SLICE_X13Y113_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y113_SLICE_X13Y113_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y113_SLICE_X13Y113_DO6),
.Q(CLBLM_L_X10Y113_SLICE_X13Y113_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffa5550bbba1110)
  ) CLBLM_L_X10Y113_SLICE_X13Y113_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y114_SLICE_X11Y114_B5Q),
.I2(CLBLM_L_X10Y113_SLICE_X13Y113_DQ),
.I3(CLBLM_R_X7Y108_SLICE_X9Y108_AQ),
.I4(CLBLM_R_X13Y113_SLICE_X18Y113_CQ),
.I5(CLBLM_L_X10Y104_SLICE_X12Y104_BO6),
.O5(CLBLM_L_X10Y113_SLICE_X13Y113_DO5),
.O6(CLBLM_L_X10Y113_SLICE_X13Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hb1a0b1a0faff5055)
  ) CLBLM_L_X10Y113_SLICE_X13Y113_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y113_SLICE_X13Y113_CQ),
.I2(CLBLM_L_X8Y113_SLICE_X10Y113_DQ),
.I3(RIOB33_X105Y119_IOB_X1Y119_I),
.I4(CLBLM_R_X5Y109_SLICE_X7Y109_BQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y113_SLICE_X13Y113_CO5),
.O6(CLBLM_L_X10Y113_SLICE_X13Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffc000c0ffcc00cc)
  ) CLBLM_L_X10Y113_SLICE_X13Y113_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y113_SLICE_X13Y113_BQ),
.I2(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y113_SLICE_X13Y113_C5Q),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_L_X10Y113_SLICE_X13Y113_BO5),
.O6(CLBLM_L_X10Y113_SLICE_X13Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffeeffe000ee00e0)
  ) CLBLM_L_X10Y113_SLICE_X13Y113_ALUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.I2(CLBLM_L_X10Y113_SLICE_X13Y113_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y113_SLICE_X13Y113_C5Q),
.I5(CLBLM_L_X10Y113_SLICE_X12Y113_CQ),
.O5(CLBLM_L_X10Y113_SLICE_X13Y113_AO5),
.O6(CLBLM_L_X10Y113_SLICE_X13Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y114_SLICE_X12Y114_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y114_SLICE_X12Y114_AO6),
.Q(CLBLM_L_X10Y114_SLICE_X12Y114_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y114_SLICE_X12Y114_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y114_SLICE_X12Y114_BO6),
.Q(CLBLM_L_X10Y114_SLICE_X12Y114_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y114_SLICE_X12Y114_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y114_SLICE_X12Y114_CO6),
.Q(CLBLM_L_X10Y114_SLICE_X12Y114_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y114_SLICE_X12Y114_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y114_SLICE_X12Y114_DO6),
.Q(CLBLM_L_X10Y114_SLICE_X12Y114_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfeaa5400feaa5400)
  ) CLBLM_L_X10Y114_SLICE_X12Y114_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y114_SLICE_X12Y114_AQ),
.I2(CLBLM_L_X10Y114_SLICE_X12Y114_DQ),
.I3(CLBLM_R_X7Y115_SLICE_X9Y115_DO6),
.I4(CLBLM_L_X8Y108_SLICE_X10Y108_DQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y114_SLICE_X12Y114_DO5),
.O6(CLBLM_L_X10Y114_SLICE_X12Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haafe0054aafe0054)
  ) CLBLM_L_X10Y114_SLICE_X12Y114_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y114_SLICE_X12Y114_CQ),
.I2(CLBLM_R_X11Y113_SLICE_X15Y113_DQ),
.I3(CLBLM_R_X5Y115_SLICE_X7Y115_CO6),
.I4(CLBLM_R_X5Y115_SLICE_X6Y115_BQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y114_SLICE_X12Y114_CO5),
.O6(CLBLM_L_X10Y114_SLICE_X12Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fcf0f3000c0003)
  ) CLBLM_L_X10Y114_SLICE_X12Y114_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y108_SLICE_X10Y108_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_L_X10Y113_SLICE_X12Y113_DO5),
.I5(CLBLM_L_X10Y116_SLICE_X12Y116_BQ),
.O5(CLBLM_L_X10Y114_SLICE_X12Y114_BO5),
.O6(CLBLM_L_X10Y114_SLICE_X12Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haafcaafcaa00aa00)
  ) CLBLM_L_X10Y114_SLICE_X12Y114_ALUT (
.I0(CLBLM_R_X7Y115_SLICE_X8Y115_B5Q),
.I1(CLBLM_L_X12Y114_SLICE_X16Y114_AQ),
.I2(CLBLM_L_X10Y114_SLICE_X12Y114_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLM_R_X7Y115_SLICE_X9Y115_DO6),
.O5(CLBLM_L_X10Y114_SLICE_X12Y114_AO5),
.O6(CLBLM_L_X10Y114_SLICE_X12Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y114_SLICE_X13Y114_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y114_SLICE_X13Y114_AO6),
.Q(CLBLM_L_X10Y114_SLICE_X13Y114_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y114_SLICE_X13Y114_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y114_SLICE_X13Y114_BO6),
.Q(CLBLM_L_X10Y114_SLICE_X13Y114_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y114_SLICE_X13Y114_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y114_SLICE_X13Y114_CO6),
.Q(CLBLM_L_X10Y114_SLICE_X13Y114_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffc)
  ) CLBLM_L_X10Y114_SLICE_X13Y114_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y112_SLICE_X7Y112_CQ),
.I2(CLBLM_L_X10Y115_SLICE_X13Y115_DO6),
.I3(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I4(CLBLM_R_X11Y114_SLICE_X14Y114_CQ),
.I5(CLBLM_L_X8Y108_SLICE_X10Y108_BQ),
.O5(CLBLM_L_X10Y114_SLICE_X13Y114_DO5),
.O6(CLBLM_L_X10Y114_SLICE_X13Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0f5a0f5a0e4a0e4)
  ) CLBLM_L_X10Y114_SLICE_X13Y114_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y114_SLICE_X13Y114_CQ),
.I2(CLBLM_L_X10Y114_SLICE_X13Y114_BQ),
.I3(CLBLM_R_X5Y115_SLICE_X7Y115_CO6),
.I4(1'b1),
.I5(CLBLM_L_X10Y109_SLICE_X12Y109_AQ),
.O5(CLBLM_L_X10Y114_SLICE_X13Y114_CO5),
.O6(CLBLM_L_X10Y114_SLICE_X13Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcacacacacac0cac0)
  ) CLBLM_L_X10Y114_SLICE_X13Y114_BLUT (
.I0(CLBLL_L_X4Y116_SLICE_X4Y116_BO6),
.I1(CLBLM_R_X11Y115_SLICE_X15Y115_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X12Y112_SLICE_X17Y112_BQ),
.I4(1'b1),
.I5(CLBLM_L_X10Y114_SLICE_X13Y114_BQ),
.O5(CLBLM_L_X10Y114_SLICE_X13Y114_BO5),
.O6(CLBLM_L_X10Y114_SLICE_X13Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdfc3130ddcc1100)
  ) CLBLM_L_X10Y114_SLICE_X13Y114_ALUT (
.I0(CLBLM_L_X10Y114_SLICE_X13Y114_DO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y114_SLICE_X13Y114_AQ),
.I3(CLBLM_L_X8Y115_SLICE_X11Y115_CO6),
.I4(CLBLM_L_X12Y114_SLICE_X16Y114_AQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X10Y114_SLICE_X13Y114_AO5),
.O6(CLBLM_L_X10Y114_SLICE_X13Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y115_SLICE_X12Y115_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y115_SLICE_X12Y115_AO6),
.Q(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y115_SLICE_X12Y115_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y115_SLICE_X12Y115_BO6),
.Q(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y115_SLICE_X12Y115_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y115_SLICE_X12Y115_CO6),
.Q(CLBLM_L_X10Y115_SLICE_X12Y115_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y115_SLICE_X12Y115_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y115_SLICE_X12Y115_DO5),
.O6(CLBLM_L_X10Y115_SLICE_X12Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaeeaaee00440044)
  ) CLBLM_L_X10Y115_SLICE_X12Y115_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y115_SLICE_X12Y115_AQ),
.I2(1'b1),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(1'b1),
.I5(CLBLM_L_X10Y114_SLICE_X12Y114_BQ),
.O5(CLBLM_L_X10Y115_SLICE_X12Y115_CO5),
.O6(CLBLM_L_X10Y115_SLICE_X12Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f3f0fc0003000c)
  ) CLBLM_L_X10Y115_SLICE_X12Y115_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y114_SLICE_X11Y114_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X11Y112_SLICE_X14Y112_AO5),
.I5(CLBLM_L_X8Y116_SLICE_X11Y116_AQ),
.O5(CLBLM_L_X10Y115_SLICE_X12Y115_BO5),
.O6(CLBLM_L_X10Y115_SLICE_X12Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0afa0afa0)
  ) CLBLM_L_X10Y115_SLICE_X12Y115_ALUT (
.I0(CLBLM_R_X11Y116_SLICE_X14Y116_AQ),
.I1(1'b1),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y115_SLICE_X9Y115_A5Q),
.I4(1'b1),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X10Y115_SLICE_X12Y115_AO5),
.O6(CLBLM_L_X10Y115_SLICE_X12Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y115_SLICE_X13Y115_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y115_SLICE_X13Y115_AO6),
.Q(CLBLM_L_X10Y115_SLICE_X13Y115_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y115_SLICE_X13Y115_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y115_SLICE_X13Y115_BO6),
.Q(CLBLM_L_X10Y115_SLICE_X13Y115_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y115_SLICE_X13Y115_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y115_SLICE_X13Y115_CO6),
.Q(CLBLM_L_X10Y115_SLICE_X13Y115_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffeffff33330000)
  ) CLBLM_L_X10Y115_SLICE_X13Y115_DLUT (
.I0(CLBLM_R_X11Y110_SLICE_X15Y110_BQ),
.I1(RIOB33_X105Y121_IOB_X1Y121_I),
.I2(CLBLM_R_X11Y115_SLICE_X15Y115_AQ),
.I3(CLBLM_L_X12Y110_SLICE_X17Y110_CQ),
.I4(CLBLM_R_X11Y113_SLICE_X14Y113_CQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y115_SLICE_X13Y115_DO5),
.O6(CLBLM_L_X10Y115_SLICE_X13Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefefefa54545450)
  ) CLBLM_L_X10Y115_SLICE_X13Y115_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y117_SLICE_X13Y117_AO5),
.I2(CLBLM_L_X10Y116_SLICE_X13Y116_DO6),
.I3(CLBLM_L_X10Y113_SLICE_X13Y113_CQ),
.I4(CLBLM_R_X5Y108_SLICE_X6Y108_BO6),
.I5(CLBLM_L_X10Y114_SLICE_X13Y114_CQ),
.O5(CLBLM_L_X10Y115_SLICE_X13Y115_CO5),
.O6(CLBLM_L_X10Y115_SLICE_X13Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefe0e0ef0f00000)
  ) CLBLM_L_X10Y115_SLICE_X13Y115_BLUT (
.I0(CLBLM_L_X12Y113_SLICE_X17Y113_DO6),
.I1(CLBLM_L_X10Y115_SLICE_X13Y115_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(CLBLM_R_X7Y117_SLICE_X9Y117_A5Q),
.I5(CLBLM_R_X7Y115_SLICE_X9Y115_DO6),
.O5(CLBLM_L_X10Y115_SLICE_X13Y115_BO5),
.O6(CLBLM_L_X10Y115_SLICE_X13Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heefaeefaeefaeeaa)
  ) CLBLM_L_X10Y115_SLICE_X13Y115_ALUT (
.I0(CLBLM_R_X7Y112_SLICE_X9Y112_DO6),
.I1(CLBLM_R_X5Y114_SLICE_X7Y114_BQ),
.I2(CLBLM_L_X10Y115_SLICE_X13Y115_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.O5(CLBLM_L_X10Y115_SLICE_X13Y115_AO5),
.O6(CLBLM_L_X10Y115_SLICE_X13Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y116_SLICE_X12Y116_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y116_SLICE_X12Y116_AO6),
.Q(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y116_SLICE_X12Y116_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y116_SLICE_X12Y116_BO6),
.Q(CLBLM_L_X10Y116_SLICE_X12Y116_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y116_SLICE_X12Y116_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y116_SLICE_X12Y116_CO6),
.Q(CLBLM_L_X10Y116_SLICE_X12Y116_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00cd00cd0000fffe)
  ) CLBLM_L_X10Y116_SLICE_X12Y116_DLUT (
.I0(CLBLM_L_X10Y119_SLICE_X12Y119_AQ),
.I1(CLBLM_R_X7Y114_SLICE_X8Y114_A5Q),
.I2(CLBLM_R_X7Y118_SLICE_X8Y118_CQ),
.I3(CLBLM_L_X8Y118_SLICE_X10Y118_AQ),
.I4(CLBLM_L_X10Y117_SLICE_X13Y117_CO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y116_SLICE_X12Y116_DO5),
.O6(CLBLM_L_X10Y116_SLICE_X12Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hafaa0500efea4540)
  ) CLBLM_L_X10Y116_SLICE_X12Y116_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y116_SLICE_X12Y116_CQ),
.I2(CLBLM_R_X7Y118_SLICE_X8Y118_DO6),
.I3(CLBLM_L_X8Y116_SLICE_X10Y116_CQ),
.I4(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.I5(CLBLM_L_X10Y117_SLICE_X13Y117_AO5),
.O5(CLBLM_L_X10Y116_SLICE_X12Y116_CO5),
.O6(CLBLM_L_X10Y116_SLICE_X12Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf505f000fd0df808)
  ) CLBLM_L_X10Y116_SLICE_X12Y116_BLUT (
.I0(CLBLM_R_X7Y118_SLICE_X8Y118_DO6),
.I1(CLBLM_L_X10Y116_SLICE_X12Y116_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X5Y115_SLICE_X7Y115_BQ),
.I4(CLBLM_L_X10Y116_SLICE_X12Y116_CQ),
.I5(CLBLM_L_X10Y117_SLICE_X13Y117_AO5),
.O5(CLBLM_L_X10Y116_SLICE_X12Y116_BO5),
.O6(CLBLM_L_X10Y116_SLICE_X12Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hddcc1100fdec3120)
  ) CLBLM_L_X10Y116_SLICE_X12Y116_ALUT (
.I0(CLBLM_R_X7Y118_SLICE_X8Y118_DO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I3(CLBLM_R_X11Y116_SLICE_X14Y116_AQ),
.I4(CLBLM_R_X7Y111_SLICE_X9Y111_AQ),
.I5(CLBLM_L_X10Y117_SLICE_X13Y117_AO5),
.O5(CLBLM_L_X10Y116_SLICE_X12Y116_AO5),
.O6(CLBLM_L_X10Y116_SLICE_X12Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y116_SLICE_X13Y116_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y116_SLICE_X13Y116_AO6),
.Q(CLBLM_L_X10Y116_SLICE_X13Y116_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y116_SLICE_X13Y116_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y116_SLICE_X13Y116_BO6),
.Q(CLBLM_L_X10Y116_SLICE_X13Y116_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y116_SLICE_X13Y116_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y116_SLICE_X13Y116_CO6),
.Q(CLBLM_L_X10Y116_SLICE_X13Y116_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3232cccc3232ccc8)
  ) CLBLM_L_X10Y116_SLICE_X13Y116_DLUT (
.I0(CLBLM_L_X10Y119_SLICE_X12Y119_AQ),
.I1(CLBLM_L_X10Y115_SLICE_X13Y115_CQ),
.I2(CLBLM_R_X7Y118_SLICE_X8Y118_CQ),
.I3(CLBLM_R_X7Y114_SLICE_X8Y114_A5Q),
.I4(CLBLM_R_X7Y118_SLICE_X9Y118_BO5),
.I5(CLBLM_L_X8Y118_SLICE_X10Y118_AQ),
.O5(CLBLM_L_X10Y116_SLICE_X13Y116_DO5),
.O6(CLBLM_L_X10Y116_SLICE_X13Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000ff90ff90)
  ) CLBLM_L_X10Y116_SLICE_X13Y116_CLUT (
.I0(CLBLM_R_X11Y117_SLICE_X14Y117_AO6),
.I1(CLBLM_L_X10Y116_SLICE_X13Y116_CQ),
.I2(CLBLM_L_X10Y116_SLICE_X12Y116_DO5),
.I3(CLBLM_L_X10Y118_SLICE_X13Y118_CO6),
.I4(CLBLM_L_X12Y110_SLICE_X17Y110_DQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y116_SLICE_X13Y116_CO5),
.O6(CLBLM_L_X10Y116_SLICE_X13Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff00ffff540054)
  ) CLBLM_L_X10Y116_SLICE_X13Y116_BLUT (
.I0(CLBLM_R_X7Y118_SLICE_X8Y118_DO6),
.I1(CLBLM_L_X10Y116_SLICE_X13Y116_BQ),
.I2(CLBLM_L_X10Y116_SLICE_X13Y116_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLL_L_X4Y114_SLICE_X4Y114_BQ),
.I5(CLBLM_L_X10Y117_SLICE_X13Y117_AO5),
.O5(CLBLM_L_X10Y116_SLICE_X13Y116_BO5),
.O6(CLBLM_L_X10Y116_SLICE_X13Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hddccfdec11003120)
  ) CLBLM_L_X10Y116_SLICE_X13Y116_ALUT (
.I0(CLBLM_R_X7Y118_SLICE_X8Y118_DO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y116_SLICE_X13Y116_AQ),
.I3(CLBLM_L_X10Y116_SLICE_X12Y116_BQ),
.I4(CLBLM_L_X10Y117_SLICE_X13Y117_AO5),
.I5(CLBLM_L_X10Y111_SLICE_X13Y111_CQ),
.O5(CLBLM_L_X10Y116_SLICE_X13Y116_AO5),
.O6(CLBLM_L_X10Y116_SLICE_X13Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y117_SLICE_X12Y117_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y117_SLICE_X12Y117_AO5),
.Q(CLBLM_L_X10Y117_SLICE_X12Y117_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y117_SLICE_X12Y117_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y117_SLICE_X12Y117_AO6),
.Q(CLBLM_L_X10Y117_SLICE_X12Y117_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y117_SLICE_X12Y117_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y117_SLICE_X12Y117_BO6),
.Q(CLBLM_L_X10Y117_SLICE_X12Y117_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f3f3f3f3f3f2f3f)
  ) CLBLM_L_X10Y117_SLICE_X12Y117_DLUT (
.I0(CLBLM_L_X10Y119_SLICE_X12Y119_AQ),
.I1(CLBLM_R_X11Y117_SLICE_X15Y117_AQ),
.I2(CLBLM_R_X7Y118_SLICE_X9Y118_BO5),
.I3(CLBLM_L_X8Y118_SLICE_X10Y118_AQ),
.I4(CLBLM_R_X7Y118_SLICE_X8Y118_CQ),
.I5(CLBLM_R_X7Y114_SLICE_X8Y114_A5Q),
.O5(CLBLM_L_X10Y117_SLICE_X12Y117_DO5),
.O6(CLBLM_L_X10Y117_SLICE_X12Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0004ffff4444)
  ) CLBLM_L_X10Y117_SLICE_X12Y117_CLUT (
.I0(CLBLM_L_X8Y116_SLICE_X11Y116_CO6),
.I1(CLBLM_L_X8Y116_SLICE_X10Y116_CQ),
.I2(CLBLM_L_X10Y116_SLICE_X13Y116_CQ),
.I3(CLBLM_L_X10Y119_SLICE_X12Y119_CO6),
.I4(CLBLM_L_X10Y117_SLICE_X12Y117_DO6),
.I5(CLBLM_L_X10Y119_SLICE_X12Y119_BO6),
.O5(CLBLM_L_X10Y117_SLICE_X12Y117_CO5),
.O6(CLBLM_L_X10Y117_SLICE_X12Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfb0bfa0afe0efa0a)
  ) CLBLM_L_X10Y117_SLICE_X12Y117_BLUT (
.I0(CLBLM_L_X10Y118_SLICE_X13Y118_CO6),
.I1(CLBLM_L_X10Y117_SLICE_X12Y117_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y115_SLICE_X8Y115_DQ),
.I4(CLBLM_L_X10Y116_SLICE_X12Y116_DO5),
.I5(CLBLM_L_X10Y117_SLICE_X12Y117_CO6),
.O5(CLBLM_L_X10Y117_SLICE_X12Y117_BO5),
.O6(CLBLM_L_X10Y117_SLICE_X12Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa0afa0acacacaca)
  ) CLBLM_L_X10Y117_SLICE_X12Y117_ALUT (
.I0(RIOB33_X105Y143_IOB_X1Y144_I),
.I1(CLBLM_L_X10Y116_SLICE_X13Y116_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X3Y114_SLICE_X2Y114_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y117_SLICE_X12Y117_AO5),
.O6(CLBLM_L_X10Y117_SLICE_X12Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff77ffffffffffff)
  ) CLBLM_L_X10Y117_SLICE_X13Y117_DLUT (
.I0(CLBLM_R_X11Y116_SLICE_X14Y116_BQ),
.I1(CLBLM_L_X12Y117_SLICE_X17Y117_BQ),
.I2(1'b1),
.I3(CLBLM_R_X11Y117_SLICE_X14Y117_DO6),
.I4(CLBLM_L_X10Y116_SLICE_X13Y116_CQ),
.I5(CLBLM_L_X10Y117_SLICE_X12Y117_BQ),
.O5(CLBLM_L_X10Y117_SLICE_X13Y117_DO5),
.O6(CLBLM_L_X10Y117_SLICE_X13Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h005080d000008080)
  ) CLBLM_L_X10Y117_SLICE_X13Y117_CLUT (
.I0(CLBLM_R_X11Y117_SLICE_X15Y117_DQ),
.I1(CLBLM_R_X11Y117_SLICE_X15Y117_CQ),
.I2(CLBLM_R_X7Y118_SLICE_X9Y118_CO5),
.I3(CLBLM_L_X10Y119_SLICE_X12Y119_CO6),
.I4(CLBLM_L_X10Y117_SLICE_X13Y117_DO6),
.I5(CLBLM_L_X10Y117_SLICE_X13Y117_BO5),
.O5(CLBLM_L_X10Y117_SLICE_X13Y117_CO5),
.O6(CLBLM_L_X10Y117_SLICE_X13Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffa00010001)
  ) CLBLM_L_X10Y117_SLICE_X13Y117_BLUT (
.I0(CLBLM_L_X10Y116_SLICE_X13Y116_CQ),
.I1(CLBLM_R_X11Y117_SLICE_X15Y117_CQ),
.I2(CLBLM_L_X12Y117_SLICE_X17Y117_BQ),
.I3(CLBLM_L_X10Y117_SLICE_X12Y117_BQ),
.I4(CLBLM_L_X10Y119_SLICE_X12Y119_CO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y117_SLICE_X13Y117_BO5),
.O6(CLBLM_L_X10Y117_SLICE_X13Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000020000000003)
  ) CLBLM_L_X10Y117_SLICE_X13Y117_ALUT (
.I0(CLBLM_R_X7Y118_SLICE_X9Y118_BO5),
.I1(CLBLM_R_X7Y114_SLICE_X8Y114_A5Q),
.I2(CLBLM_R_X7Y118_SLICE_X8Y118_CQ),
.I3(CLBLM_L_X8Y118_SLICE_X10Y118_AQ),
.I4(CLBLM_L_X10Y119_SLICE_X12Y119_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y117_SLICE_X13Y117_AO5),
.O6(CLBLM_L_X10Y117_SLICE_X13Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y118_SLICE_X12Y118_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y118_SLICE_X12Y118_AO6),
.Q(CLBLM_L_X10Y118_SLICE_X12Y118_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y118_SLICE_X12Y118_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y118_SLICE_X12Y118_BO6),
.Q(CLBLM_L_X10Y118_SLICE_X12Y118_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000febfffff)
  ) CLBLM_L_X10Y118_SLICE_X12Y118_DLUT (
.I0(CLBLM_L_X8Y116_SLICE_X11Y116_CO6),
.I1(CLBLM_L_X10Y118_SLICE_X12Y118_AQ),
.I2(CLBLM_L_X10Y118_SLICE_X13Y118_AQ),
.I3(CLBLM_L_X8Y118_SLICE_X10Y118_CO5),
.I4(CLBLM_L_X8Y116_SLICE_X10Y116_BQ),
.I5(CLBLM_L_X10Y117_SLICE_X12Y117_DO6),
.O5(CLBLM_L_X10Y118_SLICE_X12Y118_DO5),
.O6(CLBLM_L_X10Y118_SLICE_X12Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc69cc33cc33cc33)
  ) CLBLM_L_X10Y118_SLICE_X12Y118_CLUT (
.I0(CLBLM_L_X10Y118_SLICE_X13Y118_AQ),
.I1(CLBLM_L_X10Y118_SLICE_X12Y118_AQ),
.I2(CLBLM_L_X8Y118_SLICE_X10Y118_CO5),
.I3(CLBLM_L_X10Y117_SLICE_X12Y117_DO6),
.I4(CLBLM_L_X8Y117_SLICE_X10Y117_AQ),
.I5(CLBLM_R_X7Y118_SLICE_X9Y118_CO5),
.O5(CLBLM_L_X10Y118_SLICE_X12Y118_CO5),
.O6(CLBLM_L_X10Y118_SLICE_X12Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00f8f8f4f4)
  ) CLBLM_L_X10Y118_SLICE_X12Y118_BLUT (
.I0(CLBLM_L_X10Y118_SLICE_X12Y118_DO6),
.I1(CLBLM_L_X10Y116_SLICE_X12Y116_DO5),
.I2(CLBLM_L_X10Y118_SLICE_X13Y118_CO6),
.I3(CLBLM_L_X8Y118_SLICE_X10Y118_BQ),
.I4(CLBLM_L_X10Y118_SLICE_X12Y118_BQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y118_SLICE_X12Y118_BO5),
.O6(CLBLM_L_X10Y118_SLICE_X12Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfc3030fffc3330)
  ) CLBLM_L_X10Y118_SLICE_X12Y118_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y118_SLICE_X13Y118_CO6),
.I3(CLBLM_L_X10Y116_SLICE_X12Y116_DO5),
.I4(CLBLM_R_X7Y105_SLICE_X8Y105_AQ),
.I5(CLBLM_L_X10Y118_SLICE_X12Y118_CO6),
.O5(CLBLM_L_X10Y118_SLICE_X12Y118_AO5),
.O6(CLBLM_L_X10Y118_SLICE_X12Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y118_SLICE_X13Y118_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y118_SLICE_X13Y118_AO6),
.Q(CLBLM_L_X10Y118_SLICE_X13Y118_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h22dd000033cc0000)
  ) CLBLM_L_X10Y118_SLICE_X13Y118_DLUT (
.I0(CLBLM_L_X8Y116_SLICE_X11Y116_CO6),
.I1(CLBLM_L_X10Y117_SLICE_X12Y117_DO6),
.I2(1'b1),
.I3(CLBLM_L_X10Y118_SLICE_X13Y118_AQ),
.I4(CLBLM_L_X10Y116_SLICE_X12Y116_DO5),
.I5(CLBLM_L_X10Y116_SLICE_X13Y116_BQ),
.O5(CLBLM_L_X10Y118_SLICE_X13Y118_DO5),
.O6(CLBLM_L_X10Y118_SLICE_X13Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcb004100ca00ca00)
  ) CLBLM_L_X10Y118_SLICE_X13Y118_CLUT (
.I0(CLBLM_L_X8Y118_SLICE_X10Y118_AQ),
.I1(CLBLM_L_X10Y119_SLICE_X12Y119_AQ),
.I2(CLBLM_R_X7Y118_SLICE_X8Y118_CQ),
.I3(CLBLM_L_X10Y117_SLICE_X13Y117_CO6),
.I4(CLBLM_R_X11Y117_SLICE_X15Y117_AQ),
.I5(CLBLM_R_X7Y114_SLICE_X8Y114_A5Q),
.O5(CLBLM_L_X10Y118_SLICE_X13Y118_CO5),
.O6(CLBLM_L_X10Y118_SLICE_X13Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0033233333333333)
  ) CLBLM_L_X10Y118_SLICE_X13Y118_BLUT (
.I0(CLBLM_L_X10Y119_SLICE_X12Y119_BO6),
.I1(CLBLM_L_X10Y117_SLICE_X12Y117_DO6),
.I2(CLBLM_L_X10Y117_SLICE_X12Y117_BQ),
.I3(CLBLM_R_X7Y118_SLICE_X9Y118_CO5),
.I4(CLBLM_L_X10Y119_SLICE_X13Y119_AO6),
.I5(CLBLM_L_X10Y116_SLICE_X12Y116_CQ),
.O5(CLBLM_L_X10Y118_SLICE_X13Y118_BO5),
.O6(CLBLM_L_X10Y118_SLICE_X13Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff00ffffaa00aa)
  ) CLBLM_L_X10Y118_SLICE_X13Y118_ALUT (
.I0(CLBLM_L_X10Y118_SLICE_X13Y118_DO6),
.I1(1'b1),
.I2(1'b1),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y113_SLICE_X13Y113_DQ),
.I5(CLBLM_L_X10Y118_SLICE_X13Y118_CO6),
.O5(CLBLM_L_X10Y118_SLICE_X13Y118_AO5),
.O6(CLBLM_L_X10Y118_SLICE_X13Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y119_SLICE_X12Y119_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y119_SLICE_X12Y119_AO6),
.Q(CLBLM_L_X10Y119_SLICE_X12Y119_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y119_SLICE_X12Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y119_SLICE_X12Y119_DO5),
.O6(CLBLM_L_X10Y119_SLICE_X12Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffffbb)
  ) CLBLM_L_X10Y119_SLICE_X12Y119_CLUT (
.I0(CLBLM_R_X11Y116_SLICE_X14Y116_BQ),
.I1(CLBLM_L_X8Y118_SLICE_X10Y118_CO5),
.I2(1'b1),
.I3(CLBLM_L_X10Y118_SLICE_X12Y118_AQ),
.I4(CLBLM_L_X10Y118_SLICE_X13Y118_AQ),
.I5(CLBLM_L_X10Y118_SLICE_X12Y118_BQ),
.O5(CLBLM_L_X10Y119_SLICE_X12Y119_CO5),
.O6(CLBLM_L_X10Y119_SLICE_X12Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff7fffffff)
  ) CLBLM_L_X10Y119_SLICE_X12Y119_BLUT (
.I0(CLBLM_L_X10Y118_SLICE_X12Y118_AQ),
.I1(CLBLM_L_X10Y116_SLICE_X13Y116_CQ),
.I2(CLBLM_L_X10Y118_SLICE_X13Y118_AQ),
.I3(CLBLM_L_X10Y118_SLICE_X12Y118_BQ),
.I4(CLBLM_R_X11Y116_SLICE_X14Y116_BQ),
.I5(CLBLM_L_X8Y118_SLICE_X10Y118_CO5),
.O5(CLBLM_L_X10Y119_SLICE_X12Y119_BO5),
.O6(CLBLM_L_X10Y119_SLICE_X12Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd8d8888d88d8888)
  ) CLBLM_L_X10Y119_SLICE_X12Y119_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y114_SLICE_X12Y114_AQ),
.I2(CLBLM_L_X10Y119_SLICE_X12Y119_AQ),
.I3(CLBLM_L_X8Y118_SLICE_X10Y118_DO6),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(CLBLM_L_X10Y117_SLICE_X13Y117_AO5),
.O5(CLBLM_L_X10Y119_SLICE_X12Y119_AO5),
.O6(CLBLM_L_X10Y119_SLICE_X12Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y119_SLICE_X13Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y119_SLICE_X13Y119_DO5),
.O6(CLBLM_L_X10Y119_SLICE_X13Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y119_SLICE_X13Y119_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y119_SLICE_X13Y119_CO5),
.O6(CLBLM_L_X10Y119_SLICE_X13Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y119_SLICE_X13Y119_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y119_SLICE_X13Y119_BO5),
.O6(CLBLM_L_X10Y119_SLICE_X13Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0003000300030003)
  ) CLBLM_L_X10Y119_SLICE_X13Y119_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y117_SLICE_X12Y117_BQ),
.I2(CLBLM_L_X10Y119_SLICE_X12Y119_CO6),
.I3(CLBLM_L_X10Y116_SLICE_X13Y116_CQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y119_SLICE_X13Y119_AO5),
.O6(CLBLM_L_X10Y119_SLICE_X13Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y148_SLICE_X12Y148_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y148_SLICE_X12Y148_DO5),
.O6(CLBLM_L_X10Y148_SLICE_X12Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y148_SLICE_X12Y148_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y148_SLICE_X12Y148_CO5),
.O6(CLBLM_L_X10Y148_SLICE_X12Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y148_SLICE_X12Y148_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y148_SLICE_X12Y148_BO5),
.O6(CLBLM_L_X10Y148_SLICE_X12Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555555555555555)
  ) CLBLM_L_X10Y148_SLICE_X12Y148_ALUT (
.I0(CLBLM_L_X10Y110_SLICE_X12Y110_B5Q),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y148_SLICE_X12Y148_AO5),
.O6(CLBLM_L_X10Y148_SLICE_X12Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y148_SLICE_X13Y148_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y148_SLICE_X13Y148_DO5),
.O6(CLBLM_L_X10Y148_SLICE_X13Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y148_SLICE_X13Y148_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y148_SLICE_X13Y148_CO5),
.O6(CLBLM_L_X10Y148_SLICE_X13Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y148_SLICE_X13Y148_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y148_SLICE_X13Y148_BO5),
.O6(CLBLM_L_X10Y148_SLICE_X13Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y148_SLICE_X13Y148_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y148_SLICE_X13Y148_AO5),
.O6(CLBLM_L_X10Y148_SLICE_X13Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y105_SLICE_X16Y105_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y105_SLICE_X16Y105_AO6),
.Q(CLBLM_L_X12Y105_SLICE_X16Y105_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y105_SLICE_X16Y105_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y105_SLICE_X16Y105_DO5),
.O6(CLBLM_L_X12Y105_SLICE_X16Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0fbf0fff30003000)
  ) CLBLM_L_X12Y105_SLICE_X16Y105_CLUT (
.I0(CLBLM_R_X13Y108_SLICE_X18Y108_BO5),
.I1(CLBLM_L_X12Y105_SLICE_X16Y105_AQ),
.I2(CLBLM_R_X11Y106_SLICE_X15Y106_DO5),
.I3(CLBLM_R_X11Y105_SLICE_X15Y105_BQ),
.I4(CLBLM_L_X12Y107_SLICE_X17Y107_BQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y105_SLICE_X16Y105_CO5),
.O6(CLBLM_L_X12Y105_SLICE_X16Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000500040000)
  ) CLBLM_L_X12Y105_SLICE_X16Y105_BLUT (
.I0(CLBLM_R_X13Y109_SLICE_X19Y109_BQ),
.I1(CLBLM_R_X11Y106_SLICE_X15Y106_DO5),
.I2(CLBLM_L_X12Y105_SLICE_X16Y105_AQ),
.I3(CLBLM_R_X13Y113_SLICE_X18Y113_BQ),
.I4(CLBLM_L_X12Y107_SLICE_X17Y107_BQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y105_SLICE_X16Y105_BO5),
.O6(CLBLM_L_X12Y105_SLICE_X16Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff120012ff030003)
  ) CLBLM_L_X12Y105_SLICE_X16Y105_ALUT (
.I0(CLBLM_L_X12Y107_SLICE_X17Y107_DO6),
.I1(RIOB33_X105Y121_IOB_X1Y121_I),
.I2(CLBLM_L_X12Y105_SLICE_X16Y105_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y106_SLICE_X8Y106_CQ),
.I5(CLBLM_L_X12Y105_SLICE_X16Y105_CO6),
.O5(CLBLM_L_X12Y105_SLICE_X16Y105_AO5),
.O6(CLBLM_L_X12Y105_SLICE_X16Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y105_SLICE_X17Y105_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y105_SLICE_X17Y105_DO5),
.O6(CLBLM_L_X12Y105_SLICE_X17Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h33323333ffffffff)
  ) CLBLM_L_X12Y105_SLICE_X17Y105_CLUT (
.I0(CLBLM_L_X12Y105_SLICE_X16Y105_AQ),
.I1(CLBLM_R_X11Y105_SLICE_X15Y105_BQ),
.I2(CLBLM_R_X13Y109_SLICE_X19Y109_BQ),
.I3(CLBLM_R_X13Y113_SLICE_X18Y113_BQ),
.I4(CLBLM_L_X12Y107_SLICE_X17Y107_BQ),
.I5(CLBLM_R_X11Y106_SLICE_X15Y106_DO5),
.O5(CLBLM_L_X12Y105_SLICE_X17Y105_CO5),
.O6(CLBLM_L_X12Y105_SLICE_X17Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hd033dd33cc88cc88)
  ) CLBLM_L_X12Y105_SLICE_X17Y105_BLUT (
.I0(CLBLM_R_X13Y109_SLICE_X19Y109_BQ),
.I1(CLBLM_R_X13Y113_SLICE_X18Y113_BQ),
.I2(CLBLM_R_X11Y105_SLICE_X15Y105_BQ),
.I3(CLBLM_L_X12Y107_SLICE_X17Y107_BQ),
.I4(CLBLM_L_X12Y105_SLICE_X16Y105_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y105_SLICE_X17Y105_BO5),
.O6(CLBLM_L_X12Y105_SLICE_X17Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000555503ff13ff)
  ) CLBLM_L_X12Y105_SLICE_X17Y105_ALUT (
.I0(CLBLM_R_X13Y109_SLICE_X19Y109_BQ),
.I1(CLBLM_L_X12Y107_SLICE_X17Y107_DO5),
.I2(CLBLM_R_X11Y105_SLICE_X14Y105_DQ),
.I3(CLBLM_R_X11Y106_SLICE_X15Y106_DO5),
.I4(CLBLM_R_X13Y113_SLICE_X18Y113_BQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y105_SLICE_X17Y105_AO5),
.O6(CLBLM_L_X12Y105_SLICE_X17Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y106_SLICE_X16Y106_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y106_SLICE_X16Y106_AO6),
.Q(CLBLM_L_X12Y106_SLICE_X16Y106_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f4f1f0f0f0f0f0)
  ) CLBLM_L_X12Y106_SLICE_X16Y106_DLUT (
.I0(CLBLM_L_X12Y105_SLICE_X17Y105_AO5),
.I1(CLBLM_R_X13Y108_SLICE_X19Y108_BQ),
.I2(CLBLM_L_X12Y105_SLICE_X17Y105_CO6),
.I3(CLBLM_L_X12Y105_SLICE_X17Y105_BO5),
.I4(CLBLM_L_X12Y108_SLICE_X16Y108_BQ),
.I5(CLBLM_R_X11Y105_SLICE_X15Y105_CQ),
.O5(CLBLM_L_X12Y106_SLICE_X16Y106_DO5),
.O6(CLBLM_L_X12Y106_SLICE_X16Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h55555555aa56aaaa)
  ) CLBLM_L_X12Y106_SLICE_X16Y106_CLUT (
.I0(CLBLM_L_X12Y107_SLICE_X16Y107_AQ),
.I1(CLBLM_L_X12Y106_SLICE_X17Y106_CO6),
.I2(CLBLM_L_X12Y106_SLICE_X17Y106_DO6),
.I3(CLBLM_L_X12Y105_SLICE_X17Y105_AO5),
.I4(CLBLM_R_X11Y106_SLICE_X14Y106_CQ),
.I5(CLBLM_L_X12Y105_SLICE_X17Y105_CO6),
.O5(CLBLM_L_X12Y106_SLICE_X16Y106_CO5),
.O6(CLBLM_L_X12Y106_SLICE_X16Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5a5a595a5a5a565a)
  ) CLBLM_L_X12Y106_SLICE_X16Y106_BLUT (
.I0(CLBLM_L_X12Y108_SLICE_X16Y108_BQ),
.I1(CLBLM_R_X13Y108_SLICE_X19Y108_BQ),
.I2(CLBLM_L_X12Y105_SLICE_X17Y105_CO6),
.I3(CLBLM_L_X12Y108_SLICE_X17Y108_BQ),
.I4(CLBLM_L_X12Y105_SLICE_X17Y105_AO5),
.I5(CLBLM_L_X12Y105_SLICE_X17Y105_BO5),
.O5(CLBLM_L_X12Y106_SLICE_X16Y106_BO5),
.O6(CLBLM_L_X12Y106_SLICE_X16Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00ccf0cc00ccf5)
  ) CLBLM_L_X12Y106_SLICE_X16Y106_ALUT (
.I0(CLBLM_R_X13Y109_SLICE_X19Y109_BQ),
.I1(CLBLM_R_X11Y105_SLICE_X15Y105_BQ),
.I2(CLBLM_L_X12Y105_SLICE_X16Y105_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X12Y107_SLICE_X17Y107_BQ),
.I5(CLBLM_R_X13Y113_SLICE_X18Y113_BQ),
.O5(CLBLM_L_X12Y106_SLICE_X16Y106_AO5),
.O6(CLBLM_L_X12Y106_SLICE_X16Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y106_SLICE_X17Y106_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y106_SLICE_X17Y106_AO6),
.Q(CLBLM_L_X12Y106_SLICE_X17Y106_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h2000000000000000)
  ) CLBLM_L_X12Y106_SLICE_X17Y106_DLUT (
.I0(CLBLM_R_X13Y107_SLICE_X19Y107_AQ),
.I1(CLBLM_L_X12Y105_SLICE_X17Y105_BO5),
.I2(CLBLM_L_X12Y108_SLICE_X16Y108_BQ),
.I3(CLBLM_R_X13Y108_SLICE_X19Y108_BQ),
.I4(CLBLM_L_X12Y107_SLICE_X16Y107_BQ),
.I5(CLBLM_R_X13Y107_SLICE_X19Y107_BQ),
.O5(CLBLM_L_X12Y106_SLICE_X17Y106_DO5),
.O6(CLBLM_L_X12Y106_SLICE_X17Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000004)
  ) CLBLM_L_X12Y106_SLICE_X17Y106_CLUT (
.I0(CLBLM_R_X13Y107_SLICE_X19Y107_AQ),
.I1(CLBLM_L_X12Y105_SLICE_X17Y105_BO5),
.I2(CLBLM_L_X12Y108_SLICE_X16Y108_BQ),
.I3(CLBLM_R_X13Y108_SLICE_X19Y108_BQ),
.I4(CLBLM_L_X12Y107_SLICE_X16Y107_BQ),
.I5(CLBLM_R_X13Y107_SLICE_X19Y107_BQ),
.O5(CLBLM_L_X12Y106_SLICE_X17Y106_CO5),
.O6(CLBLM_L_X12Y106_SLICE_X17Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff08ff0cff08ff00)
  ) CLBLM_L_X12Y106_SLICE_X17Y106_BLUT (
.I0(CLBLM_L_X12Y106_SLICE_X17Y106_DO6),
.I1(CLBLM_L_X12Y107_SLICE_X16Y107_CQ),
.I2(CLBLM_L_X12Y105_SLICE_X17Y105_AO5),
.I3(CLBLM_L_X12Y105_SLICE_X17Y105_CO6),
.I4(CLBLM_L_X12Y107_SLICE_X16Y107_AQ),
.I5(CLBLM_L_X12Y106_SLICE_X17Y106_CO6),
.O5(CLBLM_L_X12Y106_SLICE_X17Y106_BO5),
.O6(CLBLM_L_X12Y106_SLICE_X17Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccfc0030ccfc0030)
  ) CLBLM_L_X12Y106_SLICE_X17Y106_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X12Y106_SLICE_X17Y106_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X13Y107_SLICE_X18Y107_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y106_SLICE_X17Y106_AO5),
.O6(CLBLM_L_X12Y106_SLICE_X17Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y107_SLICE_X16Y107_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y107_SLICE_X16Y107_AO6),
.Q(CLBLM_L_X12Y107_SLICE_X16Y107_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y107_SLICE_X16Y107_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y107_SLICE_X16Y107_BO6),
.Q(CLBLM_L_X12Y107_SLICE_X16Y107_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y107_SLICE_X16Y107_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y107_SLICE_X16Y107_CO6),
.Q(CLBLM_L_X12Y107_SLICE_X16Y107_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y107_SLICE_X16Y107_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y107_SLICE_X16Y107_DO6),
.Q(CLBLM_L_X12Y107_SLICE_X16Y107_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff00003b083b08)
  ) CLBLM_L_X12Y107_SLICE_X16Y107_DLUT (
.I0(CLBLM_L_X12Y107_SLICE_X16Y107_DQ),
.I1(CLBLM_L_X12Y105_SLICE_X16Y105_CO5),
.I2(CLBLM_L_X12Y105_SLICE_X16Y105_BO6),
.I3(CLBLM_L_X12Y108_SLICE_X16Y108_CQ),
.I4(CLBLM_L_X10Y110_SLICE_X13Y110_DQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X12Y107_SLICE_X16Y107_DO5),
.O6(CLBLM_L_X12Y107_SLICE_X16Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf505fd0df000f808)
  ) CLBLM_L_X12Y107_SLICE_X16Y107_CLUT (
.I0(CLBLM_L_X12Y105_SLICE_X16Y105_CO5),
.I1(CLBLM_L_X12Y107_SLICE_X16Y107_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y113_SLICE_X10Y113_CQ),
.I4(CLBLM_L_X12Y105_SLICE_X16Y105_BO6),
.I5(CLBLM_R_X11Y106_SLICE_X14Y106_CQ),
.O5(CLBLM_L_X12Y107_SLICE_X16Y107_CO5),
.O6(CLBLM_L_X12Y107_SLICE_X16Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000aaaaf3fc)
  ) CLBLM_L_X12Y107_SLICE_X16Y107_BLUT (
.I0(CLBLM_L_X10Y118_SLICE_X13Y118_AQ),
.I1(CLBLM_L_X12Y107_SLICE_X16Y107_BQ),
.I2(CLBLM_L_X12Y107_SLICE_X17Y107_CO5),
.I3(CLBLM_L_X12Y106_SLICE_X16Y106_DO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X12Y108_SLICE_X17Y108_CO5),
.O5(CLBLM_L_X12Y107_SLICE_X16Y107_BO5),
.O6(CLBLM_L_X12Y107_SLICE_X16Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000fffc00fc)
  ) CLBLM_L_X12Y107_SLICE_X16Y107_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X12Y106_SLICE_X16Y106_CO6),
.I2(CLBLM_L_X12Y107_SLICE_X17Y107_CO5),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y107_SLICE_X9Y107_BQ),
.I5(CLBLM_L_X12Y108_SLICE_X17Y108_CO5),
.O5(CLBLM_L_X12Y107_SLICE_X16Y107_AO5),
.O6(CLBLM_L_X12Y107_SLICE_X16Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y107_SLICE_X17Y107_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y107_SLICE_X17Y107_AO6),
.Q(CLBLM_L_X12Y107_SLICE_X17Y107_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y107_SLICE_X17Y107_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y107_SLICE_X17Y107_BO6),
.Q(CLBLM_L_X12Y107_SLICE_X17Y107_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000200030003000)
  ) CLBLM_L_X12Y107_SLICE_X17Y107_DLUT (
.I0(CLBLM_R_X13Y108_SLICE_X18Y108_BO6),
.I1(CLBLM_R_X11Y105_SLICE_X15Y105_BQ),
.I2(CLBLM_L_X12Y107_SLICE_X17Y107_BQ),
.I3(CLBLM_L_X12Y105_SLICE_X16Y105_AQ),
.I4(CLBLM_L_X12Y107_SLICE_X17Y107_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y107_SLICE_X17Y107_DO5),
.O6(CLBLM_L_X12Y107_SLICE_X17Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h33000005c4a5f5a0)
  ) CLBLM_L_X12Y107_SLICE_X17Y107_CLUT (
.I0(CLBLM_R_X13Y113_SLICE_X18Y113_BQ),
.I1(CLBLM_R_X11Y105_SLICE_X15Y105_BQ),
.I2(CLBLM_R_X13Y109_SLICE_X19Y109_BQ),
.I3(CLBLM_L_X12Y107_SLICE_X17Y107_BQ),
.I4(CLBLM_L_X12Y105_SLICE_X16Y105_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y107_SLICE_X17Y107_CO5),
.O6(CLBLM_L_X12Y107_SLICE_X17Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0e4f5a0a0b1a0)
  ) CLBLM_L_X12Y107_SLICE_X17Y107_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X12Y105_SLICE_X17Y105_BO6),
.I2(CLBLM_R_X13Y113_SLICE_X18Y113_AQ),
.I3(CLBLM_R_X13Y108_SLICE_X18Y108_BO6),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(CLBLM_L_X12Y107_SLICE_X17Y107_BQ),
.O5(CLBLM_L_X12Y107_SLICE_X17Y107_BO5),
.O6(CLBLM_L_X12Y107_SLICE_X17Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00eaeaff00fafa)
  ) CLBLM_L_X12Y107_SLICE_X17Y107_ALUT (
.I0(CLBLM_L_X12Y107_SLICE_X17Y107_DO6),
.I1(CLBLM_L_X12Y108_SLICE_X17Y108_CO5),
.I2(CLBLM_L_X12Y107_SLICE_X17Y107_AQ),
.I3(CLBLM_L_X8Y109_SLICE_X10Y109_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X12Y107_SLICE_X17Y107_CO6),
.O5(CLBLM_L_X12Y107_SLICE_X17Y107_AO5),
.O6(CLBLM_L_X12Y107_SLICE_X17Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y108_SLICE_X16Y108_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y108_SLICE_X16Y108_AO6),
.Q(CLBLM_L_X12Y108_SLICE_X16Y108_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y108_SLICE_X16Y108_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y108_SLICE_X16Y108_BO6),
.Q(CLBLM_L_X12Y108_SLICE_X16Y108_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y108_SLICE_X16Y108_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y108_SLICE_X16Y108_CO6),
.Q(CLBLM_L_X12Y108_SLICE_X16Y108_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y108_SLICE_X16Y108_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y108_SLICE_X16Y108_DO6),
.Q(CLBLM_L_X12Y108_SLICE_X16Y108_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaccaaffaaccaafc)
  ) CLBLM_L_X12Y108_SLICE_X16Y108_DLUT (
.I0(CLBLM_L_X8Y116_SLICE_X10Y116_DQ),
.I1(CLBLM_L_X12Y105_SLICE_X16Y105_BO6),
.I2(CLBLM_L_X12Y108_SLICE_X16Y108_DQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X12Y105_SLICE_X16Y105_CO5),
.I5(CLBLM_R_X11Y108_SLICE_X14Y108_AQ),
.O5(CLBLM_L_X12Y108_SLICE_X16Y108_DO5),
.O6(CLBLM_L_X12Y108_SLICE_X16Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haeaeffaa04045500)
  ) CLBLM_L_X12Y108_SLICE_X16Y108_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X12Y108_SLICE_X16Y108_CQ),
.I2(CLBLM_L_X12Y105_SLICE_X16Y105_BO6),
.I3(CLBLM_R_X11Y105_SLICE_X15Y105_CQ),
.I4(CLBLM_L_X12Y105_SLICE_X16Y105_CO5),
.I5(CLBLM_R_X7Y109_SLICE_X9Y109_BQ),
.O5(CLBLM_L_X12Y108_SLICE_X16Y108_CO5),
.O6(CLBLM_L_X12Y108_SLICE_X16Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc0fcc0fcc0fcc00)
  ) CLBLM_L_X12Y108_SLICE_X16Y108_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X12Y112_SLICE_X16Y112_AQ),
.I2(CLBLM_L_X12Y108_SLICE_X17Y108_CO5),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X12Y106_SLICE_X16Y106_BO6),
.I5(CLBLM_L_X12Y107_SLICE_X17Y107_CO5),
.O5(CLBLM_L_X12Y108_SLICE_X16Y108_BO5),
.O6(CLBLM_L_X12Y108_SLICE_X16Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00ccaa000f0000)
  ) CLBLM_L_X12Y108_SLICE_X16Y108_ALUT (
.I0(CLBLM_L_X10Y115_SLICE_X12Y115_CQ),
.I1(CLBLM_L_X12Y109_SLICE_X17Y109_BQ),
.I2(CLBLM_R_X7Y115_SLICE_X8Y115_DQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_L_X12Y108_SLICE_X16Y108_AO5),
.O6(CLBLM_L_X12Y108_SLICE_X16Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y108_SLICE_X17Y108_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y108_SLICE_X17Y108_AO6),
.Q(CLBLM_L_X12Y108_SLICE_X17Y108_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y108_SLICE_X17Y108_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y108_SLICE_X17Y108_BO6),
.Q(CLBLM_L_X12Y108_SLICE_X17Y108_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3033303bffffffff)
  ) CLBLM_L_X12Y108_SLICE_X17Y108_DLUT (
.I0(CLBLM_R_X11Y105_SLICE_X15Y105_BQ),
.I1(CLBLM_L_X12Y107_SLICE_X17Y107_BQ),
.I2(CLBLM_L_X12Y105_SLICE_X16Y105_AQ),
.I3(CLBLM_R_X13Y113_SLICE_X18Y113_BQ),
.I4(CLBLM_R_X13Y109_SLICE_X19Y109_BQ),
.I5(CLBLM_L_X12Y109_SLICE_X17Y109_BQ),
.O5(CLBLM_L_X12Y108_SLICE_X17Y108_DO5),
.O6(CLBLM_L_X12Y108_SLICE_X17Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5050515100ff00fe)
  ) CLBLM_L_X12Y108_SLICE_X17Y108_CLUT (
.I0(CLBLM_L_X12Y107_SLICE_X17Y107_BQ),
.I1(CLBLM_R_X13Y113_SLICE_X18Y113_BQ),
.I2(CLBLM_L_X12Y105_SLICE_X16Y105_AQ),
.I3(CLBLM_R_X13Y108_SLICE_X18Y108_BO5),
.I4(CLBLM_R_X13Y109_SLICE_X19Y109_BQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y108_SLICE_X17Y108_CO5),
.O6(CLBLM_L_X12Y108_SLICE_X17Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfeeccee03220022)
  ) CLBLM_L_X12Y108_SLICE_X17Y108_BLUT (
.I0(CLBLM_L_X12Y108_SLICE_X16Y108_DQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X12Y105_SLICE_X16Y105_BO6),
.I3(CLBLM_L_X12Y105_SLICE_X16Y105_CO5),
.I4(CLBLM_L_X12Y108_SLICE_X17Y108_BQ),
.I5(CLBLM_L_X12Y109_SLICE_X17Y109_CQ),
.O5(CLBLM_L_X12Y108_SLICE_X17Y108_BO5),
.O6(CLBLM_L_X12Y108_SLICE_X17Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc50ff5000)
  ) CLBLM_L_X12Y108_SLICE_X17Y108_ALUT (
.I0(CLBLM_L_X12Y105_SLICE_X16Y105_BO6),
.I1(CLBLM_R_X7Y109_SLICE_X8Y109_BQ),
.I2(CLBLM_L_X12Y108_SLICE_X17Y108_AQ),
.I3(CLBLM_L_X12Y105_SLICE_X16Y105_CO5),
.I4(CLBLM_L_X12Y107_SLICE_X16Y107_CQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X12Y108_SLICE_X17Y108_AO5),
.O6(CLBLM_L_X12Y108_SLICE_X17Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y109_SLICE_X16Y109_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y109_SLICE_X16Y109_DO5),
.Q(CLBLM_L_X12Y109_SLICE_X16Y109_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y109_SLICE_X16Y109_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y109_SLICE_X16Y109_AO6),
.Q(CLBLM_L_X12Y109_SLICE_X16Y109_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y109_SLICE_X16Y109_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y109_SLICE_X16Y109_BO6),
.Q(CLBLM_L_X12Y109_SLICE_X16Y109_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y109_SLICE_X16Y109_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y109_SLICE_X16Y109_CO6),
.Q(CLBLM_L_X12Y109_SLICE_X16Y109_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y109_SLICE_X16Y109_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y109_SLICE_X16Y109_DO6),
.Q(CLBLM_L_X12Y109_SLICE_X16Y109_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc30fc30bbbb8888)
  ) CLBLM_L_X12Y109_SLICE_X16Y109_DLUT (
.I0(CLBLM_L_X12Y109_SLICE_X16Y109_BQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X12Y112_SLICE_X17Y112_B5Q),
.I3(CLBLM_L_X10Y105_SLICE_X12Y105_AQ),
.I4(CLBLM_R_X13Y109_SLICE_X18Y109_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y109_SLICE_X16Y109_DO5),
.O6(CLBLM_L_X12Y109_SLICE_X16Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hafacafacafacafac)
  ) CLBLM_L_X12Y109_SLICE_X16Y109_CLUT (
.I0(CLBLM_L_X8Y106_SLICE_X11Y106_A5Q),
.I1(CLBLM_L_X12Y108_SLICE_X17Y108_CO6),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X12Y112_SLICE_X16Y112_CQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y109_SLICE_X16Y109_CO5),
.O6(CLBLM_L_X12Y109_SLICE_X16Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff8aa88aa88aa8)
  ) CLBLM_L_X12Y109_SLICE_X16Y109_BLUT (
.I0(CLBLM_L_X12Y117_SLICE_X16Y117_AO6),
.I1(CLBLM_L_X12Y109_SLICE_X16Y109_BQ),
.I2(CLBLM_R_X11Y108_SLICE_X14Y108_BO6),
.I3(CLBLM_R_X11Y109_SLICE_X15Y109_CO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X12Y109_SLICE_X16Y109_DQ),
.O5(CLBLM_L_X12Y109_SLICE_X16Y109_BO5),
.O6(CLBLM_L_X12Y109_SLICE_X16Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfeaafc00faaaf000)
  ) CLBLM_L_X12Y109_SLICE_X16Y109_ALUT (
.I0(CLBLM_R_X13Y110_SLICE_X18Y110_AQ),
.I1(CLBLM_L_X12Y110_SLICE_X17Y110_BQ),
.I2(CLBLM_L_X12Y109_SLICE_X16Y109_AQ),
.I3(CLBLM_L_X12Y108_SLICE_X16Y108_AO5),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X12Y110_SLICE_X16Y110_CO5),
.O5(CLBLM_L_X12Y109_SLICE_X16Y109_AO5),
.O6(CLBLM_L_X12Y109_SLICE_X16Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y109_SLICE_X17Y109_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y109_SLICE_X17Y109_AO6),
.Q(CLBLM_L_X12Y109_SLICE_X17Y109_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y109_SLICE_X17Y109_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y109_SLICE_X17Y109_BO6),
.Q(CLBLM_L_X12Y109_SLICE_X17Y109_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y109_SLICE_X17Y109_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y109_SLICE_X17Y109_CO6),
.Q(CLBLM_L_X12Y109_SLICE_X17Y109_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y109_SLICE_X17Y109_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y109_SLICE_X17Y109_DO6),
.Q(CLBLM_L_X12Y109_SLICE_X17Y109_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaeeea00004440)
  ) CLBLM_L_X12Y109_SLICE_X17Y109_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.I2(CLBLM_L_X12Y109_SLICE_X17Y109_DQ),
.I3(CLBLM_R_X7Y109_SLICE_X8Y109_DO6),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLM_R_X11Y112_SLICE_X14Y112_BQ),
.O5(CLBLM_L_X12Y109_SLICE_X17Y109_DO5),
.O6(CLBLM_L_X12Y109_SLICE_X17Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc5500cccc5500)
  ) CLBLM_L_X12Y109_SLICE_X17Y109_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X10Y111_SLICE_X13Y111_BQ),
.I2(1'b1),
.I3(CLBLM_R_X7Y115_SLICE_X8Y115_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_L_X12Y109_SLICE_X17Y109_CO5),
.O6(CLBLM_L_X12Y109_SLICE_X17Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8888d8d88888d8d8)
  ) CLBLM_L_X12Y109_SLICE_X17Y109_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y107_SLICE_X7Y107_BQ),
.I2(CLBLM_L_X12Y109_SLICE_X17Y109_AQ),
.I3(1'b1),
.I4(CLBLM_L_X12Y108_SLICE_X17Y108_CO6),
.I5(1'b1),
.O5(CLBLM_L_X12Y109_SLICE_X17Y109_BO5),
.O6(CLBLM_L_X12Y109_SLICE_X17Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hafa5afa4a0a0a0a0)
  ) CLBLM_L_X12Y109_SLICE_X17Y109_ALUT (
.I0(CLBLM_L_X12Y105_SLICE_X16Y105_AQ),
.I1(CLBLM_R_X13Y113_SLICE_X18Y113_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X12Y107_SLICE_X17Y107_BQ),
.I4(CLBLM_R_X13Y109_SLICE_X19Y109_BQ),
.I5(CLBLM_L_X12Y109_SLICE_X16Y109_CQ),
.O5(CLBLM_L_X12Y109_SLICE_X17Y109_AO5),
.O6(CLBLM_L_X12Y109_SLICE_X17Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y110_SLICE_X16Y110_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y77_IOB_X0Y77_I),
.D(CLBLM_L_X12Y107_SLICE_X16Y107_CQ),
.Q(CLBLM_L_X12Y110_SLICE_X16Y110_AQ),
.R(CLBLM_L_X12Y117_SLICE_X16Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf8f0f0f088000000)
  ) CLBLM_L_X12Y110_SLICE_X16Y110_DLUT (
.I0(CLBLM_L_X12Y109_SLICE_X16Y109_AQ),
.I1(CLBLM_L_X12Y110_SLICE_X17Y110_BQ),
.I2(CLBLM_L_X10Y106_SLICE_X12Y106_BO6),
.I3(CLBLM_R_X11Y110_SLICE_X15Y110_AQ),
.I4(CLBLM_R_X13Y110_SLICE_X19Y110_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y110_SLICE_X16Y110_DO5),
.O6(CLBLM_L_X12Y110_SLICE_X16Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h070f000007000000)
  ) CLBLM_L_X12Y110_SLICE_X16Y110_CLUT (
.I0(CLBLM_L_X12Y109_SLICE_X16Y109_AQ),
.I1(CLBLM_L_X12Y110_SLICE_X17Y110_BQ),
.I2(CLBLM_L_X10Y106_SLICE_X12Y106_BO6),
.I3(CLBLM_R_X11Y110_SLICE_X15Y110_AQ),
.I4(CLBLM_R_X13Y110_SLICE_X19Y110_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y110_SLICE_X16Y110_CO5),
.O6(CLBLM_L_X12Y110_SLICE_X16Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaafc00fc00fc00)
  ) CLBLM_L_X12Y110_SLICE_X16Y110_BLUT (
.I0(CLBLL_L_X4Y117_SLICE_X4Y117_CQ),
.I1(CLBLM_R_X11Y112_SLICE_X14Y112_BQ),
.I2(CLBLM_L_X10Y110_SLICE_X13Y110_CQ),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_L_X12Y110_SLICE_X16Y110_BO5),
.O6(CLBLM_L_X12Y110_SLICE_X16Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfecc3200fa00fa00)
  ) CLBLM_L_X12Y110_SLICE_X16Y110_ALUT (
.I0(CLBLM_L_X8Y109_SLICE_X10Y109_DQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X8Y112_SLICE_X10Y112_A5Q),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(CLBLM_L_X12Y110_SLICE_X17Y110_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y110_SLICE_X16Y110_AO5),
.O6(CLBLM_L_X12Y110_SLICE_X16Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y110_SLICE_X17Y110_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y110_SLICE_X17Y110_AO6),
.Q(CLBLM_L_X12Y110_SLICE_X17Y110_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y110_SLICE_X17Y110_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y110_SLICE_X17Y110_BO6),
.Q(CLBLM_L_X12Y110_SLICE_X17Y110_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y110_SLICE_X17Y110_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y110_SLICE_X17Y110_CO6),
.Q(CLBLM_L_X12Y110_SLICE_X17Y110_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y110_SLICE_X17Y110_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y110_SLICE_X17Y110_DO6),
.Q(CLBLM_L_X12Y110_SLICE_X17Y110_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbbbbb88b8b8b888)
  ) CLBLM_L_X12Y110_SLICE_X17Y110_DLUT (
.I0(CLBLM_L_X8Y109_SLICE_X11Y109_CQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X12Y110_SLICE_X17Y110_DQ),
.I3(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLM_L_X10Y109_SLICE_X13Y109_CO6),
.O5(CLBLM_L_X12Y110_SLICE_X17Y110_DO5),
.O6(CLBLM_L_X12Y110_SLICE_X17Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcddccddc01100110)
  ) CLBLM_L_X12Y110_SLICE_X17Y110_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X12Y110_SLICE_X16Y110_BO5),
.I3(CLBLM_L_X8Y115_SLICE_X10Y115_CQ),
.I4(1'b1),
.I5(CLBLM_L_X12Y108_SLICE_X16Y108_BQ),
.O5(CLBLM_L_X12Y110_SLICE_X17Y110_CO5),
.O6(CLBLM_L_X12Y110_SLICE_X17Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff2800000028)
  ) CLBLM_L_X12Y110_SLICE_X17Y110_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X12Y110_SLICE_X17Y110_BQ),
.I2(CLBLM_L_X12Y110_SLICE_X16Y110_CO5),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y115_SLICE_X8Y115_DQ),
.I5(CLBLM_L_X12Y108_SLICE_X16Y108_AQ),
.O5(CLBLM_L_X12Y110_SLICE_X17Y110_BO5),
.O6(CLBLM_L_X12Y110_SLICE_X17Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdddcdddc11101110)
  ) CLBLM_L_X12Y110_SLICE_X17Y110_ALUT (
.I0(CLBLM_R_X5Y115_SLICE_X7Y115_CO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X12Y110_SLICE_X17Y110_AQ),
.I3(CLBLM_R_X11Y110_SLICE_X14Y110_CQ),
.I4(1'b1),
.I5(CLBLM_L_X8Y115_SLICE_X10Y115_CQ),
.O5(CLBLM_L_X12Y110_SLICE_X17Y110_AO5),
.O6(CLBLM_L_X12Y110_SLICE_X17Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y111_SLICE_X16Y111_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y111_SLICE_X16Y111_AO6),
.Q(CLBLM_L_X12Y111_SLICE_X16Y111_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y111_SLICE_X16Y111_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y111_SLICE_X16Y111_BO6),
.Q(CLBLM_L_X12Y111_SLICE_X16Y111_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y111_SLICE_X16Y111_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y111_SLICE_X16Y111_CO6),
.Q(CLBLM_L_X12Y111_SLICE_X16Y111_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y111_SLICE_X16Y111_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y111_SLICE_X16Y111_DO6),
.Q(CLBLM_L_X12Y111_SLICE_X16Y111_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf044f044f044f044)
  ) CLBLM_L_X12Y111_SLICE_X16Y111_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X12Y111_SLICE_X16Y111_CQ),
.I2(CLBLM_R_X11Y108_SLICE_X15Y108_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y111_SLICE_X16Y111_DO5),
.O6(CLBLM_L_X12Y111_SLICE_X16Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf088f088f088f088)
  ) CLBLM_L_X12Y111_SLICE_X16Y111_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X8Y111_SLICE_X11Y111_CQ),
.I2(CLBLM_R_X11Y107_SLICE_X15Y107_CQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y111_SLICE_X16Y111_CO5),
.O6(CLBLM_L_X12Y111_SLICE_X16Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa0af808fa0af808)
  ) CLBLM_L_X12Y111_SLICE_X16Y111_BLUT (
.I0(CLBLM_R_X7Y115_SLICE_X9Y115_DO6),
.I1(CLBLM_L_X12Y111_SLICE_X16Y111_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X12Y108_SLICE_X16Y108_CQ),
.I4(CLBLM_L_X12Y112_SLICE_X16Y112_DQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y111_SLICE_X16Y111_BO5),
.O6(CLBLM_L_X12Y111_SLICE_X16Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00f0f0ff00fcfc)
  ) CLBLM_L_X12Y111_SLICE_X16Y111_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y141_IOB_X1Y142_I),
.I2(CLBLM_L_X12Y111_SLICE_X16Y111_AQ),
.I3(CLBLM_L_X10Y113_SLICE_X12Y113_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y119_SLICE_X10Y119_AQ),
.O5(CLBLM_L_X12Y111_SLICE_X16Y111_AO5),
.O6(CLBLM_L_X12Y111_SLICE_X16Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y111_SLICE_X17Y111_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y111_SLICE_X17Y111_DO5),
.O6(CLBLM_L_X12Y111_SLICE_X17Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y111_SLICE_X17Y111_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y111_SLICE_X17Y111_CO5),
.O6(CLBLM_L_X12Y111_SLICE_X17Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y111_SLICE_X17Y111_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y111_SLICE_X17Y111_BO5),
.O6(CLBLM_L_X12Y111_SLICE_X17Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y111_SLICE_X17Y111_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y111_SLICE_X17Y111_AO5),
.O6(CLBLM_L_X12Y111_SLICE_X17Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y112_SLICE_X16Y112_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y112_SLICE_X14Y112_AO6),
.Q(CLBLM_L_X12Y112_SLICE_X16Y112_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y112_SLICE_X16Y112_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y112_SLICE_X16Y112_BO5),
.Q(CLBLM_L_X12Y112_SLICE_X16Y112_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y112_SLICE_X16Y112_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y112_SLICE_X16Y112_AO6),
.Q(CLBLM_L_X12Y112_SLICE_X16Y112_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y112_SLICE_X16Y112_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y112_SLICE_X16Y112_BO6),
.Q(CLBLM_L_X12Y112_SLICE_X16Y112_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y112_SLICE_X16Y112_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y112_SLICE_X16Y112_CO6),
.Q(CLBLM_L_X12Y112_SLICE_X16Y112_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y112_SLICE_X16Y112_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y112_SLICE_X16Y112_DO6),
.Q(CLBLM_L_X12Y112_SLICE_X16Y112_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffcff0000fc0000)
  ) CLBLM_L_X12Y112_SLICE_X16Y112_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X12Y113_SLICE_X16Y113_CQ),
.I2(CLBLM_L_X12Y112_SLICE_X16Y112_DQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y115_SLICE_X9Y115_DO6),
.I5(CLBLM_L_X8Y105_SLICE_X11Y105_BQ),
.O5(CLBLM_L_X12Y112_SLICE_X16Y112_DO5),
.O6(CLBLM_L_X12Y112_SLICE_X16Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000ffaa00aa)
  ) CLBLM_L_X12Y112_SLICE_X16Y112_CLUT (
.I0(CLBLM_L_X12Y112_SLICE_X16Y112_BQ),
.I1(1'b1),
.I2(1'b1),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X11Y114_SLICE_X14Y114_CQ),
.I5(CLBLM_L_X12Y108_SLICE_X17Y108_CO6),
.O5(CLBLM_L_X12Y112_SLICE_X16Y112_CO5),
.O6(CLBLM_L_X12Y112_SLICE_X16Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0afa0a0cacacaca)
  ) CLBLM_L_X12Y112_SLICE_X16Y112_BLUT (
.I0(CLBLM_R_X11Y116_SLICE_X14Y116_A5Q),
.I1(CLBLM_L_X10Y112_SLICE_X12Y112_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X12Y108_SLICE_X17Y108_CO6),
.I4(CLBLM_L_X12Y109_SLICE_X17Y109_BQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y112_SLICE_X16Y112_BO5),
.O6(CLBLM_L_X12Y112_SLICE_X16Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdcc3100fccc3000)
  ) CLBLM_L_X12Y112_SLICE_X16Y112_ALUT (
.I0(RIOB33_X105Y121_IOB_X1Y121_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X12Y112_SLICE_X16Y112_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X11Y113_SLICE_X15Y113_AQ),
.I5(CLBLM_R_X11Y113_SLICE_X14Y113_CQ),
.O5(CLBLM_L_X12Y112_SLICE_X16Y112_AO5),
.O6(CLBLM_L_X12Y112_SLICE_X16Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y112_SLICE_X17Y112_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y110_SLICE_X16Y110_AO6),
.Q(CLBLM_L_X12Y112_SLICE_X17Y112_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y112_SLICE_X17Y112_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y112_SLICE_X17Y112_CO6),
.Q(CLBLM_L_X12Y112_SLICE_X17Y112_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y112_SLICE_X17Y112_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y112_SLICE_X17Y112_AO6),
.Q(CLBLM_L_X12Y112_SLICE_X17Y112_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y112_SLICE_X17Y112_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y112_SLICE_X17Y112_BO6),
.Q(CLBLM_L_X12Y112_SLICE_X17Y112_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffafffffffa)
  ) CLBLM_L_X12Y112_SLICE_X17Y112_DLUT (
.I0(CLBLM_R_X11Y111_SLICE_X15Y111_BQ),
.I1(1'b1),
.I2(CLBLM_R_X7Y115_SLICE_X8Y115_CQ),
.I3(CLBLM_L_X12Y111_SLICE_X16Y111_CQ),
.I4(CLBLM_L_X12Y109_SLICE_X17Y109_CQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y112_SLICE_X17Y112_DO5),
.O6(CLBLM_L_X12Y112_SLICE_X17Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaf0aac0f0f0c0c0)
  ) CLBLM_L_X12Y112_SLICE_X17Y112_CLUT (
.I0(CLBLM_R_X13Y110_SLICE_X18Y110_BQ),
.I1(CLBLM_R_X11Y111_SLICE_X15Y111_BQ),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X12Y110_SLICE_X17Y110_DQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y112_SLICE_X17Y112_CO5),
.O6(CLBLM_L_X12Y112_SLICE_X17Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0011112222)
  ) CLBLM_L_X12Y112_SLICE_X17Y112_BLUT (
.I0(CLBLM_R_X5Y112_SLICE_X7Y112_CQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(1'b1),
.I3(CLBLM_L_X12Y109_SLICE_X16Y109_CQ),
.I4(CLBLM_L_X12Y112_SLICE_X17Y112_CO5),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X12Y112_SLICE_X17Y112_BO5),
.O6(CLBLM_L_X12Y112_SLICE_X17Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaaffaaffaa3f)
  ) CLBLM_L_X12Y112_SLICE_X17Y112_ALUT (
.I0(CLBLM_L_X12Y112_SLICE_X17Y112_B5Q),
.I1(RIOB33_X105Y135_IOB_X1Y135_I),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X13Y113_SLICE_X18Y113_DO6),
.I5(RIOB33_X105Y135_IOB_X1Y136_I),
.O5(CLBLM_L_X12Y112_SLICE_X17Y112_AO5),
.O6(CLBLM_L_X12Y112_SLICE_X17Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y113_SLICE_X16Y113_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y113_SLICE_X16Y113_AO6),
.Q(CLBLM_L_X12Y113_SLICE_X16Y113_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y113_SLICE_X16Y113_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y113_SLICE_X16Y113_BO6),
.Q(CLBLM_L_X12Y113_SLICE_X16Y113_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y113_SLICE_X16Y113_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y113_SLICE_X16Y113_CO6),
.Q(CLBLM_L_X12Y113_SLICE_X16Y113_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffefefefe)
  ) CLBLM_L_X12Y113_SLICE_X16Y113_DLUT (
.I0(CLBLM_L_X8Y115_SLICE_X10Y115_AQ),
.I1(CLBLM_L_X12Y113_SLICE_X16Y113_CQ),
.I2(CLBLM_L_X8Y115_SLICE_X11Y115_BQ),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X10Y115_SLICE_X13Y115_BQ),
.O5(CLBLM_L_X12Y113_SLICE_X16Y113_DO5),
.O6(CLBLM_L_X12Y113_SLICE_X16Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5a0a0e4e4a0a0)
  ) CLBLM_L_X12Y113_SLICE_X16Y113_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X12Y113_SLICE_X16Y113_CQ),
.I2(CLBLM_L_X12Y113_SLICE_X16Y113_BQ),
.I3(1'b1),
.I4(CLBLM_R_X7Y115_SLICE_X9Y115_DO6),
.I5(CLBLM_R_X11Y113_SLICE_X15Y113_AQ),
.O5(CLBLM_L_X12Y113_SLICE_X16Y113_CO5),
.O6(CLBLM_L_X12Y113_SLICE_X16Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000ff00eeee)
  ) CLBLM_L_X12Y113_SLICE_X16Y113_BLUT (
.I0(CLBLM_R_X11Y114_SLICE_X14Y114_DQ),
.I1(CLBLM_L_X12Y113_SLICE_X16Y113_BQ),
.I2(1'b1),
.I3(CLBLM_L_X12Y112_SLICE_X16Y112_DQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X5Y115_SLICE_X7Y115_CO6),
.O5(CLBLM_L_X12Y113_SLICE_X16Y113_BO5),
.O6(CLBLM_L_X12Y113_SLICE_X16Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffa50ea40)
  ) CLBLM_L_X12Y113_SLICE_X16Y113_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_L_X12Y113_SLICE_X16Y113_AQ),
.I3(CLBLM_L_X12Y113_SLICE_X16Y113_CQ),
.I4(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.I5(CLBLM_R_X7Y112_SLICE_X9Y112_CO6),
.O5(CLBLM_L_X12Y113_SLICE_X16Y113_AO5),
.O6(CLBLM_L_X12Y113_SLICE_X16Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y113_SLICE_X17Y113_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y113_SLICE_X17Y113_BO5),
.Q(CLBLM_L_X12Y113_SLICE_X17Y113_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y113_SLICE_X17Y113_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y113_SLICE_X17Y113_AO6),
.Q(CLBLM_L_X12Y113_SLICE_X17Y113_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y113_SLICE_X17Y113_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y113_SLICE_X17Y113_BO6),
.Q(CLBLM_L_X12Y113_SLICE_X17Y113_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y113_SLICE_X17Y113_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y113_SLICE_X17Y113_CO6),
.Q(CLBLM_L_X12Y113_SLICE_X17Y113_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ffffffff000a)
  ) CLBLM_L_X12Y113_SLICE_X17Y113_DLUT (
.I0(CLBLM_R_X11Y109_SLICE_X15Y109_DO6),
.I1(1'b1),
.I2(CLBLM_L_X12Y114_SLICE_X17Y114_CO6),
.I3(CLBLM_L_X12Y113_SLICE_X16Y113_DO6),
.I4(CLBLM_R_X13Y113_SLICE_X18Y113_CQ),
.I5(CLBLM_L_X12Y114_SLICE_X17Y114_BQ),
.O5(CLBLM_L_X12Y113_SLICE_X17Y113_DO5),
.O6(CLBLM_L_X12Y113_SLICE_X17Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff0ffccfff0ff88)
  ) CLBLM_L_X12Y113_SLICE_X17Y113_CLUT (
.I0(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.I1(CLBLM_L_X12Y113_SLICE_X17Y113_CQ),
.I2(CLBLM_R_X13Y113_SLICE_X19Y113_AQ),
.I3(CLBLM_R_X7Y110_SLICE_X9Y110_CO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_L_X12Y113_SLICE_X17Y113_CO5),
.O6(CLBLM_L_X12Y113_SLICE_X17Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff000f0f022f022)
  ) CLBLM_L_X12Y113_SLICE_X17Y113_BLUT (
.I0(CLBLM_L_X12Y113_SLICE_X17Y113_B5Q),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_L_X12Y112_SLICE_X17Y112_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X11Y115_SLICE_X15Y115_B5Q),
.I5(1'b1),
.O5(CLBLM_L_X12Y113_SLICE_X17Y113_BO5),
.O6(CLBLM_L_X12Y113_SLICE_X17Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5f5f5f5b1f5f5)
  ) CLBLM_L_X12Y113_SLICE_X17Y113_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(CLBLM_L_X12Y109_SLICE_X17Y109_AQ),
.I3(RIOB33_X105Y135_IOB_X1Y135_I),
.I4(RIOB33_X105Y135_IOB_X1Y136_I),
.I5(CLBLM_R_X13Y113_SLICE_X18Y113_DO6),
.O5(CLBLM_L_X12Y113_SLICE_X17Y113_AO5),
.O6(CLBLM_L_X12Y113_SLICE_X17Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y114_SLICE_X16Y114_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y114_SLICE_X16Y114_AO6),
.Q(CLBLM_L_X12Y114_SLICE_X16Y114_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y114_SLICE_X16Y114_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y114_SLICE_X16Y114_BO6),
.Q(CLBLM_L_X12Y114_SLICE_X16Y114_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y114_SLICE_X16Y114_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y114_SLICE_X16Y114_CO6),
.Q(CLBLM_L_X12Y114_SLICE_X16Y114_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5544554455555050)
  ) CLBLM_L_X12Y114_SLICE_X16Y114_DLUT (
.I0(CLBLM_L_X10Y113_SLICE_X13Y113_CQ),
.I1(CLBLM_L_X12Y114_SLICE_X16Y114_CQ),
.I2(CLBLM_L_X10Y110_SLICE_X13Y110_DQ),
.I3(CLBLM_L_X8Y115_SLICE_X11Y115_AQ),
.I4(CLBLM_L_X12Y113_SLICE_X16Y113_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y114_SLICE_X16Y114_DO5),
.O6(CLBLM_L_X12Y114_SLICE_X16Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f055004400)
  ) CLBLM_L_X12Y114_SLICE_X16Y114_CLUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_L_X12Y114_SLICE_X16Y114_CQ),
.I2(CLBLM_L_X12Y117_SLICE_X17Y117_BQ),
.I3(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.I4(CLBLM_L_X10Y111_SLICE_X13Y111_DO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X12Y114_SLICE_X16Y114_CO5),
.O6(CLBLM_L_X12Y114_SLICE_X16Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0eff0e000e000e)
  ) CLBLM_L_X12Y114_SLICE_X16Y114_BLUT (
.I0(CLBLM_R_X11Y115_SLICE_X15Y115_CQ),
.I1(CLBLM_L_X12Y114_SLICE_X16Y114_BQ),
.I2(CLBLM_R_X5Y115_SLICE_X7Y115_CO6),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLM_R_X11Y114_SLICE_X14Y114_DQ),
.O5(CLBLM_L_X12Y114_SLICE_X16Y114_BO5),
.O6(CLBLM_L_X12Y114_SLICE_X16Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f3c0c0f3c0c0c0)
  ) CLBLM_L_X12Y114_SLICE_X16Y114_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X11Y111_SLICE_X15Y111_CQ),
.I3(CLBLM_L_X12Y114_SLICE_X16Y114_AQ),
.I4(CLBLM_R_X7Y115_SLICE_X9Y115_DO6),
.I5(CLBLM_L_X8Y114_SLICE_X10Y114_BQ),
.O5(CLBLM_L_X12Y114_SLICE_X16Y114_AO5),
.O6(CLBLM_L_X12Y114_SLICE_X16Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y114_SLICE_X17Y114_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y114_SLICE_X17Y114_AO6),
.Q(CLBLM_L_X12Y114_SLICE_X17Y114_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y114_SLICE_X17Y114_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y114_SLICE_X17Y114_BO6),
.Q(CLBLM_L_X12Y114_SLICE_X17Y114_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y114_SLICE_X17Y114_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y114_SLICE_X17Y114_DO5),
.O6(CLBLM_L_X12Y114_SLICE_X17Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffeeeeffffeeee)
  ) CLBLM_L_X12Y114_SLICE_X17Y114_CLUT (
.I0(CLBLM_L_X12Y112_SLICE_X16Y112_DQ),
.I1(CLBLM_L_X12Y114_SLICE_X17Y114_AQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_L_X12Y111_SLICE_X16Y111_BQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y114_SLICE_X17Y114_CO5),
.O6(CLBLM_L_X12Y114_SLICE_X17Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00aafcaafc)
  ) CLBLM_L_X12Y114_SLICE_X17Y114_BLUT (
.I0(CLBLM_R_X11Y115_SLICE_X15Y115_AQ),
.I1(CLBLM_L_X12Y114_SLICE_X17Y114_BQ),
.I2(CLBLM_L_X12Y114_SLICE_X17Y114_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLM_R_X5Y115_SLICE_X7Y115_CO6),
.O5(CLBLM_L_X12Y114_SLICE_X17Y114_BO5),
.O6(CLBLM_L_X12Y114_SLICE_X17Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa33aa33aa30aa30)
  ) CLBLM_L_X12Y114_SLICE_X17Y114_ALUT (
.I0(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.I1(CLBLM_R_X5Y115_SLICE_X7Y115_CO6),
.I2(CLBLM_L_X12Y114_SLICE_X17Y114_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLM_L_X12Y111_SLICE_X16Y111_BQ),
.O5(CLBLM_L_X12Y114_SLICE_X17Y114_AO5),
.O6(CLBLM_L_X12Y114_SLICE_X17Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y115_SLICE_X16Y115_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y115_SLICE_X14Y115_BO6),
.Q(CLBLM_L_X12Y115_SLICE_X16Y115_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y115_SLICE_X16Y115_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y115_SLICE_X16Y115_DO5),
.O6(CLBLM_L_X12Y115_SLICE_X16Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y115_SLICE_X16Y115_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y115_SLICE_X16Y115_CO5),
.O6(CLBLM_L_X12Y115_SLICE_X16Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y115_SLICE_X16Y115_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y115_SLICE_X16Y115_BO5),
.O6(CLBLM_L_X12Y115_SLICE_X16Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y115_SLICE_X16Y115_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y115_SLICE_X16Y115_AO5),
.O6(CLBLM_L_X12Y115_SLICE_X16Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y115_SLICE_X17Y115_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y115_SLICE_X17Y115_DO5),
.O6(CLBLM_L_X12Y115_SLICE_X17Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y115_SLICE_X17Y115_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y115_SLICE_X17Y115_CO5),
.O6(CLBLM_L_X12Y115_SLICE_X17Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y115_SLICE_X17Y115_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y115_SLICE_X17Y115_BO5),
.O6(CLBLM_L_X12Y115_SLICE_X17Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y115_SLICE_X17Y115_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y115_SLICE_X17Y115_AO5),
.O6(CLBLM_L_X12Y115_SLICE_X17Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y117_SLICE_X16Y117_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y77_IOB_X0Y77_I),
.D(CLBLM_R_X13Y109_SLICE_X19Y109_BQ),
.Q(CLBLM_L_X12Y117_SLICE_X16Y117_AQ),
.R(CLBLM_L_X12Y117_SLICE_X16Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y117_SLICE_X16Y117_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y117_SLICE_X16Y117_DO5),
.O6(CLBLM_L_X12Y117_SLICE_X16Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y117_SLICE_X16Y117_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y117_SLICE_X16Y117_CO5),
.O6(CLBLM_L_X12Y117_SLICE_X16Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y117_SLICE_X16Y117_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y117_SLICE_X16Y117_BO5),
.O6(CLBLM_L_X12Y117_SLICE_X16Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000ccffccff)
  ) CLBLM_L_X12Y117_SLICE_X16Y117_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y119_SLICE_X10Y119_AQ),
.I2(1'b1),
.I3(RIOB33_X105Y141_IOB_X1Y142_I),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X12Y117_SLICE_X16Y117_AO5),
.O6(CLBLM_L_X12Y117_SLICE_X16Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y117_SLICE_X17Y117_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y117_SLICE_X17Y117_AO6),
.Q(CLBLM_L_X12Y117_SLICE_X17Y117_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y117_SLICE_X17Y117_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y117_SLICE_X17Y117_BO6),
.Q(CLBLM_L_X12Y117_SLICE_X17Y117_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y117_SLICE_X17Y117_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y117_SLICE_X17Y117_DO5),
.O6(CLBLM_L_X12Y117_SLICE_X17Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y117_SLICE_X17Y117_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y117_SLICE_X17Y117_CO5),
.O6(CLBLM_L_X12Y117_SLICE_X17Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaffffc030)
  ) CLBLM_L_X12Y117_SLICE_X17Y117_BLUT (
.I0(CLBLM_L_X12Y107_SLICE_X17Y107_AQ),
.I1(CLBLM_L_X12Y117_SLICE_X17Y117_BQ),
.I2(CLBLM_L_X10Y116_SLICE_X12Y116_DO5),
.I3(CLBLM_L_X10Y118_SLICE_X13Y118_BO6),
.I4(CLBLM_L_X10Y118_SLICE_X13Y118_CO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X12Y117_SLICE_X17Y117_BO5),
.O6(CLBLM_L_X12Y117_SLICE_X17Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00f0f0fcfc)
  ) CLBLM_L_X12Y117_SLICE_X17Y117_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y141_IOB_X1Y142_I),
.I2(CLBLM_L_X12Y117_SLICE_X17Y117_AQ),
.I3(CLBLM_R_X11Y117_SLICE_X15Y117_CQ),
.I4(CLBLM_L_X8Y119_SLICE_X10Y119_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X12Y117_SLICE_X17Y117_AO5),
.O6(CLBLM_L_X12Y117_SLICE_X17Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y118_SLICE_X16Y118_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y77_IOB_X0Y77_I),
.D(CLBLM_R_X11Y117_SLICE_X15Y117_AQ),
.Q(CLBLM_L_X12Y118_SLICE_X16Y118_AQ),
.R(CLBLM_L_X12Y117_SLICE_X16Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y118_SLICE_X16Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y118_SLICE_X16Y118_DO5),
.O6(CLBLM_L_X12Y118_SLICE_X16Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y118_SLICE_X16Y118_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y118_SLICE_X16Y118_CO5),
.O6(CLBLM_L_X12Y118_SLICE_X16Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y118_SLICE_X16Y118_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y118_SLICE_X16Y118_BO5),
.O6(CLBLM_L_X12Y118_SLICE_X16Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y118_SLICE_X16Y118_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y118_SLICE_X16Y118_AO5),
.O6(CLBLM_L_X12Y118_SLICE_X16Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y118_SLICE_X17Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y118_SLICE_X17Y118_DO5),
.O6(CLBLM_L_X12Y118_SLICE_X17Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y118_SLICE_X17Y118_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y118_SLICE_X17Y118_CO5),
.O6(CLBLM_L_X12Y118_SLICE_X17Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y118_SLICE_X17Y118_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y118_SLICE_X17Y118_BO5),
.O6(CLBLM_L_X12Y118_SLICE_X17Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y118_SLICE_X17Y118_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y118_SLICE_X17Y118_AO5),
.O6(CLBLM_L_X12Y118_SLICE_X17Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y106_SLICE_X2Y106_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y106_SLICE_X2Y106_DO5),
.O6(CLBLM_R_X3Y106_SLICE_X2Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffaaee00cc)
  ) CLBLM_R_X3Y106_SLICE_X2Y106_CLUT (
.I0(LIOB33_X0Y53_IOB_X0Y53_I),
.I1(LIOB33_X0Y51_IOB_X0Y51_I),
.I2(1'b1),
.I3(CLBLL_L_X2Y110_SLICE_X1Y110_DO6),
.I4(CLBLM_R_X3Y111_SLICE_X2Y111_CO6),
.I5(CLBLM_R_X3Y109_SLICE_X2Y109_DO6),
.O5(CLBLM_R_X3Y106_SLICE_X2Y106_CO5),
.O6(CLBLM_R_X3Y106_SLICE_X2Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h33333333bfffbfff)
  ) CLBLM_R_X3Y106_SLICE_X2Y106_BLUT (
.I0(CLBLM_R_X3Y109_SLICE_X2Y109_AQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X3Y110_SLICE_X3Y110_AO6),
.I3(CLBLL_L_X4Y113_SLICE_X4Y113_BQ),
.I4(1'b1),
.I5(CLBLM_R_X3Y106_SLICE_X2Y106_CO6),
.O5(CLBLM_R_X3Y106_SLICE_X2Y106_BO5),
.O6(CLBLM_R_X3Y106_SLICE_X2Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000cccc8ccccccc)
  ) CLBLM_R_X3Y106_SLICE_X2Y106_ALUT (
.I0(CLBLM_R_X3Y109_SLICE_X2Y109_AQ),
.I1(CLBLM_R_X5Y106_SLICE_X7Y106_CO6),
.I2(CLBLM_R_X3Y110_SLICE_X3Y110_AO6),
.I3(CLBLL_L_X4Y113_SLICE_X4Y113_BQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X3Y106_SLICE_X2Y106_CO6),
.O5(CLBLM_R_X3Y106_SLICE_X2Y106_AO5),
.O6(CLBLM_R_X3Y106_SLICE_X2Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y106_SLICE_X3Y106_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y106_SLICE_X3Y106_DO5),
.O6(CLBLM_R_X3Y106_SLICE_X3Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y106_SLICE_X3Y106_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y106_SLICE_X3Y106_CO5),
.O6(CLBLM_R_X3Y106_SLICE_X3Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y106_SLICE_X3Y106_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y106_SLICE_X3Y106_BO5),
.O6(CLBLM_R_X3Y106_SLICE_X3Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y106_SLICE_X3Y106_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y106_SLICE_X3Y106_AO5),
.O6(CLBLM_R_X3Y106_SLICE_X3Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f000f000f000f00)
  ) CLBLM_R_X3Y107_SLICE_X2Y107_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLL_L_X2Y108_SLICE_X1Y108_AO6),
.I3(CLBLM_R_X7Y106_SLICE_X8Y106_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y107_SLICE_X2Y107_DO5),
.O6(CLBLM_R_X3Y107_SLICE_X2Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000040000)
  ) CLBLM_R_X3Y107_SLICE_X2Y107_CLUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(RIOB33_X105Y133_IOB_X1Y134_I),
.I2(RIOB33_X105Y133_IOB_X1Y133_I),
.I3(RIOB33_X105Y131_IOB_X1Y132_I),
.I4(CLBLM_R_X5Y107_SLICE_X6Y107_DQ),
.I5(CLBLL_L_X2Y114_SLICE_X0Y114_AO6),
.O5(CLBLM_R_X3Y107_SLICE_X2Y107_CO5),
.O6(CLBLM_R_X3Y107_SLICE_X2Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000200000000000)
  ) CLBLM_R_X3Y107_SLICE_X2Y107_BLUT (
.I0(RIOB33_X105Y133_IOB_X1Y133_I),
.I1(CLBLL_L_X2Y114_SLICE_X0Y114_AO6),
.I2(RIOB33_X105Y133_IOB_X1Y134_I),
.I3(CLBLM_R_X5Y107_SLICE_X6Y107_BQ),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(RIOB33_X105Y131_IOB_X1Y132_I),
.O5(CLBLM_R_X3Y107_SLICE_X2Y107_BO5),
.O6(CLBLM_R_X3Y107_SLICE_X2Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h2000000000000000)
  ) CLBLM_R_X3Y107_SLICE_X2Y107_ALUT (
.I0(RIOB33_X105Y133_IOB_X1Y133_I),
.I1(CLBLL_L_X2Y114_SLICE_X0Y114_AO6),
.I2(CLBLM_R_X5Y109_SLICE_X6Y109_AQ),
.I3(RIOB33_X105Y133_IOB_X1Y134_I),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(RIOB33_X105Y131_IOB_X1Y132_I),
.O5(CLBLM_R_X3Y107_SLICE_X2Y107_AO5),
.O6(CLBLM_R_X3Y107_SLICE_X2Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y107_SLICE_X3Y107_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y107_SLICE_X3Y107_AO6),
.Q(CLBLM_R_X3Y107_SLICE_X3Y107_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y107_SLICE_X3Y107_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y107_SLICE_X3Y107_DO5),
.O6(CLBLM_R_X3Y107_SLICE_X3Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000001)
  ) CLBLM_R_X3Y107_SLICE_X3Y107_CLUT (
.I0(CLBLM_R_X3Y108_SLICE_X3Y108_AO6),
.I1(CLBLL_L_X2Y111_SLICE_X1Y111_CO6),
.I2(CLBLM_R_X3Y110_SLICE_X2Y110_DO6),
.I3(CLBLM_R_X3Y109_SLICE_X2Y109_CO6),
.I4(CLBLM_R_X3Y111_SLICE_X2Y111_CO6),
.I5(CLBLM_R_X3Y110_SLICE_X3Y110_AO6),
.O5(CLBLM_R_X3Y107_SLICE_X3Y107_CO5),
.O6(CLBLM_R_X3Y107_SLICE_X3Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffaffc0ccc0cc)
  ) CLBLM_R_X3Y107_SLICE_X3Y107_BLUT (
.I0(RIOB33_X105Y127_IOB_X1Y128_I),
.I1(CLBLM_R_X5Y107_SLICE_X7Y107_BQ),
.I2(RIOB33_X105Y129_IOB_X1Y129_I),
.I3(RIOB33_X105Y137_IOB_X1Y137_I),
.I4(CLBLM_R_X3Y110_SLICE_X3Y110_AO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y107_SLICE_X3Y107_BO5),
.O6(CLBLM_R_X3Y107_SLICE_X3Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccca5a5aaa5)
  ) CLBLM_R_X3Y107_SLICE_X3Y107_ALUT (
.I0(CLBLL_L_X4Y107_SLICE_X5Y107_DO6),
.I1(CLBLM_L_X10Y112_SLICE_X13Y112_AQ),
.I2(CLBLM_R_X3Y107_SLICE_X3Y107_AQ),
.I3(RIOB33_X105Y137_IOB_X1Y137_I),
.I4(RIOB33_X105Y129_IOB_X1Y129_I),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X3Y107_SLICE_X3Y107_AO5),
.O6(CLBLM_R_X3Y107_SLICE_X3Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffffba)
  ) CLBLM_R_X3Y108_SLICE_X2Y108_DLUT (
.I0(CLBLL_L_X4Y108_SLICE_X5Y108_BO6),
.I1(CLBLL_L_X2Y110_SLICE_X1Y110_CO6),
.I2(CLBLL_L_X2Y108_SLICE_X1Y108_AO5),
.I3(CLBLM_R_X3Y108_SLICE_X3Y108_DO6),
.I4(CLBLL_L_X2Y109_SLICE_X1Y109_DO6),
.I5(CLBLM_R_X3Y107_SLICE_X2Y107_DO6),
.O5(CLBLM_R_X3Y108_SLICE_X2Y108_DO5),
.O6(CLBLM_R_X3Y108_SLICE_X2Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffafffe)
  ) CLBLM_R_X3Y108_SLICE_X2Y108_CLUT (
.I0(CLBLM_R_X3Y108_SLICE_X2Y108_AO6),
.I1(CLBLM_R_X7Y106_SLICE_X8Y106_AQ),
.I2(CLBLL_L_X2Y109_SLICE_X0Y109_DO6),
.I3(CLBLM_R_X3Y107_SLICE_X2Y107_AO6),
.I4(CLBLL_L_X2Y108_SLICE_X1Y108_AO6),
.I5(CLBLM_R_X3Y111_SLICE_X3Y111_AO6),
.O5(CLBLM_R_X3Y108_SLICE_X2Y108_CO5),
.O6(CLBLM_R_X3Y108_SLICE_X2Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000300000001)
  ) CLBLM_R_X3Y108_SLICE_X2Y108_BLUT (
.I0(CLBLL_L_X2Y108_SLICE_X1Y108_AO5),
.I1(CLBLM_R_X3Y108_SLICE_X3Y108_DO6),
.I2(CLBLL_L_X4Y108_SLICE_X5Y108_BO6),
.I3(CLBLL_L_X2Y108_SLICE_X1Y108_CO6),
.I4(CLBLM_L_X10Y112_SLICE_X12Y112_DO6),
.I5(CLBLL_L_X2Y110_SLICE_X1Y110_CO6),
.O5(CLBLM_R_X3Y108_SLICE_X2Y108_BO5),
.O6(CLBLM_R_X3Y108_SLICE_X2Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000040000000000)
  ) CLBLM_R_X3Y108_SLICE_X2Y108_ALUT (
.I0(RIOB33_X105Y133_IOB_X1Y133_I),
.I1(CLBLM_R_X7Y109_SLICE_X9Y109_AQ),
.I2(CLBLM_R_X3Y116_SLICE_X3Y116_AO6),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(RIOB33_X105Y131_IOB_X1Y132_I),
.I5(RIOB33_X105Y133_IOB_X1Y134_I),
.O5(CLBLM_R_X3Y108_SLICE_X2Y108_AO5),
.O6(CLBLM_R_X3Y108_SLICE_X2Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0c0cffff0c0c0c0c)
  ) CLBLM_R_X3Y108_SLICE_X3Y108_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y109_SLICE_X6Y109_AQ),
.I2(CLBLM_R_X3Y112_SLICE_X2Y112_AO5),
.I3(1'b1),
.I4(CLBLL_L_X2Y110_SLICE_X0Y110_BO5),
.I5(CLBLM_R_X7Y109_SLICE_X9Y109_AQ),
.O5(CLBLM_R_X3Y108_SLICE_X3Y108_DO5),
.O6(CLBLM_R_X3Y108_SLICE_X3Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0e10f0f0f0f)
  ) CLBLM_R_X3Y108_SLICE_X3Y108_CLUT (
.I0(CLBLL_L_X4Y108_SLICE_X5Y108_BO6),
.I1(CLBLM_R_X3Y108_SLICE_X2Y108_CO6),
.I2(CLBLM_R_X5Y107_SLICE_X7Y107_AQ),
.I3(CLBLM_L_X10Y112_SLICE_X12Y112_DO6),
.I4(CLBLL_L_X2Y109_SLICE_X1Y109_AO6),
.I5(CLBLM_R_X11Y110_SLICE_X14Y110_AQ),
.O5(CLBLM_R_X3Y108_SLICE_X3Y108_CO5),
.O6(CLBLM_R_X3Y108_SLICE_X3Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000004000)
  ) CLBLM_R_X3Y108_SLICE_X3Y108_BLUT (
.I0(RIOB33_X105Y133_IOB_X1Y133_I),
.I1(RIOB33_X105Y133_IOB_X1Y134_I),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(CLBLL_L_X4Y112_SLICE_X4Y112_BQ),
.I4(CLBLM_R_X3Y116_SLICE_X3Y116_AO6),
.I5(RIOB33_X105Y131_IOB_X1Y132_I),
.O5(CLBLM_R_X3Y108_SLICE_X3Y108_BO5),
.O6(CLBLM_R_X3Y108_SLICE_X3Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffeffffffff)
  ) CLBLM_R_X3Y108_SLICE_X3Y108_ALUT (
.I0(CLBLL_L_X2Y109_SLICE_X1Y109_AO6),
.I1(CLBLM_R_X3Y109_SLICE_X3Y109_AO6),
.I2(CLBLM_R_X3Y108_SLICE_X2Y108_CO6),
.I3(CLBLL_L_X4Y108_SLICE_X5Y108_BO6),
.I4(CLBLL_L_X4Y109_SLICE_X4Y109_DO6),
.I5(CLBLL_L_X2Y109_SLICE_X1Y109_CO6),
.O5(CLBLM_R_X3Y108_SLICE_X3Y108_AO5),
.O6(CLBLM_R_X3Y108_SLICE_X3Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y109_SLICE_X2Y109_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y109_SLICE_X2Y109_AO5),
.Q(CLBLM_R_X3Y109_SLICE_X2Y109_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y109_SLICE_X2Y109_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y109_SLICE_X2Y109_AO6),
.Q(CLBLM_R_X3Y109_SLICE_X2Y109_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0ea00aac0c00000)
  ) CLBLM_R_X3Y109_SLICE_X2Y109_DLUT (
.I0(CLBLM_R_X3Y109_SLICE_X2Y109_CO6),
.I1(CLBLL_L_X4Y113_SLICE_X5Y113_B5Q),
.I2(CLBLM_R_X3Y110_SLICE_X2Y110_DO6),
.I3(CLBLM_R_X3Y109_SLICE_X2Y109_A5Q),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X3Y115_SLICE_X2Y115_AQ),
.O5(CLBLM_R_X3Y109_SLICE_X2Y109_DO5),
.O6(CLBLM_R_X3Y109_SLICE_X2Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffcfcfffffdfc)
  ) CLBLM_R_X3Y109_SLICE_X2Y109_CLUT (
.I0(CLBLL_L_X2Y110_SLICE_X1Y110_CO6),
.I1(CLBLM_R_X3Y110_SLICE_X3Y110_CO6),
.I2(CLBLL_L_X4Y109_SLICE_X5Y109_DO6),
.I3(CLBLL_L_X2Y109_SLICE_X0Y109_BO5),
.I4(CLBLL_L_X4Y112_SLICE_X4Y112_DO6),
.I5(CLBLL_L_X2Y112_SLICE_X1Y112_AO6),
.O5(CLBLM_R_X3Y109_SLICE_X2Y109_CO5),
.O6(CLBLM_R_X3Y109_SLICE_X2Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000008)
  ) CLBLM_R_X3Y109_SLICE_X2Y109_BLUT (
.I0(RIOB33_X105Y133_IOB_X1Y133_I),
.I1(CLBLM_R_X5Y115_SLICE_X6Y115_AQ),
.I2(RIOB33_X105Y133_IOB_X1Y134_I),
.I3(CLBLM_R_X3Y116_SLICE_X3Y116_AO6),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(RIOB33_X105Y131_IOB_X1Y132_I),
.O5(CLBLM_R_X3Y109_SLICE_X2Y109_BO5),
.O6(CLBLM_R_X3Y109_SLICE_X2Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5a0f5a0eeee4444)
  ) CLBLM_R_X3Y109_SLICE_X2Y109_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X3Y115_SLICE_X2Y115_AQ),
.I2(CLBLL_L_X4Y109_SLICE_X4Y109_BQ),
.I3(CLBLL_L_X4Y113_SLICE_X4Y113_BQ),
.I4(CLBLM_R_X3Y107_SLICE_X3Y107_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y109_SLICE_X2Y109_AO5),
.O6(CLBLM_R_X3Y109_SLICE_X2Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55ff00fff5fff0)
  ) CLBLM_R_X3Y109_SLICE_X3Y109_DLUT (
.I0(CLBLL_L_X2Y109_SLICE_X0Y109_AO6),
.I1(1'b1),
.I2(CLBLL_L_X4Y112_SLICE_X4Y112_BQ),
.I3(CLBLM_R_X3Y109_SLICE_X3Y109_CO6),
.I4(LIOB33_X0Y65_IOB_X0Y66_I),
.I5(CLBLL_L_X2Y110_SLICE_X0Y110_BO5),
.O5(CLBLM_R_X3Y109_SLICE_X3Y109_DO5),
.O6(CLBLM_R_X3Y109_SLICE_X3Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbbfbbbb000f0000)
  ) CLBLM_R_X3Y109_SLICE_X3Y109_CLUT (
.I0(RIOB33_X105Y129_IOB_X1Y129_I),
.I1(RIOB33_X105Y137_IOB_X1Y137_I),
.I2(CLBLL_L_X2Y114_SLICE_X0Y114_AO5),
.I3(CLBLL_L_X2Y112_SLICE_X0Y112_AO5),
.I4(CLBLM_R_X5Y112_SLICE_X7Y112_DQ),
.I5(CLBLM_R_X5Y107_SLICE_X7Y107_BQ),
.O5(CLBLM_R_X3Y109_SLICE_X3Y109_CO5),
.O6(CLBLM_R_X3Y109_SLICE_X3Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hababbbabaaaabbaa)
  ) CLBLM_R_X3Y109_SLICE_X3Y109_BLUT (
.I0(CLBLM_R_X3Y107_SLICE_X3Y107_BO5),
.I1(CLBLL_L_X2Y114_SLICE_X0Y114_AO5),
.I2(CLBLL_L_X2Y112_SLICE_X0Y112_AO5),
.I3(LIOB33_X0Y65_IOB_X0Y66_I),
.I4(CLBLL_L_X2Y112_SLICE_X0Y112_AO6),
.I5(CLBLM_R_X5Y112_SLICE_X7Y112_DQ),
.O5(CLBLM_R_X3Y109_SLICE_X3Y109_BO5),
.O6(CLBLM_R_X3Y109_SLICE_X3Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffefffefffffffe)
  ) CLBLM_R_X3Y109_SLICE_X3Y109_ALUT (
.I0(CLBLM_R_X3Y112_SLICE_X3Y112_CO6),
.I1(CLBLM_R_X3Y109_SLICE_X2Y109_BO6),
.I2(CLBLM_R_X3Y108_SLICE_X3Y108_BO6),
.I3(CLBLM_R_X3Y109_SLICE_X3Y109_BO6),
.I4(RIOB33_X105Y111_IOB_X1Y111_I),
.I5(CLBLL_L_X2Y111_SLICE_X1Y111_BO5),
.O5(CLBLM_R_X3Y109_SLICE_X3Y109_AO5),
.O6(CLBLM_R_X3Y109_SLICE_X3Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffeeeeeefe)
  ) CLBLM_R_X3Y110_SLICE_X2Y110_DLUT (
.I0(CLBLL_L_X4Y109_SLICE_X5Y109_BO6),
.I1(CLBLM_R_X3Y111_SLICE_X2Y111_DO6),
.I2(CLBLL_L_X2Y111_SLICE_X1Y111_AO5),
.I3(CLBLL_L_X2Y110_SLICE_X1Y110_CO6),
.I4(CLBLM_R_X3Y112_SLICE_X2Y112_DO6),
.I5(CLBLL_L_X4Y110_SLICE_X5Y110_DO6),
.O5(CLBLM_R_X3Y110_SLICE_X2Y110_DO5),
.O6(CLBLM_R_X3Y110_SLICE_X2Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffdfffffff)
  ) CLBLM_R_X3Y110_SLICE_X2Y110_CLUT (
.I0(CLBLM_R_X3Y110_SLICE_X2Y110_AO6),
.I1(CLBLL_L_X2Y110_SLICE_X1Y110_CO6),
.I2(CLBLM_R_X3Y112_SLICE_X3Y112_BO5),
.I3(CLBLL_L_X2Y108_SLICE_X1Y108_AO5),
.I4(CLBLL_L_X2Y111_SLICE_X1Y111_AO5),
.I5(CLBLL_L_X2Y112_SLICE_X1Y112_AO6),
.O5(CLBLM_R_X3Y110_SLICE_X2Y110_CO5),
.O6(CLBLM_R_X3Y110_SLICE_X2Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_R_X3Y110_SLICE_X2Y110_BLUT (
.I0(CLBLL_L_X2Y111_SLICE_X1Y111_DO6),
.I1(CLBLM_R_X3Y108_SLICE_X2Y108_DO6),
.I2(CLBLM_R_X3Y110_SLICE_X3Y110_DO6),
.I3(CLBLM_R_X3Y110_SLICE_X2Y110_DO6),
.I4(CLBLL_L_X2Y112_SLICE_X1Y112_BO6),
.I5(CLBLM_R_X3Y109_SLICE_X2Y109_CO6),
.O5(CLBLM_R_X3Y110_SLICE_X2Y110_BO5),
.O6(CLBLM_R_X3Y110_SLICE_X2Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffeffffffffffffb)
  ) CLBLM_R_X3Y110_SLICE_X2Y110_ALUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(RIOB33_X105Y133_IOB_X1Y134_I),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(CLBLL_L_X2Y114_SLICE_X0Y114_AO6),
.I4(RIOB33_X105Y133_IOB_X1Y133_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y110_SLICE_X2Y110_AO5),
.O6(CLBLM_R_X3Y110_SLICE_X2Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffff3fffffffb)
  ) CLBLM_R_X3Y110_SLICE_X3Y110_DLUT (
.I0(CLBLM_R_X5Y115_SLICE_X6Y115_AQ),
.I1(CLBLL_L_X2Y109_SLICE_X1Y109_CO6),
.I2(CLBLM_R_X3Y109_SLICE_X3Y109_DO6),
.I3(CLBLL_L_X4Y109_SLICE_X4Y109_DO6),
.I4(CLBLM_R_X3Y111_SLICE_X3Y111_DO6),
.I5(CLBLL_L_X2Y110_SLICE_X0Y110_CO5),
.O5(CLBLM_R_X3Y110_SLICE_X3Y110_DO5),
.O6(CLBLM_R_X3Y110_SLICE_X3Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffff3fbf0fa)
  ) CLBLM_R_X3Y110_SLICE_X3Y110_CLUT (
.I0(CLBLM_R_X7Y109_SLICE_X8Y109_BQ),
.I1(CLBLM_R_X3Y112_SLICE_X3Y112_BO6),
.I2(CLBLM_R_X3Y111_SLICE_X3Y111_CO6),
.I3(CLBLL_L_X2Y110_SLICE_X0Y110_BO6),
.I4(CLBLM_R_X5Y114_SLICE_X7Y114_AQ),
.I5(CLBLM_R_X3Y110_SLICE_X3Y110_BO6),
.O5(CLBLM_R_X3Y110_SLICE_X3Y110_CO5),
.O6(CLBLM_R_X3Y110_SLICE_X3Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000110020203120)
  ) CLBLM_R_X3Y110_SLICE_X3Y110_BLUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(CLBLL_L_X2Y110_SLICE_X0Y110_AO5),
.I2(RIOB33_X105Y109_IOB_X1Y110_I),
.I3(CLBLM_R_X5Y109_SLICE_X6Y109_BQ),
.I4(CLBLM_R_X3Y116_SLICE_X3Y116_AO6),
.I5(CLBLL_L_X2Y114_SLICE_X0Y114_AO6),
.O5(CLBLM_R_X3Y110_SLICE_X3Y110_BO5),
.O6(CLBLM_R_X3Y110_SLICE_X3Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffcfffffffe)
  ) CLBLM_R_X3Y110_SLICE_X3Y110_ALUT (
.I0(CLBLL_L_X2Y109_SLICE_X1Y109_BO6),
.I1(CLBLL_L_X4Y110_SLICE_X5Y110_CO6),
.I2(CLBLL_L_X4Y110_SLICE_X4Y110_DO6),
.I3(CLBLM_R_X3Y114_SLICE_X3Y114_AO6),
.I4(CLBLL_L_X4Y110_SLICE_X5Y110_BO6),
.I5(CLBLM_R_X3Y112_SLICE_X2Y112_DO6),
.O5(CLBLM_R_X3Y110_SLICE_X3Y110_AO5),
.O6(CLBLM_R_X3Y110_SLICE_X3Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_R_X3Y111_SLICE_X2Y111_DLUT (
.I0(CLBLL_L_X2Y111_SLICE_X0Y111_CO6),
.I1(CLBLM_R_X3Y107_SLICE_X2Y107_BO6),
.I2(CLBLM_R_X3Y112_SLICE_X2Y112_BO6),
.I3(CLBLM_R_X3Y107_SLICE_X2Y107_CO6),
.I4(CLBLM_R_X3Y113_SLICE_X2Y113_DO6),
.I5(CLBLM_R_X3Y115_SLICE_X2Y115_DO6),
.O5(CLBLM_R_X3Y111_SLICE_X2Y111_DO5),
.O6(CLBLM_R_X3Y111_SLICE_X2Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffaaffffffae)
  ) CLBLM_R_X3Y111_SLICE_X2Y111_CLUT (
.I0(CLBLM_R_X3Y115_SLICE_X2Y115_CO6),
.I1(CLBLL_L_X2Y111_SLICE_X1Y111_AO5),
.I2(CLBLM_R_X3Y112_SLICE_X2Y112_DO6),
.I3(CLBLL_L_X4Y111_SLICE_X5Y111_DO6),
.I4(CLBLL_L_X4Y111_SLICE_X4Y111_DO6),
.I5(CLBLL_L_X2Y110_SLICE_X1Y110_CO6),
.O5(CLBLM_R_X3Y111_SLICE_X2Y111_CO5),
.O6(CLBLM_R_X3Y111_SLICE_X2Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffddfffdffccfffc)
  ) CLBLM_R_X3Y111_SLICE_X2Y111_BLUT (
.I0(CLBLM_R_X3Y112_SLICE_X2Y112_AO5),
.I1(CLBLM_R_X3Y111_SLICE_X3Y111_BO6),
.I2(CLBLM_R_X5Y113_SLICE_X7Y113_AQ),
.I3(CLBLL_L_X2Y111_SLICE_X0Y111_AO6),
.I4(CLBLL_L_X2Y110_SLICE_X0Y110_BO5),
.I5(CLBLL_L_X4Y108_SLICE_X4Y108_AQ),
.O5(CLBLM_R_X3Y111_SLICE_X2Y111_BO5),
.O6(CLBLM_R_X3Y111_SLICE_X2Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0caeffff0cae0cae)
  ) CLBLM_R_X3Y111_SLICE_X2Y111_ALUT (
.I0(CLBLM_R_X5Y106_SLICE_X7Y106_AQ),
.I1(RIOB33_X105Y113_IOB_X1Y113_I),
.I2(CLBLL_L_X2Y111_SLICE_X1Y111_BO5),
.I3(CLBLL_L_X2Y108_SLICE_X1Y108_AO5),
.I4(CLBLL_L_X2Y110_SLICE_X0Y110_BO6),
.I5(CLBLL_L_X4Y111_SLICE_X4Y111_BQ),
.O5(CLBLM_R_X3Y111_SLICE_X2Y111_AO5),
.O6(CLBLM_R_X3Y111_SLICE_X2Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h77335500f7f3f5f0)
  ) CLBLM_R_X3Y111_SLICE_X3Y111_DLUT (
.I0(CLBLM_R_X3Y110_SLICE_X2Y110_AO5),
.I1(CLBLL_L_X2Y111_SLICE_X1Y111_BO5),
.I2(CLBLM_R_X5Y112_SLICE_X6Y112_BQ),
.I3(CLBLM_R_X5Y110_SLICE_X6Y110_CQ),
.I4(RIOB33_X105Y111_IOB_X1Y111_I),
.I5(CLBLL_L_X2Y111_SLICE_X1Y111_AO6),
.O5(CLBLM_R_X3Y111_SLICE_X3Y111_DO5),
.O6(CLBLM_R_X3Y111_SLICE_X3Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000100000)
  ) CLBLM_R_X3Y111_SLICE_X3Y111_CLUT (
.I0(CLBLM_R_X3Y116_SLICE_X3Y116_AO6),
.I1(RIOB33_X105Y133_IOB_X1Y134_I),
.I2(RIOB33_X105Y133_IOB_X1Y133_I),
.I3(RIOB33_X105Y131_IOB_X1Y132_I),
.I4(CLBLM_L_X8Y110_SLICE_X11Y110_AQ),
.I5(RIOB33_X105Y131_IOB_X1Y131_I),
.O5(CLBLM_R_X3Y111_SLICE_X3Y111_CO5),
.O6(CLBLM_R_X3Y111_SLICE_X3Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000ff101010)
  ) CLBLM_R_X3Y111_SLICE_X3Y111_BLUT (
.I0(CLBLL_L_X2Y114_SLICE_X0Y114_AO5),
.I1(CLBLM_R_X3Y115_SLICE_X3Y115_AO6),
.I2(CLBLM_R_X5Y114_SLICE_X6Y114_AQ),
.I3(CLBLL_L_X4Y110_SLICE_X4Y110_C5Q),
.I4(CLBLL_L_X2Y107_SLICE_X1Y107_AO6),
.I5(RIOB33_X105Y131_IOB_X1Y132_I),
.O5(CLBLM_R_X3Y111_SLICE_X3Y111_BO5),
.O6(CLBLM_R_X3Y111_SLICE_X3Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0c0d5c0c0)
  ) CLBLM_R_X3Y111_SLICE_X3Y111_ALUT (
.I0(CLBLL_L_X2Y114_SLICE_X0Y114_AO5),
.I1(CLBLL_L_X4Y110_SLICE_X4Y110_CQ),
.I2(CLBLL_L_X2Y107_SLICE_X1Y107_AO6),
.I3(CLBLM_R_X3Y115_SLICE_X3Y115_AO6),
.I4(CLBLM_R_X5Y115_SLICE_X7Y115_BQ),
.I5(RIOB33_X105Y131_IOB_X1Y132_I),
.O5(CLBLM_R_X3Y111_SLICE_X3Y111_AO5),
.O6(CLBLM_R_X3Y111_SLICE_X3Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f2f0f2fffffffff)
  ) CLBLM_R_X3Y112_SLICE_X2Y112_DLUT (
.I0(RIOB33_X105Y135_IOB_X1Y136_I),
.I1(CLBLL_L_X26Y136_SLICE_X38Y136_AO6),
.I2(CLBLM_R_X3Y112_SLICE_X3Y112_BO5),
.I3(CLBLL_L_X2Y109_SLICE_X0Y109_AO5),
.I4(1'b1),
.I5(CLBLL_L_X2Y108_SLICE_X1Y108_AO5),
.O5(CLBLM_R_X3Y112_SLICE_X2Y112_DO5),
.O6(CLBLM_R_X3Y112_SLICE_X2Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0fff00ffafffaa)
  ) CLBLM_R_X3Y112_SLICE_X2Y112_CLUT (
.I0(CLBLM_R_X5Y106_SLICE_X7Y106_AQ),
.I1(1'b1),
.I2(CLBLM_R_X3Y112_SLICE_X3Y112_BO6),
.I3(CLBLM_R_X3Y113_SLICE_X2Y113_AO6),
.I4(CLBLM_R_X7Y115_SLICE_X9Y115_AQ),
.I5(CLBLL_L_X2Y108_SLICE_X1Y108_AO5),
.O5(CLBLM_R_X3Y112_SLICE_X2Y112_CO5),
.O6(CLBLM_R_X3Y112_SLICE_X2Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000005410)
  ) CLBLM_R_X3Y112_SLICE_X2Y112_BLUT (
.I0(RIOB33_X105Y135_IOB_X1Y135_I),
.I1(RIOB33_X105Y135_IOB_X1Y136_I),
.I2(CLBLM_L_X8Y109_SLICE_X10Y109_AQ),
.I3(RIOB33_X105Y109_IOB_X1Y109_I),
.I4(CLBLL_L_X26Y136_SLICE_X38Y136_AO6),
.I5(CLBLL_L_X2Y112_SLICE_X0Y112_AO6),
.O5(CLBLM_R_X3Y112_SLICE_X2Y112_BO5),
.O6(CLBLM_R_X3Y112_SLICE_X2Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hafffffffdfffffff)
  ) CLBLM_R_X3Y112_SLICE_X2Y112_ALUT (
.I0(RIOB33_X105Y131_IOB_X1Y132_I),
.I1(CLBLL_L_X2Y114_SLICE_X0Y114_AO6),
.I2(RIOB33_X105Y133_IOB_X1Y134_I),
.I3(RIOB33_X105Y133_IOB_X1Y133_I),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y112_SLICE_X2Y112_AO5),
.O6(CLBLM_R_X3Y112_SLICE_X2Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y112_SLICE_X3Y112_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y112_SLICE_X3Y112_AO6),
.Q(CLBLM_R_X3Y112_SLICE_X3Y112_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y112_SLICE_X3Y112_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y112_SLICE_X3Y112_DO5),
.O6(CLBLM_R_X3Y112_SLICE_X3Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000c0000000a)
  ) CLBLM_R_X3Y112_SLICE_X3Y112_CLUT (
.I0(CLBLM_R_X5Y112_SLICE_X6Y112_BQ),
.I1(CLBLM_R_X5Y110_SLICE_X6Y110_CQ),
.I2(RIOB33_X105Y135_IOB_X1Y135_I),
.I3(CLBLL_L_X26Y136_SLICE_X38Y136_AO6),
.I4(CLBLL_L_X2Y112_SLICE_X0Y112_AO5),
.I5(RIOB33_X105Y135_IOB_X1Y136_I),
.O5(CLBLM_R_X3Y112_SLICE_X3Y112_CO5),
.O6(CLBLM_R_X3Y112_SLICE_X3Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffff7ffffffdf)
  ) CLBLM_R_X3Y112_SLICE_X3Y112_BLUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(RIOB33_X105Y133_IOB_X1Y133_I),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(RIOB33_X105Y133_IOB_X1Y134_I),
.I4(CLBLM_R_X3Y116_SLICE_X3Y116_AO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y112_SLICE_X3Y112_BO5),
.O6(CLBLM_R_X3Y112_SLICE_X3Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00fcf0fcf0)
  ) CLBLM_R_X3Y112_SLICE_X3Y112_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X3Y112_SLICE_X3Y112_AQ),
.I3(CLBLM_R_X11Y105_SLICE_X14Y105_CQ),
.I4(1'b1),
.I5(CLBLL_L_X4Y108_SLICE_X4Y108_CO6),
.O5(CLBLM_R_X3Y112_SLICE_X3Y112_AO5),
.O6(CLBLM_R_X3Y112_SLICE_X3Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0002000233330002)
  ) CLBLM_R_X3Y113_SLICE_X2Y113_DLUT (
.I0(CLBLM_R_X3Y112_SLICE_X3Y112_AQ),
.I1(CLBLL_L_X2Y114_SLICE_X0Y114_AO5),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(CLBLM_R_X3Y115_SLICE_X3Y115_AO5),
.I4(LIOB33_X0Y63_IOB_X0Y63_I),
.I5(CLBLL_L_X2Y112_SLICE_X0Y112_AO6),
.O5(CLBLM_R_X3Y113_SLICE_X2Y113_DO5),
.O6(CLBLM_R_X3Y113_SLICE_X2Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0002000200030000)
  ) CLBLM_R_X3Y113_SLICE_X2Y113_CLUT (
.I0(CLBLM_R_X3Y113_SLICE_X3Y113_AQ),
.I1(CLBLL_L_X2Y114_SLICE_X0Y114_AO5),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(CLBLL_L_X2Y112_SLICE_X1Y112_DO6),
.I4(CLBLM_R_X5Y110_SLICE_X6Y110_DQ),
.I5(RIOB33_X105Y131_IOB_X1Y131_I),
.O5(CLBLM_R_X3Y113_SLICE_X2Y113_CO5),
.O6(CLBLM_R_X3Y113_SLICE_X2Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff04ff0404)
  ) CLBLM_R_X3Y113_SLICE_X2Y113_BLUT (
.I0(CLBLL_L_X2Y114_SLICE_X0Y114_AO5),
.I1(CLBLL_L_X4Y114_SLICE_X4Y114_AQ),
.I2(CLBLM_R_X3Y112_SLICE_X2Y112_AO6),
.I3(CLBLL_L_X2Y110_SLICE_X0Y110_AO5),
.I4(CLBLL_L_X2Y113_SLICE_X1Y113_BO6),
.I5(CLBLM_R_X3Y114_SLICE_X2Y114_CO6),
.O5(CLBLM_R_X3Y113_SLICE_X2Y113_BO5),
.O6(CLBLM_R_X3Y113_SLICE_X2Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000003100000020)
  ) CLBLM_R_X3Y113_SLICE_X2Y113_ALUT (
.I0(RIOB33_X105Y135_IOB_X1Y136_I),
.I1(CLBLL_L_X26Y136_SLICE_X38Y136_AO6),
.I2(RIOB33_X105Y113_IOB_X1Y113_I),
.I3(CLBLL_L_X2Y112_SLICE_X0Y112_AO6),
.I4(RIOB33_X105Y135_IOB_X1Y135_I),
.I5(CLBLL_L_X4Y111_SLICE_X4Y111_BQ),
.O5(CLBLM_R_X3Y113_SLICE_X2Y113_AO5),
.O6(CLBLM_R_X3Y113_SLICE_X2Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y113_SLICE_X3Y113_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y113_SLICE_X3Y113_AO6),
.Q(CLBLM_R_X3Y113_SLICE_X3Y113_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffdfffc)
  ) CLBLM_R_X3Y113_SLICE_X3Y113_DLUT (
.I0(CLBLM_R_X3Y110_SLICE_X2Y110_AO5),
.I1(CLBLL_L_X4Y113_SLICE_X4Y113_DO6),
.I2(CLBLM_R_X5Y113_SLICE_X6Y113_DO6),
.I3(CLBLM_R_X3Y113_SLICE_X3Y113_CO6),
.I4(CLBLM_R_X5Y113_SLICE_X6Y113_CQ),
.I5(CLBLM_R_X3Y113_SLICE_X3Y113_BO6),
.O5(CLBLM_R_X3Y113_SLICE_X3Y113_DO5),
.O6(CLBLM_R_X3Y113_SLICE_X3Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0100010033330100)
  ) CLBLM_R_X3Y113_SLICE_X3Y113_CLUT (
.I0(CLBLM_R_X3Y115_SLICE_X3Y115_AO6),
.I1(CLBLL_L_X2Y114_SLICE_X0Y114_AO6),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(CLBLM_R_X5Y109_SLICE_X7Y109_B5Q),
.I4(RIOB33_X105Y105_IOB_X1Y106_I),
.I5(CLBLL_L_X2Y112_SLICE_X0Y112_AO6),
.O5(CLBLM_R_X3Y113_SLICE_X3Y113_CO5),
.O6(CLBLM_R_X3Y113_SLICE_X3Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0404040404ff0404)
  ) CLBLM_R_X3Y113_SLICE_X3Y113_BLUT (
.I0(CLBLL_L_X2Y112_SLICE_X0Y112_AO5),
.I1(CLBLM_R_X5Y112_SLICE_X7Y112_BQ),
.I2(CLBLM_R_X3Y116_SLICE_X3Y116_AO6),
.I3(CLBLL_L_X2Y114_SLICE_X0Y114_AO6),
.I4(RIOB33_X105Y113_IOB_X1Y114_I),
.I5(CLBLL_L_X2Y109_SLICE_X0Y109_AO5),
.O5(CLBLM_R_X3Y113_SLICE_X3Y113_BO5),
.O6(CLBLM_R_X3Y113_SLICE_X3Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdecc1200fccc3000)
  ) CLBLM_R_X3Y113_SLICE_X3Y113_ALUT (
.I0(CLBLM_R_X3Y114_SLICE_X2Y114_BQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X3Y113_SLICE_X3Y113_AQ),
.I3(CLBLL_L_X4Y113_SLICE_X4Y113_CO6),
.I4(CLBLM_R_X3Y112_SLICE_X3Y112_AQ),
.I5(CLBLL_L_X4Y111_SLICE_X5Y111_BO6),
.O5(CLBLM_R_X3Y113_SLICE_X3Y113_AO5),
.O6(CLBLM_R_X3Y113_SLICE_X3Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y114_SLICE_X2Y114_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y114_SLICE_X2Y114_AO6),
.Q(CLBLM_R_X3Y114_SLICE_X2Y114_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y114_SLICE_X2Y114_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y114_SLICE_X2Y114_BO6),
.Q(CLBLM_R_X3Y114_SLICE_X2Y114_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaeeaaaafafe)
  ) CLBLM_R_X3Y114_SLICE_X2Y114_DLUT (
.I0(CLBLM_R_X3Y114_SLICE_X2Y114_CO5),
.I1(CLBLL_L_X4Y114_SLICE_X4Y114_CQ),
.I2(LIOB33_X0Y65_IOB_X0Y65_I),
.I3(CLBLL_L_X2Y112_SLICE_X0Y112_AO5),
.I4(CLBLL_L_X2Y114_SLICE_X0Y114_AO5),
.I5(CLBLL_L_X2Y112_SLICE_X0Y112_AO6),
.O5(CLBLM_R_X3Y114_SLICE_X2Y114_DO5),
.O6(CLBLM_R_X3Y114_SLICE_X2Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbbb0000b0b0b0b0)
  ) CLBLM_R_X3Y114_SLICE_X2Y114_CLUT (
.I0(RIOB33_X105Y129_IOB_X1Y129_I),
.I1(RIOB33_X105Y137_IOB_X1Y137_I),
.I2(CLBLL_L_X4Y115_SLICE_X5Y115_A5Q),
.I3(1'b1),
.I4(CLBLL_L_X4Y110_SLICE_X5Y110_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y114_SLICE_X2Y114_CO5),
.O6(CLBLM_R_X3Y114_SLICE_X2Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hb1a0b1a0e4a0e4a0)
  ) CLBLM_R_X3Y114_SLICE_X2Y114_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLL_L_X4Y111_SLICE_X5Y111_BO6),
.I2(CLBLM_R_X3Y114_SLICE_X2Y114_AQ),
.I3(CLBLL_L_X4Y113_SLICE_X4Y113_CO6),
.I4(1'b1),
.I5(CLBLM_R_X3Y114_SLICE_X2Y114_BQ),
.O5(CLBLM_R_X3Y114_SLICE_X2Y114_BO5),
.O6(CLBLM_R_X3Y114_SLICE_X2Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc5500ccccf000)
  ) CLBLM_R_X3Y114_SLICE_X2Y114_ALUT (
.I0(CLBLM_R_X3Y115_SLICE_X2Y115_AO5),
.I1(CLBLM_R_X7Y106_SLICE_X9Y106_BQ),
.I2(CLBLM_R_X3Y114_SLICE_X2Y114_AQ),
.I3(CLBLL_L_X4Y113_SLICE_X4Y113_CO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLL_L_X4Y114_SLICE_X5Y114_BO6),
.O5(CLBLM_R_X3Y114_SLICE_X2Y114_AO5),
.O6(CLBLM_R_X3Y114_SLICE_X2Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000005050dcdc)
  ) CLBLM_R_X3Y114_SLICE_X3Y114_DLUT (
.I0(CLBLL_L_X2Y109_SLICE_X0Y109_AO5),
.I1(CLBLM_R_X7Y106_SLICE_X9Y106_CQ),
.I2(RIOB33_X105Y115_IOB_X1Y116_I),
.I3(1'b1),
.I4(CLBLL_L_X2Y112_SLICE_X0Y112_AO5),
.I5(CLBLL_L_X2Y114_SLICE_X0Y114_AO6),
.O5(CLBLM_R_X3Y114_SLICE_X3Y114_DO5),
.O6(CLBLM_R_X3Y114_SLICE_X3Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000f000c0c0f0c)
  ) CLBLM_R_X3Y114_SLICE_X3Y114_CLUT (
.I0(1'b1),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLL_L_X2Y114_SLICE_X0Y114_AO5),
.I3(CLBLL_L_X4Y115_SLICE_X5Y115_CQ),
.I4(CLBLL_L_X2Y112_SLICE_X0Y112_AO5),
.I5(CLBLL_L_X2Y112_SLICE_X0Y112_AO6),
.O5(CLBLM_R_X3Y114_SLICE_X3Y114_CO5),
.O6(CLBLM_R_X3Y114_SLICE_X3Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000200000000000)
  ) CLBLM_R_X3Y114_SLICE_X3Y114_BLUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(CLBLL_L_X2Y114_SLICE_X0Y114_AO6),
.I2(RIOB33_X105Y133_IOB_X1Y133_I),
.I3(RIOB33_X105Y107_IOB_X1Y108_I),
.I4(RIOB33_X105Y133_IOB_X1Y134_I),
.I5(RIOB33_X105Y131_IOB_X1Y132_I),
.O5(CLBLM_R_X3Y114_SLICE_X3Y114_BO5),
.O6(CLBLM_R_X3Y114_SLICE_X3Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_R_X3Y114_SLICE_X3Y114_ALUT (
.I0(CLBLM_R_X3Y114_SLICE_X3Y114_DO6),
.I1(CLBLM_R_X3Y115_SLICE_X3Y115_DO6),
.I2(CLBLM_R_X3Y115_SLICE_X3Y115_CO6),
.I3(CLBLM_R_X3Y114_SLICE_X3Y114_BO6),
.I4(CLBLM_R_X3Y114_SLICE_X3Y114_CO6),
.I5(CLBLL_L_X4Y114_SLICE_X4Y114_DO6),
.O5(CLBLM_R_X3Y114_SLICE_X3Y114_AO5),
.O6(CLBLM_R_X3Y114_SLICE_X3Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y115_SLICE_X2Y115_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y115_SLICE_X2Y115_AO6),
.Q(CLBLM_R_X3Y115_SLICE_X2Y115_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000200020002)
  ) CLBLM_R_X3Y115_SLICE_X2Y115_DLUT (
.I0(CLBLM_R_X3Y114_SLICE_X2Y114_AQ),
.I1(CLBLM_R_X3Y115_SLICE_X3Y115_AO6),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(CLBLL_L_X2Y114_SLICE_X0Y114_AO5),
.I4(CLBLL_L_X4Y115_SLICE_X5Y115_AQ),
.I5(CLBLL_L_X2Y107_SLICE_X1Y107_AO6),
.O5(CLBLM_R_X3Y115_SLICE_X2Y115_DO5),
.O6(CLBLM_R_X3Y115_SLICE_X2Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_R_X3Y115_SLICE_X2Y115_CLUT (
.I0(CLBLL_L_X4Y115_SLICE_X4Y115_AO6),
.I1(CLBLL_L_X2Y114_SLICE_X0Y114_BO6),
.I2(CLBLM_R_X3Y115_SLICE_X3Y115_BO6),
.I3(CLBLM_R_X3Y113_SLICE_X2Y113_CO6),
.I4(CLBLM_R_X3Y116_SLICE_X2Y116_AO6),
.I5(CLBLM_R_X3Y115_SLICE_X2Y115_BO6),
.O5(CLBLM_R_X3Y115_SLICE_X2Y115_CO5),
.O6(CLBLM_R_X3Y115_SLICE_X2Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0080000000000000)
  ) CLBLM_R_X3Y115_SLICE_X2Y115_BLUT (
.I0(RIOB33_X105Y131_IOB_X1Y132_I),
.I1(RIOB33_X105Y133_IOB_X1Y133_I),
.I2(RIOB33_X105Y133_IOB_X1Y134_I),
.I3(CLBLL_L_X2Y114_SLICE_X0Y114_AO6),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(CLBLL_L_X4Y111_SLICE_X4Y111_CQ),
.O5(CLBLM_R_X3Y115_SLICE_X2Y115_BO5),
.O6(CLBLM_R_X3Y115_SLICE_X2Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heaaa0000c0000000)
  ) CLBLM_R_X3Y115_SLICE_X2Y115_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X3Y114_SLICE_X2Y114_BQ),
.I2(CLBLM_R_X3Y114_SLICE_X2Y114_AQ),
.I3(CLBLM_R_X3Y113_SLICE_X3Y113_AQ),
.I4(CLBLL_L_X4Y114_SLICE_X5Y114_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y115_SLICE_X2Y115_AO5),
.O6(CLBLM_R_X3Y115_SLICE_X2Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000050d0000000c)
  ) CLBLM_R_X3Y115_SLICE_X3Y115_DLUT (
.I0(CLBLM_R_X3Y115_SLICE_X3Y115_AO6),
.I1(CLBLL_L_X4Y116_SLICE_X5Y116_A5Q),
.I2(CLBLL_L_X2Y114_SLICE_X0Y114_AO5),
.I3(CLBLM_R_X3Y115_SLICE_X3Y115_AO5),
.I4(RIOB33_X105Y131_IOB_X1Y132_I),
.I5(CLBLL_L_X4Y114_SLICE_X5Y114_AQ),
.O5(CLBLM_R_X3Y115_SLICE_X3Y115_DO5),
.O6(CLBLM_R_X3Y115_SLICE_X3Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccec000000a0)
  ) CLBLM_R_X3Y115_SLICE_X3Y115_CLUT (
.I0(LIOB33_X0Y57_IOB_X0Y57_I),
.I1(CLBLM_R_X7Y114_SLICE_X8Y114_AQ),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(CLBLL_L_X2Y114_SLICE_X0Y114_AO5),
.I4(CLBLM_R_X3Y115_SLICE_X3Y115_AO6),
.I5(CLBLL_L_X2Y107_SLICE_X1Y107_AO6),
.O5(CLBLM_R_X3Y115_SLICE_X3Y115_CO5),
.O6(CLBLM_R_X3Y115_SLICE_X3Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000ff040404)
  ) CLBLM_R_X3Y115_SLICE_X3Y115_BLUT (
.I0(RIOB33_X105Y131_IOB_X1Y132_I),
.I1(CLBLM_R_X5Y112_SLICE_X6Y112_AQ),
.I2(CLBLL_L_X2Y114_SLICE_X0Y114_AO5),
.I3(CLBLL_L_X2Y107_SLICE_X1Y107_AO6),
.I4(CLBLM_L_X8Y111_SLICE_X10Y111_A5Q),
.I5(CLBLM_R_X3Y115_SLICE_X3Y115_AO5),
.O5(CLBLM_R_X3Y115_SLICE_X3Y115_BO5),
.O6(CLBLM_R_X3Y115_SLICE_X3Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff33ffff33ffffff)
  ) CLBLM_R_X3Y115_SLICE_X3Y115_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(1'b1),
.I3(RIOB33_X105Y133_IOB_X1Y133_I),
.I4(RIOB33_X105Y133_IOB_X1Y134_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y115_SLICE_X3Y115_AO5),
.O6(CLBLM_R_X3Y115_SLICE_X3Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y116_SLICE_X2Y116_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y116_SLICE_X2Y116_DO5),
.O6(CLBLM_R_X3Y116_SLICE_X2Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y116_SLICE_X2Y116_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y116_SLICE_X2Y116_CO5),
.O6(CLBLM_R_X3Y116_SLICE_X2Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y116_SLICE_X2Y116_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y116_SLICE_X2Y116_BO5),
.O6(CLBLM_R_X3Y116_SLICE_X2Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000008000000)
  ) CLBLM_R_X3Y116_SLICE_X2Y116_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y61_I),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(CLBLL_L_X2Y114_SLICE_X0Y114_AO5),
.I3(RIOB33_X105Y131_IOB_X1Y132_I),
.I4(RIOB33_X105Y133_IOB_X1Y133_I),
.I5(RIOB33_X105Y133_IOB_X1Y134_I),
.O5(CLBLM_R_X3Y116_SLICE_X2Y116_AO5),
.O6(CLBLM_R_X3Y116_SLICE_X2Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y116_SLICE_X3Y116_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y116_SLICE_X3Y116_DO5),
.O6(CLBLM_R_X3Y116_SLICE_X3Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y116_SLICE_X3Y116_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y116_SLICE_X3Y116_CO5),
.O6(CLBLM_R_X3Y116_SLICE_X3Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y116_SLICE_X3Y116_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y116_SLICE_X3Y116_BO5),
.O6(CLBLM_R_X3Y116_SLICE_X3Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffefffffffef)
  ) CLBLM_R_X3Y116_SLICE_X3Y116_ALUT (
.I0(RIOB33_X105Y135_IOB_X1Y135_I),
.I1(RIOB33_X105Y135_IOB_X1Y136_I),
.I2(RIOB33_X105Y137_IOB_X1Y137_I),
.I3(RIOB33_X105Y129_IOB_X1Y130_I),
.I4(RIOB33_X105Y129_IOB_X1Y129_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y116_SLICE_X3Y116_AO5),
.O6(CLBLM_R_X3Y116_SLICE_X3Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y118_SLICE_X2Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y118_SLICE_X2Y118_DO5),
.O6(CLBLM_R_X3Y118_SLICE_X2Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y118_SLICE_X2Y118_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y118_SLICE_X2Y118_CO5),
.O6(CLBLM_R_X3Y118_SLICE_X2Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y118_SLICE_X2Y118_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y118_SLICE_X2Y118_BO5),
.O6(CLBLM_R_X3Y118_SLICE_X2Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y118_SLICE_X2Y118_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y118_SLICE_X2Y118_AO5),
.O6(CLBLM_R_X3Y118_SLICE_X2Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y118_SLICE_X3Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y118_SLICE_X3Y118_DO5),
.O6(CLBLM_R_X3Y118_SLICE_X3Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y118_SLICE_X3Y118_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y118_SLICE_X3Y118_CO5),
.O6(CLBLM_R_X3Y118_SLICE_X3Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y118_SLICE_X3Y118_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y118_SLICE_X3Y118_BO5),
.O6(CLBLM_R_X3Y118_SLICE_X3Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_R_X3Y118_SLICE_X3Y118_ALUT (
.I0(CLBLL_L_X4Y118_SLICE_X4Y118_A5Q),
.I1(CLBLL_L_X4Y117_SLICE_X4Y117_AQ),
.I2(CLBLL_L_X4Y118_SLICE_X4Y118_AQ),
.I3(CLBLL_L_X4Y116_SLICE_X5Y116_AQ),
.I4(CLBLL_L_X4Y117_SLICE_X4Y117_DQ),
.I5(CLBLL_L_X4Y117_SLICE_X5Y117_AQ),
.O5(CLBLM_R_X3Y118_SLICE_X3Y118_AO5),
.O6(CLBLM_R_X3Y118_SLICE_X3Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y105_SLICE_X6Y105_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y105_SLICE_X6Y105_AO6),
.Q(CLBLM_R_X5Y105_SLICE_X6Y105_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y105_SLICE_X6Y105_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y105_SLICE_X6Y105_BO6),
.Q(CLBLM_R_X5Y105_SLICE_X6Y105_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y105_SLICE_X6Y105_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y105_SLICE_X6Y105_DO5),
.O6(CLBLM_R_X5Y105_SLICE_X6Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y105_SLICE_X6Y105_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y105_SLICE_X6Y105_CO5),
.O6(CLBLM_R_X5Y105_SLICE_X6Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haeaeaeae04040404)
  ) CLBLM_R_X5Y105_SLICE_X6Y105_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLL_L_X4Y106_SLICE_X5Y106_BQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X5Y107_SLICE_X6Y107_BQ),
.O5(CLBLM_R_X5Y105_SLICE_X6Y105_BO5),
.O6(CLBLM_R_X5Y105_SLICE_X6Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccff00ccccfa50)
  ) CLBLM_R_X5Y105_SLICE_X6Y105_ALUT (
.I0(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.I1(CLBLM_R_X5Y107_SLICE_X7Y107_AQ),
.I2(CLBLM_R_X5Y105_SLICE_X6Y105_AQ),
.I3(CLBLL_L_X4Y107_SLICE_X4Y107_DQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_R_X5Y105_SLICE_X6Y105_AO5),
.O6(CLBLM_R_X5Y105_SLICE_X6Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y105_SLICE_X7Y105_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y105_SLICE_X7Y105_AO6),
.Q(CLBLM_R_X5Y105_SLICE_X7Y105_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y105_SLICE_X7Y105_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y105_SLICE_X7Y105_BO6),
.Q(CLBLM_R_X5Y105_SLICE_X7Y105_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y105_SLICE_X7Y105_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y105_SLICE_X7Y105_DO5),
.O6(CLBLM_R_X5Y105_SLICE_X7Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y105_SLICE_X7Y105_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y105_SLICE_X7Y105_CO5),
.O6(CLBLM_R_X5Y105_SLICE_X7Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa000faaaa000c)
  ) CLBLM_R_X5Y105_SLICE_X7Y105_BLUT (
.I0(CLBLM_R_X7Y105_SLICE_X8Y105_CQ),
.I1(CLBLM_R_X5Y105_SLICE_X7Y105_BQ),
.I2(CLBLM_R_X5Y106_SLICE_X7Y106_BO5),
.I3(CLBLM_L_X10Y113_SLICE_X13Y113_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X5Y107_SLICE_X7Y107_DO6),
.O5(CLBLM_R_X5Y105_SLICE_X7Y105_BO5),
.O6(CLBLM_R_X5Y105_SLICE_X7Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff005454ff005454)
  ) CLBLM_R_X5Y105_SLICE_X7Y105_ALUT (
.I0(CLBLL_L_X4Y112_SLICE_X4Y112_CO5),
.I1(CLBLL_L_X4Y106_SLICE_X5Y106_BQ),
.I2(CLBLM_R_X5Y105_SLICE_X7Y105_AQ),
.I3(CLBLM_R_X7Y105_SLICE_X9Y105_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y105_SLICE_X7Y105_AO5),
.O6(CLBLM_R_X5Y105_SLICE_X7Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y106_SLICE_X6Y106_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y106_SLICE_X6Y106_AO6),
.Q(CLBLM_R_X5Y106_SLICE_X6Y106_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y106_SLICE_X6Y106_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y106_SLICE_X6Y106_BO6),
.Q(CLBLM_R_X5Y106_SLICE_X6Y106_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y106_SLICE_X6Y106_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y106_SLICE_X6Y106_CO6),
.Q(CLBLM_R_X5Y106_SLICE_X6Y106_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y106_SLICE_X6Y106_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y106_SLICE_X6Y106_DO6),
.Q(CLBLM_R_X5Y106_SLICE_X6Y106_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc00ffcccc0000)
  ) CLBLM_R_X5Y106_SLICE_X6Y106_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y106_SLICE_X6Y106_AQ),
.I2(1'b1),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y107_SLICE_X9Y107_CQ),
.O5(CLBLM_R_X5Y106_SLICE_X6Y106_DO5),
.O6(CLBLM_R_X5Y106_SLICE_X6Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff060006ff060006)
  ) CLBLM_R_X5Y106_SLICE_X6Y106_CLUT (
.I0(CLBLM_R_X5Y106_SLICE_X7Y106_BO6),
.I1(CLBLM_R_X5Y106_SLICE_X6Y106_CQ),
.I2(CLBLM_L_X10Y113_SLICE_X13Y113_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLL_L_X4Y111_SLICE_X4Y111_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y106_SLICE_X6Y106_CO5),
.O6(CLBLM_R_X5Y106_SLICE_X6Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f055f000f044)
  ) CLBLM_R_X5Y106_SLICE_X6Y106_BLUT (
.I0(CLBLM_L_X10Y113_SLICE_X13Y113_AQ),
.I1(CLBLM_R_X5Y106_SLICE_X6Y106_BQ),
.I2(CLBLM_R_X7Y109_SLICE_X9Y109_CQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X5Y106_SLICE_X7Y106_BO6),
.I5(CLBLM_R_X5Y106_SLICE_X7Y106_BO5),
.O5(CLBLM_R_X5Y106_SLICE_X6Y106_BO5),
.O6(CLBLM_R_X5Y106_SLICE_X6Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccaaf0aaf0)
  ) CLBLM_R_X5Y106_SLICE_X6Y106_ALUT (
.I0(CLBLM_R_X7Y108_SLICE_X8Y108_CQ),
.I1(CLBLM_R_X7Y110_SLICE_X8Y110_BQ),
.I2(CLBLM_R_X5Y106_SLICE_X6Y106_AQ),
.I3(CLBLL_L_X4Y112_SLICE_X4Y112_CO5),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X5Y106_SLICE_X6Y106_AO5),
.O6(CLBLM_R_X5Y106_SLICE_X6Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y106_SLICE_X7Y106_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y106_SLICE_X7Y106_AO6),
.Q(CLBLM_R_X5Y106_SLICE_X7Y106_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff757575ff303030)
  ) CLBLM_R_X5Y106_SLICE_X7Y106_DLUT (
.I0(CLBLM_L_X8Y104_SLICE_X11Y104_AQ),
.I1(CLBLM_R_X5Y107_SLICE_X7Y107_CO5),
.I2(CLBLM_R_X3Y109_SLICE_X2Y109_CO6),
.I3(CLBLL_L_X4Y117_SLICE_X4Y117_CQ),
.I4(CLBLL_L_X2Y111_SLICE_X1Y111_DO6),
.I5(CLBLM_R_X3Y110_SLICE_X3Y110_DO6),
.O5(CLBLM_R_X5Y106_SLICE_X7Y106_DO5),
.O6(CLBLM_R_X5Y106_SLICE_X7Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h505572775055faff)
  ) CLBLM_R_X5Y106_SLICE_X7Y106_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X8Y106_SLICE_X11Y106_A5Q),
.I2(CLBLL_L_X4Y107_SLICE_X4Y107_BO5),
.I3(CLBLM_R_X3Y108_SLICE_X2Y108_DO6),
.I4(CLBLM_R_X5Y106_SLICE_X7Y106_DO6),
.I5(CLBLM_R_X3Y110_SLICE_X2Y110_DO6),
.O5(CLBLM_R_X5Y106_SLICE_X7Y106_CO5),
.O6(CLBLM_R_X5Y106_SLICE_X7Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000080800000)
  ) CLBLM_R_X5Y106_SLICE_X7Y106_BLUT (
.I0(CLBLM_R_X7Y105_SLICE_X9Y105_CQ),
.I1(CLBLM_R_X5Y105_SLICE_X7Y105_BQ),
.I2(CLBLM_R_X7Y107_SLICE_X8Y107_DO6),
.I3(CLBLM_R_X5Y106_SLICE_X6Y106_BQ),
.I4(CLBLM_L_X8Y106_SLICE_X10Y106_BQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y106_SLICE_X7Y106_BO5),
.O6(CLBLM_R_X5Y106_SLICE_X7Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffcc00ccf5cca0)
  ) CLBLM_R_X5Y106_SLICE_X7Y106_ALUT (
.I0(CLBLM_L_X8Y114_SLICE_X11Y114_B5Q),
.I1(CLBLM_L_X10Y106_SLICE_X13Y106_CQ),
.I2(CLBLM_R_X5Y106_SLICE_X7Y106_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y106_SLICE_X9Y106_AQ),
.I5(CLBLM_L_X10Y104_SLICE_X12Y104_BO6),
.O5(CLBLM_R_X5Y106_SLICE_X7Y106_AO5),
.O6(CLBLM_R_X5Y106_SLICE_X7Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y107_SLICE_X6Y107_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y107_SLICE_X6Y107_AO6),
.Q(CLBLM_R_X5Y107_SLICE_X6Y107_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y107_SLICE_X6Y107_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y107_SLICE_X6Y107_BO6),
.Q(CLBLM_R_X5Y107_SLICE_X6Y107_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y107_SLICE_X6Y107_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y107_SLICE_X6Y107_CO6),
.Q(CLBLM_R_X5Y107_SLICE_X6Y107_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y107_SLICE_X6Y107_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y107_SLICE_X6Y107_DO6),
.Q(CLBLM_R_X5Y107_SLICE_X6Y107_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffc8fffa00c800fa)
  ) CLBLM_R_X5Y107_SLICE_X6Y107_DLUT (
.I0(CLBLM_L_X8Y106_SLICE_X10Y106_BQ),
.I1(CLBLM_L_X10Y104_SLICE_X12Y104_BO6),
.I2(CLBLM_R_X5Y107_SLICE_X6Y107_DQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y114_SLICE_X11Y114_B5Q),
.I5(CLBLM_R_X5Y105_SLICE_X7Y105_BQ),
.O5(CLBLM_R_X5Y107_SLICE_X6Y107_DO5),
.O6(CLBLM_R_X5Y107_SLICE_X6Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff5a0000005a)
  ) CLBLM_R_X5Y107_SLICE_X6Y107_CLUT (
.I0(CLBLM_R_X7Y111_SLICE_X9Y111_DO6),
.I1(1'b1),
.I2(CLBLM_R_X7Y111_SLICE_X8Y111_DQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLL_L_X4Y107_SLICE_X4Y107_DQ),
.O5(CLBLM_R_X5Y107_SLICE_X6Y107_CO5),
.O6(CLBLM_R_X5Y107_SLICE_X6Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00dfdf8080)
  ) CLBLM_R_X5Y107_SLICE_X6Y107_BLUT (
.I0(CLBLM_R_X7Y105_SLICE_X8Y105_CQ),
.I1(CLBLM_R_X5Y107_SLICE_X6Y107_BQ),
.I2(CLBLL_L_X4Y110_SLICE_X4Y110_AQ),
.I3(CLBLL_L_X4Y109_SLICE_X5Y109_AQ),
.I4(CLBLM_L_X8Y106_SLICE_X10Y106_BQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X5Y107_SLICE_X6Y107_BO5),
.O6(CLBLM_R_X5Y107_SLICE_X6Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc55f0ccccf0f0)
  ) CLBLM_R_X5Y107_SLICE_X6Y107_ALUT (
.I0(CLBLL_L_X4Y108_SLICE_X5Y108_AO6),
.I1(CLBLL_L_X4Y110_SLICE_X4Y110_AQ),
.I2(CLBLM_R_X5Y107_SLICE_X6Y107_AQ),
.I3(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_R_X5Y107_SLICE_X6Y107_AO5),
.O6(CLBLM_R_X5Y107_SLICE_X6Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y107_SLICE_X7Y107_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y107_SLICE_X7Y107_BO5),
.Q(CLBLM_R_X5Y107_SLICE_X7Y107_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y107_SLICE_X7Y107_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y107_SLICE_X7Y107_AO6),
.Q(CLBLM_R_X5Y107_SLICE_X7Y107_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y107_SLICE_X7Y107_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y107_SLICE_X7Y107_BO6),
.Q(CLBLM_R_X5Y107_SLICE_X7Y107_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c000003333ffff)
  ) CLBLM_R_X5Y107_SLICE_X7Y107_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y105_SLICE_X9Y105_CQ),
.I2(CLBLM_R_X7Y107_SLICE_X8Y107_DO6),
.I3(1'b1),
.I4(CLBLM_L_X8Y106_SLICE_X10Y106_BQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y107_SLICE_X7Y107_DO5),
.O6(CLBLM_R_X5Y107_SLICE_X7Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hbaff0000cfcfffff)
  ) CLBLM_R_X5Y107_SLICE_X7Y107_CLUT (
.I0(CLBLM_L_X8Y106_SLICE_X11Y106_A5Q),
.I1(CLBLM_L_X8Y109_SLICE_X10Y109_CQ),
.I2(CLBLM_R_X5Y109_SLICE_X6Y109_CQ),
.I3(CLBLM_R_X7Y115_SLICE_X8Y115_DQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y107_SLICE_X7Y107_CO5),
.O6(CLBLM_R_X5Y107_SLICE_X7Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'heeee4444ffa0ffa0)
  ) CLBLM_R_X5Y107_SLICE_X7Y107_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X3Y110_SLICE_X3Y110_DO6),
.I2(CLBLM_R_X5Y105_SLICE_X7Y105_AQ),
.I3(CLBLM_R_X5Y108_SLICE_X7Y108_CO6),
.I4(CLBLM_L_X8Y107_SLICE_X10Y107_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y107_SLICE_X7Y107_BO5),
.O6(CLBLM_R_X5Y107_SLICE_X7Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffac80000fac8)
  ) CLBLM_R_X5Y107_SLICE_X7Y107_ALUT (
.I0(CLBLM_R_X7Y107_SLICE_X8Y107_CQ),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_R_X5Y107_SLICE_X7Y107_AQ),
.I3(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLL_L_X4Y116_SLICE_X5Y116_B5Q),
.O5(CLBLM_R_X5Y107_SLICE_X7Y107_AO5),
.O6(CLBLM_R_X5Y107_SLICE_X7Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffcfffffffc)
  ) CLBLM_R_X5Y108_SLICE_X6Y108_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y106_SLICE_X6Y106_DQ),
.I2(CLBLM_R_X7Y111_SLICE_X8Y111_DQ),
.I3(CLBLM_R_X5Y107_SLICE_X6Y107_CQ),
.I4(CLBLM_R_X5Y113_SLICE_X7Y113_BQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y108_SLICE_X6Y108_DO5),
.O6(CLBLM_R_X5Y108_SLICE_X6Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h4cff4c4cffff4c4c)
  ) CLBLM_R_X5Y108_SLICE_X6Y108_CLUT (
.I0(CLBLM_R_X5Y105_SLICE_X7Y105_BQ),
.I1(CLBLM_R_X5Y107_SLICE_X7Y107_DO5),
.I2(CLBLM_R_X5Y106_SLICE_X6Y106_BQ),
.I3(CLBLM_L_X8Y110_SLICE_X10Y110_BQ),
.I4(CLBLM_R_X7Y108_SLICE_X9Y108_BO5),
.I5(CLBLM_R_X7Y108_SLICE_X9Y108_AQ),
.O5(CLBLM_R_X5Y108_SLICE_X6Y108_CO5),
.O6(CLBLM_R_X5Y108_SLICE_X6Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbffabaf00000000)
  ) CLBLM_R_X5Y108_SLICE_X6Y108_BLUT (
.I0(CLBLL_L_X4Y108_SLICE_X5Y108_AO5),
.I1(CLBLM_R_X3Y110_SLICE_X3Y110_AO6),
.I2(CLBLM_R_X3Y111_SLICE_X2Y111_CO6),
.I3(CLBLM_R_X3Y110_SLICE_X2Y110_DO6),
.I4(CLBLL_L_X2Y110_SLICE_X1Y110_DO6),
.I5(CLBLM_R_X5Y108_SLICE_X6Y108_CO6),
.O5(CLBLM_R_X5Y108_SLICE_X6Y108_BO5),
.O6(CLBLM_R_X5Y108_SLICE_X6Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hefffffffffffffff)
  ) CLBLM_R_X5Y108_SLICE_X6Y108_ALUT (
.I0(CLBLM_R_X7Y108_SLICE_X9Y108_BO5),
.I1(CLBLM_R_X5Y107_SLICE_X7Y107_DO5),
.I2(CLBLM_L_X8Y110_SLICE_X10Y110_BQ),
.I3(CLBLM_R_X5Y106_SLICE_X6Y106_BQ),
.I4(CLBLM_L_X10Y113_SLICE_X13Y113_CQ),
.I5(CLBLM_R_X5Y106_SLICE_X6Y106_CQ),
.O5(CLBLM_R_X5Y108_SLICE_X6Y108_AO5),
.O6(CLBLM_R_X5Y108_SLICE_X6Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y108_SLICE_X7Y108_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y108_SLICE_X7Y108_AO6),
.Q(CLBLM_R_X5Y108_SLICE_X7Y108_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0008000000000000)
  ) CLBLM_R_X5Y108_SLICE_X7Y108_DLUT (
.I0(CLBLM_L_X10Y108_SLICE_X12Y108_CQ),
.I1(CLBLM_R_X7Y107_SLICE_X9Y107_CQ),
.I2(CLBLM_R_X5Y108_SLICE_X6Y108_DO6),
.I3(CLBLL_L_X4Y112_SLICE_X5Y112_DO6),
.I4(CLBLM_R_X5Y108_SLICE_X7Y108_AQ),
.I5(CLBLM_R_X5Y105_SLICE_X6Y105_BQ),
.O5(CLBLM_R_X5Y108_SLICE_X7Y108_DO5),
.O6(CLBLM_R_X5Y108_SLICE_X7Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000f078f0f0)
  ) CLBLM_R_X5Y108_SLICE_X7Y108_CLUT (
.I0(CLBLM_R_X5Y109_SLICE_X7Y109_BQ),
.I1(CLBLM_R_X5Y109_SLICE_X7Y109_DQ),
.I2(CLBLM_R_X5Y107_SLICE_X7Y107_B5Q),
.I3(CLBLM_L_X10Y104_SLICE_X12Y104_BO6),
.I4(CLBLM_R_X5Y109_SLICE_X7Y109_B5Q),
.I5(CLBLM_R_X5Y108_SLICE_X7Y108_BO6),
.O5(CLBLM_R_X5Y108_SLICE_X7Y108_CO5),
.O6(CLBLM_R_X5Y108_SLICE_X7Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff3b33ffff3b3b)
  ) CLBLM_R_X5Y108_SLICE_X7Y108_BLUT (
.I0(CLBLM_R_X7Y115_SLICE_X8Y115_DQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_L_X8Y106_SLICE_X11Y106_A5Q),
.I3(CLBLM_L_X8Y109_SLICE_X10Y109_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X5Y109_SLICE_X6Y109_CQ),
.O5(CLBLM_R_X5Y108_SLICE_X7Y108_BO5),
.O6(CLBLM_R_X5Y108_SLICE_X7Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa000faaaa0f00)
  ) CLBLM_R_X5Y108_SLICE_X7Y108_ALUT (
.I0(CLBLM_R_X5Y110_SLICE_X6Y110_B5Q),
.I1(1'b1),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X7Y108_SLICE_X8Y108_DO5),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X5Y107_SLICE_X6Y107_CQ),
.O5(CLBLM_R_X5Y108_SLICE_X7Y108_AO5),
.O6(CLBLM_R_X5Y108_SLICE_X7Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y109_SLICE_X6Y109_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y109_SLICE_X6Y109_AO6),
.Q(CLBLM_R_X5Y109_SLICE_X6Y109_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y109_SLICE_X6Y109_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y109_SLICE_X6Y109_BO6),
.Q(CLBLM_R_X5Y109_SLICE_X6Y109_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y109_SLICE_X6Y109_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y109_SLICE_X6Y109_CO6),
.Q(CLBLM_R_X5Y109_SLICE_X6Y109_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y109_SLICE_X6Y109_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y109_SLICE_X6Y109_DO6),
.Q(CLBLM_R_X5Y109_SLICE_X6Y109_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hacaca0a0acaca0a0)
  ) CLBLM_R_X5Y109_SLICE_X6Y109_DLUT (
.I0(CLBLL_L_X4Y108_SLICE_X4Y108_AQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(CLBLM_R_X7Y110_SLICE_X8Y110_BQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y109_SLICE_X6Y109_DO5),
.O6(CLBLM_R_X5Y109_SLICE_X6Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haac0aa00aa00aa00)
  ) CLBLM_R_X5Y109_SLICE_X6Y109_CLUT (
.I0(CLBLM_R_X7Y112_SLICE_X8Y112_C5Q),
.I1(CLBLM_R_X5Y107_SLICE_X7Y107_B5Q),
.I2(CLBLM_R_X5Y109_SLICE_X7Y109_B5Q),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X5Y109_SLICE_X7Y109_DQ),
.I5(CLBLM_R_X5Y109_SLICE_X7Y109_BQ),
.O5(CLBLM_R_X5Y109_SLICE_X6Y109_CO5),
.O6(CLBLM_R_X5Y109_SLICE_X6Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ccaaf0f0ccaa)
  ) CLBLM_R_X5Y109_SLICE_X6Y109_BLUT (
.I0(CLBLM_R_X5Y106_SLICE_X6Y106_DQ),
.I1(CLBLM_R_X5Y109_SLICE_X6Y109_BQ),
.I2(CLBLM_R_X11Y105_SLICE_X14Y105_C5Q),
.I3(CLBLL_L_X4Y112_SLICE_X4Y112_CO5),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y109_SLICE_X6Y109_BO5),
.O6(CLBLM_R_X5Y109_SLICE_X6Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8888bbb8bbb8bbb8)
  ) CLBLM_R_X5Y109_SLICE_X6Y109_ALUT (
.I0(CLBLM_R_X11Y117_SLICE_X15Y117_DQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X5Y109_SLICE_X6Y109_AQ),
.I3(CLBLM_R_X7Y109_SLICE_X9Y109_CQ),
.I4(CLBLL_L_X4Y110_SLICE_X4Y110_AQ),
.I5(CLBLM_R_X7Y105_SLICE_X8Y105_CQ),
.O5(CLBLM_R_X5Y109_SLICE_X6Y109_AO5),
.O6(CLBLM_R_X5Y109_SLICE_X6Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y109_SLICE_X7Y109_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y106_SLICE_X9Y106_DO5),
.Q(CLBLM_R_X5Y109_SLICE_X7Y109_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y109_SLICE_X7Y109_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y109_SLICE_X7Y109_CO6),
.Q(CLBLM_R_X5Y109_SLICE_X7Y109_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y109_SLICE_X7Y109_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y109_SLICE_X7Y109_AO6),
.Q(CLBLM_R_X5Y109_SLICE_X7Y109_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y109_SLICE_X7Y109_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y109_SLICE_X7Y109_BO6),
.Q(CLBLM_R_X5Y109_SLICE_X7Y109_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y109_SLICE_X7Y109_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y109_SLICE_X7Y109_DO6),
.Q(CLBLM_R_X5Y109_SLICE_X7Y109_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff840084ffc000c0)
  ) CLBLM_R_X5Y109_SLICE_X7Y109_DLUT (
.I0(CLBLM_R_X5Y109_SLICE_X7Y109_CO5),
.I1(CLBLM_R_X5Y107_SLICE_X7Y107_CO6),
.I2(CLBLM_R_X5Y109_SLICE_X7Y109_DQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y111_SLICE_X13Y111_AQ),
.I5(CLBLM_R_X5Y109_SLICE_X7Y109_BQ),
.O5(CLBLM_R_X5Y109_SLICE_X7Y109_DO5),
.O6(CLBLM_R_X5Y109_SLICE_X7Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0eac0d5aaaaffff)
  ) CLBLM_R_X5Y109_SLICE_X7Y109_CLUT (
.I0(CLBLM_L_X10Y104_SLICE_X12Y104_BO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X5Y114_SLICE_X7Y114_B5Q),
.I3(CLBLM_R_X5Y108_SLICE_X7Y108_BO6),
.I4(CLBLM_R_X5Y109_SLICE_X7Y109_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X5Y109_SLICE_X7Y109_CO5),
.O6(CLBLM_R_X5Y109_SLICE_X7Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc0cf303f000f000)
  ) CLBLM_R_X5Y109_SLICE_X7Y109_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y109_SLICE_X7Y109_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y109_SLICE_X10Y109_BQ),
.I4(CLBLM_R_X5Y109_SLICE_X7Y109_CO5),
.I5(CLBLM_R_X5Y107_SLICE_X7Y107_CO6),
.O5(CLBLM_R_X5Y109_SLICE_X7Y109_BO5),
.O6(CLBLM_R_X5Y109_SLICE_X7Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf101f101f202f202)
  ) CLBLM_R_X5Y109_SLICE_X7Y109_ALUT (
.I0(CLBLM_R_X7Y109_SLICE_X8Y109_CO6),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLL_L_X4Y106_SLICE_X5Y106_BQ),
.I4(1'b1),
.I5(CLBLM_R_X5Y113_SLICE_X7Y113_BQ),
.O5(CLBLM_R_X5Y109_SLICE_X7Y109_AO5),
.O6(CLBLM_R_X5Y109_SLICE_X7Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y110_SLICE_X6Y110_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y110_SLICE_X6Y110_BO5),
.Q(CLBLM_R_X5Y110_SLICE_X6Y110_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y110_SLICE_X6Y110_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y110_SLICE_X6Y110_AO6),
.Q(CLBLM_R_X5Y110_SLICE_X6Y110_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y110_SLICE_X6Y110_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y110_SLICE_X6Y110_BO6),
.Q(CLBLM_R_X5Y110_SLICE_X6Y110_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y110_SLICE_X6Y110_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y110_SLICE_X6Y110_CO6),
.Q(CLBLM_R_X5Y110_SLICE_X6Y110_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y110_SLICE_X6Y110_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y110_SLICE_X6Y110_DO6),
.Q(CLBLM_R_X5Y110_SLICE_X6Y110_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hd8ddd888d8ddd888)
  ) CLBLM_R_X5Y110_SLICE_X6Y110_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X13Y107_SLICE_X19Y107_BQ),
.I2(CLBLM_R_X5Y110_SLICE_X6Y110_DQ),
.I3(CLBLL_L_X4Y113_SLICE_X5Y113_DO6),
.I4(CLBLL_L_X4Y116_SLICE_X5Y116_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X5Y110_SLICE_X6Y110_DO5),
.O6(CLBLM_R_X5Y110_SLICE_X6Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffaf8c0000af8c)
  ) CLBLM_R_X5Y110_SLICE_X6Y110_CLUT (
.I0(CLBLM_L_X10Y104_SLICE_X12Y104_BO6),
.I1(CLBLM_R_X5Y110_SLICE_X6Y110_CQ),
.I2(CLBLM_L_X8Y114_SLICE_X11Y114_B5Q),
.I3(CLBLM_R_X5Y106_SLICE_X6Y106_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y119_SLICE_X10Y119_AQ),
.O5(CLBLM_R_X5Y110_SLICE_X6Y110_CO5),
.O6(CLBLM_R_X5Y110_SLICE_X6Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hafa0afa0cfcfc0c0)
  ) CLBLM_R_X5Y110_SLICE_X6Y110_BLUT (
.I0(CLBLM_R_X5Y110_SLICE_X6Y110_CQ),
.I1(CLBLM_R_X5Y117_SLICE_X7Y117_AQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X5Y115_SLICE_X6Y115_BQ),
.I4(CLBLL_L_X4Y107_SLICE_X4Y107_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y110_SLICE_X6Y110_BO5),
.O6(CLBLM_R_X5Y110_SLICE_X6Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0c0c0cac0)
  ) CLBLM_R_X5Y110_SLICE_X6Y110_ALUT (
.I0(CLBLM_R_X5Y105_SLICE_X7Y105_BQ),
.I1(CLBLM_R_X5Y110_SLICE_X6Y110_DQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y113_SLICE_X10Y113_D5Q),
.I4(CLBLM_R_X5Y108_SLICE_X6Y108_AO6),
.I5(CLBLM_R_X7Y108_SLICE_X9Y108_AQ),
.O5(CLBLM_R_X5Y110_SLICE_X6Y110_AO5),
.O6(CLBLM_R_X5Y110_SLICE_X6Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y110_SLICE_X7Y110_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y110_SLICE_X7Y110_BO5),
.Q(CLBLM_R_X5Y110_SLICE_X7Y110_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y110_SLICE_X7Y110_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y110_SLICE_X7Y110_AO6),
.Q(CLBLM_R_X5Y110_SLICE_X7Y110_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y110_SLICE_X7Y110_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y110_SLICE_X7Y110_BO6),
.Q(CLBLM_R_X5Y110_SLICE_X7Y110_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000fdff0000ffff)
  ) CLBLM_R_X5Y110_SLICE_X7Y110_DLUT (
.I0(CLBLM_R_X5Y111_SLICE_X7Y111_AQ),
.I1(CLBLM_R_X3Y107_SLICE_X3Y107_CO6),
.I2(CLBLM_R_X5Y115_SLICE_X7Y115_DO6),
.I3(CLBLM_R_X5Y110_SLICE_X7Y110_BQ),
.I4(CLBLM_R_X5Y110_SLICE_X7Y110_B5Q),
.I5(CLBLL_L_X4Y113_SLICE_X5Y113_BQ),
.O5(CLBLM_R_X5Y110_SLICE_X7Y110_DO5),
.O6(CLBLM_R_X5Y110_SLICE_X7Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff002000ff0000)
  ) CLBLM_R_X5Y110_SLICE_X7Y110_CLUT (
.I0(CLBLM_R_X5Y111_SLICE_X7Y111_AQ),
.I1(CLBLM_R_X5Y115_SLICE_X7Y115_CO6),
.I2(CLBLM_R_X5Y110_SLICE_X7Y110_BQ),
.I3(CLBLM_L_X8Y110_SLICE_X11Y110_BO5),
.I4(CLBLM_R_X5Y110_SLICE_X7Y110_B5Q),
.I5(CLBLL_L_X4Y113_SLICE_X5Y113_BQ),
.O5(CLBLM_R_X5Y110_SLICE_X7Y110_CO5),
.O6(CLBLM_R_X5Y110_SLICE_X7Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffa0ffa0ffffc0c0)
  ) CLBLM_R_X5Y110_SLICE_X7Y110_BLUT (
.I0(CLBLL_L_X4Y115_SLICE_X5Y115_CQ),
.I1(CLBLM_R_X5Y111_SLICE_X7Y111_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLL_L_X4Y110_SLICE_X5Y110_AO6),
.I4(CLBLM_R_X5Y110_SLICE_X7Y110_CO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y110_SLICE_X7Y110_BO5),
.O6(CLBLM_R_X5Y110_SLICE_X7Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccf0f0ccccaaaa)
  ) CLBLM_R_X5Y110_SLICE_X7Y110_ALUT (
.I0(CLBLM_R_X5Y114_SLICE_X7Y114_B5Q),
.I1(CLBLM_R_X11Y111_SLICE_X15Y111_BQ),
.I2(CLBLM_R_X5Y110_SLICE_X7Y110_AQ),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLL_L_X4Y113_SLICE_X5Y113_DO6),
.O5(CLBLM_R_X5Y110_SLICE_X7Y110_AO5),
.O6(CLBLM_R_X5Y110_SLICE_X7Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y111_SLICE_X6Y111_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y111_SLICE_X6Y111_AO6),
.Q(CLBLM_R_X5Y111_SLICE_X6Y111_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y111_SLICE_X6Y111_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y111_SLICE_X6Y111_BO6),
.Q(CLBLM_R_X5Y111_SLICE_X6Y111_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y111_SLICE_X6Y111_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y111_SLICE_X6Y111_CO6),
.Q(CLBLM_R_X5Y111_SLICE_X6Y111_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h77ff77ffffffffff)
  ) CLBLM_R_X5Y111_SLICE_X6Y111_DLUT (
.I0(CLBLM_R_X5Y111_SLICE_X7Y111_AQ),
.I1(CLBLL_L_X4Y113_SLICE_X5Y113_BQ),
.I2(1'b1),
.I3(CLBLM_R_X5Y110_SLICE_X7Y110_B5Q),
.I4(1'b1),
.I5(CLBLM_R_X5Y110_SLICE_X7Y110_BQ),
.O5(CLBLM_R_X5Y111_SLICE_X6Y111_DO5),
.O6(CLBLM_R_X5Y111_SLICE_X6Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0c03aaaa0c03)
  ) CLBLM_R_X5Y111_SLICE_X6Y111_CLUT (
.I0(CLBLM_R_X5Y109_SLICE_X6Y109_AQ),
.I1(CLBLM_R_X7Y111_SLICE_X9Y111_DO5),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_L_X10Y111_SLICE_X12Y111_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y111_SLICE_X6Y111_CO5),
.O6(CLBLM_R_X5Y111_SLICE_X6Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00fe000e00fe000e)
  ) CLBLM_R_X5Y111_SLICE_X6Y111_BLUT (
.I0(CLBLM_R_X7Y111_SLICE_X8Y111_DQ),
.I1(CLBLM_R_X5Y111_SLICE_X6Y111_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLL_L_X4Y112_SLICE_X4Y112_CO6),
.I4(CLBLL_L_X4Y116_SLICE_X4Y116_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y111_SLICE_X6Y111_BO5),
.O6(CLBLM_R_X5Y111_SLICE_X6Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaf0ccaaaacccc)
  ) CLBLM_R_X5Y111_SLICE_X6Y111_ALUT (
.I0(CLBLM_R_X5Y116_SLICE_X6Y116_CQ),
.I1(CLBLM_R_X7Y108_SLICE_X9Y108_AQ),
.I2(CLBLM_R_X5Y111_SLICE_X6Y111_AQ),
.I3(CLBLM_R_X7Y105_SLICE_X8Y105_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLL_L_X4Y110_SLICE_X4Y110_AQ),
.O5(CLBLM_R_X5Y111_SLICE_X6Y111_AO5),
.O6(CLBLM_R_X5Y111_SLICE_X6Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y111_SLICE_X7Y111_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y111_SLICE_X7Y111_AO6),
.Q(CLBLM_R_X5Y111_SLICE_X7Y111_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y111_SLICE_X7Y111_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y111_SLICE_X7Y111_BO6),
.Q(CLBLM_R_X5Y111_SLICE_X7Y111_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y111_SLICE_X7Y111_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y111_SLICE_X7Y111_CO6),
.Q(CLBLM_R_X5Y111_SLICE_X7Y111_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf7ffffffffffffff)
  ) CLBLM_R_X5Y111_SLICE_X7Y111_DLUT (
.I0(CLBLM_L_X10Y111_SLICE_X12Y111_AQ),
.I1(CLBLM_R_X7Y109_SLICE_X9Y109_DQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X5Y111_SLICE_X6Y111_CQ),
.I4(CLBLM_R_X5Y109_SLICE_X7Y109_AQ),
.I5(CLBLL_L_X4Y106_SLICE_X5Y106_BQ),
.O5(CLBLM_R_X5Y111_SLICE_X7Y111_DO5),
.O6(CLBLM_R_X5Y111_SLICE_X7Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffaaac0000aaac)
  ) CLBLM_R_X5Y111_SLICE_X7Y111_CLUT (
.I0(CLBLM_L_X8Y111_SLICE_X10Y111_DO6),
.I1(CLBLM_R_X5Y111_SLICE_X7Y111_CQ),
.I2(RIOB33_X105Y117_IOB_X1Y118_I),
.I3(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X5Y106_SLICE_X7Y106_AQ),
.O5(CLBLM_R_X5Y111_SLICE_X7Y111_CO5),
.O6(CLBLM_R_X5Y111_SLICE_X7Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff005d5dff000c0c)
  ) CLBLM_R_X5Y111_SLICE_X7Y111_BLUT (
.I0(CLBLM_R_X5Y111_SLICE_X7Y111_DO6),
.I1(CLBLM_R_X5Y111_SLICE_X7Y111_BQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_L_X12Y109_SLICE_X16Y109_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X5Y108_SLICE_X7Y108_DO6),
.O5(CLBLM_R_X5Y111_SLICE_X7Y111_BO5),
.O6(CLBLM_R_X5Y111_SLICE_X7Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00ebc3aa00fbf3)
  ) CLBLM_R_X5Y111_SLICE_X7Y111_ALUT (
.I0(CLBLM_R_X7Y118_SLICE_X8Y118_AQ),
.I1(CLBLM_R_X5Y115_SLICE_X7Y115_CO6),
.I2(CLBLM_R_X5Y111_SLICE_X7Y111_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y110_SLICE_X11Y110_BO5),
.I5(CLBLM_R_X5Y111_SLICE_X6Y111_DO6),
.O5(CLBLM_R_X5Y111_SLICE_X7Y111_AO5),
.O6(CLBLM_R_X5Y111_SLICE_X7Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y112_SLICE_X6Y112_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y112_SLICE_X6Y112_AO6),
.Q(CLBLM_R_X5Y112_SLICE_X6Y112_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y112_SLICE_X6Y112_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y112_SLICE_X6Y112_BO6),
.Q(CLBLM_R_X5Y112_SLICE_X6Y112_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y112_SLICE_X6Y112_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y112_SLICE_X6Y112_CO6),
.Q(CLBLM_R_X5Y112_SLICE_X6Y112_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00002f2200002f22)
  ) CLBLM_R_X5Y112_SLICE_X6Y112_DLUT (
.I0(CLBLM_R_X7Y114_SLICE_X9Y114_BQ),
.I1(CLBLL_L_X2Y109_SLICE_X0Y109_AO5),
.I2(CLBLL_L_X2Y112_SLICE_X0Y112_AO5),
.I3(CLBLM_R_X7Y113_SLICE_X8Y113_AQ),
.I4(CLBLM_R_X3Y116_SLICE_X3Y116_AO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y112_SLICE_X6Y112_DO5),
.O6(CLBLM_R_X5Y112_SLICE_X6Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haafaaaea00500040)
  ) CLBLM_R_X5Y112_SLICE_X6Y112_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y112_SLICE_X6Y112_CQ),
.I2(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_R_X11Y114_SLICE_X14Y114_BQ),
.I5(CLBLL_L_X4Y112_SLICE_X5Y112_AQ),
.O5(CLBLM_R_X5Y112_SLICE_X6Y112_CO5),
.O6(CLBLM_R_X5Y112_SLICE_X6Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefefcfcaaaa0000)
  ) CLBLM_R_X5Y112_SLICE_X6Y112_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y112_SLICE_X6Y112_BQ),
.I2(CLBLM_L_X8Y113_SLICE_X11Y113_AQ),
.I3(1'b1),
.I4(CLBLM_R_X13Y112_SLICE_X18Y112_AQ),
.I5(CLBLL_L_X4Y112_SLICE_X4Y112_CO6),
.O5(CLBLM_R_X5Y112_SLICE_X6Y112_BO5),
.O6(CLBLM_R_X5Y112_SLICE_X6Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff505050ff505050)
  ) CLBLM_R_X5Y112_SLICE_X6Y112_ALUT (
.I0(CLBLL_L_X4Y108_SLICE_X4Y108_CO6),
.I1(1'b1),
.I2(CLBLM_R_X5Y112_SLICE_X6Y112_AQ),
.I3(CLBLM_R_X5Y112_SLICE_X6Y112_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y112_SLICE_X6Y112_AO5),
.O6(CLBLM_R_X5Y112_SLICE_X6Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y112_SLICE_X7Y112_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y112_SLICE_X7Y112_AO6),
.Q(CLBLM_R_X5Y112_SLICE_X7Y112_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y112_SLICE_X7Y112_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y112_SLICE_X7Y112_BO6),
.Q(CLBLM_R_X5Y112_SLICE_X7Y112_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y112_SLICE_X7Y112_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y112_SLICE_X7Y112_CO6),
.Q(CLBLM_R_X5Y112_SLICE_X7Y112_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y112_SLICE_X7Y112_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y112_SLICE_X7Y112_DO6),
.Q(CLBLM_R_X5Y112_SLICE_X7Y112_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbbbbaba11111010)
  ) CLBLM_R_X5Y112_SLICE_X7Y112_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLL_L_X4Y113_SLICE_X5Y113_DO6),
.I2(CLBLM_R_X5Y112_SLICE_X7Y112_DQ),
.I3(1'b1),
.I4(CLBLM_R_X7Y115_SLICE_X8Y115_B5Q),
.I5(CLBLM_L_X12Y108_SLICE_X16Y108_DQ),
.O5(CLBLM_R_X5Y112_SLICE_X7Y112_DO5),
.O6(CLBLM_R_X5Y112_SLICE_X7Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0b1a0b1b1a0b1a0)
  ) CLBLM_R_X5Y112_SLICE_X7Y112_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X7Y112_SLICE_X8Y112_DQ),
.I3(CLBLM_R_X11Y110_SLICE_X14Y110_BO5),
.I4(1'b1),
.I5(CLBLM_R_X11Y114_SLICE_X14Y114_CQ),
.O5(CLBLM_R_X5Y112_SLICE_X7Y112_CO5),
.O6(CLBLM_R_X5Y112_SLICE_X7Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00f000ff00f000cc)
  ) CLBLM_R_X5Y112_SLICE_X7Y112_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y112_SLICE_X7Y112_BQ),
.I2(CLBLM_R_X5Y112_SLICE_X7Y112_AQ),
.I3(CLBLL_L_X4Y112_SLICE_X4Y112_CO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y111_SLICE_X9Y111_CQ),
.O5(CLBLM_R_X5Y112_SLICE_X7Y112_BO5),
.O6(CLBLM_R_X5Y112_SLICE_X7Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff005050ff00d8d8)
  ) CLBLM_R_X5Y112_SLICE_X7Y112_ALUT (
.I0(CLBLM_R_X7Y105_SLICE_X8Y105_BO5),
.I1(CLBLM_R_X3Y110_SLICE_X3Y110_AO6),
.I2(CLBLM_R_X5Y112_SLICE_X7Y112_AQ),
.I3(CLBLM_L_X10Y119_SLICE_X12Y119_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X5Y112_SLICE_X7Y112_AO5),
.O6(CLBLM_R_X5Y112_SLICE_X7Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y113_SLICE_X6Y113_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y113_SLICE_X6Y113_AO6),
.Q(CLBLM_R_X5Y113_SLICE_X6Y113_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y113_SLICE_X6Y113_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y113_SLICE_X6Y113_BO6),
.Q(CLBLM_R_X5Y113_SLICE_X6Y113_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y113_SLICE_X6Y113_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y113_SLICE_X6Y113_CO6),
.Q(CLBLM_R_X5Y113_SLICE_X6Y113_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000c0000000a0)
  ) CLBLM_R_X5Y113_SLICE_X6Y113_DLUT (
.I0(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.I1(CLBLM_R_X5Y116_SLICE_X6Y116_BQ),
.I2(RIOB33_X105Y133_IOB_X1Y133_I),
.I3(CLBLM_R_X5Y114_SLICE_X6Y114_BO6),
.I4(RIOB33_X105Y133_IOB_X1Y134_I),
.I5(RIOB33_X105Y131_IOB_X1Y131_I),
.O5(CLBLM_R_X5Y113_SLICE_X6Y113_DO5),
.O6(CLBLM_R_X5Y113_SLICE_X6Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfaeefafa50445050)
  ) CLBLM_R_X5Y113_SLICE_X6Y113_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y113_SLICE_X6Y113_CQ),
.I2(CLBLM_L_X8Y110_SLICE_X10Y110_BQ),
.I3(CLBLM_L_X10Y104_SLICE_X12Y104_BO6),
.I4(CLBLM_L_X8Y114_SLICE_X11Y114_B5Q),
.I5(CLBLL_L_X4Y116_SLICE_X5Y116_A5Q),
.O5(CLBLM_R_X5Y113_SLICE_X6Y113_CO5),
.O6(CLBLM_R_X5Y113_SLICE_X6Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf1f1f2f201010202)
  ) CLBLM_R_X5Y113_SLICE_X6Y113_BLUT (
.I0(CLBLM_R_X7Y113_SLICE_X9Y113_DO6),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(CLBLM_R_X7Y112_SLICE_X9Y112_AQ),
.I5(CLBLM_R_X5Y114_SLICE_X7Y114_C5Q),
.O5(CLBLM_R_X5Y113_SLICE_X6Y113_BO5),
.O6(CLBLM_R_X5Y113_SLICE_X6Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccff00ccccaaaa)
  ) CLBLM_R_X5Y113_SLICE_X6Y113_ALUT (
.I0(CLBLM_R_X5Y113_SLICE_X6Y113_AQ),
.I1(CLBLM_R_X11Y113_SLICE_X14Y113_DQ),
.I2(1'b1),
.I3(CLBLM_L_X10Y111_SLICE_X12Y111_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLL_L_X4Y112_SLICE_X4Y112_CO5),
.O5(CLBLM_R_X5Y113_SLICE_X6Y113_AO5),
.O6(CLBLM_R_X5Y113_SLICE_X6Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y113_SLICE_X7Y113_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y113_SLICE_X7Y113_AO6),
.Q(CLBLM_R_X5Y113_SLICE_X7Y113_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y113_SLICE_X7Y113_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y113_SLICE_X7Y113_BO6),
.Q(CLBLM_R_X5Y113_SLICE_X7Y113_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8800880000000000)
  ) CLBLM_R_X5Y113_SLICE_X7Y113_DLUT (
.I0(CLBLM_R_X7Y115_SLICE_X9Y115_A5Q),
.I1(CLBLM_R_X5Y109_SLICE_X7Y109_A5Q),
.I2(1'b1),
.I3(CLBLM_R_X7Y114_SLICE_X8Y114_CQ),
.I4(1'b1),
.I5(CLBLM_L_X8Y113_SLICE_X11Y113_AQ),
.O5(CLBLM_R_X5Y113_SLICE_X7Y113_DO5),
.O6(CLBLM_R_X5Y113_SLICE_X7Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000e200000000)
  ) CLBLM_R_X5Y113_SLICE_X7Y113_CLUT (
.I0(CLBLM_L_X10Y113_SLICE_X12Y113_AQ),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(CLBLM_L_X8Y114_SLICE_X11Y114_AQ),
.I3(CLBLM_R_X5Y114_SLICE_X6Y114_BO6),
.I4(RIOB33_X105Y133_IOB_X1Y134_I),
.I5(RIOB33_X105Y133_IOB_X1Y133_I),
.O5(CLBLM_R_X5Y113_SLICE_X7Y113_CO5),
.O6(CLBLM_R_X5Y113_SLICE_X7Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00066f0f00066)
  ) CLBLM_R_X5Y113_SLICE_X7Y113_BLUT (
.I0(CLBLM_R_X7Y109_SLICE_X9Y109_DQ),
.I1(CLBLM_R_X7Y113_SLICE_X9Y113_BO6),
.I2(CLBLM_R_X5Y113_SLICE_X7Y113_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y113_SLICE_X7Y113_BO5),
.O6(CLBLM_R_X5Y113_SLICE_X7Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00fcfcff003030)
  ) CLBLM_R_X5Y113_SLICE_X7Y113_ALUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y112_SLICE_X4Y112_CO5),
.I2(CLBLM_R_X5Y113_SLICE_X7Y113_AQ),
.I3(CLBLM_L_X12Y113_SLICE_X17Y113_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y114_SLICE_X8Y114_CQ),
.O5(CLBLM_R_X5Y113_SLICE_X7Y113_AO5),
.O6(CLBLM_R_X5Y113_SLICE_X7Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y114_SLICE_X6Y114_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y114_SLICE_X6Y114_AO6),
.Q(CLBLM_R_X5Y114_SLICE_X6Y114_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffc)
  ) CLBLM_R_X5Y114_SLICE_X6Y114_DLUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y116_SLICE_X4Y116_A5Q),
.I2(CLBLM_R_X5Y114_SLICE_X7Y114_B5Q),
.I3(CLBLL_L_X4Y116_SLICE_X5Y116_B5Q),
.I4(CLBLM_R_X5Y110_SLICE_X6Y110_BQ),
.I5(CLBLM_R_X7Y113_SLICE_X9Y113_A5Q),
.O5(CLBLM_R_X5Y114_SLICE_X6Y114_DO5),
.O6(CLBLM_R_X5Y114_SLICE_X6Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h020202020202ff02)
  ) CLBLM_R_X5Y114_SLICE_X6Y114_CLUT (
.I0(CLBLM_L_X8Y114_SLICE_X10Y114_AQ),
.I1(CLBLL_L_X2Y112_SLICE_X0Y112_AO5),
.I2(CLBLM_R_X3Y116_SLICE_X3Y116_AO6),
.I3(RIOB33_X105Y117_IOB_X1Y117_I),
.I4(CLBLL_L_X2Y114_SLICE_X0Y114_AO6),
.I5(CLBLL_L_X2Y109_SLICE_X0Y109_AO5),
.O5(CLBLM_R_X5Y114_SLICE_X6Y114_CO5),
.O6(CLBLM_R_X5Y114_SLICE_X6Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffeff)
  ) CLBLM_R_X5Y114_SLICE_X6Y114_BLUT (
.I0(RIOB33_X105Y135_IOB_X1Y135_I),
.I1(RIOB33_X105Y129_IOB_X1Y130_I),
.I2(RIOB33_X105Y135_IOB_X1Y136_I),
.I3(RIOB33_X105Y137_IOB_X1Y137_I),
.I4(RIOB33_X105Y129_IOB_X1Y129_I),
.I5(RIOB33_X105Y131_IOB_X1Y132_I),
.O5(CLBLM_R_X5Y114_SLICE_X6Y114_BO5),
.O6(CLBLM_R_X5Y114_SLICE_X6Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaafcfcaaaa0000)
  ) CLBLM_R_X5Y114_SLICE_X6Y114_ALUT (
.I0(CLBLM_R_X5Y113_SLICE_X6Y113_AQ),
.I1(CLBLM_R_X7Y115_SLICE_X9Y115_B5Q),
.I2(CLBLM_R_X5Y114_SLICE_X6Y114_AQ),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLL_L_X4Y113_SLICE_X5Y113_DO6),
.O5(CLBLM_R_X5Y114_SLICE_X6Y114_AO5),
.O6(CLBLM_R_X5Y114_SLICE_X6Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y114_SLICE_X7Y114_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y114_SLICE_X7Y114_BO5),
.Q(CLBLM_R_X5Y114_SLICE_X7Y114_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y114_SLICE_X7Y114_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y114_SLICE_X7Y114_CO5),
.Q(CLBLM_R_X5Y114_SLICE_X7Y114_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y114_SLICE_X7Y114_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y114_SLICE_X7Y114_AO6),
.Q(CLBLM_R_X5Y114_SLICE_X7Y114_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y114_SLICE_X7Y114_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y114_SLICE_X7Y114_BO6),
.Q(CLBLM_R_X5Y114_SLICE_X7Y114_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y114_SLICE_X7Y114_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y114_SLICE_X7Y114_CO6),
.Q(CLBLM_R_X5Y114_SLICE_X7Y114_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_R_X5Y114_SLICE_X7Y114_DLUT (
.I0(CLBLM_R_X7Y115_SLICE_X8Y115_D5Q),
.I1(CLBLL_L_X4Y116_SLICE_X5Y116_B5Q),
.I2(CLBLM_R_X5Y110_SLICE_X6Y110_BQ),
.I3(CLBLL_L_X4Y116_SLICE_X4Y116_A5Q),
.I4(CLBLM_R_X5Y114_SLICE_X7Y114_B5Q),
.I5(CLBLM_R_X5Y116_SLICE_X6Y116_D5Q),
.O5(CLBLM_R_X5Y114_SLICE_X7Y114_DO5),
.O6(CLBLM_R_X5Y114_SLICE_X7Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hd8d8d8d8fafa5050)
  ) CLBLM_R_X5Y114_SLICE_X7Y114_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y114_SLICE_X8Y114_CQ),
.I2(RIOB33_X105Y101_IOB_X1Y102_I),
.I3(1'b1),
.I4(CLBLM_R_X7Y110_SLICE_X8Y110_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y114_SLICE_X7Y114_CO5),
.O6(CLBLM_R_X5Y114_SLICE_X7Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc5c5c0c0fc0cfc0c)
  ) CLBLM_R_X5Y114_SLICE_X7Y114_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X7Y116_SLICE_X9Y116_AQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X5Y113_SLICE_X6Y113_CQ),
.I4(CLBLM_L_X8Y114_SLICE_X10Y114_DQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y114_SLICE_X7Y114_BO5),
.O6(CLBLM_R_X5Y114_SLICE_X7Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hee44fa50ee44fa50)
  ) CLBLM_R_X5Y114_SLICE_X7Y114_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X11Y114_SLICE_X14Y114_CQ),
.I2(CLBLM_R_X5Y114_SLICE_X7Y114_AQ),
.I3(CLBLM_R_X5Y116_SLICE_X7Y116_AQ),
.I4(CLBLL_L_X4Y116_SLICE_X4Y116_BO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y114_SLICE_X7Y114_AO5),
.O6(CLBLM_R_X5Y114_SLICE_X7Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y115_SLICE_X6Y115_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y115_SLICE_X6Y115_AO6),
.Q(CLBLM_R_X5Y115_SLICE_X6Y115_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y115_SLICE_X6Y115_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y115_SLICE_X6Y115_BO6),
.Q(CLBLM_R_X5Y115_SLICE_X6Y115_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y115_SLICE_X6Y115_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y115_SLICE_X6Y115_CO6),
.Q(CLBLM_R_X5Y115_SLICE_X6Y115_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffddffdfdddddddd)
  ) CLBLM_R_X5Y115_SLICE_X6Y115_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X7Y115_SLICE_X9Y115_B5Q),
.I2(CLBLL_L_X4Y107_SLICE_X5Y107_BO6),
.I3(CLBLM_R_X5Y114_SLICE_X6Y114_DO6),
.I4(CLBLM_R_X3Y110_SLICE_X2Y110_BO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y115_SLICE_X6Y115_DO5),
.O6(CLBLM_R_X5Y115_SLICE_X6Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'he4e4e4e4f5a0f5a0)
  ) CLBLM_R_X5Y115_SLICE_X6Y115_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y115_SLICE_X6Y115_CQ),
.I2(CLBLM_R_X13Y117_SLICE_X18Y117_BQ),
.I3(CLBLM_R_X7Y115_SLICE_X8Y115_D5Q),
.I4(1'b1),
.I5(CLBLL_L_X4Y113_SLICE_X5Y113_DO6),
.O5(CLBLM_R_X5Y115_SLICE_X6Y115_CO5),
.O6(CLBLM_R_X5Y115_SLICE_X6Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf6f66666f0f00000)
  ) CLBLM_R_X5Y115_SLICE_X6Y115_BLUT (
.I0(CLBLM_R_X7Y116_SLICE_X9Y116_BO5),
.I1(CLBLM_R_X5Y115_SLICE_X6Y115_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(CLBLL_L_X4Y113_SLICE_X5Y113_AQ),
.I5(CLBLM_R_X7Y115_SLICE_X9Y115_CO6),
.O5(CLBLM_R_X5Y115_SLICE_X6Y115_BO5),
.O6(CLBLM_R_X5Y115_SLICE_X6Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55aa00fa50aa00)
  ) CLBLM_R_X5Y115_SLICE_X6Y115_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(1'b1),
.I2(CLBLM_R_X5Y115_SLICE_X6Y115_AQ),
.I3(CLBLL_L_X4Y115_SLICE_X5Y115_AQ),
.I4(CLBLL_L_X4Y116_SLICE_X4Y116_BO6),
.I5(CLBLM_L_X8Y116_SLICE_X11Y116_BQ),
.O5(CLBLM_R_X5Y115_SLICE_X6Y115_AO5),
.O6(CLBLM_R_X5Y115_SLICE_X6Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y115_SLICE_X7Y115_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y115_SLICE_X7Y115_AO6),
.Q(CLBLM_R_X5Y115_SLICE_X7Y115_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y115_SLICE_X7Y115_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y115_SLICE_X7Y115_BO6),
.Q(CLBLM_R_X5Y115_SLICE_X7Y115_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffdfd)
  ) CLBLM_R_X5Y115_SLICE_X7Y115_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X7Y115_SLICE_X9Y115_B5Q),
.I2(CLBLM_R_X7Y115_SLICE_X8Y115_B5Q),
.I3(1'b1),
.I4(CLBLM_R_X5Y114_SLICE_X7Y114_DO6),
.I5(CLBLM_R_X7Y113_SLICE_X9Y113_A5Q),
.O5(CLBLM_R_X5Y115_SLICE_X7Y115_DO5),
.O6(CLBLM_R_X5Y115_SLICE_X7Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffafb)
  ) CLBLM_R_X5Y115_SLICE_X7Y115_CLUT (
.I0(CLBLM_R_X5Y115_SLICE_X6Y115_DO5),
.I1(CLBLM_R_X3Y110_SLICE_X2Y110_BO6),
.I2(CLBLM_R_X7Y115_SLICE_X8Y115_B5Q),
.I3(CLBLL_L_X4Y107_SLICE_X5Y107_BO6),
.I4(CLBLM_R_X5Y114_SLICE_X7Y114_DO6),
.I5(CLBLM_R_X7Y113_SLICE_X9Y113_A5Q),
.O5(CLBLM_R_X5Y115_SLICE_X7Y115_CO5),
.O6(CLBLM_R_X5Y115_SLICE_X7Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000fe0efe0e)
  ) CLBLM_R_X5Y115_SLICE_X7Y115_BLUT (
.I0(CLBLM_R_X5Y116_SLICE_X6Y116_D5Q),
.I1(CLBLM_R_X5Y115_SLICE_X7Y115_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y117_SLICE_X10Y117_BQ),
.I4(1'b1),
.I5(CLBLL_L_X4Y113_SLICE_X5Y113_DO6),
.O5(CLBLM_R_X5Y115_SLICE_X7Y115_BO5),
.O6(CLBLM_R_X5Y115_SLICE_X7Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdecc5a00fcccf000)
  ) CLBLM_R_X5Y115_SLICE_X7Y115_ALUT (
.I0(CLBLM_R_X5Y116_SLICE_X7Y116_DO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X5Y115_SLICE_X7Y115_AQ),
.I3(CLBLM_R_X7Y115_SLICE_X9Y115_CO6),
.I4(CLBLM_R_X5Y109_SLICE_X7Y109_AQ),
.I5(CLBLM_R_X5Y116_SLICE_X6Y116_CQ),
.O5(CLBLM_R_X5Y115_SLICE_X7Y115_AO5),
.O6(CLBLM_R_X5Y115_SLICE_X7Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y116_SLICE_X6Y116_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y116_SLICE_X6Y116_DO5),
.Q(CLBLM_R_X5Y116_SLICE_X6Y116_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y116_SLICE_X6Y116_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y116_SLICE_X6Y116_BO6),
.Q(CLBLM_R_X5Y116_SLICE_X6Y116_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y116_SLICE_X6Y116_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y116_SLICE_X6Y116_CO6),
.Q(CLBLM_R_X5Y116_SLICE_X6Y116_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y116_SLICE_X6Y116_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y116_SLICE_X6Y116_DO6),
.Q(CLBLM_R_X5Y116_SLICE_X6Y116_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'heeee4444f5a0f5a0)
  ) CLBLM_R_X5Y116_SLICE_X6Y116_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y113_SLICE_X13Y113_AQ),
.I2(CLBLM_R_X5Y116_SLICE_X6Y116_DQ),
.I3(CLBLM_R_X7Y117_SLICE_X9Y117_AQ),
.I4(CLBLM_R_X3Y115_SLICE_X2Y115_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y116_SLICE_X6Y116_DO5),
.O6(CLBLM_R_X5Y116_SLICE_X6Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff282828282828)
  ) CLBLM_R_X5Y116_SLICE_X6Y116_CLUT (
.I0(CLBLM_R_X7Y115_SLICE_X9Y115_CO6),
.I1(CLBLM_R_X5Y116_SLICE_X6Y116_CQ),
.I2(CLBLM_R_X5Y116_SLICE_X7Y116_DO6),
.I3(1'b1),
.I4(CLBLM_R_X5Y116_SLICE_X6Y116_BQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X5Y116_SLICE_X6Y116_CO5),
.O6(CLBLM_R_X5Y116_SLICE_X6Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hacacafafacaca0a0)
  ) CLBLM_R_X5Y116_SLICE_X6Y116_BLUT (
.I0(CLBLM_R_X7Y117_SLICE_X8Y117_AQ),
.I1(CLBLM_R_X5Y116_SLICE_X6Y116_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(CLBLL_L_X4Y116_SLICE_X4Y116_BO6),
.I5(CLBLM_R_X13Y117_SLICE_X18Y117_BQ),
.O5(CLBLM_R_X5Y116_SLICE_X6Y116_BO5),
.O6(CLBLM_R_X5Y116_SLICE_X6Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0c0c0c0000aaaa)
  ) CLBLM_R_X5Y116_SLICE_X6Y116_ALUT (
.I0(RIOB33_X105Y121_IOB_X1Y121_I),
.I1(CLBLL_L_X4Y116_SLICE_X5Y116_A5Q),
.I2(CLBLL_L_X4Y108_SLICE_X4Y108_CO6),
.I3(CLBLM_L_X8Y116_SLICE_X10Y116_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y116_SLICE_X6Y116_AO5),
.O6(CLBLM_R_X5Y116_SLICE_X6Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y116_SLICE_X7Y116_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y116_SLICE_X7Y116_CO6),
.Q(CLBLM_R_X5Y116_SLICE_X7Y116_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y116_SLICE_X7Y116_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y116_SLICE_X7Y116_AO6),
.Q(CLBLM_R_X5Y116_SLICE_X7Y116_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y116_SLICE_X7Y116_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y116_SLICE_X7Y116_BO6),
.Q(CLBLM_R_X5Y116_SLICE_X7Y116_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_R_X5Y116_SLICE_X7Y116_DLUT (
.I0(CLBLM_R_X7Y117_SLICE_X9Y117_AQ),
.I1(CLBLM_R_X7Y117_SLICE_X9Y117_A5Q),
.I2(CLBLM_R_X7Y116_SLICE_X9Y116_AQ),
.I3(CLBLM_R_X7Y117_SLICE_X9Y117_BQ),
.I4(CLBLM_R_X5Y116_SLICE_X7Y116_AQ),
.I5(CLBLM_R_X5Y115_SLICE_X6Y115_BQ),
.O5(CLBLM_R_X5Y116_SLICE_X7Y116_DO5),
.O6(CLBLM_R_X5Y116_SLICE_X7Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hacacacacaa000000)
  ) CLBLM_R_X5Y116_SLICE_X7Y116_CLUT (
.I0(CLBLM_R_X5Y115_SLICE_X7Y115_AQ),
.I1(RIOB33_X105Y127_IOB_X1Y127_I),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X5Y116_SLICE_X6Y116_CQ),
.I4(CLBLM_R_X5Y116_SLICE_X7Y116_DO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y116_SLICE_X7Y116_CO5),
.O6(CLBLM_R_X5Y116_SLICE_X7Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f0fcf03300cc00)
  ) CLBLM_R_X5Y116_SLICE_X7Y116_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y116_SLICE_X7Y116_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y115_SLICE_X9Y115_CO6),
.I4(CLBLM_R_X5Y116_SLICE_X7Y116_CO5),
.I5(CLBLM_R_X5Y106_SLICE_X6Y106_CQ),
.O5(CLBLM_R_X5Y116_SLICE_X7Y116_BO5),
.O6(CLBLM_R_X5Y116_SLICE_X7Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbafa30f0eaaac000)
  ) CLBLM_R_X5Y116_SLICE_X7Y116_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y117_SLICE_X9Y117_A5Q),
.I2(CLBLM_R_X7Y115_SLICE_X9Y115_CO6),
.I3(CLBLM_R_X7Y117_SLICE_X9Y117_AQ),
.I4(CLBLM_R_X5Y111_SLICE_X6Y111_AQ),
.I5(CLBLM_R_X5Y116_SLICE_X7Y116_AQ),
.O5(CLBLM_R_X5Y116_SLICE_X7Y116_AO5),
.O6(CLBLM_R_X5Y116_SLICE_X7Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y117_SLICE_X6Y117_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y117_SLICE_X6Y117_DO5),
.O6(CLBLM_R_X5Y117_SLICE_X6Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y117_SLICE_X6Y117_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y117_SLICE_X6Y117_CO5),
.O6(CLBLM_R_X5Y117_SLICE_X6Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y117_SLICE_X6Y117_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y117_SLICE_X6Y117_BO5),
.O6(CLBLM_R_X5Y117_SLICE_X6Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y117_SLICE_X6Y117_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y117_SLICE_X6Y117_AO5),
.O6(CLBLM_R_X5Y117_SLICE_X6Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y117_SLICE_X7Y117_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y117_SLICE_X7Y117_AO6),
.Q(CLBLM_R_X5Y117_SLICE_X7Y117_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y117_SLICE_X7Y117_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y117_SLICE_X7Y117_DO5),
.O6(CLBLM_R_X5Y117_SLICE_X7Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y117_SLICE_X7Y117_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y117_SLICE_X7Y117_CO5),
.O6(CLBLM_R_X5Y117_SLICE_X7Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y117_SLICE_X7Y117_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y117_SLICE_X7Y117_BO5),
.O6(CLBLM_R_X5Y117_SLICE_X7Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000ffee5544)
  ) CLBLM_R_X5Y117_SLICE_X7Y117_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(1'b1),
.I3(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.I4(CLBLL_L_X4Y117_SLICE_X4Y117_BQ),
.I5(CLBLM_L_X8Y114_SLICE_X11Y114_DO6),
.O5(CLBLM_R_X5Y117_SLICE_X7Y117_AO5),
.O6(CLBLM_R_X5Y117_SLICE_X7Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y105_SLICE_X8Y105_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y105_SLICE_X8Y105_BO6),
.Q(CLBLM_R_X7Y105_SLICE_X8Y105_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y105_SLICE_X8Y105_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y105_SLICE_X8Y105_AO6),
.Q(CLBLM_R_X7Y105_SLICE_X8Y105_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y105_SLICE_X8Y105_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y105_SLICE_X8Y105_CO6),
.Q(CLBLM_R_X7Y105_SLICE_X8Y105_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00cf00cf00ef00ef)
  ) CLBLM_R_X7Y105_SLICE_X8Y105_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X7Y116_SLICE_X8Y116_CQ),
.I2(CLBLM_L_X10Y104_SLICE_X12Y104_AQ),
.I3(CLBLM_R_X7Y105_SLICE_X8Y105_A5Q),
.I4(1'b1),
.I5(CLBLM_R_X3Y110_SLICE_X2Y110_DO6),
.O5(CLBLM_R_X7Y105_SLICE_X8Y105_DO5),
.O6(CLBLM_R_X7Y105_SLICE_X8Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'heeeeaaee44440044)
  ) CLBLM_R_X7Y105_SLICE_X8Y105_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y105_SLICE_X8Y105_CQ),
.I2(1'b1),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.I5(CLBLM_R_X7Y105_SLICE_X9Y105_BQ),
.O5(CLBLM_R_X7Y105_SLICE_X8Y105_CO5),
.O6(CLBLM_R_X7Y105_SLICE_X8Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff100010c0c0c0c0)
  ) CLBLM_R_X7Y105_SLICE_X8Y105_BLUT (
.I0(CLBLM_R_X7Y105_SLICE_X8Y105_DO6),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y104_SLICE_X11Y104_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y105_SLICE_X8Y105_BO5),
.O6(CLBLM_R_X7Y105_SLICE_X8Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffafa0000fafa)
  ) CLBLM_R_X7Y105_SLICE_X8Y105_ALUT (
.I0(CLBLM_R_X7Y115_SLICE_X8Y115_DQ),
.I1(1'b1),
.I2(CLBLM_R_X7Y105_SLICE_X8Y105_AQ),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(LIOB33_X0Y79_IOB_X0Y79_I),
.O5(CLBLM_R_X7Y105_SLICE_X8Y105_AO5),
.O6(CLBLM_R_X7Y105_SLICE_X8Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y105_SLICE_X9Y105_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y105_SLICE_X9Y105_AO6),
.Q(CLBLM_R_X7Y105_SLICE_X9Y105_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y105_SLICE_X9Y105_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y105_SLICE_X9Y105_BO6),
.Q(CLBLM_R_X7Y105_SLICE_X9Y105_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y105_SLICE_X9Y105_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y105_SLICE_X9Y105_CO6),
.Q(CLBLM_R_X7Y105_SLICE_X9Y105_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000323200003333)
  ) CLBLM_R_X7Y105_SLICE_X9Y105_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X7Y116_SLICE_X8Y116_CQ),
.I2(CLBLM_L_X10Y104_SLICE_X12Y104_AQ),
.I3(1'b1),
.I4(CLBLM_R_X7Y105_SLICE_X9Y105_AQ),
.I5(CLBLM_R_X3Y110_SLICE_X3Y110_AO6),
.O5(CLBLM_R_X7Y105_SLICE_X9Y105_DO5),
.O6(CLBLM_R_X7Y105_SLICE_X9Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaabebe00001414)
  ) CLBLM_R_X7Y105_SLICE_X9Y105_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y105_SLICE_X9Y105_CQ),
.I2(CLBLM_R_X7Y107_SLICE_X8Y107_DO6),
.I3(1'b1),
.I4(CLBLM_L_X10Y113_SLICE_X13Y113_AQ),
.I5(CLBLM_L_X8Y105_SLICE_X11Y105_AQ),
.O5(CLBLM_R_X7Y105_SLICE_X9Y105_CO5),
.O6(CLBLM_R_X7Y105_SLICE_X9Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hacaca0a0afa0afa0)
  ) CLBLM_R_X7Y105_SLICE_X9Y105_BLUT (
.I0(CLBLM_R_X5Y107_SLICE_X6Y107_AQ),
.I1(CLBLM_R_X7Y105_SLICE_X9Y105_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y105_SLICE_X11Y105_AQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_L_X10Y106_SLICE_X12Y106_BO6),
.O5(CLBLM_R_X7Y105_SLICE_X9Y105_BO5),
.O6(CLBLM_R_X7Y105_SLICE_X9Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcd01cc000000f0f0)
  ) CLBLM_R_X7Y105_SLICE_X9Y105_ALUT (
.I0(CLBLM_R_X7Y105_SLICE_X9Y105_DO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(RIOB33_X105Y117_IOB_X1Y118_I),
.I3(CLBLM_R_X5Y113_SLICE_X6Y113_BQ),
.I4(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y105_SLICE_X9Y105_AO5),
.O6(CLBLM_R_X7Y105_SLICE_X9Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y106_SLICE_X8Y106_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y106_SLICE_X8Y106_AO6),
.Q(CLBLM_R_X7Y106_SLICE_X8Y106_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y106_SLICE_X8Y106_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y106_SLICE_X8Y106_BO6),
.Q(CLBLM_R_X7Y106_SLICE_X8Y106_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y106_SLICE_X8Y106_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y106_SLICE_X8Y106_CO6),
.Q(CLBLM_R_X7Y106_SLICE_X8Y106_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y106_SLICE_X8Y106_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y106_SLICE_X8Y106_DO5),
.O6(CLBLM_R_X7Y106_SLICE_X8Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafaeaea50504040)
  ) CLBLM_R_X7Y106_SLICE_X8Y106_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y106_SLICE_X8Y106_CQ),
.I2(CLBLM_L_X8Y104_SLICE_X10Y104_AO6),
.I3(1'b1),
.I4(CLBLM_R_X7Y109_SLICE_X9Y109_CQ),
.I5(CLBLM_R_X7Y109_SLICE_X8Y109_AQ),
.O5(CLBLM_R_X7Y106_SLICE_X8Y106_CO5),
.O6(CLBLM_R_X7Y106_SLICE_X8Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hafacafaca0a0a0a0)
  ) CLBLM_R_X7Y106_SLICE_X8Y106_BLUT (
.I0(CLBLM_L_X8Y109_SLICE_X10Y109_CQ),
.I1(CLBLM_R_X7Y106_SLICE_X8Y106_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X5Y105_SLICE_X7Y105_BQ),
.I4(1'b1),
.I5(CLBLM_L_X8Y104_SLICE_X10Y104_AO6),
.O5(CLBLM_R_X7Y106_SLICE_X8Y106_BO5),
.O6(CLBLM_R_X7Y106_SLICE_X8Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa33aaffaa30aaf0)
  ) CLBLM_R_X7Y106_SLICE_X8Y106_ALUT (
.I0(CLBLM_L_X12Y107_SLICE_X16Y107_DQ),
.I1(CLBLM_R_X7Y105_SLICE_X8Y105_CQ),
.I2(CLBLM_R_X7Y106_SLICE_X8Y106_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLL_L_X4Y110_SLICE_X4Y110_AQ),
.I5(CLBLM_R_X5Y106_SLICE_X6Y106_CQ),
.O5(CLBLM_R_X7Y106_SLICE_X8Y106_AO5),
.O6(CLBLM_R_X7Y106_SLICE_X8Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y106_SLICE_X9Y106_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y106_SLICE_X9Y106_AO6),
.Q(CLBLM_R_X7Y106_SLICE_X9Y106_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y106_SLICE_X9Y106_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y106_SLICE_X9Y106_BO6),
.Q(CLBLM_R_X7Y106_SLICE_X9Y106_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y106_SLICE_X9Y106_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y106_SLICE_X9Y106_CO6),
.Q(CLBLM_R_X7Y106_SLICE_X9Y106_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h11110000aa00fa50)
  ) CLBLM_R_X7Y106_SLICE_X9Y106_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y111_SLICE_X12Y111_CQ),
.I2(CLBLM_R_X7Y111_SLICE_X8Y111_BQ),
.I3(CLBLL_L_X4Y107_SLICE_X4Y107_CQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y106_SLICE_X9Y106_DO5),
.O6(CLBLM_R_X7Y106_SLICE_X9Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffeeaaaa55440000)
  ) CLBLM_R_X7Y106_SLICE_X9Y106_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y106_SLICE_X9Y106_CQ),
.I2(1'b1),
.I3(CLBLM_R_X7Y105_SLICE_X9Y105_CQ),
.I4(CLBLM_L_X8Y104_SLICE_X10Y104_AO6),
.I5(CLBLM_R_X7Y112_SLICE_X8Y112_BQ),
.O5(CLBLM_R_X7Y106_SLICE_X9Y106_CO5),
.O6(CLBLM_R_X7Y106_SLICE_X9Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000ff00e0e0)
  ) CLBLM_R_X7Y106_SLICE_X9Y106_BLUT (
.I0(CLBLM_R_X11Y107_SLICE_X15Y107_BQ),
.I1(CLBLM_R_X7Y106_SLICE_X9Y106_BQ),
.I2(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.I3(CLBLL_L_X4Y113_SLICE_X4Y113_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_R_X7Y106_SLICE_X9Y106_BO5),
.O6(CLBLM_R_X7Y106_SLICE_X9Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc05505050)
  ) CLBLM_R_X7Y106_SLICE_X9Y106_ALUT (
.I0(CLBLM_L_X10Y113_SLICE_X13Y113_AQ),
.I1(CLBLM_L_X12Y109_SLICE_X16Y109_D5Q),
.I2(CLBLM_R_X7Y106_SLICE_X9Y106_AQ),
.I3(CLBLM_R_X7Y105_SLICE_X9Y105_AO5),
.I4(CLBLM_R_X7Y109_SLICE_X9Y109_CQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X7Y106_SLICE_X9Y106_AO5),
.O6(CLBLM_R_X7Y106_SLICE_X9Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y107_SLICE_X8Y107_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y107_SLICE_X8Y107_AO6),
.Q(CLBLM_R_X7Y107_SLICE_X8Y107_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y107_SLICE_X8Y107_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y107_SLICE_X8Y107_BO6),
.Q(CLBLM_R_X7Y107_SLICE_X8Y107_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y107_SLICE_X8Y107_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y107_SLICE_X8Y107_CO6),
.Q(CLBLM_R_X7Y107_SLICE_X8Y107_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000800000000000)
  ) CLBLM_R_X7Y107_SLICE_X8Y107_DLUT (
.I0(CLBLM_R_X7Y106_SLICE_X9Y106_AQ),
.I1(CLBLM_R_X7Y108_SLICE_X9Y108_AQ),
.I2(CLBLM_L_X8Y110_SLICE_X10Y110_BQ),
.I3(CLBLM_R_X7Y109_SLICE_X9Y109_CQ),
.I4(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_R_X7Y107_SLICE_X8Y107_DO5),
.O6(CLBLM_R_X7Y107_SLICE_X8Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00aafcaa00)
  ) CLBLM_R_X7Y107_SLICE_X8Y107_CLUT (
.I0(CLBLM_R_X7Y113_SLICE_X9Y113_AQ),
.I1(CLBLM_R_X7Y107_SLICE_X8Y107_CQ),
.I2(CLBLM_L_X8Y107_SLICE_X10Y107_CQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_R_X7Y107_SLICE_X8Y107_CO5),
.O6(CLBLM_R_X7Y107_SLICE_X8Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff00f00fef40e04)
  ) CLBLM_R_X7Y107_SLICE_X8Y107_BLUT (
.I0(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.I1(CLBLM_R_X7Y107_SLICE_X8Y107_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y107_SLICE_X9Y107_BQ),
.I4(CLBLM_R_X5Y110_SLICE_X7Y110_AQ),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_R_X7Y107_SLICE_X8Y107_BO5),
.O6(CLBLM_R_X7Y107_SLICE_X8Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00e4e4cccc)
  ) CLBLM_R_X7Y107_SLICE_X8Y107_ALUT (
.I0(CLBLM_R_X7Y105_SLICE_X8Y105_CQ),
.I1(CLBLM_L_X8Y110_SLICE_X10Y110_BQ),
.I2(CLBLM_R_X7Y107_SLICE_X8Y107_AQ),
.I3(CLBLM_L_X12Y106_SLICE_X17Y106_AQ),
.I4(CLBLL_L_X4Y110_SLICE_X4Y110_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X7Y107_SLICE_X8Y107_AO5),
.O6(CLBLM_R_X7Y107_SLICE_X8Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y107_SLICE_X9Y107_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y107_SLICE_X9Y107_CO5),
.Q(CLBLM_R_X7Y107_SLICE_X9Y107_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y107_SLICE_X9Y107_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y107_SLICE_X9Y107_AO6),
.Q(CLBLM_R_X7Y107_SLICE_X9Y107_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y107_SLICE_X9Y107_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y107_SLICE_X9Y107_BO6),
.Q(CLBLM_R_X7Y107_SLICE_X9Y107_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y107_SLICE_X9Y107_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y107_SLICE_X9Y107_CO6),
.Q(CLBLM_R_X7Y107_SLICE_X9Y107_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h2424424242422424)
  ) CLBLM_R_X7Y107_SLICE_X9Y107_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X7Y107_SLICE_X9Y107_CQ),
.I2(CLBLM_R_X7Y108_SLICE_X8Y108_CQ),
.I3(1'b1),
.I4(CLBLM_L_X10Y108_SLICE_X12Y108_CQ),
.I5(CLBLM_R_X5Y105_SLICE_X6Y105_BQ),
.O5(CLBLM_R_X7Y107_SLICE_X9Y107_DO5),
.O6(CLBLM_R_X7Y107_SLICE_X9Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hdddd8888fa50fa50)
  ) CLBLM_R_X7Y107_SLICE_X9Y107_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y110_SLICE_X9Y110_AQ),
.I2(CLBLM_L_X8Y108_SLICE_X10Y108_AQ),
.I3(CLBLM_R_X7Y107_SLICE_X9Y107_AQ),
.I4(CLBLM_R_X7Y107_SLICE_X9Y107_DO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y107_SLICE_X9Y107_CO5),
.O6(CLBLM_R_X7Y107_SLICE_X9Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff00a8000000a8)
  ) CLBLM_R_X7Y107_SLICE_X9Y107_BLUT (
.I0(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.I1(CLBLM_R_X7Y107_SLICE_X9Y107_BQ),
.I2(CLBLM_R_X7Y107_SLICE_X9Y107_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X5Y116_SLICE_X6Y116_D5Q),
.O5(CLBLM_R_X7Y107_SLICE_X9Y107_BO5),
.O6(CLBLM_R_X7Y107_SLICE_X9Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f05555f0f01111)
  ) CLBLM_R_X7Y107_SLICE_X9Y107_ALUT (
.I0(CLBLM_R_X7Y108_SLICE_X9Y108_DO6),
.I1(RIOB33_X105Y141_IOB_X1Y142_I),
.I2(CLBLM_R_X7Y107_SLICE_X9Y107_CQ),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y119_SLICE_X10Y119_AQ),
.O5(CLBLM_R_X7Y107_SLICE_X9Y107_AO5),
.O6(CLBLM_R_X7Y107_SLICE_X9Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y108_SLICE_X8Y108_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y108_SLICE_X8Y108_AO6),
.Q(CLBLM_R_X7Y108_SLICE_X8Y108_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y108_SLICE_X8Y108_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y108_SLICE_X8Y108_BO6),
.Q(CLBLM_R_X7Y108_SLICE_X8Y108_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y108_SLICE_X8Y108_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y108_SLICE_X8Y108_CO6),
.Q(CLBLM_R_X7Y108_SLICE_X8Y108_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h1111fffff000ffff)
  ) CLBLM_R_X7Y108_SLICE_X8Y108_DLUT (
.I0(CLBLM_L_X8Y109_SLICE_X11Y109_AQ),
.I1(CLBLM_R_X11Y111_SLICE_X15Y111_BQ),
.I2(CLBLM_R_X5Y111_SLICE_X7Y111_CQ),
.I3(CLBLM_R_X7Y115_SLICE_X8Y115_CQ),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y108_SLICE_X8Y108_DO5),
.O6(CLBLM_R_X7Y108_SLICE_X8Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h88d8888d88d8888d)
  ) CLBLM_R_X7Y108_SLICE_X8Y108_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y112_SLICE_X10Y112_A5Q),
.I2(CLBLM_L_X10Y108_SLICE_X12Y108_CQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X7Y108_SLICE_X8Y108_DO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y108_SLICE_X8Y108_CO5),
.O6(CLBLM_R_X7Y108_SLICE_X8Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccf5f5a0a0)
  ) CLBLM_R_X7Y108_SLICE_X8Y108_BLUT (
.I0(CLBLL_L_X4Y112_SLICE_X4Y112_CO5),
.I1(CLBLM_R_X7Y107_SLICE_X8Y107_AQ),
.I2(CLBLM_R_X7Y109_SLICE_X9Y109_DQ),
.I3(1'b1),
.I4(CLBLM_R_X7Y108_SLICE_X8Y108_BQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X7Y108_SLICE_X8Y108_BO5),
.O6(CLBLM_R_X7Y108_SLICE_X8Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa00fcfcfc)
  ) CLBLM_R_X7Y108_SLICE_X8Y108_ALUT (
.I0(CLBLM_L_X8Y113_SLICE_X10Y113_D5Q),
.I1(CLBLM_R_X5Y106_SLICE_X6Y106_BQ),
.I2(CLBLM_R_X7Y108_SLICE_X8Y108_AQ),
.I3(CLBLM_R_X7Y105_SLICE_X8Y105_CQ),
.I4(CLBLL_L_X4Y110_SLICE_X4Y110_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X7Y108_SLICE_X8Y108_AO5),
.O6(CLBLM_R_X7Y108_SLICE_X8Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y108_SLICE_X9Y108_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y108_SLICE_X9Y108_AO6),
.Q(CLBLM_R_X7Y108_SLICE_X9Y108_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000000fcc0f33)
  ) CLBLM_R_X7Y108_SLICE_X9Y108_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y109_SLICE_X11Y109_CQ),
.I2(CLBLM_R_X7Y107_SLICE_X9Y107_C5Q),
.I3(CLBLM_R_X5Y115_SLICE_X7Y115_CO6),
.I4(CLBLM_L_X10Y109_SLICE_X13Y109_BO5),
.I5(CLBLM_R_X7Y107_SLICE_X9Y107_AQ),
.O5(CLBLM_R_X7Y108_SLICE_X9Y108_DO5),
.O6(CLBLM_R_X7Y108_SLICE_X9Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbfffbffffffffff)
  ) CLBLM_R_X7Y108_SLICE_X9Y108_CLUT (
.I0(CLBLL_L_X4Y107_SLICE_X5Y107_BO6),
.I1(CLBLL_L_X4Y108_SLICE_X5Y108_AO6),
.I2(CLBLM_L_X10Y112_SLICE_X12Y112_DO6),
.I3(CLBLL_L_X2Y110_SLICE_X1Y110_DO6),
.I4(1'b1),
.I5(CLBLM_R_X3Y110_SLICE_X2Y110_DO6),
.O5(CLBLM_R_X7Y108_SLICE_X9Y108_CO5),
.O6(CLBLM_R_X7Y108_SLICE_X9Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h300000000f0fffff)
  ) CLBLM_R_X7Y108_SLICE_X9Y108_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.I2(CLBLM_R_X7Y106_SLICE_X9Y106_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_R_X7Y109_SLICE_X9Y109_CQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y108_SLICE_X9Y108_BO5),
.O6(CLBLM_R_X7Y108_SLICE_X9Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000aaaa3cf0)
  ) CLBLM_R_X7Y108_SLICE_X9Y108_ALUT (
.I0(CLBLM_R_X7Y115_SLICE_X8Y115_CQ),
.I1(CLBLM_L_X8Y110_SLICE_X10Y110_BQ),
.I2(CLBLM_R_X7Y108_SLICE_X9Y108_AQ),
.I3(CLBLM_R_X7Y108_SLICE_X9Y108_BO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X10Y113_SLICE_X13Y113_AQ),
.O5(CLBLM_R_X7Y108_SLICE_X9Y108_AO5),
.O6(CLBLM_R_X7Y108_SLICE_X9Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y109_SLICE_X8Y109_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y109_SLICE_X8Y109_AO6),
.Q(CLBLM_R_X7Y109_SLICE_X8Y109_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y109_SLICE_X8Y109_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y109_SLICE_X8Y109_BO6),
.Q(CLBLM_R_X7Y109_SLICE_X8Y109_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffae0400005555)
  ) CLBLM_R_X7Y109_SLICE_X8Y109_DLUT (
.I0(CLBLM_L_X10Y104_SLICE_X12Y104_AQ),
.I1(CLBLL_L_X2Y111_SLICE_X1Y111_DO6),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X7Y109_SLICE_X8Y109_CO6),
.I4(CLBLM_R_X7Y116_SLICE_X8Y116_CQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y109_SLICE_X8Y109_DO5),
.O6(CLBLM_R_X7Y109_SLICE_X8Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff00000eeee0000)
  ) CLBLM_R_X7Y109_SLICE_X8Y109_CLUT (
.I0(CLBLM_R_X7Y113_SLICE_X9Y113_AQ),
.I1(CLBLM_R_X5Y109_SLICE_X6Y109_DQ),
.I2(CLBLL_L_X4Y109_SLICE_X5Y109_AQ),
.I3(CLBLM_L_X8Y112_SLICE_X10Y112_A5Q),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y109_SLICE_X8Y109_CO5),
.O6(CLBLM_R_X7Y109_SLICE_X8Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffa8a8a8a8a8a8)
  ) CLBLM_R_X7Y109_SLICE_X8Y109_BLUT (
.I0(CLBLL_L_X4Y112_SLICE_X4Y112_CO6),
.I1(CLBLM_R_X7Y109_SLICE_X8Y109_BQ),
.I2(CLBLM_R_X5Y108_SLICE_X7Y108_AQ),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y111_SLICE_X9Y111_BQ),
.O5(CLBLM_R_X7Y109_SLICE_X8Y109_BO5),
.O6(CLBLM_R_X7Y109_SLICE_X8Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcff3033fccc3000)
  ) CLBLM_R_X7Y109_SLICE_X8Y109_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X7Y109_SLICE_X8Y109_AQ),
.I3(CLBLL_L_X4Y116_SLICE_X4Y116_BO6),
.I4(CLBLM_R_X5Y109_SLICE_X6Y109_DQ),
.I5(CLBLM_L_X8Y114_SLICE_X11Y114_CQ),
.O5(CLBLM_R_X7Y109_SLICE_X8Y109_AO5),
.O6(CLBLM_R_X7Y109_SLICE_X8Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y109_SLICE_X9Y109_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y109_SLICE_X9Y109_AO6),
.Q(CLBLM_R_X7Y109_SLICE_X9Y109_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y109_SLICE_X9Y109_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y109_SLICE_X9Y109_BO6),
.Q(CLBLM_R_X7Y109_SLICE_X9Y109_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y109_SLICE_X9Y109_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y109_SLICE_X9Y109_CO6),
.Q(CLBLM_R_X7Y109_SLICE_X9Y109_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y109_SLICE_X9Y109_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y109_SLICE_X9Y109_DO6),
.Q(CLBLM_R_X7Y109_SLICE_X9Y109_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf044f044f011f011)
  ) CLBLM_R_X7Y109_SLICE_X9Y109_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X8Y109_SLICE_X11Y109_DO6),
.I2(CLBLM_L_X12Y112_SLICE_X16Y112_B5Q),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLM_R_X5Y106_SLICE_X6Y106_DQ),
.O5(CLBLM_R_X7Y109_SLICE_X9Y109_DO5),
.O6(CLBLM_R_X7Y109_SLICE_X9Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55ff55eb41ee44)
  ) CLBLM_R_X7Y109_SLICE_X9Y109_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y109_SLICE_X9Y109_CQ),
.I2(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.I3(CLBLM_L_X8Y114_SLICE_X11Y114_CQ),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLM_L_X10Y113_SLICE_X13Y113_AQ),
.O5(CLBLM_R_X7Y109_SLICE_X9Y109_CO5),
.O6(CLBLM_R_X7Y109_SLICE_X9Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfe0ef404fe0ef404)
  ) CLBLM_R_X7Y109_SLICE_X9Y109_BLUT (
.I0(CLBLL_L_X4Y112_SLICE_X4Y112_CO5),
.I1(CLBLM_R_X7Y109_SLICE_X9Y109_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y108_SLICE_X12Y108_CQ),
.I4(CLBLM_L_X12Y108_SLICE_X16Y108_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y109_SLICE_X9Y109_BO5),
.O6(CLBLM_R_X7Y109_SLICE_X9Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefefcfcaaaa0000)
  ) CLBLM_R_X7Y109_SLICE_X9Y109_ALUT (
.I0(CLBLM_R_X7Y110_SLICE_X9Y110_BQ),
.I1(CLBLM_R_X7Y111_SLICE_X8Y111_BQ),
.I2(CLBLM_R_X7Y109_SLICE_X9Y109_AQ),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLL_L_X4Y112_SLICE_X4Y112_CO6),
.O5(CLBLM_R_X7Y109_SLICE_X9Y109_AO5),
.O6(CLBLM_R_X7Y109_SLICE_X9Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y110_SLICE_X8Y110_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y110_SLICE_X8Y110_AO6),
.Q(CLBLM_R_X7Y110_SLICE_X8Y110_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y110_SLICE_X8Y110_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y110_SLICE_X8Y110_BO6),
.Q(CLBLM_R_X7Y110_SLICE_X8Y110_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y110_SLICE_X8Y110_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y110_SLICE_X8Y110_CO6),
.Q(CLBLM_R_X7Y110_SLICE_X8Y110_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hb1b1b1b10000ccff)
  ) CLBLM_R_X7Y110_SLICE_X8Y110_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLL_L_X2Y110_SLICE_X1Y110_DO6),
.I2(CLBLM_L_X8Y106_SLICE_X11Y106_AQ),
.I3(CLBLM_R_X5Y106_SLICE_X6Y106_CQ),
.I4(CLBLM_L_X10Y113_SLICE_X13Y113_CQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y110_SLICE_X8Y110_DO5),
.O6(CLBLM_R_X7Y110_SLICE_X8Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa0faa0faa0caa0c)
  ) CLBLM_R_X7Y110_SLICE_X8Y110_CLUT (
.I0(CLBLM_R_X7Y112_SLICE_X8Y112_AQ),
.I1(CLBLM_R_X7Y110_SLICE_X8Y110_CQ),
.I2(CLBLM_R_X5Y115_SLICE_X7Y115_CO6),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLM_L_X8Y109_SLICE_X11Y109_CQ),
.O5(CLBLM_R_X7Y110_SLICE_X8Y110_CO5),
.O6(CLBLM_R_X7Y110_SLICE_X8Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0cacac0c0caca)
  ) CLBLM_R_X7Y110_SLICE_X8Y110_BLUT (
.I0(CLBLM_R_X5Y114_SLICE_X7Y114_BQ),
.I1(CLBLM_R_X7Y105_SLICE_X8Y105_A5Q),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y110_SLICE_X8Y110_BO5),
.O6(CLBLM_R_X7Y110_SLICE_X8Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaf0cccccc)
  ) CLBLM_R_X7Y110_SLICE_X8Y110_ALUT (
.I0(CLBLM_R_X11Y110_SLICE_X14Y110_A5Q),
.I1(CLBLM_R_X7Y105_SLICE_X9Y105_CQ),
.I2(CLBLM_R_X7Y110_SLICE_X8Y110_AQ),
.I3(CLBLM_R_X7Y105_SLICE_X8Y105_CQ),
.I4(CLBLL_L_X4Y110_SLICE_X4Y110_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X7Y110_SLICE_X8Y110_AO5),
.O6(CLBLM_R_X7Y110_SLICE_X8Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y110_SLICE_X9Y110_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y110_SLICE_X9Y110_AO6),
.Q(CLBLM_R_X7Y110_SLICE_X9Y110_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y110_SLICE_X9Y110_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y110_SLICE_X9Y110_BO6),
.Q(CLBLM_R_X7Y110_SLICE_X9Y110_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haa88a080aacca0c0)
  ) CLBLM_R_X7Y110_SLICE_X9Y110_DLUT (
.I0(CLBLM_R_X7Y109_SLICE_X8Y109_CO5),
.I1(CLBLM_L_X10Y104_SLICE_X12Y104_AQ),
.I2(RIOB33_X105Y117_IOB_X1Y118_I),
.I3(CLBLM_R_X7Y116_SLICE_X8Y116_CQ),
.I4(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.I5(CLBLL_L_X4Y108_SLICE_X5Y108_AO6),
.O5(CLBLM_R_X7Y110_SLICE_X9Y110_DO5),
.O6(CLBLM_R_X7Y110_SLICE_X9Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0300010033003300)
  ) CLBLM_R_X7Y110_SLICE_X9Y110_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X7Y116_SLICE_X8Y116_CQ),
.I3(CLBLM_L_X8Y110_SLICE_X10Y110_DO6),
.I4(CLBLM_R_X3Y110_SLICE_X3Y110_DO6),
.I5(CLBLM_R_X7Y111_SLICE_X9Y111_DO5),
.O5(CLBLM_R_X7Y110_SLICE_X9Y110_CO5),
.O6(CLBLM_R_X7Y110_SLICE_X9Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffff0ccf088)
  ) CLBLM_R_X7Y110_SLICE_X9Y110_BLUT (
.I0(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.I1(CLBLM_R_X7Y110_SLICE_X9Y110_BQ),
.I2(CLBLM_R_X7Y113_SLICE_X8Y113_C5Q),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLM_R_X7Y110_SLICE_X9Y110_CO6),
.O5(CLBLM_R_X7Y110_SLICE_X9Y110_BO5),
.O6(CLBLM_R_X7Y110_SLICE_X9Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fa000af0f50005)
  ) CLBLM_R_X7Y110_SLICE_X9Y110_ALUT (
.I0(CLBLM_L_X8Y113_SLICE_X10Y113_CQ),
.I1(1'b1),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X11Y110_SLICE_X14Y110_AQ),
.I5(CLBLM_L_X8Y112_SLICE_X10Y112_BO6),
.O5(CLBLM_R_X7Y110_SLICE_X9Y110_AO5),
.O6(CLBLM_R_X7Y110_SLICE_X9Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y111_SLICE_X8Y111_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y111_SLICE_X8Y111_AO6),
.Q(CLBLM_R_X7Y111_SLICE_X8Y111_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y111_SLICE_X8Y111_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y111_SLICE_X8Y111_BO6),
.Q(CLBLM_R_X7Y111_SLICE_X8Y111_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y111_SLICE_X8Y111_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y111_SLICE_X8Y111_CO6),
.Q(CLBLM_R_X7Y111_SLICE_X8Y111_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y111_SLICE_X8Y111_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y111_SLICE_X8Y111_DO6),
.Q(CLBLM_R_X7Y111_SLICE_X8Y111_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haabbaaee00110044)
  ) CLBLM_R_X7Y111_SLICE_X8Y111_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y111_SLICE_X6Y111_CQ),
.I2(1'b1),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X7Y109_SLICE_X8Y109_CO5),
.I5(CLBLM_L_X10Y113_SLICE_X13Y113_CQ),
.O5(CLBLM_R_X7Y111_SLICE_X8Y111_DO5),
.O6(CLBLM_R_X7Y111_SLICE_X8Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0e4a0a0a0e4a0)
  ) CLBLM_R_X7Y111_SLICE_X8Y111_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y111_SLICE_X8Y111_CQ),
.I2(CLBLM_R_X7Y111_SLICE_X8Y111_DQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X7Y112_SLICE_X8Y112_CQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y111_SLICE_X8Y111_CO5),
.O6(CLBLM_R_X7Y111_SLICE_X8Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0c0cfcfc0)
  ) CLBLM_R_X7Y111_SLICE_X8Y111_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y107_SLICE_X8Y107_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y114_SLICE_X8Y114_CQ),
.I4(CLBLM_L_X8Y111_SLICE_X10Y111_DO6),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X7Y111_SLICE_X8Y111_BO5),
.O6(CLBLM_R_X7Y111_SLICE_X8Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcffecee30332022)
  ) CLBLM_R_X7Y111_SLICE_X8Y111_ALUT (
.I0(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X7Y111_SLICE_X8Y111_AQ),
.I3(CLBLM_L_X8Y112_SLICE_X10Y112_BO6),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLL_L_X4Y116_SLICE_X4Y116_A5Q),
.O5(CLBLM_R_X7Y111_SLICE_X8Y111_AO5),
.O6(CLBLM_R_X7Y111_SLICE_X8Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y111_SLICE_X9Y111_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y111_SLICE_X9Y111_AO6),
.Q(CLBLM_R_X7Y111_SLICE_X9Y111_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y111_SLICE_X9Y111_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y111_SLICE_X9Y111_BO6),
.Q(CLBLM_R_X7Y111_SLICE_X9Y111_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y111_SLICE_X9Y111_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y111_SLICE_X9Y111_CO6),
.Q(CLBLM_R_X7Y111_SLICE_X9Y111_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff33cc0037373737)
  ) CLBLM_R_X7Y111_SLICE_X9Y111_DLUT (
.I0(CLBLM_R_X7Y111_SLICE_X8Y111_AQ),
.I1(RIOB33_X105Y121_IOB_X1Y121_I),
.I2(CLBLM_R_X5Y114_SLICE_X7Y114_BQ),
.I3(CLBLM_R_X11Y112_SLICE_X14Y112_CQ),
.I4(CLBLM_L_X8Y113_SLICE_X11Y113_BQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y111_SLICE_X9Y111_DO5),
.O6(CLBLM_R_X7Y111_SLICE_X9Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haabb0011bbaa1100)
  ) CLBLM_R_X7Y111_SLICE_X9Y111_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(1'b1),
.I3(CLBLM_L_X8Y112_SLICE_X10Y112_CO6),
.I4(CLBLM_R_X5Y105_SLICE_X6Y105_AQ),
.I5(CLBLM_R_X7Y110_SLICE_X9Y110_AQ),
.O5(CLBLM_R_X7Y111_SLICE_X9Y111_CO5),
.O6(CLBLM_R_X7Y111_SLICE_X9Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffeca0a0ffeca0a0)
  ) CLBLM_R_X7Y111_SLICE_X9Y111_BLUT (
.I0(CLBLM_L_X12Y111_SLICE_X16Y111_CQ),
.I1(CLBLM_R_X7Y111_SLICE_X9Y111_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y110_SLICE_X9Y110_AQ),
.I4(CLBLL_L_X4Y112_SLICE_X4Y112_CO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y111_SLICE_X9Y111_BO5),
.O6(CLBLM_R_X7Y111_SLICE_X9Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffcec0000fcec)
  ) CLBLM_R_X7Y111_SLICE_X9Y111_ALUT (
.I0(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.I1(CLBLM_R_X7Y110_SLICE_X9Y110_DO6),
.I2(CLBLM_R_X7Y111_SLICE_X9Y111_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLL_L_X4Y113_SLICE_X5Y113_BQ),
.O5(CLBLM_R_X7Y111_SLICE_X9Y111_AO5),
.O6(CLBLM_R_X7Y111_SLICE_X9Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y112_SLICE_X8Y112_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y112_SLICE_X8Y112_CO5),
.Q(CLBLM_R_X7Y112_SLICE_X8Y112_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y112_SLICE_X8Y112_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y112_SLICE_X8Y112_AO6),
.Q(CLBLM_R_X7Y112_SLICE_X8Y112_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y112_SLICE_X8Y112_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y112_SLICE_X8Y112_BO6),
.Q(CLBLM_R_X7Y112_SLICE_X8Y112_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y112_SLICE_X8Y112_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y112_SLICE_X8Y112_CO6),
.Q(CLBLM_R_X7Y112_SLICE_X8Y112_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y112_SLICE_X8Y112_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y112_SLICE_X8Y112_DO6),
.Q(CLBLM_R_X7Y112_SLICE_X8Y112_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000bbb0bbb0)
  ) CLBLM_R_X7Y112_SLICE_X8Y112_DLUT (
.I0(CLBLM_L_X10Y104_SLICE_X12Y104_BO6),
.I1(CLBLM_L_X8Y114_SLICE_X11Y114_B5Q),
.I2(CLBLM_R_X7Y112_SLICE_X8Y112_DQ),
.I3(CLBLM_R_X5Y106_SLICE_X6Y106_CQ),
.I4(CLBLM_R_X7Y113_SLICE_X8Y113_DQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X7Y112_SLICE_X8Y112_DO5),
.O6(CLBLM_R_X7Y112_SLICE_X8Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcc33008b8b8888)
  ) CLBLM_R_X7Y112_SLICE_X8Y112_CLUT (
.I0(CLBLL_L_X4Y107_SLICE_X5Y107_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_L_X10Y112_SLICE_X12Y112_AQ),
.I4(CLBLM_R_X11Y112_SLICE_X14Y112_CQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y112_SLICE_X8Y112_CO5),
.O6(CLBLM_R_X7Y112_SLICE_X8Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000c0cff000c0c)
  ) CLBLM_R_X7Y112_SLICE_X8Y112_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y112_SLICE_X8Y112_BQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X7Y113_SLICE_X8Y113_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y112_SLICE_X8Y112_BO5),
.O6(CLBLM_R_X7Y112_SLICE_X8Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffbaba0000baba)
  ) CLBLM_R_X7Y112_SLICE_X8Y112_ALUT (
.I0(CLBLM_R_X7Y114_SLICE_X8Y114_DO6),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X7Y112_SLICE_X8Y112_AQ),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X10Y112_SLICE_X12Y112_AQ),
.O5(CLBLM_R_X7Y112_SLICE_X8Y112_AO5),
.O6(CLBLM_R_X7Y112_SLICE_X8Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y112_SLICE_X9Y112_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y112_SLICE_X9Y112_AO6),
.Q(CLBLM_R_X7Y112_SLICE_X9Y112_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y112_SLICE_X9Y112_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y112_SLICE_X9Y112_BO6),
.Q(CLBLM_R_X7Y112_SLICE_X9Y112_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0b0b0b0a0a0a0a)
  ) CLBLM_R_X7Y112_SLICE_X9Y112_DLUT (
.I0(CLBLM_R_X7Y109_SLICE_X8Y109_DO5),
.I1(RIOB33_X105Y121_IOB_X1Y121_I),
.I2(CLBLM_R_X7Y113_SLICE_X9Y113_CO6),
.I3(CLBLM_R_X7Y115_SLICE_X8Y115_CQ),
.I4(CLBLM_R_X5Y111_SLICE_X7Y111_CQ),
.I5(CLBLM_R_X3Y110_SLICE_X3Y110_AO6),
.O5(CLBLM_R_X7Y112_SLICE_X9Y112_DO5),
.O6(CLBLM_R_X7Y112_SLICE_X9Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0b0a0a0e0a0a0a)
  ) CLBLM_R_X7Y112_SLICE_X9Y112_CLUT (
.I0(CLBLM_R_X7Y109_SLICE_X8Y109_DO5),
.I1(RIOB33_X105Y121_IOB_X1Y121_I),
.I2(CLBLM_R_X7Y113_SLICE_X9Y113_CO6),
.I3(CLBLM_R_X11Y112_SLICE_X14Y112_CQ),
.I4(CLBLM_R_X3Y110_SLICE_X2Y110_DO6),
.I5(CLBLM_L_X8Y113_SLICE_X11Y113_BQ),
.O5(CLBLM_R_X7Y112_SLICE_X9Y112_CO5),
.O6(CLBLM_R_X7Y112_SLICE_X9Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0afafa0a0a0a0)
  ) CLBLM_R_X7Y112_SLICE_X9Y112_BLUT (
.I0(CLBLM_R_X5Y112_SLICE_X7Y112_DQ),
.I1(1'b1),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_L_X10Y111_SLICE_X13Y111_C5Q),
.O5(CLBLM_R_X7Y112_SLICE_X9Y112_BO5),
.O6(CLBLM_R_X7Y112_SLICE_X9Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f5f5f000050500)
  ) CLBLM_R_X7Y112_SLICE_X9Y112_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(1'b1),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y112_SLICE_X11Y112_DO6),
.I4(CLBLM_L_X8Y113_SLICE_X11Y113_AQ),
.I5(CLBLM_R_X7Y108_SLICE_X8Y108_CQ),
.O5(CLBLM_R_X7Y112_SLICE_X9Y112_AO5),
.O6(CLBLM_R_X7Y112_SLICE_X9Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y113_SLICE_X8Y113_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y113_SLICE_X8Y113_CO5),
.Q(CLBLM_R_X7Y113_SLICE_X8Y113_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y113_SLICE_X8Y113_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y113_SLICE_X8Y113_AO6),
.Q(CLBLM_R_X7Y113_SLICE_X8Y113_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y113_SLICE_X8Y113_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y113_SLICE_X8Y113_BO6),
.Q(CLBLM_R_X7Y113_SLICE_X8Y113_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y113_SLICE_X8Y113_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y113_SLICE_X8Y113_CO6),
.Q(CLBLM_R_X7Y113_SLICE_X8Y113_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y113_SLICE_X8Y113_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y113_SLICE_X8Y113_DO6),
.Q(CLBLM_R_X7Y113_SLICE_X8Y113_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000fafa5050)
  ) CLBLM_R_X7Y113_SLICE_X8Y113_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(1'b1),
.I2(CLBLM_R_X7Y113_SLICE_X8Y113_DQ),
.I3(1'b1),
.I4(CLBLM_L_X8Y113_SLICE_X11Y113_AQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X7Y113_SLICE_X8Y113_DO5),
.O6(CLBLM_R_X7Y113_SLICE_X8Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5a0a0ff55aa00)
  ) CLBLM_R_X7Y113_SLICE_X8Y113_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(1'b1),
.I2(CLBLM_R_X7Y107_SLICE_X8Y107_CQ),
.I3(CLBLM_R_X7Y113_SLICE_X8Y113_BQ),
.I4(RIOB33_X105Y101_IOB_X1Y101_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y113_SLICE_X8Y113_CO5),
.O6(CLBLM_R_X7Y113_SLICE_X8Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa0afa0afc0cfc0c)
  ) CLBLM_R_X7Y113_SLICE_X8Y113_BLUT (
.I0(CLBLM_R_X5Y109_SLICE_X7Y109_AQ),
.I1(CLBLM_R_X7Y113_SLICE_X8Y113_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y117_SLICE_X12Y117_A5Q),
.I4(1'b1),
.I5(CLBLL_L_X4Y112_SLICE_X4Y112_CO5),
.O5(CLBLM_R_X7Y113_SLICE_X8Y113_BO5),
.O6(CLBLM_R_X7Y113_SLICE_X8Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00aaaaff00f0f0)
  ) CLBLM_R_X7Y113_SLICE_X8Y113_ALUT (
.I0(CLBLM_L_X8Y113_SLICE_X10Y113_CQ),
.I1(1'b1),
.I2(CLBLM_R_X7Y113_SLICE_X8Y113_AQ),
.I3(CLBLM_R_X7Y114_SLICE_X8Y114_A5Q),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLL_L_X4Y112_SLICE_X4Y112_CO5),
.O5(CLBLM_R_X7Y113_SLICE_X8Y113_AO5),
.O6(CLBLM_R_X7Y113_SLICE_X8Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y113_SLICE_X9Y113_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y113_SLICE_X9Y113_BO5),
.Q(CLBLM_R_X7Y113_SLICE_X9Y113_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y113_SLICE_X9Y113_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y113_SLICE_X9Y113_AO6),
.Q(CLBLM_R_X7Y113_SLICE_X9Y113_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hee44eb41ee44eb41)
  ) CLBLM_R_X7Y113_SLICE_X9Y113_DLUT (
.I0(RIOB33_X105Y121_IOB_X1Y121_I),
.I1(CLBLM_L_X8Y109_SLICE_X10Y109_BQ),
.I2(CLBLM_R_X7Y114_SLICE_X9Y114_AO5),
.I3(CLBLM_R_X5Y114_SLICE_X7Y114_BQ),
.I4(CLBLM_R_X7Y117_SLICE_X9Y117_DQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y113_SLICE_X9Y113_DO5),
.O6(CLBLM_R_X7Y113_SLICE_X9Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffffae)
  ) CLBLM_R_X7Y113_SLICE_X9Y113_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y104_SLICE_X12Y104_AQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X7Y116_SLICE_X8Y116_CQ),
.I4(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_R_X7Y113_SLICE_X9Y113_CO5),
.O6(CLBLM_R_X7Y113_SLICE_X9Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfc0000f0aaf0aa)
  ) CLBLM_R_X7Y113_SLICE_X9Y113_BLUT (
.I0(CLBLM_R_X5Y116_SLICE_X6Y116_CQ),
.I1(CLBLM_L_X10Y111_SLICE_X13Y111_C5Q),
.I2(CLBLM_L_X8Y111_SLICE_X11Y111_BQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y113_SLICE_X9Y113_BO5),
.O6(CLBLM_R_X7Y113_SLICE_X9Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffcffa800fc00a8)
  ) CLBLM_R_X7Y113_SLICE_X9Y113_ALUT (
.I0(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.I1(CLBLM_L_X8Y112_SLICE_X10Y112_CO6),
.I2(CLBLM_R_X7Y113_SLICE_X9Y113_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLM_L_X10Y116_SLICE_X12Y116_CQ),
.O5(CLBLM_R_X7Y113_SLICE_X9Y113_AO5),
.O6(CLBLM_R_X7Y113_SLICE_X9Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y114_SLICE_X8Y114_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y114_SLICE_X8Y114_AO5),
.Q(CLBLM_R_X7Y114_SLICE_X8Y114_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y114_SLICE_X8Y114_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y114_SLICE_X8Y114_AO6),
.Q(CLBLM_R_X7Y114_SLICE_X8Y114_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y114_SLICE_X8Y114_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y114_SLICE_X8Y114_BO6),
.Q(CLBLM_R_X7Y114_SLICE_X8Y114_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y114_SLICE_X8Y114_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y114_SLICE_X8Y114_CO6),
.Q(CLBLM_R_X7Y114_SLICE_X8Y114_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000500000000)
  ) CLBLM_R_X7Y114_SLICE_X8Y114_DLUT (
.I0(CLBLL_L_X4Y110_SLICE_X4Y110_BQ),
.I1(1'b1),
.I2(CLBLM_R_X7Y114_SLICE_X9Y114_DO6),
.I3(CLBLM_L_X12Y108_SLICE_X16Y108_AQ),
.I4(CLBLM_L_X8Y115_SLICE_X10Y115_DO6),
.I5(CLBLM_R_X5Y113_SLICE_X7Y113_DO6),
.O5(CLBLM_R_X7Y114_SLICE_X8Y114_DO5),
.O6(CLBLM_R_X7Y114_SLICE_X8Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f01144f0f01144)
  ) CLBLM_R_X7Y114_SLICE_X8Y114_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X7Y111_SLICE_X9Y111_CQ),
.I2(CLBLM_R_X7Y117_SLICE_X9Y117_BQ),
.I3(CLBLM_L_X8Y113_SLICE_X11Y113_CO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y114_SLICE_X8Y114_CO5),
.O6(CLBLM_R_X7Y114_SLICE_X8Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hefef4545eaea4040)
  ) CLBLM_R_X7Y114_SLICE_X8Y114_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y114_SLICE_X8Y114_BQ),
.I2(CLBLL_L_X4Y112_SLICE_X4Y112_CO5),
.I3(1'b1),
.I4(CLBLM_R_X5Y113_SLICE_X7Y113_BQ),
.I5(CLBLM_L_X10Y115_SLICE_X12Y115_CQ),
.O5(CLBLM_R_X7Y114_SLICE_X8Y114_BO5),
.O6(CLBLM_R_X7Y114_SLICE_X8Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccff00fafaaaaa)
  ) CLBLM_R_X7Y114_SLICE_X8Y114_ALUT (
.I0(CLBLM_R_X7Y116_SLICE_X8Y116_DO6),
.I1(CLBLM_L_X10Y104_SLICE_X12Y104_AQ),
.I2(CLBLM_R_X5Y114_SLICE_X6Y114_AQ),
.I3(CLBLM_R_X3Y110_SLICE_X3Y110_AO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y114_SLICE_X8Y114_AO5),
.O6(CLBLM_R_X7Y114_SLICE_X8Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y114_SLICE_X9Y114_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y114_SLICE_X9Y114_BO6),
.Q(CLBLM_R_X7Y114_SLICE_X9Y114_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3ffffffffffffff)
  ) CLBLM_R_X7Y114_SLICE_X9Y114_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y113_SLICE_X10Y113_CQ),
.I2(CLBLM_R_X7Y111_SLICE_X8Y111_BQ),
.I3(CLBLM_R_X7Y112_SLICE_X9Y112_AQ),
.I4(CLBLM_R_X7Y110_SLICE_X9Y110_AQ),
.I5(CLBLM_R_X5Y113_SLICE_X6Y113_BQ),
.O5(CLBLM_R_X7Y114_SLICE_X9Y114_DO5),
.O6(CLBLM_R_X7Y114_SLICE_X9Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffefffafffafff)
  ) CLBLM_R_X7Y114_SLICE_X9Y114_CLUT (
.I0(CLBLM_R_X7Y114_SLICE_X9Y114_AO6),
.I1(CLBLM_L_X10Y114_SLICE_X13Y114_BQ),
.I2(CLBLM_R_X5Y116_SLICE_X6Y116_CQ),
.I3(CLBLM_R_X5Y116_SLICE_X7Y116_DO6),
.I4(CLBLM_L_X12Y112_SLICE_X17Y112_BQ),
.I5(CLBLL_L_X4Y116_SLICE_X4Y116_BO6),
.O5(CLBLM_R_X7Y114_SLICE_X9Y114_CO5),
.O6(CLBLM_R_X7Y114_SLICE_X9Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00fe54aa00fe54)
  ) CLBLM_R_X7Y114_SLICE_X9Y114_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y114_SLICE_X9Y114_BQ),
.I2(CLBLM_R_X5Y113_SLICE_X7Y113_BQ),
.I3(CLBLM_R_X11Y115_SLICE_X14Y115_AQ),
.I4(CLBLL_L_X4Y112_SLICE_X4Y112_CO5),
.I5(1'b1),
.O5(CLBLM_R_X7Y114_SLICE_X9Y114_BO5),
.O6(CLBLM_R_X7Y114_SLICE_X9Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfb04ff00ffffdddd)
  ) CLBLM_R_X7Y114_SLICE_X9Y114_ALUT (
.I0(CLBLM_R_X7Y111_SLICE_X8Y111_CQ),
.I1(CLBLM_L_X8Y114_SLICE_X10Y114_CQ),
.I2(CLBLM_R_X7Y117_SLICE_X9Y117_DQ),
.I3(CLBLM_R_X7Y115_SLICE_X8Y115_BQ),
.I4(CLBLM_L_X10Y112_SLICE_X12Y112_BQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y114_SLICE_X9Y114_AO5),
.O6(CLBLM_R_X7Y114_SLICE_X9Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y115_SLICE_X8Y115_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y115_SLICE_X8Y115_BO5),
.Q(CLBLM_R_X7Y115_SLICE_X8Y115_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y115_SLICE_X8Y115_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y115_SLICE_X8Y115_DO5),
.Q(CLBLM_R_X7Y115_SLICE_X8Y115_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y115_SLICE_X8Y115_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y115_SLICE_X8Y115_AO6),
.Q(CLBLM_R_X7Y115_SLICE_X8Y115_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y115_SLICE_X8Y115_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y115_SLICE_X8Y115_BO6),
.Q(CLBLM_R_X7Y115_SLICE_X8Y115_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y115_SLICE_X8Y115_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y115_SLICE_X8Y115_CO6),
.Q(CLBLM_R_X7Y115_SLICE_X8Y115_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y115_SLICE_X8Y115_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y115_SLICE_X8Y115_DO6),
.Q(CLBLM_R_X7Y115_SLICE_X8Y115_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfc0c0cafa0afa0)
  ) CLBLM_R_X7Y115_SLICE_X8Y115_DLUT (
.I0(CLBLM_R_X11Y114_SLICE_X14Y114_BQ),
.I1(CLBLM_L_X12Y113_SLICE_X17Y113_AQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X5Y116_SLICE_X7Y116_AQ),
.I4(CLBLM_L_X8Y118_SLICE_X10Y118_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y115_SLICE_X8Y115_DO5),
.O6(CLBLM_R_X7Y115_SLICE_X8Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00a0a0ff00a0a0)
  ) CLBLM_R_X7Y115_SLICE_X8Y115_CLUT (
.I0(CLBLM_R_X7Y112_SLICE_X8Y112_C5Q),
.I1(1'b1),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X7Y116_SLICE_X8Y116_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y115_SLICE_X8Y115_CO5),
.O6(CLBLM_R_X7Y115_SLICE_X8Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fc000ccacacaca)
  ) CLBLM_R_X7Y115_SLICE_X8Y115_BLUT (
.I0(CLBLM_R_X5Y115_SLICE_X7Y115_AQ),
.I1(CLBLM_R_X7Y115_SLICE_X8Y115_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X5Y115_SLICE_X6Y115_CQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y115_SLICE_X8Y115_BO5),
.O6(CLBLM_R_X7Y115_SLICE_X8Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0f0fcccc0005)
  ) CLBLM_R_X7Y115_SLICE_X8Y115_ALUT (
.I0(CLBLM_R_X7Y118_SLICE_X8Y118_CQ),
.I1(CLBLM_R_X3Y109_SLICE_X2Y109_AQ),
.I2(CLBLM_L_X8Y118_SLICE_X10Y118_AQ),
.I3(CLBLM_L_X10Y119_SLICE_X12Y119_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y114_SLICE_X8Y114_A5Q),
.O5(CLBLM_R_X7Y115_SLICE_X8Y115_AO5),
.O6(CLBLM_R_X7Y115_SLICE_X8Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y115_SLICE_X9Y115_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y115_SLICE_X9Y115_CO5),
.Q(CLBLM_R_X7Y115_SLICE_X9Y115_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y115_SLICE_X9Y115_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y115_SLICE_X9Y115_BO5),
.Q(CLBLM_R_X7Y115_SLICE_X9Y115_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y115_SLICE_X9Y115_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y115_SLICE_X9Y115_AO6),
.Q(CLBLM_R_X7Y115_SLICE_X9Y115_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y115_SLICE_X9Y115_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y115_SLICE_X9Y115_BO6),
.Q(CLBLM_R_X7Y115_SLICE_X9Y115_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000505)
  ) CLBLM_R_X7Y115_SLICE_X9Y115_DLUT (
.I0(CLBLM_R_X7Y115_SLICE_X8Y115_D5Q),
.I1(1'b1),
.I2(CLBLM_R_X7Y115_SLICE_X8Y115_B5Q),
.I3(1'b1),
.I4(CLBLM_R_X5Y115_SLICE_X6Y115_DO6),
.I5(CLBLM_R_X5Y116_SLICE_X6Y116_D5Q),
.O5(CLBLM_R_X7Y115_SLICE_X9Y115_DO5),
.O6(CLBLM_R_X7Y115_SLICE_X9Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0c000000f202f202)
  ) CLBLM_R_X7Y115_SLICE_X9Y115_CLUT (
.I0(CLBLL_L_X4Y110_SLICE_X4Y110_BQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y112_SLICE_X12Y112_C5Q),
.I4(CLBLM_L_X12Y112_SLICE_X16Y112_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X7Y115_SLICE_X9Y115_CO5),
.O6(CLBLM_R_X7Y115_SLICE_X9Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f03300ff00aaaa)
  ) CLBLM_R_X7Y115_SLICE_X9Y115_BLUT (
.I0(CLBLM_R_X7Y117_SLICE_X9Y117_A5Q),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X7Y109_SLICE_X9Y109_DQ),
.I3(CLBLM_L_X12Y112_SLICE_X17Y112_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y115_SLICE_X9Y115_BO5),
.O6(CLBLM_R_X7Y115_SLICE_X9Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfaff5055faaa5000)
  ) CLBLM_R_X7Y115_SLICE_X9Y115_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(1'b1),
.I2(CLBLM_R_X7Y115_SLICE_X9Y115_AQ),
.I3(CLBLL_L_X4Y116_SLICE_X4Y116_BO6),
.I4(CLBLM_R_X7Y115_SLICE_X8Y115_AQ),
.I5(CLBLM_L_X10Y114_SLICE_X12Y114_BQ),
.O5(CLBLM_R_X7Y115_SLICE_X9Y115_AO5),
.O6(CLBLM_R_X7Y115_SLICE_X9Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y116_SLICE_X8Y116_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y116_SLICE_X8Y116_AO6),
.Q(CLBLM_R_X7Y116_SLICE_X8Y116_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y116_SLICE_X8Y116_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y116_SLICE_X8Y116_BO6),
.Q(CLBLM_R_X7Y116_SLICE_X8Y116_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y116_SLICE_X8Y116_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y116_SLICE_X8Y116_CO6),
.Q(CLBLM_R_X7Y116_SLICE_X8Y116_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h2288aa000288aa00)
  ) CLBLM_R_X7Y116_SLICE_X8Y116_DLUT (
.I0(CLBLM_R_X5Y116_SLICE_X6Y116_AO5),
.I1(CLBLM_R_X11Y117_SLICE_X15Y117_AQ),
.I2(CLBLM_L_X8Y118_SLICE_X10Y118_AQ),
.I3(CLBLM_R_X7Y114_SLICE_X8Y114_A5Q),
.I4(CLBLM_R_X7Y118_SLICE_X9Y118_BO5),
.I5(CLBLM_L_X10Y117_SLICE_X13Y117_CO6),
.O5(CLBLM_R_X7Y116_SLICE_X8Y116_DO5),
.O6(CLBLM_R_X7Y116_SLICE_X8Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00fefeff000404)
  ) CLBLM_R_X7Y116_SLICE_X8Y116_CLUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_R_X7Y116_SLICE_X8Y116_CQ),
.I2(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.I3(CLBLL_L_X4Y118_SLICE_X4Y118_A5Q),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X10Y113_SLICE_X13Y113_AQ),
.O5(CLBLM_R_X7Y116_SLICE_X8Y116_CO5),
.O6(CLBLM_R_X7Y116_SLICE_X8Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000fafa5050)
  ) CLBLM_R_X7Y116_SLICE_X8Y116_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(1'b1),
.I2(CLBLM_R_X7Y116_SLICE_X8Y116_AQ),
.I3(1'b1),
.I4(CLBLM_L_X10Y113_SLICE_X12Y113_AQ),
.I5(CLBLM_L_X10Y116_SLICE_X12Y116_DO6),
.O5(CLBLM_R_X7Y116_SLICE_X8Y116_BO5),
.O6(CLBLM_R_X7Y116_SLICE_X8Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0f5a0f5a0a0a0a0)
  ) CLBLM_R_X7Y116_SLICE_X8Y116_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(1'b1),
.I2(CLBLM_L_X8Y115_SLICE_X11Y115_BQ),
.I3(CLBLM_L_X10Y116_SLICE_X12Y116_DO6),
.I4(1'b1),
.I5(CLBLM_R_X7Y117_SLICE_X8Y117_AQ),
.O5(CLBLM_R_X7Y116_SLICE_X8Y116_AO5),
.O6(CLBLM_R_X7Y116_SLICE_X8Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y116_SLICE_X9Y116_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y116_SLICE_X9Y116_AO6),
.Q(CLBLM_R_X7Y116_SLICE_X9Y116_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h55555fff5fff5fff)
  ) CLBLM_R_X7Y116_SLICE_X9Y116_DLUT (
.I0(CLBLM_R_X5Y116_SLICE_X7Y116_BQ),
.I1(1'b1),
.I2(CLBLM_R_X5Y115_SLICE_X7Y115_AQ),
.I3(CLBLM_R_X5Y116_SLICE_X6Y116_CQ),
.I4(CLBLM_R_X7Y116_SLICE_X9Y116_AQ),
.I5(CLBLM_R_X5Y115_SLICE_X6Y115_BQ),
.O5(CLBLM_R_X7Y116_SLICE_X9Y116_DO5),
.O6(CLBLM_R_X7Y116_SLICE_X9Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha556aa56a566aa66)
  ) CLBLM_R_X7Y116_SLICE_X9Y116_CLUT (
.I0(CLBLL_L_X4Y108_SLICE_X5Y108_AO6),
.I1(CLBLM_R_X7Y114_SLICE_X8Y114_A5Q),
.I2(CLBLM_L_X8Y118_SLICE_X10Y118_AQ),
.I3(CLBLM_L_X10Y115_SLICE_X13Y115_CQ),
.I4(CLBLM_R_X7Y118_SLICE_X8Y118_CQ),
.I5(CLBLM_L_X10Y119_SLICE_X12Y119_AQ),
.O5(CLBLM_R_X7Y116_SLICE_X9Y116_CO5),
.O6(CLBLM_R_X7Y116_SLICE_X9Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haabfbfbfc0000000)
  ) CLBLM_R_X7Y116_SLICE_X9Y116_BLUT (
.I0(CLBLM_R_X7Y116_SLICE_X9Y116_DO6),
.I1(CLBLM_R_X7Y117_SLICE_X9Y117_A5Q),
.I2(CLBLM_R_X7Y117_SLICE_X9Y117_AQ),
.I3(CLBLM_R_X7Y117_SLICE_X9Y117_BQ),
.I4(CLBLM_R_X5Y116_SLICE_X7Y116_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y116_SLICE_X9Y116_BO5),
.O6(CLBLM_R_X7Y116_SLICE_X9Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff7800000078)
  ) CLBLM_R_X7Y116_SLICE_X9Y116_ALUT (
.I0(CLBLM_R_X7Y116_SLICE_X9Y116_BO5),
.I1(CLBLM_R_X5Y115_SLICE_X6Y115_BQ),
.I2(CLBLM_R_X7Y116_SLICE_X9Y116_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y132_SLICE_X9Y132_AO6),
.I5(CLBLM_L_X8Y112_SLICE_X10Y112_AQ),
.O5(CLBLM_R_X7Y116_SLICE_X9Y116_AO5),
.O6(CLBLM_R_X7Y116_SLICE_X9Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y117_SLICE_X8Y117_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y117_SLICE_X8Y117_AO6),
.Q(CLBLM_R_X7Y117_SLICE_X8Y117_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y117_SLICE_X8Y117_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y117_SLICE_X8Y117_BO6),
.Q(CLBLM_R_X7Y117_SLICE_X8Y117_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y117_SLICE_X8Y117_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y117_SLICE_X8Y117_DO5),
.O6(CLBLM_R_X7Y117_SLICE_X8Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y117_SLICE_X8Y117_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y117_SLICE_X8Y117_CO5),
.O6(CLBLM_R_X7Y117_SLICE_X8Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haf05aa00af05aa00)
  ) CLBLM_R_X7Y117_SLICE_X8Y117_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(1'b1),
.I2(CLBLM_L_X10Y116_SLICE_X12Y116_DO6),
.I3(CLBLL_L_X4Y115_SLICE_X5Y115_BQ),
.I4(CLBLM_L_X8Y116_SLICE_X11Y116_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y117_SLICE_X8Y117_BO5),
.O6(CLBLM_R_X7Y117_SLICE_X8Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaafcfcaaaafcfc)
  ) CLBLM_R_X7Y117_SLICE_X8Y117_ALUT (
.I0(CLBLM_L_X8Y111_SLICE_X10Y111_A5Q),
.I1(CLBLM_R_X7Y117_SLICE_X8Y117_BQ),
.I2(CLBLM_L_X10Y116_SLICE_X12Y116_DO6),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y117_SLICE_X8Y117_AO5),
.O6(CLBLM_R_X7Y117_SLICE_X8Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y117_SLICE_X9Y117_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y117_SLICE_X9Y117_CO6),
.Q(CLBLM_R_X7Y117_SLICE_X9Y117_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y117_SLICE_X9Y117_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y117_SLICE_X9Y117_AO6),
.Q(CLBLM_R_X7Y117_SLICE_X9Y117_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y117_SLICE_X9Y117_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y117_SLICE_X9Y117_BO6),
.Q(CLBLM_R_X7Y117_SLICE_X9Y117_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y117_SLICE_X9Y117_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y117_SLICE_X9Y117_DO6),
.Q(CLBLM_R_X7Y117_SLICE_X9Y117_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hbabaaaaa10100000)
  ) CLBLM_R_X7Y117_SLICE_X9Y117_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y112_SLICE_X8Y112_CQ),
.I2(CLBLM_R_X7Y117_SLICE_X9Y117_DQ),
.I3(1'b1),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLL_L_X4Y117_SLICE_X4Y117_AQ),
.O5(CLBLM_R_X7Y117_SLICE_X9Y117_DO5),
.O6(CLBLM_R_X7Y117_SLICE_X9Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcacfcfcaff000000)
  ) CLBLM_R_X7Y117_SLICE_X9Y117_CLUT (
.I0(CLBLM_R_X7Y132_SLICE_X9Y132_AO6),
.I1(CLBLM_L_X8Y110_SLICE_X11Y110_DQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y117_SLICE_X9Y117_A5Q),
.I4(CLBLM_R_X7Y117_SLICE_X9Y117_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y117_SLICE_X9Y117_CO5),
.O6(CLBLM_R_X7Y117_SLICE_X9Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'habaeaeae01040404)
  ) CLBLM_R_X7Y117_SLICE_X9Y117_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y117_SLICE_X9Y117_BQ),
.I2(CLBLM_R_X7Y132_SLICE_X9Y132_AO6),
.I3(CLBLM_R_X5Y116_SLICE_X7Y116_AQ),
.I4(CLBLM_R_X7Y117_SLICE_X9Y117_CO5),
.I5(CLBLM_R_X7Y112_SLICE_X8Y112_CQ),
.O5(CLBLM_R_X7Y117_SLICE_X9Y117_BO5),
.O6(CLBLM_R_X7Y117_SLICE_X9Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff7fffff007f00ff)
  ) CLBLM_R_X7Y117_SLICE_X9Y117_ALUT (
.I0(CLBLM_L_X10Y112_SLICE_X12Y112_C5Q),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X7Y117_SLICE_X9Y117_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X12Y112_SLICE_X16Y112_B5Q),
.I5(CLBLM_L_X8Y109_SLICE_X11Y109_BQ),
.O5(CLBLM_R_X7Y117_SLICE_X9Y117_AO5),
.O6(CLBLM_R_X7Y117_SLICE_X9Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y118_SLICE_X8Y118_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y118_SLICE_X8Y118_AO6),
.Q(CLBLM_R_X7Y118_SLICE_X8Y118_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y118_SLICE_X8Y118_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y118_SLICE_X8Y118_BO6),
.Q(CLBLM_R_X7Y118_SLICE_X8Y118_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y118_SLICE_X8Y118_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y118_SLICE_X8Y118_CO6),
.Q(CLBLM_R_X7Y118_SLICE_X8Y118_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000008)
  ) CLBLM_R_X7Y118_SLICE_X8Y118_DLUT (
.I0(CLBLM_R_X7Y117_SLICE_X8Y117_BQ),
.I1(CLBLM_R_X11Y117_SLICE_X15Y117_AQ),
.I2(CLBLM_R_X7Y118_SLICE_X8Y118_BQ),
.I3(CLBLM_R_X7Y118_SLICE_X9Y118_AQ),
.I4(CLBLM_R_X7Y118_SLICE_X8Y118_AQ),
.I5(CLBLM_R_X7Y114_SLICE_X8Y114_A5Q),
.O5(CLBLM_R_X7Y118_SLICE_X8Y118_DO5),
.O6(CLBLM_R_X7Y118_SLICE_X8Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000ff00e4e4)
  ) CLBLM_R_X7Y118_SLICE_X8Y118_CLUT (
.I0(CLBLM_L_X10Y117_SLICE_X13Y117_CO6),
.I1(CLBLM_R_X7Y118_SLICE_X8Y118_CQ),
.I2(CLBLM_L_X10Y119_SLICE_X12Y119_AQ),
.I3(CLBLL_L_X4Y118_SLICE_X4Y118_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y121_IOB_X1Y121_I),
.O5(CLBLM_R_X7Y118_SLICE_X8Y118_CO5),
.O6(CLBLM_R_X7Y118_SLICE_X8Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0e4e4e4e4a0a0)
  ) CLBLM_R_X7Y118_SLICE_X8Y118_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y118_SLICE_X9Y118_BO6),
.I2(CLBLM_R_X7Y114_SLICE_X8Y114_BQ),
.I3(1'b1),
.I4(CLBLM_R_X7Y117_SLICE_X8Y117_BQ),
.I5(CLBLM_R_X7Y118_SLICE_X8Y118_BQ),
.O5(CLBLM_R_X7Y118_SLICE_X8Y118_BO5),
.O6(CLBLM_R_X7Y118_SLICE_X8Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'he4a0e4a0a0e4e4a0)
  ) CLBLM_R_X7Y118_SLICE_X8Y118_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y118_SLICE_X9Y118_BO6),
.I2(CLBLM_L_X8Y113_SLICE_X10Y113_AQ),
.I3(CLBLM_R_X7Y118_SLICE_X8Y118_AQ),
.I4(CLBLM_R_X7Y117_SLICE_X8Y117_BQ),
.I5(CLBLM_R_X7Y118_SLICE_X8Y118_BQ),
.O5(CLBLM_R_X7Y118_SLICE_X8Y118_AO5),
.O6(CLBLM_R_X7Y118_SLICE_X8Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y118_SLICE_X9Y118_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y118_SLICE_X9Y118_AO6),
.Q(CLBLM_R_X7Y118_SLICE_X9Y118_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y118_SLICE_X9Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y118_SLICE_X9Y118_DO5),
.O6(CLBLM_R_X7Y118_SLICE_X9Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000f0000000100)
  ) CLBLM_R_X7Y118_SLICE_X9Y118_CLUT (
.I0(CLBLM_L_X8Y116_SLICE_X11Y116_CO6),
.I1(CLBLM_R_X7Y118_SLICE_X9Y118_AQ),
.I2(CLBLM_R_X7Y118_SLICE_X8Y118_AQ),
.I3(CLBLM_R_X7Y117_SLICE_X8Y117_BQ),
.I4(CLBLM_R_X7Y118_SLICE_X8Y118_BQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y118_SLICE_X9Y118_CO5),
.O6(CLBLM_R_X7Y118_SLICE_X9Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0d00000022)
  ) CLBLM_R_X7Y118_SLICE_X9Y118_BLUT (
.I0(CLBLM_R_X7Y117_SLICE_X8Y117_BQ),
.I1(CLBLM_R_X7Y118_SLICE_X8Y118_AQ),
.I2(CLBLM_L_X10Y117_SLICE_X13Y117_AO5),
.I3(CLBLM_R_X7Y118_SLICE_X8Y118_BQ),
.I4(CLBLM_R_X7Y118_SLICE_X9Y118_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y118_SLICE_X9Y118_BO5),
.O6(CLBLM_R_X7Y118_SLICE_X9Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdddd8d8dddddd8d8)
  ) CLBLM_R_X7Y118_SLICE_X9Y118_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y111_SLICE_X8Y111_BQ),
.I2(CLBLM_R_X7Y118_SLICE_X9Y118_AQ),
.I3(1'b1),
.I4(CLBLM_L_X10Y117_SLICE_X13Y117_AO5),
.I5(CLBLM_R_X7Y118_SLICE_X9Y118_CO6),
.O5(CLBLM_R_X7Y118_SLICE_X9Y118_AO5),
.O6(CLBLM_R_X7Y118_SLICE_X9Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y132_SLICE_X8Y132_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y132_SLICE_X8Y132_DO5),
.O6(CLBLM_R_X7Y132_SLICE_X8Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y132_SLICE_X8Y132_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y132_SLICE_X8Y132_CO5),
.O6(CLBLM_R_X7Y132_SLICE_X8Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y132_SLICE_X8Y132_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y132_SLICE_X8Y132_BO5),
.O6(CLBLM_R_X7Y132_SLICE_X8Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y132_SLICE_X8Y132_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y132_SLICE_X8Y132_AO5),
.O6(CLBLM_R_X7Y132_SLICE_X8Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y132_SLICE_X9Y132_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y132_SLICE_X9Y132_DO5),
.O6(CLBLM_R_X7Y132_SLICE_X9Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y132_SLICE_X9Y132_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y132_SLICE_X9Y132_CO5),
.O6(CLBLM_R_X7Y132_SLICE_X9Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y132_SLICE_X9Y132_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y132_SLICE_X9Y132_BO5),
.O6(CLBLM_R_X7Y132_SLICE_X9Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5f5fffffcc000000)
  ) CLBLM_R_X7Y132_SLICE_X9Y132_ALUT (
.I0(CLBLM_L_X10Y112_SLICE_X12Y112_C5Q),
.I1(RIOB33_X105Y139_IOB_X1Y140_I),
.I2(CLBLM_L_X12Y112_SLICE_X16Y112_B5Q),
.I3(RIOB33_X105Y141_IOB_X1Y141_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y132_SLICE_X9Y132_AO5),
.O6(CLBLM_R_X7Y132_SLICE_X9Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y105_SLICE_X14Y105_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y105_SLICE_X14Y105_CO5),
.Q(CLBLM_R_X11Y105_SLICE_X14Y105_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y105_SLICE_X14Y105_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y105_SLICE_X14Y105_AO6),
.Q(CLBLM_R_X11Y105_SLICE_X14Y105_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y105_SLICE_X14Y105_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y105_SLICE_X14Y105_BO6),
.Q(CLBLM_R_X11Y105_SLICE_X14Y105_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y105_SLICE_X14Y105_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y105_SLICE_X14Y105_CO6),
.Q(CLBLM_R_X11Y105_SLICE_X14Y105_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y105_SLICE_X14Y105_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y105_SLICE_X14Y105_DO6),
.Q(CLBLM_R_X11Y105_SLICE_X14Y105_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffbaffbe55105514)
  ) CLBLM_R_X11Y105_SLICE_X14Y105_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X11Y106_SLICE_X15Y106_DO5),
.I2(CLBLM_R_X11Y105_SLICE_X14Y105_DQ),
.I3(CLBLM_L_X12Y105_SLICE_X16Y105_BO6),
.I4(CLBLM_L_X12Y105_SLICE_X17Y105_AO6),
.I5(CLBLL_L_X4Y107_SLICE_X4Y107_AQ),
.O5(CLBLM_R_X11Y105_SLICE_X14Y105_DO5),
.O6(CLBLM_R_X11Y105_SLICE_X14Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaaff00f8f8f8f8)
  ) CLBLM_R_X11Y105_SLICE_X14Y105_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLL_L_X4Y112_SLICE_X4Y112_BQ),
.I2(CLBLM_L_X10Y105_SLICE_X13Y105_AO6),
.I3(CLBLM_L_X10Y105_SLICE_X13Y105_BO6),
.I4(CLBLM_R_X13Y107_SLICE_X19Y107_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y105_SLICE_X14Y105_CO5),
.O6(CLBLM_R_X11Y105_SLICE_X14Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff88f0000088f0)
  ) CLBLM_R_X11Y105_SLICE_X14Y105_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X11Y105_SLICE_X14Y105_BQ),
.I2(CLBLM_L_X10Y111_SLICE_X13Y111_BQ),
.I3(CLBLM_L_X10Y106_SLICE_X12Y106_BO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X13Y112_SLICE_X18Y112_BQ),
.O5(CLBLM_R_X11Y105_SLICE_X14Y105_BO5),
.O6(CLBLM_R_X11Y105_SLICE_X14Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hecffeccc20332000)
  ) CLBLM_R_X11Y105_SLICE_X14Y105_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X11Y105_SLICE_X14Y105_AQ),
.I3(CLBLM_L_X10Y106_SLICE_X12Y106_BO6),
.I4(CLBLM_L_X10Y105_SLICE_X12Y105_BQ),
.I5(CLBLM_R_X11Y105_SLICE_X15Y105_CQ),
.O5(CLBLM_R_X11Y105_SLICE_X14Y105_AO5),
.O6(CLBLM_R_X11Y105_SLICE_X14Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y105_SLICE_X15Y105_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y105_SLICE_X15Y105_DO6),
.Q(CLBLM_R_X11Y105_SLICE_X15Y105_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y105_SLICE_X15Y105_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y105_SLICE_X15Y105_AO6),
.Q(CLBLM_R_X11Y105_SLICE_X15Y105_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y105_SLICE_X15Y105_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y105_SLICE_X15Y105_BO6),
.Q(CLBLM_R_X11Y105_SLICE_X15Y105_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y105_SLICE_X15Y105_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y105_SLICE_X15Y105_CO6),
.Q(CLBLM_R_X11Y105_SLICE_X15Y105_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'heffe455400f000f0)
  ) CLBLM_R_X11Y105_SLICE_X15Y105_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X12Y105_SLICE_X16Y105_BO6),
.I2(CLBLM_L_X12Y112_SLICE_X16Y112_CQ),
.I3(CLBLM_R_X11Y105_SLICE_X15Y105_A5Q),
.I4(CLBLM_L_X10Y111_SLICE_X12Y111_BQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y105_SLICE_X15Y105_DO5),
.O6(CLBLM_R_X11Y105_SLICE_X15Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hafef0545aaea0040)
  ) CLBLM_R_X11Y105_SLICE_X15Y105_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X11Y105_SLICE_X15Y105_CQ),
.I2(CLBLM_L_X12Y105_SLICE_X16Y105_CO5),
.I3(CLBLM_L_X12Y105_SLICE_X16Y105_BO6),
.I4(CLBLM_R_X7Y105_SLICE_X9Y105_CQ),
.I5(CLBLM_L_X12Y108_SLICE_X17Y108_BQ),
.O5(CLBLM_R_X11Y105_SLICE_X15Y105_CO5),
.O6(CLBLM_R_X11Y105_SLICE_X15Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff030003ff0e000e)
  ) CLBLM_R_X11Y105_SLICE_X15Y105_BLUT (
.I0(CLBLM_L_X12Y105_SLICE_X16Y105_BO5),
.I1(CLBLM_R_X11Y105_SLICE_X15Y105_BQ),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X11Y112_SLICE_X15Y112_AQ),
.I5(CLBLM_R_X11Y106_SLICE_X15Y106_CO6),
.O5(CLBLM_R_X11Y105_SLICE_X15Y105_BO5),
.O6(CLBLM_R_X11Y105_SLICE_X15Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0000cccc0550)
  ) CLBLM_R_X11Y105_SLICE_X15Y105_ALUT (
.I0(CLBLM_R_X11Y106_SLICE_X15Y106_DO5),
.I1(CLBLM_R_X11Y115_SLICE_X14Y115_BQ),
.I2(CLBLM_R_X11Y105_SLICE_X15Y105_AQ),
.I3(CLBLM_R_X11Y105_SLICE_X15Y105_DO5),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X12Y105_SLICE_X16Y105_BO6),
.O5(CLBLM_R_X11Y105_SLICE_X15Y105_AO5),
.O6(CLBLM_R_X11Y105_SLICE_X15Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y106_SLICE_X14Y106_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y106_SLICE_X14Y106_AO6),
.Q(CLBLM_R_X11Y106_SLICE_X14Y106_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y106_SLICE_X14Y106_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y106_SLICE_X14Y106_BO6),
.Q(CLBLM_R_X11Y106_SLICE_X14Y106_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y106_SLICE_X14Y106_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y106_SLICE_X14Y106_CO6),
.Q(CLBLM_R_X11Y106_SLICE_X14Y106_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y106_SLICE_X14Y106_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y106_SLICE_X14Y106_DO6),
.Q(CLBLM_R_X11Y106_SLICE_X14Y106_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ffa8000000a8)
  ) CLBLM_R_X11Y106_SLICE_X14Y106_DLUT (
.I0(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.I1(CLBLM_R_X11Y109_SLICE_X14Y109_AQ),
.I2(CLBLM_R_X11Y106_SLICE_X14Y106_DQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLM_R_X11Y105_SLICE_X14Y105_BQ),
.O5(CLBLM_R_X11Y106_SLICE_X14Y106_DO5),
.O6(CLBLM_R_X11Y106_SLICE_X14Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf505f000fd0df808)
  ) CLBLM_R_X11Y106_SLICE_X14Y106_CLUT (
.I0(CLBLM_L_X12Y105_SLICE_X16Y105_CO5),
.I1(CLBLM_R_X11Y106_SLICE_X14Y106_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X3Y113_SLICE_X3Y113_AQ),
.I4(CLBLM_L_X12Y107_SLICE_X16Y107_DQ),
.I5(CLBLM_L_X12Y105_SLICE_X16Y105_BO6),
.O5(CLBLM_R_X11Y106_SLICE_X14Y106_CO5),
.O6(CLBLM_R_X11Y106_SLICE_X14Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00f3f3ff00fcfc)
  ) CLBLM_R_X11Y106_SLICE_X14Y106_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y106_SLICE_X14Y106_BQ),
.I2(CLBLM_L_X12Y105_SLICE_X16Y105_BO6),
.I3(CLBLM_R_X7Y106_SLICE_X8Y106_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X11Y106_SLICE_X15Y106_DO6),
.O5(CLBLM_R_X11Y106_SLICE_X14Y106_BO5),
.O6(CLBLM_R_X11Y106_SLICE_X14Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000ccd8ccd8)
  ) CLBLM_R_X11Y106_SLICE_X14Y106_ALUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_R_X11Y106_SLICE_X14Y106_DQ),
.I2(CLBLM_R_X11Y106_SLICE_X14Y106_AQ),
.I3(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.I4(CLBLM_L_X12Y111_SLICE_X16Y111_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y106_SLICE_X14Y106_AO5),
.O6(CLBLM_R_X11Y106_SLICE_X14Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y106_SLICE_X15Y106_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y106_SLICE_X15Y106_AO6),
.Q(CLBLM_R_X11Y106_SLICE_X15Y106_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000110000000100)
  ) CLBLM_R_X11Y106_SLICE_X15Y106_DLUT (
.I0(CLBLM_R_X11Y105_SLICE_X15Y105_A5Q),
.I1(CLBLM_R_X11Y105_SLICE_X15Y105_AQ),
.I2(CLBLM_R_X11Y106_SLICE_X14Y106_BQ),
.I3(CLBLM_L_X12Y112_SLICE_X16Y112_CQ),
.I4(CLBLM_R_X11Y106_SLICE_X15Y106_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y106_SLICE_X15Y106_DO5),
.O6(CLBLM_R_X11Y106_SLICE_X15Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ff005050cccc)
  ) CLBLM_R_X11Y106_SLICE_X15Y106_CLUT (
.I0(CLBLM_L_X12Y105_SLICE_X16Y105_BO6),
.I1(CLBLM_L_X12Y108_SLICE_X17Y108_BQ),
.I2(CLBLM_R_X11Y105_SLICE_X15Y105_CQ),
.I3(CLBLM_R_X11Y108_SLICE_X14Y108_AQ),
.I4(CLBLM_L_X12Y105_SLICE_X16Y105_CO5),
.I5(1'b1),
.O5(CLBLM_R_X11Y106_SLICE_X15Y106_CO5),
.O6(CLBLM_R_X11Y106_SLICE_X15Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccaaaa00300030)
  ) CLBLM_R_X11Y106_SLICE_X15Y106_BLUT (
.I0(CLBLM_L_X10Y111_SLICE_X12Y111_A5Q),
.I1(CLBLM_R_X11Y105_SLICE_X15Y105_AQ),
.I2(CLBLM_L_X12Y112_SLICE_X16Y112_CQ),
.I3(CLBLM_R_X11Y105_SLICE_X15Y105_A5Q),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y106_SLICE_X15Y106_BO5),
.O6(CLBLM_R_X11Y106_SLICE_X15Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff001212ff001010)
  ) CLBLM_R_X11Y106_SLICE_X15Y106_ALUT (
.I0(CLBLM_R_X11Y106_SLICE_X15Y106_BO5),
.I1(CLBLM_L_X12Y105_SLICE_X16Y105_BO6),
.I2(CLBLM_R_X11Y106_SLICE_X15Y106_AQ),
.I3(CLBLM_R_X11Y106_SLICE_X14Y106_DQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X11Y106_SLICE_X14Y106_BQ),
.O5(CLBLM_R_X11Y106_SLICE_X15Y106_AO5),
.O6(CLBLM_R_X11Y106_SLICE_X15Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hbb88bb88bb88aaaa)
  ) CLBLM_R_X11Y107_SLICE_X14Y107_DLUT (
.I0(CLBLM_L_X8Y109_SLICE_X10Y109_C5Q),
.I1(CLBLM_R_X5Y115_SLICE_X7Y115_DO6),
.I2(1'b1),
.I3(CLBLM_R_X11Y107_SLICE_X14Y107_CO6),
.I4(CLBLM_R_X3Y110_SLICE_X2Y110_BO6),
.I5(CLBLL_L_X4Y107_SLICE_X5Y107_BO6),
.O5(CLBLM_R_X11Y107_SLICE_X14Y107_DO5),
.O6(CLBLM_R_X11Y107_SLICE_X14Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdfd0202ffff0000)
  ) CLBLM_R_X11Y107_SLICE_X14Y107_CLUT (
.I0(CLBLM_R_X11Y105_SLICE_X14Y105_C5Q),
.I1(CLBLM_R_X11Y105_SLICE_X14Y105_CQ),
.I2(CLBLM_L_X10Y106_SLICE_X12Y106_AQ),
.I3(1'b1),
.I4(CLBLM_R_X11Y110_SLICE_X14Y110_CQ),
.I5(CLBLM_L_X10Y105_SLICE_X12Y105_AQ),
.O5(CLBLM_R_X11Y107_SLICE_X14Y107_CO5),
.O6(CLBLM_R_X11Y107_SLICE_X14Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffdfffffffdd)
  ) CLBLM_R_X11Y107_SLICE_X14Y107_BLUT (
.I0(RIOB33_X105Y137_IOB_X1Y137_I),
.I1(RIOB33_X105Y129_IOB_X1Y129_I),
.I2(CLBLM_L_X8Y107_SLICE_X11Y107_BQ),
.I3(CLBLM_L_X12Y109_SLICE_X16Y109_AQ),
.I4(CLBLM_L_X10Y116_SLICE_X13Y116_AQ),
.I5(CLBLM_L_X8Y107_SLICE_X11Y107_B5Q),
.O5(CLBLM_R_X11Y107_SLICE_X14Y107_BO5),
.O6(CLBLM_R_X11Y107_SLICE_X14Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0000fe01ff00)
  ) CLBLM_R_X11Y107_SLICE_X14Y107_ALUT (
.I0(CLBLM_R_X11Y105_SLICE_X14Y105_CQ),
.I1(CLBLM_L_X10Y105_SLICE_X12Y105_AQ),
.I2(CLBLM_L_X10Y106_SLICE_X12Y106_AQ),
.I3(CLBLM_L_X8Y115_SLICE_X11Y115_BQ),
.I4(CLBLM_R_X11Y105_SLICE_X14Y105_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X11Y107_SLICE_X14Y107_AO5),
.O6(CLBLM_R_X11Y107_SLICE_X14Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y107_SLICE_X15Y107_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y107_SLICE_X15Y107_AO6),
.Q(CLBLM_R_X11Y107_SLICE_X15Y107_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y107_SLICE_X15Y107_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y107_SLICE_X15Y107_BO6),
.Q(CLBLM_R_X11Y107_SLICE_X15Y107_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y107_SLICE_X15Y107_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y107_SLICE_X15Y107_CO6),
.Q(CLBLM_R_X11Y107_SLICE_X15Y107_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0053005c0050005f)
  ) CLBLM_R_X11Y107_SLICE_X15Y107_DLUT (
.I0(CLBLM_L_X8Y109_SLICE_X10Y109_C5Q),
.I1(CLBLM_R_X11Y108_SLICE_X15Y108_AO5),
.I2(CLBLM_R_X5Y115_SLICE_X7Y115_CO6),
.I3(CLBLM_R_X11Y107_SLICE_X15Y107_AQ),
.I4(CLBLM_R_X11Y110_SLICE_X14Y110_CQ),
.I5(CLBLM_R_X11Y107_SLICE_X14Y107_AO6),
.O5(CLBLM_R_X11Y107_SLICE_X15Y107_DO5),
.O6(CLBLM_R_X11Y107_SLICE_X15Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hafae0504aaaa0000)
  ) CLBLM_R_X11Y107_SLICE_X15Y107_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X11Y107_SLICE_X15Y107_CQ),
.I2(RIOB33_X105Y117_IOB_X1Y118_I),
.I3(CLBLM_L_X10Y107_SLICE_X12Y107_DO6),
.I4(CLBLM_L_X8Y108_SLICE_X11Y108_AQ),
.I5(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.O5(CLBLM_R_X11Y107_SLICE_X15Y107_CO5),
.O6(CLBLM_R_X11Y107_SLICE_X15Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0ff000ff0f30003)
  ) CLBLM_R_X11Y107_SLICE_X15Y107_BLUT (
.I0(1'b1),
.I1(RIOB33_X105Y141_IOB_X1Y142_I),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X11Y109_SLICE_X15Y109_BO6),
.I4(CLBLM_L_X10Y105_SLICE_X12Y105_BQ),
.I5(CLBLM_L_X8Y119_SLICE_X10Y119_AQ),
.O5(CLBLM_R_X11Y107_SLICE_X15Y107_BO5),
.O6(CLBLM_R_X11Y107_SLICE_X15Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f05555f0f01111)
  ) CLBLM_R_X11Y107_SLICE_X15Y107_ALUT (
.I0(CLBLM_R_X11Y107_SLICE_X15Y107_DO6),
.I1(RIOB33_X105Y141_IOB_X1Y142_I),
.I2(CLBLM_L_X8Y114_SLICE_X11Y114_B5Q),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y119_SLICE_X10Y119_AQ),
.O5(CLBLM_R_X11Y107_SLICE_X15Y107_AO5),
.O6(CLBLM_R_X11Y107_SLICE_X15Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y108_SLICE_X14Y108_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y108_SLICE_X14Y108_AO6),
.Q(CLBLM_R_X11Y108_SLICE_X14Y108_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000abab5454ffff)
  ) CLBLM_R_X11Y108_SLICE_X14Y108_DLUT (
.I0(CLBLM_R_X5Y115_SLICE_X7Y115_DO6),
.I1(CLBLM_R_X3Y110_SLICE_X2Y110_BO6),
.I2(CLBLL_L_X4Y107_SLICE_X5Y107_BO6),
.I3(1'b1),
.I4(CLBLM_R_X13Y117_SLICE_X18Y117_AQ),
.I5(CLBLM_L_X10Y108_SLICE_X12Y108_AO6),
.O5(CLBLM_R_X11Y108_SLICE_X14Y108_DO5),
.O6(CLBLM_R_X11Y108_SLICE_X14Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333cccc27728dd8)
  ) CLBLM_R_X11Y108_SLICE_X14Y108_CLUT (
.I0(CLBLM_R_X5Y115_SLICE_X7Y115_DO6),
.I1(CLBLM_R_X13Y112_SLICE_X18Y112_A5Q),
.I2(CLBLM_R_X11Y108_SLICE_X15Y108_BO6),
.I3(CLBLM_R_X11Y107_SLICE_X14Y107_AO5),
.I4(CLBLM_L_X8Y112_SLICE_X10Y112_AQ),
.I5(CLBLM_R_X3Y107_SLICE_X3Y107_CO6),
.O5(CLBLM_R_X11Y108_SLICE_X14Y108_CO5),
.O6(CLBLM_R_X11Y108_SLICE_X14Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h9669699669969669)
  ) CLBLM_R_X11Y108_SLICE_X14Y108_BLUT (
.I0(CLBLM_R_X11Y108_SLICE_X14Y108_DO6),
.I1(CLBLM_L_X10Y109_SLICE_X13Y109_DO6),
.I2(CLBLM_R_X11Y108_SLICE_X15Y108_CO6),
.I3(CLBLM_R_X11Y107_SLICE_X14Y107_DO6),
.I4(CLBLM_L_X10Y108_SLICE_X13Y108_DO6),
.I5(CLBLM_R_X11Y108_SLICE_X14Y108_CO6),
.O5(CLBLM_R_X11Y108_SLICE_X14Y108_BO5),
.O6(CLBLM_R_X11Y108_SLICE_X14Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haafaeeee00504444)
  ) CLBLM_R_X11Y108_SLICE_X14Y108_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X12Y108_SLICE_X17Y108_AQ),
.I2(CLBLM_R_X11Y108_SLICE_X14Y108_AQ),
.I3(CLBLM_L_X12Y105_SLICE_X16Y105_BO6),
.I4(CLBLM_L_X12Y105_SLICE_X16Y105_CO5),
.I5(CLBLM_L_X8Y116_SLICE_X10Y116_BQ),
.O5(CLBLM_R_X11Y108_SLICE_X14Y108_AO5),
.O6(CLBLM_R_X11Y108_SLICE_X14Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y108_SLICE_X15Y108_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y106_SLICE_X15Y106_BO6),
.Q(CLBLM_R_X11Y108_SLICE_X15Y108_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000333301003233)
  ) CLBLM_R_X11Y108_SLICE_X15Y108_DLUT (
.I0(CLBLM_R_X11Y105_SLICE_X14Y105_CQ),
.I1(CLBLM_L_X12Y109_SLICE_X16Y109_DQ),
.I2(CLBLM_R_X11Y105_SLICE_X14Y105_C5Q),
.I3(CLBLM_L_X10Y105_SLICE_X12Y105_AQ),
.I4(CLBLM_L_X12Y113_SLICE_X17Y113_DO6),
.I5(CLBLM_L_X10Y106_SLICE_X12Y106_AQ),
.O5(CLBLM_R_X11Y108_SLICE_X15Y108_DO5),
.O6(CLBLM_R_X11Y108_SLICE_X15Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h33cc33cc33cc5a5a)
  ) CLBLM_R_X11Y108_SLICE_X15Y108_CLUT (
.I0(CLBLM_R_X11Y108_SLICE_X15Y108_AO6),
.I1(CLBLM_R_X11Y111_SLICE_X15Y111_CQ),
.I2(CLBLM_R_X11Y109_SLICE_X15Y109_AO5),
.I3(CLBLM_R_X11Y108_SLICE_X15Y108_AQ),
.I4(CLBLM_R_X5Y115_SLICE_X7Y115_DO6),
.I5(CLBLM_R_X3Y107_SLICE_X3Y107_CO6),
.O5(CLBLM_R_X11Y108_SLICE_X15Y108_CO5),
.O6(CLBLM_R_X11Y108_SLICE_X15Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00f708fcfcffff)
  ) CLBLM_R_X11Y108_SLICE_X15Y108_BLUT (
.I0(CLBLM_L_X10Y105_SLICE_X12Y105_AQ),
.I1(CLBLM_L_X10Y106_SLICE_X12Y106_AQ),
.I2(CLBLM_R_X11Y105_SLICE_X14Y105_C5Q),
.I3(CLBLM_L_X10Y110_SLICE_X12Y110_AQ),
.I4(CLBLM_R_X11Y105_SLICE_X14Y105_CQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y108_SLICE_X15Y108_BO5),
.O6(CLBLM_R_X11Y108_SLICE_X15Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hefff1000ff55ff55)
  ) CLBLM_R_X11Y108_SLICE_X15Y108_ALUT (
.I0(CLBLM_L_X10Y105_SLICE_X12Y105_AQ),
.I1(CLBLM_L_X10Y106_SLICE_X12Y106_AQ),
.I2(CLBLM_R_X11Y105_SLICE_X14Y105_C5Q),
.I3(CLBLM_R_X11Y105_SLICE_X14Y105_CQ),
.I4(CLBLM_L_X12Y110_SLICE_X17Y110_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y108_SLICE_X15Y108_AO5),
.O6(CLBLM_R_X11Y108_SLICE_X15Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y109_SLICE_X14Y109_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y109_SLICE_X14Y109_AO6),
.Q(CLBLM_R_X11Y109_SLICE_X14Y109_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y109_SLICE_X14Y109_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y109_SLICE_X14Y109_BO6),
.Q(CLBLM_R_X11Y109_SLICE_X14Y109_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0011331100213321)
  ) CLBLM_R_X11Y109_SLICE_X14Y109_DLUT (
.I0(CLBLM_L_X8Y115_SLICE_X10Y115_AQ),
.I1(CLBLM_R_X11Y109_SLICE_X14Y109_AQ),
.I2(CLBLM_L_X10Y105_SLICE_X12Y105_AQ),
.I3(CLBLM_R_X5Y115_SLICE_X7Y115_CO6),
.I4(CLBLM_R_X13Y117_SLICE_X18Y117_AQ),
.I5(CLBLM_R_X11Y108_SLICE_X15Y108_BO5),
.O5(CLBLM_R_X11Y109_SLICE_X14Y109_DO5),
.O6(CLBLM_R_X11Y109_SLICE_X14Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0001050450515554)
  ) CLBLM_R_X11Y109_SLICE_X14Y109_CLUT (
.I0(CLBLM_R_X11Y109_SLICE_X14Y109_BQ),
.I1(CLBLM_L_X10Y105_SLICE_X12Y105_AQ),
.I2(CLBLM_R_X5Y115_SLICE_X7Y115_CO6),
.I3(CLBLM_R_X11Y108_SLICE_X15Y108_BO5),
.I4(CLBLM_L_X10Y115_SLICE_X13Y115_BQ),
.I5(CLBLM_R_X11Y111_SLICE_X15Y111_C5Q),
.O5(CLBLM_R_X11Y109_SLICE_X14Y109_CO5),
.O6(CLBLM_R_X11Y109_SLICE_X14Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000faff5055)
  ) CLBLM_R_X11Y109_SLICE_X14Y109_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(1'b1),
.I2(CLBLM_L_X8Y119_SLICE_X10Y119_AQ),
.I3(RIOB33_X105Y141_IOB_X1Y142_I),
.I4(CLBLM_L_X10Y109_SLICE_X12Y109_BQ),
.I5(CLBLM_R_X11Y109_SLICE_X14Y109_CO6),
.O5(CLBLM_R_X11Y109_SLICE_X14Y109_BO5),
.O6(CLBLM_R_X11Y109_SLICE_X14Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff005050ff005555)
  ) CLBLM_R_X11Y109_SLICE_X14Y109_ALUT (
.I0(CLBLM_R_X11Y109_SLICE_X14Y109_DO6),
.I1(1'b1),
.I2(CLBLM_L_X8Y119_SLICE_X10Y119_AQ),
.I3(CLBLM_R_X7Y108_SLICE_X8Y108_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y141_IOB_X1Y142_I),
.O5(CLBLM_R_X11Y109_SLICE_X14Y109_AO5),
.O6(CLBLM_R_X11Y109_SLICE_X14Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000001)
  ) CLBLM_R_X11Y109_SLICE_X15Y109_DLUT (
.I0(CLBLM_R_X11Y113_SLICE_X15Y113_AQ),
.I1(CLBLM_L_X10Y110_SLICE_X12Y110_AQ),
.I2(CLBLM_R_X11Y110_SLICE_X14Y110_CQ),
.I3(CLBLM_L_X8Y109_SLICE_X11Y109_CQ),
.I4(CLBLM_L_X12Y110_SLICE_X17Y110_AQ),
.I5(CLBLM_R_X7Y110_SLICE_X8Y110_CQ),
.O5(CLBLM_R_X11Y109_SLICE_X15Y109_DO5),
.O6(CLBLM_R_X11Y109_SLICE_X15Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaafaaafaaafaabe)
  ) CLBLM_R_X11Y109_SLICE_X15Y109_CLUT (
.I0(CLBLM_R_X5Y115_SLICE_X7Y115_CO6),
.I1(CLBLM_R_X11Y105_SLICE_X14Y105_C5Q),
.I2(CLBLM_L_X12Y113_SLICE_X17Y113_DO6),
.I3(CLBLM_L_X12Y109_SLICE_X16Y109_DQ),
.I4(CLBLM_L_X10Y106_SLICE_X12Y106_AQ),
.I5(CLBLM_R_X11Y108_SLICE_X15Y108_AO5),
.O5(CLBLM_R_X11Y109_SLICE_X15Y109_CO5),
.O6(CLBLM_R_X11Y109_SLICE_X15Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0011004100bb00eb)
  ) CLBLM_R_X11Y109_SLICE_X15Y109_BLUT (
.I0(CLBLM_R_X5Y115_SLICE_X7Y115_CO6),
.I1(CLBLM_R_X11Y113_SLICE_X15Y113_AQ),
.I2(CLBLM_R_X11Y105_SLICE_X14Y105_CQ),
.I3(CLBLM_R_X11Y107_SLICE_X15Y107_BQ),
.I4(CLBLM_R_X11Y109_SLICE_X15Y109_AO6),
.I5(CLBLM_R_X11Y111_SLICE_X15Y111_CQ),
.O5(CLBLM_R_X11Y109_SLICE_X15Y109_BO5),
.O6(CLBLM_R_X11Y109_SLICE_X15Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafafffffb04ff00)
  ) CLBLM_R_X11Y109_SLICE_X15Y109_ALUT (
.I0(CLBLM_L_X10Y105_SLICE_X12Y105_AQ),
.I1(CLBLM_R_X11Y105_SLICE_X14Y105_CQ),
.I2(CLBLM_R_X11Y105_SLICE_X14Y105_C5Q),
.I3(CLBLM_R_X11Y113_SLICE_X15Y113_AQ),
.I4(CLBLM_L_X10Y106_SLICE_X12Y106_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y109_SLICE_X15Y109_AO5),
.O6(CLBLM_R_X11Y109_SLICE_X15Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y110_SLICE_X14Y110_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y110_SLICE_X14Y110_BO6),
.Q(CLBLM_R_X11Y110_SLICE_X14Y110_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y110_SLICE_X14Y110_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y110_SLICE_X14Y110_DO5),
.Q(CLBLM_R_X11Y110_SLICE_X14Y110_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y110_SLICE_X14Y110_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y110_SLICE_X14Y110_AO6),
.Q(CLBLM_R_X11Y110_SLICE_X14Y110_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y110_SLICE_X14Y110_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y110_SLICE_X14Y110_CO6),
.Q(CLBLM_R_X11Y110_SLICE_X14Y110_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y110_SLICE_X14Y110_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y110_SLICE_X14Y110_DO6),
.Q(CLBLM_R_X11Y110_SLICE_X14Y110_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5a0a0ee44ee44)
  ) CLBLM_R_X11Y110_SLICE_X14Y110_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X11Y112_SLICE_X14Y112_C5Q),
.I2(CLBLM_R_X11Y105_SLICE_X14Y105_AQ),
.I3(CLBLM_R_X11Y109_SLICE_X14Y109_AQ),
.I4(RIOB33_X105Y103_IOB_X1Y104_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y110_SLICE_X14Y110_DO5),
.O6(CLBLM_R_X11Y110_SLICE_X14Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00fcfc0000)
  ) CLBLM_R_X11Y110_SLICE_X14Y110_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y110_SLICE_X14Y110_CQ),
.I2(CLBLM_L_X8Y115_SLICE_X11Y115_BQ),
.I3(CLBLM_R_X13Y110_SLICE_X19Y110_BQ),
.I4(CLBLM_R_X7Y115_SLICE_X9Y115_DO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y110_SLICE_X14Y110_CO5),
.O6(CLBLM_R_X11Y110_SLICE_X14Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccf0a0f0a0f0a0)
  ) CLBLM_R_X11Y110_SLICE_X14Y110_BLUT (
.I0(CLBLM_R_X13Y112_SLICE_X18Y112_CQ),
.I1(CLBLM_R_X11Y107_SLICE_X15Y107_BQ),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLM_R_X13Y110_SLICE_X19Y110_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y110_SLICE_X14Y110_BO5),
.O6(CLBLM_R_X11Y110_SLICE_X14Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffaeeea55504440)
  ) CLBLM_R_X11Y110_SLICE_X14Y110_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_R_X11Y110_SLICE_X14Y110_AQ),
.I3(CLBLM_R_X13Y110_SLICE_X18Y110_AQ),
.I4(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.I5(CLBLM_L_X10Y110_SLICE_X12Y110_B5Q),
.O5(CLBLM_R_X11Y110_SLICE_X14Y110_AO5),
.O6(CLBLM_R_X11Y110_SLICE_X14Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y110_SLICE_X15Y110_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y110_SLICE_X16Y110_BO6),
.Q(CLBLM_R_X11Y110_SLICE_X15Y110_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y110_SLICE_X15Y110_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y110_SLICE_X15Y110_AO6),
.Q(CLBLM_R_X11Y110_SLICE_X15Y110_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y110_SLICE_X15Y110_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y110_SLICE_X15Y110_BO6),
.Q(CLBLM_R_X11Y110_SLICE_X15Y110_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y110_SLICE_X15Y110_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y110_SLICE_X15Y110_CO6),
.Q(CLBLM_R_X11Y110_SLICE_X15Y110_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5faff5fa5faff5fa)
  ) CLBLM_R_X11Y110_SLICE_X15Y110_DLUT (
.I0(CLBLM_L_X8Y109_SLICE_X10Y109_C5Q),
.I1(1'b1),
.I2(CLBLM_L_X10Y114_SLICE_X13Y114_CQ),
.I3(CLBLM_L_X10Y109_SLICE_X12Y109_AQ),
.I4(CLBLM_R_X11Y108_SLICE_X15Y108_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y110_SLICE_X15Y110_DO5),
.O6(CLBLM_R_X11Y110_SLICE_X15Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000000fc00fc)
  ) CLBLM_R_X11Y110_SLICE_X15Y110_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y110_SLICE_X15Y110_CQ),
.I2(CLBLM_L_X10Y114_SLICE_X13Y114_CQ),
.I3(CLBLM_R_X5Y115_SLICE_X7Y115_CO6),
.I4(CLBLM_R_X11Y110_SLICE_X15Y110_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y110_SLICE_X15Y110_CO5),
.O6(CLBLM_R_X11Y110_SLICE_X15Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f6f0f600060006)
  ) CLBLM_R_X11Y110_SLICE_X15Y110_BLUT (
.I0(CLBLM_L_X12Y110_SLICE_X16Y110_AO5),
.I1(CLBLM_R_X11Y115_SLICE_X15Y115_AQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(1'b1),
.I5(CLBLM_L_X10Y111_SLICE_X12Y111_A5Q),
.O5(CLBLM_R_X11Y110_SLICE_X15Y110_BO5),
.O6(CLBLM_R_X11Y110_SLICE_X15Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff14ff0000140000)
  ) CLBLM_R_X11Y110_SLICE_X15Y110_ALUT (
.I0(CLBLM_R_X7Y115_SLICE_X8Y115_DQ),
.I1(CLBLM_L_X12Y110_SLICE_X16Y110_CO6),
.I2(CLBLM_R_X11Y110_SLICE_X15Y110_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_L_X8Y114_SLICE_X10Y114_CQ),
.O5(CLBLM_R_X11Y110_SLICE_X15Y110_AO5),
.O6(CLBLM_R_X11Y110_SLICE_X15Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffbbffbb)
  ) CLBLM_R_X11Y111_SLICE_X14Y111_DLUT (
.I0(CLBLM_R_X11Y113_SLICE_X15Y113_AQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(1'b1),
.I3(CLBLM_R_X7Y118_SLICE_X8Y118_CQ),
.I4(1'b1),
.I5(CLBLM_L_X8Y107_SLICE_X11Y107_B5Q),
.O5(CLBLM_R_X11Y111_SLICE_X14Y111_DO5),
.O6(CLBLM_R_X11Y111_SLICE_X14Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffeffffffffff)
  ) CLBLM_R_X11Y111_SLICE_X14Y111_CLUT (
.I0(CLBLM_L_X10Y106_SLICE_X13Y106_DO6),
.I1(CLBLM_L_X10Y110_SLICE_X12Y110_DO6),
.I2(CLBLM_L_X12Y113_SLICE_X17Y113_BQ),
.I3(RIOB33_X105Y143_IOB_X1Y143_I),
.I4(CLBLM_R_X11Y111_SLICE_X14Y111_DO6),
.I5(CLBLM_L_X8Y107_SLICE_X11Y107_BQ),
.O5(CLBLM_R_X11Y111_SLICE_X14Y111_CO5),
.O6(CLBLM_R_X11Y111_SLICE_X14Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffff0f0fcf8)
  ) CLBLM_R_X11Y111_SLICE_X14Y111_BLUT (
.I0(CLBLL_L_X4Y107_SLICE_X5Y107_BO6),
.I1(CLBLM_R_X7Y110_SLICE_X8Y110_CQ),
.I2(CLBLM_R_X11Y115_SLICE_X14Y115_CO6),
.I3(CLBLM_R_X3Y110_SLICE_X2Y110_BO6),
.I4(CLBLM_R_X5Y115_SLICE_X7Y115_DO6),
.I5(CLBLM_R_X11Y111_SLICE_X14Y111_CO6),
.O5(CLBLM_R_X11Y111_SLICE_X14Y111_BO5),
.O6(CLBLM_R_X11Y111_SLICE_X14Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000111455551114)
  ) CLBLM_R_X11Y111_SLICE_X14Y111_ALUT (
.I0(CLBLM_R_X11Y114_SLICE_X14Y114_BQ),
.I1(CLBLM_R_X7Y110_SLICE_X8Y110_CQ),
.I2(CLBLM_R_X11Y109_SLICE_X15Y109_AO6),
.I3(CLBLM_R_X11Y105_SLICE_X14Y105_CQ),
.I4(CLBLM_R_X5Y115_SLICE_X7Y115_CO6),
.I5(CLBLM_R_X11Y115_SLICE_X15Y115_BQ),
.O5(CLBLM_R_X11Y111_SLICE_X14Y111_AO5),
.O6(CLBLM_R_X11Y111_SLICE_X14Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y111_SLICE_X15Y111_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y111_SLICE_X15Y111_CO5),
.Q(CLBLM_R_X11Y111_SLICE_X15Y111_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y111_SLICE_X15Y111_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y111_SLICE_X15Y111_AO6),
.Q(CLBLM_R_X11Y111_SLICE_X15Y111_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y111_SLICE_X15Y111_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y111_SLICE_X15Y111_BO6),
.Q(CLBLM_R_X11Y111_SLICE_X15Y111_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y111_SLICE_X15Y111_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y111_SLICE_X15Y111_CO6),
.Q(CLBLM_R_X11Y111_SLICE_X15Y111_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hdfefdfeffdfefdfe)
  ) CLBLM_R_X11Y111_SLICE_X15Y111_DLUT (
.I0(CLBLM_R_X11Y110_SLICE_X15Y110_CQ),
.I1(CLBLM_R_X11Y110_SLICE_X15Y110_DO6),
.I2(CLBLM_R_X11Y114_SLICE_X14Y114_DQ),
.I3(CLBLM_R_X7Y107_SLICE_X9Y107_C5Q),
.I4(1'b1),
.I5(CLBLM_R_X11Y115_SLICE_X15Y115_BQ),
.O5(CLBLM_R_X11Y111_SLICE_X15Y111_DO5),
.O6(CLBLM_R_X11Y111_SLICE_X15Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaa00f0ccf0cc)
  ) CLBLM_R_X11Y111_SLICE_X15Y111_CLUT (
.I0(CLBLM_L_X10Y118_SLICE_X12Y118_AQ),
.I1(CLBLM_R_X11Y110_SLICE_X14Y110_A5Q),
.I2(CLBLM_R_X5Y111_SLICE_X6Y111_BQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X11Y110_SLICE_X15Y110_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X11Y111_SLICE_X15Y111_CO5),
.O6(CLBLM_R_X11Y111_SLICE_X15Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0ccf0ccf000f000)
  ) CLBLM_R_X11Y111_SLICE_X15Y111_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y112_SLICE_X15Y112_BQ),
.I2(CLBLM_R_X5Y106_SLICE_X6Y106_BQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X11Y111_SLICE_X15Y111_BO5),
.O6(CLBLM_R_X11Y111_SLICE_X15Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0e2e2e2e2)
  ) CLBLM_R_X11Y111_SLICE_X15Y111_ALUT (
.I0(CLBLM_R_X11Y112_SLICE_X14Y112_BQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y106_SLICE_X12Y106_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X11Y111_SLICE_X15Y111_AO5),
.O6(CLBLM_R_X11Y111_SLICE_X15Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y112_SLICE_X14Y112_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y112_SLICE_X14Y112_BO5),
.Q(CLBLM_R_X11Y112_SLICE_X14Y112_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y112_SLICE_X14Y112_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y112_SLICE_X14Y112_CO5),
.Q(CLBLM_R_X11Y112_SLICE_X14Y112_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y112_SLICE_X14Y112_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y112_SLICE_X14Y112_BO6),
.Q(CLBLM_R_X11Y112_SLICE_X14Y112_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y112_SLICE_X14Y112_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y112_SLICE_X14Y112_CO6),
.Q(CLBLM_R_X11Y112_SLICE_X14Y112_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffafa)
  ) CLBLM_R_X11Y112_SLICE_X14Y112_DLUT (
.I0(CLBLM_L_X8Y111_SLICE_X11Y111_CQ),
.I1(1'b1),
.I2(CLBLM_L_X8Y114_SLICE_X10Y114_DQ),
.I3(1'b1),
.I4(CLBLM_R_X11Y112_SLICE_X14Y112_B5Q),
.I5(CLBLM_R_X13Y110_SLICE_X18Y110_BQ),
.O5(CLBLM_R_X11Y112_SLICE_X14Y112_DO5),
.O6(CLBLM_R_X11Y112_SLICE_X14Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfc0c0c0fafa0a0a)
  ) CLBLM_R_X11Y112_SLICE_X14Y112_CLUT (
.I0(CLBLM_L_X10Y117_SLICE_X12Y117_AQ),
.I1(CLBLM_R_X11Y113_SLICE_X15Y113_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X11Y112_SLICE_X14Y112_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X11Y112_SLICE_X14Y112_CO5),
.O6(CLBLM_R_X11Y112_SLICE_X14Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hbaba1010b1a0b1a0)
  ) CLBLM_R_X11Y112_SLICE_X14Y112_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_L_X12Y111_SLICE_X16Y111_DQ),
.I3(CLBLM_R_X5Y109_SLICE_X6Y109_DQ),
.I4(CLBLM_L_X10Y107_SLICE_X13Y107_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y112_SLICE_X14Y112_BO5),
.O6(CLBLM_R_X11Y112_SLICE_X14Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'he4e4e4a0cccccc00)
  ) CLBLM_R_X11Y112_SLICE_X14Y112_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y121_IOB_X1Y121_I),
.I2(CLBLM_L_X10Y111_SLICE_X12Y111_C5Q),
.I3(CLBLM_R_X11Y112_SLICE_X14Y112_CQ),
.I4(CLBLM_R_X11Y112_SLICE_X15Y112_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y112_SLICE_X14Y112_AO5),
.O6(CLBLM_R_X11Y112_SLICE_X14Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y112_SLICE_X15Y112_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y112_SLICE_X15Y112_AO6),
.Q(CLBLM_R_X11Y112_SLICE_X15Y112_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y112_SLICE_X15Y112_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y112_SLICE_X15Y112_BO6),
.Q(CLBLM_R_X11Y112_SLICE_X15Y112_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000824100008241)
  ) CLBLM_R_X11Y112_SLICE_X15Y112_DLUT (
.I0(CLBLM_R_X11Y111_SLICE_X15Y111_C5Q),
.I1(CLBLM_R_X13Y117_SLICE_X18Y117_AQ),
.I2(CLBLM_R_X11Y113_SLICE_X15Y113_DQ),
.I3(CLBLM_R_X11Y113_SLICE_X15Y113_CQ),
.I4(CLBLM_R_X11Y114_SLICE_X15Y114_DO6),
.I5(1'b1),
.O5(CLBLM_R_X11Y112_SLICE_X15Y112_DO5),
.O6(CLBLM_R_X11Y112_SLICE_X15Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000080208020000)
  ) CLBLM_R_X11Y112_SLICE_X15Y112_CLUT (
.I0(CLBLM_R_X11Y112_SLICE_X15Y112_DO6),
.I1(CLBLM_L_X10Y114_SLICE_X12Y114_CQ),
.I2(CLBLM_R_X11Y111_SLICE_X15Y111_DO6),
.I3(CLBLM_R_X13Y112_SLICE_X18Y112_A5Q),
.I4(CLBLM_L_X12Y109_SLICE_X16Y109_DQ),
.I5(CLBLM_R_X11Y114_SLICE_X15Y114_BO6),
.O5(CLBLM_R_X11Y112_SLICE_X15Y112_CO5),
.O6(CLBLM_R_X11Y112_SLICE_X15Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff003333ff000000)
  ) CLBLM_R_X11Y112_SLICE_X15Y112_BLUT (
.I0(1'b1),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(1'b1),
.I3(CLBLM_L_X12Y113_SLICE_X17Y113_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X13Y112_SLICE_X18Y112_CQ),
.O5(CLBLM_R_X11Y112_SLICE_X15Y112_BO5),
.O6(CLBLM_R_X11Y112_SLICE_X15Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffa50ea40)
  ) CLBLM_R_X11Y112_SLICE_X15Y112_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_R_X11Y112_SLICE_X15Y112_AQ),
.I3(CLBLL_L_X4Y112_SLICE_X4Y112_AQ),
.I4(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.I5(CLBLM_R_X7Y112_SLICE_X9Y112_CO6),
.O5(CLBLM_R_X11Y112_SLICE_X15Y112_AO5),
.O6(CLBLM_R_X11Y112_SLICE_X15Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y113_SLICE_X14Y113_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y113_SLICE_X14Y113_AO6),
.Q(CLBLM_R_X11Y113_SLICE_X14Y113_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y113_SLICE_X14Y113_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y113_SLICE_X14Y113_BO6),
.Q(CLBLM_R_X11Y113_SLICE_X14Y113_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y113_SLICE_X14Y113_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y113_SLICE_X14Y113_CO6),
.Q(CLBLM_R_X11Y113_SLICE_X14Y113_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y113_SLICE_X14Y113_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y113_SLICE_X14Y113_DO6),
.Q(CLBLM_R_X11Y113_SLICE_X14Y113_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf1f00100f1f00100)
  ) CLBLM_R_X11Y113_SLICE_X14Y113_DLUT (
.I0(CLBLM_L_X10Y112_SLICE_X13Y112_AO6),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X13Y112_SLICE_X18Y112_BQ),
.I4(CLBLM_R_X11Y118_SLICE_X15Y118_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X11Y113_SLICE_X14Y113_DO5),
.O6(CLBLM_R_X11Y113_SLICE_X14Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0050cccc0000)
  ) CLBLM_R_X11Y113_SLICE_X14Y113_CLUT (
.I0(CLBLM_L_X10Y112_SLICE_X13Y112_AO6),
.I1(CLBLM_L_X10Y113_SLICE_X13Y113_BQ),
.I2(CLBLM_R_X11Y113_SLICE_X14Y113_BQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X13Y112_SLICE_X18Y112_BQ),
.O5(CLBLM_R_X11Y113_SLICE_X14Y113_CO5),
.O6(CLBLM_R_X11Y113_SLICE_X14Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa00fcaaaa0000)
  ) CLBLM_R_X11Y113_SLICE_X14Y113_BLUT (
.I0(CLBLM_L_X12Y113_SLICE_X17Y113_CQ),
.I1(CLBLM_R_X11Y113_SLICE_X14Y113_BQ),
.I2(CLBLM_R_X11Y113_SLICE_X14Y113_DQ),
.I3(CLBLM_R_X11Y113_SLICE_X14Y113_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X11Y113_SLICE_X14Y113_BO5),
.O6(CLBLM_R_X11Y113_SLICE_X14Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88dd888888d88888)
  ) CLBLM_R_X11Y113_SLICE_X14Y113_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X11Y113_SLICE_X14Y113_BQ),
.I2(CLBLM_R_X11Y113_SLICE_X14Y113_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.I5(CLBLM_R_X11Y107_SLICE_X15Y107_AQ),
.O5(CLBLM_R_X11Y113_SLICE_X14Y113_AO5),
.O6(CLBLM_R_X11Y113_SLICE_X14Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y113_SLICE_X15Y113_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y113_SLICE_X15Y113_AO6),
.Q(CLBLM_R_X11Y113_SLICE_X15Y113_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y113_SLICE_X15Y113_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y113_SLICE_X15Y113_BO6),
.Q(CLBLM_R_X11Y113_SLICE_X15Y113_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y113_SLICE_X15Y113_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y113_SLICE_X15Y113_CO6),
.Q(CLBLM_R_X11Y113_SLICE_X15Y113_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y113_SLICE_X15Y113_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y113_SLICE_X15Y113_DO6),
.Q(CLBLM_R_X11Y113_SLICE_X15Y113_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfeaa5400feaa5400)
  ) CLBLM_R_X11Y113_SLICE_X15Y113_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X11Y113_SLICE_X15Y113_CQ),
.I2(CLBLM_R_X11Y113_SLICE_X15Y113_DQ),
.I3(CLBLM_R_X7Y115_SLICE_X9Y115_DO6),
.I4(CLBLM_R_X11Y107_SLICE_X15Y107_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y113_SLICE_X15Y113_DO5),
.O6(CLBLM_R_X11Y113_SLICE_X15Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haca0afa0aca0afa0)
  ) CLBLM_R_X11Y113_SLICE_X15Y113_CLUT (
.I0(CLBLM_R_X7Y115_SLICE_X9Y115_AQ),
.I1(CLBLM_R_X11Y113_SLICE_X15Y113_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y115_SLICE_X9Y115_DO6),
.I4(CLBLM_R_X11Y114_SLICE_X15Y114_BO6),
.I5(1'b1),
.O5(CLBLM_R_X11Y113_SLICE_X15Y113_CO5),
.O6(CLBLM_R_X11Y113_SLICE_X15Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0f5f5a0a0e4e4)
  ) CLBLM_R_X11Y113_SLICE_X15Y113_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X11Y113_SLICE_X15Y113_BQ),
.I2(CLBLM_R_X7Y113_SLICE_X8Y113_CQ),
.I3(1'b1),
.I4(CLBLM_R_X5Y115_SLICE_X7Y115_CO6),
.I5(CLBLM_L_X10Y114_SLICE_X12Y114_DQ),
.O5(CLBLM_R_X11Y113_SLICE_X15Y113_BO5),
.O6(CLBLM_R_X11Y113_SLICE_X15Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hddddd8d888888888)
  ) CLBLM_R_X11Y113_SLICE_X15Y113_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X11Y113_SLICE_X15Y113_BQ),
.I2(CLBLM_R_X11Y113_SLICE_X15Y113_AQ),
.I3(1'b1),
.I4(CLBLM_L_X10Y110_SLICE_X12Y110_AQ),
.I5(CLBLM_R_X7Y115_SLICE_X9Y115_DO6),
.O5(CLBLM_R_X11Y113_SLICE_X15Y113_AO5),
.O6(CLBLM_R_X11Y113_SLICE_X15Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y114_SLICE_X14Y114_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y114_SLICE_X14Y114_AO6),
.Q(CLBLM_R_X11Y114_SLICE_X14Y114_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y114_SLICE_X14Y114_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y114_SLICE_X14Y114_BO6),
.Q(CLBLM_R_X11Y114_SLICE_X14Y114_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y114_SLICE_X14Y114_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y114_SLICE_X14Y114_CO6),
.Q(CLBLM_R_X11Y114_SLICE_X14Y114_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y114_SLICE_X14Y114_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y114_SLICE_X14Y114_DO6),
.Q(CLBLM_R_X11Y114_SLICE_X14Y114_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000fffa00fa)
  ) CLBLM_R_X11Y114_SLICE_X14Y114_DLUT (
.I0(CLBLM_R_X11Y110_SLICE_X15Y110_CQ),
.I1(1'b1),
.I2(CLBLM_R_X11Y114_SLICE_X14Y114_DQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I5(CLBLM_R_X5Y115_SLICE_X7Y115_CO6),
.O5(CLBLM_R_X11Y114_SLICE_X14Y114_DO5),
.O6(CLBLM_R_X11Y114_SLICE_X14Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00aa0faaf0)
  ) CLBLM_R_X11Y114_SLICE_X14Y114_CLUT (
.I0(CLBLM_R_X11Y112_SLICE_X15Y112_BQ),
.I1(1'b1),
.I2(CLBLM_R_X11Y115_SLICE_X14Y115_BO5),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X11Y114_SLICE_X14Y114_CO5),
.O6(CLBLM_R_X11Y114_SLICE_X14Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcecfcecf02030203)
  ) CLBLM_R_X11Y114_SLICE_X14Y114_BLUT (
.I0(CLBLM_L_X8Y119_SLICE_X10Y119_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X11Y111_SLICE_X14Y111_AO6),
.I3(RIOB33_X105Y141_IOB_X1Y142_I),
.I4(1'b1),
.I5(CLBLM_R_X7Y115_SLICE_X9Y115_BQ),
.O5(CLBLM_R_X11Y114_SLICE_X14Y114_BO5),
.O6(CLBLM_R_X11Y114_SLICE_X14Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbb888b8bbb888b8)
  ) CLBLM_R_X11Y114_SLICE_X14Y114_ALUT (
.I0(CLBLM_L_X12Y114_SLICE_X16Y114_CQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X11Y114_SLICE_X14Y114_AQ),
.I3(CLBLL_L_X4Y116_SLICE_X4Y116_BO6),
.I4(CLBLM_L_X10Y115_SLICE_X12Y115_BQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y114_SLICE_X14Y114_AO5),
.O6(CLBLM_R_X11Y114_SLICE_X14Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h66ff66ffff66ff66)
  ) CLBLM_R_X11Y114_SLICE_X15Y114_DLUT (
.I0(CLBLM_L_X12Y113_SLICE_X16Y113_BQ),
.I1(CLBLM_L_X8Y112_SLICE_X10Y112_AQ),
.I2(1'b1),
.I3(CLBLM_L_X8Y114_SLICE_X10Y114_BQ),
.I4(1'b1),
.I5(CLBLM_R_X11Y111_SLICE_X15Y111_CQ),
.O5(CLBLM_R_X11Y114_SLICE_X15Y114_DO5),
.O6(CLBLM_R_X11Y114_SLICE_X15Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000000000000a)
  ) CLBLM_R_X11Y114_SLICE_X15Y114_CLUT (
.I0(CLBLM_R_X11Y114_SLICE_X15Y114_AO6),
.I1(1'b1),
.I2(CLBLM_L_X10Y114_SLICE_X12Y114_CQ),
.I3(CLBLM_L_X10Y114_SLICE_X12Y114_DQ),
.I4(CLBLM_R_X11Y115_SLICE_X15Y115_DO6),
.I5(CLBLM_L_X12Y114_SLICE_X16Y114_AQ),
.O5(CLBLM_R_X11Y114_SLICE_X15Y114_CO5),
.O6(CLBLM_R_X11Y114_SLICE_X15Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5f5050505f50505f)
  ) CLBLM_R_X11Y114_SLICE_X15Y114_BLUT (
.I0(CLBLM_L_X12Y109_SLICE_X16Y109_DQ),
.I1(1'b1),
.I2(CLBLM_R_X5Y111_SLICE_X6Y111_DO6),
.I3(CLBLM_R_X11Y115_SLICE_X15Y115_CQ),
.I4(CLBLM_L_X12Y114_SLICE_X16Y114_BQ),
.I5(CLBLM_R_X11Y114_SLICE_X15Y114_CO6),
.O5(CLBLM_R_X11Y114_SLICE_X15Y114_BO5),
.O6(CLBLM_R_X11Y114_SLICE_X15Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000001)
  ) CLBLM_R_X11Y114_SLICE_X15Y114_ALUT (
.I0(CLBLM_R_X11Y114_SLICE_X14Y114_DQ),
.I1(CLBLM_L_X10Y114_SLICE_X13Y114_CQ),
.I2(CLBLM_R_X11Y110_SLICE_X15Y110_CQ),
.I3(CLBLM_L_X12Y113_SLICE_X16Y113_BQ),
.I4(CLBLM_L_X8Y114_SLICE_X10Y114_BQ),
.I5(CLBLM_L_X10Y109_SLICE_X12Y109_AQ),
.O5(CLBLM_R_X11Y114_SLICE_X15Y114_AO5),
.O6(CLBLM_R_X11Y114_SLICE_X15Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y115_SLICE_X14Y115_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y77_IOB_X0Y77_I),
.D(CLBLM_R_X11Y115_SLICE_X15Y115_CQ),
.Q(CLBLM_R_X11Y115_SLICE_X14Y115_AQ),
.R(CLBLM_L_X12Y117_SLICE_X16Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y115_SLICE_X14Y115_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y77_IOB_X0Y77_I),
.D(CLBLM_R_X11Y110_SLICE_X14Y110_DQ),
.Q(CLBLM_R_X11Y115_SLICE_X14Y115_BQ),
.R(CLBLM_L_X12Y117_SLICE_X16Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y115_SLICE_X14Y115_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y115_SLICE_X14Y115_DO5),
.O6(CLBLM_R_X11Y115_SLICE_X14Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000fadb5f5f)
  ) CLBLM_R_X11Y115_SLICE_X14Y115_CLUT (
.I0(CLBLM_L_X10Y118_SLICE_X12Y118_AQ),
.I1(CLBLM_L_X10Y119_SLICE_X12Y119_AQ),
.I2(CLBLM_L_X10Y118_SLICE_X13Y118_AQ),
.I3(CLBLM_L_X8Y118_SLICE_X10Y118_AQ),
.I4(CLBLM_R_X7Y118_SLICE_X8Y118_CQ),
.I5(CLBLM_L_X10Y117_SLICE_X12Y117_DO6),
.O5(CLBLM_R_X11Y115_SLICE_X14Y115_CO5),
.O6(CLBLM_R_X11Y115_SLICE_X14Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0cc88cc88cc88)
  ) CLBLM_R_X11Y115_SLICE_X14Y115_BLUT (
.I0(CLBLM_R_X7Y115_SLICE_X8Y115_CQ),
.I1(RIOB33_X105Y121_IOB_X1Y121_I),
.I2(CLBLM_L_X10Y110_SLICE_X13Y110_BQ),
.I3(CLBLM_L_X10Y115_SLICE_X13Y115_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y115_SLICE_X14Y115_BO5),
.O6(CLBLM_R_X11Y115_SLICE_X14Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heeea4440ccc0ccc0)
  ) CLBLM_R_X11Y115_SLICE_X14Y115_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y121_IOB_X1Y121_I),
.I2(CLBLM_L_X10Y111_SLICE_X13Y111_C5Q),
.I3(CLBLM_R_X11Y116_SLICE_X15Y116_AQ),
.I4(CLBLM_L_X10Y110_SLICE_X12Y110_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y115_SLICE_X14Y115_AO5),
.O6(CLBLM_R_X11Y115_SLICE_X14Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y115_SLICE_X15Y115_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y115_SLICE_X15Y115_BO5),
.Q(CLBLM_R_X11Y115_SLICE_X15Y115_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y115_SLICE_X15Y115_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y115_SLICE_X15Y115_AO6),
.Q(CLBLM_R_X11Y115_SLICE_X15Y115_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y115_SLICE_X15Y115_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y115_SLICE_X15Y115_BO6),
.Q(CLBLM_R_X11Y115_SLICE_X15Y115_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y115_SLICE_X15Y115_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y115_SLICE_X15Y115_CO6),
.Q(CLBLM_R_X11Y115_SLICE_X15Y115_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffeeffffffee)
  ) CLBLM_R_X11Y115_SLICE_X15Y115_DLUT (
.I0(CLBLM_R_X11Y113_SLICE_X15Y113_BQ),
.I1(CLBLM_R_X11Y113_SLICE_X15Y113_CQ),
.I2(1'b1),
.I3(CLBLM_L_X10Y114_SLICE_X12Y114_AQ),
.I4(CLBLM_R_X11Y113_SLICE_X15Y113_DQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y115_SLICE_X15Y115_DO5),
.O6(CLBLM_R_X11Y115_SLICE_X15Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000ffee00ee)
  ) CLBLM_R_X11Y115_SLICE_X15Y115_CLUT (
.I0(CLBLM_R_X11Y113_SLICE_X15Y113_BQ),
.I1(CLBLM_R_X11Y115_SLICE_X15Y115_CQ),
.I2(1'b1),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y110_SLICE_X11Y110_AQ),
.I5(CLBLM_R_X5Y115_SLICE_X7Y115_CO6),
.O5(CLBLM_R_X11Y115_SLICE_X15Y115_CO5),
.O6(CLBLM_R_X11Y115_SLICE_X15Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ccccff00aaaa)
  ) CLBLM_R_X11Y115_SLICE_X15Y115_BLUT (
.I0(RIOB33_X105Y103_IOB_X1Y103_I),
.I1(CLBLM_L_X12Y112_SLICE_X17Y112_A5Q),
.I2(CLBLM_L_X10Y113_SLICE_X13Y113_AQ),
.I3(CLBLM_L_X10Y115_SLICE_X13Y115_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y115_SLICE_X15Y115_BO5),
.O6(CLBLM_R_X11Y115_SLICE_X15Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff006600000066)
  ) CLBLM_R_X11Y115_SLICE_X15Y115_ALUT (
.I0(CLBLM_R_X11Y115_SLICE_X14Y115_AO5),
.I1(CLBLM_L_X12Y110_SLICE_X17Y110_CQ),
.I2(1'b1),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X11Y113_SLICE_X14Y113_CQ),
.O5(CLBLM_R_X11Y115_SLICE_X15Y115_AO5),
.O6(CLBLM_R_X11Y115_SLICE_X15Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y116_SLICE_X14Y116_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y117_SLICE_X15Y117_BO6),
.Q(CLBLM_R_X11Y116_SLICE_X14Y116_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y116_SLICE_X14Y116_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y116_SLICE_X14Y116_AO6),
.Q(CLBLM_R_X11Y116_SLICE_X14Y116_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y116_SLICE_X14Y116_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y116_SLICE_X14Y116_BO6),
.Q(CLBLM_R_X11Y116_SLICE_X14Y116_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0101808001808080)
  ) CLBLM_R_X11Y116_SLICE_X14Y116_DLUT (
.I0(CLBLM_L_X10Y118_SLICE_X12Y118_AQ),
.I1(CLBLM_L_X10Y118_SLICE_X12Y118_BQ),
.I2(CLBLM_L_X10Y118_SLICE_X13Y118_AQ),
.I3(CLBLM_L_X8Y118_SLICE_X10Y118_AQ),
.I4(CLBLM_R_X7Y118_SLICE_X8Y118_CQ),
.I5(CLBLM_L_X10Y119_SLICE_X12Y119_AQ),
.O5(CLBLM_R_X11Y116_SLICE_X14Y116_DO5),
.O6(CLBLM_R_X11Y116_SLICE_X14Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd77dd77fd57dd77)
  ) CLBLM_R_X11Y116_SLICE_X14Y116_CLUT (
.I0(CLBLM_L_X10Y116_SLICE_X12Y116_DO5),
.I1(CLBLM_L_X10Y117_SLICE_X12Y117_DO6),
.I2(CLBLM_R_X11Y116_SLICE_X14Y116_AQ),
.I3(CLBLM_R_X11Y116_SLICE_X14Y116_BQ),
.I4(CLBLM_R_X11Y116_SLICE_X14Y116_DO6),
.I5(CLBLM_L_X8Y116_SLICE_X11Y116_CO6),
.O5(CLBLM_R_X11Y116_SLICE_X14Y116_CO5),
.O6(CLBLM_R_X11Y116_SLICE_X14Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcacacacacfcfcfcf)
  ) CLBLM_R_X11Y116_SLICE_X14Y116_BLUT (
.I0(CLBLM_L_X10Y118_SLICE_X13Y118_CO6),
.I1(CLBLM_R_X7Y108_SLICE_X9Y108_AQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X11Y116_SLICE_X14Y116_CO6),
.O5(CLBLM_R_X11Y116_SLICE_X14Y116_BO5),
.O6(CLBLM_R_X11Y116_SLICE_X14Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdc10dc10ff33cc00)
  ) CLBLM_R_X11Y116_SLICE_X14Y116_ALUT (
.I0(CLBLM_L_X10Y117_SLICE_X13Y117_AO5),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X11Y116_SLICE_X14Y116_AQ),
.I3(CLBLM_L_X12Y114_SLICE_X16Y114_BQ),
.I4(CLBLM_L_X8Y116_SLICE_X10Y116_BQ),
.I5(CLBLM_R_X7Y118_SLICE_X8Y118_DO6),
.O5(CLBLM_R_X11Y116_SLICE_X14Y116_AO5),
.O6(CLBLM_R_X11Y116_SLICE_X14Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y116_SLICE_X15Y116_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y116_SLICE_X15Y116_AO6),
.Q(CLBLM_R_X11Y116_SLICE_X15Y116_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y116_SLICE_X15Y116_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y116_SLICE_X15Y116_DO5),
.O6(CLBLM_R_X11Y116_SLICE_X15Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y116_SLICE_X15Y116_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y116_SLICE_X15Y116_CO5),
.O6(CLBLM_R_X11Y116_SLICE_X15Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y116_SLICE_X15Y116_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y116_SLICE_X15Y116_BO5),
.O6(CLBLM_R_X11Y116_SLICE_X15Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdddddd88d8d8d888)
  ) CLBLM_R_X11Y116_SLICE_X15Y116_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X12Y114_SLICE_X17Y114_AQ),
.I2(CLBLM_R_X11Y116_SLICE_X15Y116_AQ),
.I3(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLM_L_X10Y111_SLICE_X13Y111_DO6),
.O5(CLBLM_R_X11Y116_SLICE_X15Y116_AO5),
.O6(CLBLM_R_X11Y116_SLICE_X15Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff5fffdfff5fff)
  ) CLBLM_R_X11Y117_SLICE_X14Y117_DLUT (
.I0(CLBLM_L_X10Y118_SLICE_X12Y118_AQ),
.I1(CLBLM_L_X8Y118_SLICE_X10Y118_AQ),
.I2(CLBLM_L_X10Y118_SLICE_X13Y118_AQ),
.I3(CLBLM_L_X10Y118_SLICE_X12Y118_BQ),
.I4(CLBLM_R_X7Y118_SLICE_X8Y118_CQ),
.I5(CLBLM_L_X10Y119_SLICE_X12Y119_AQ),
.O5(CLBLM_R_X11Y117_SLICE_X14Y117_DO5),
.O6(CLBLM_R_X11Y117_SLICE_X14Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff004cb300ff)
  ) CLBLM_R_X11Y117_SLICE_X14Y117_CLUT (
.I0(CLBLM_L_X10Y117_SLICE_X13Y117_BO6),
.I1(CLBLM_L_X10Y116_SLICE_X12Y116_BQ),
.I2(CLBLM_L_X10Y117_SLICE_X13Y117_DO6),
.I3(CLBLM_R_X11Y117_SLICE_X15Y117_CQ),
.I4(CLBLM_R_X7Y118_SLICE_X9Y118_CO5),
.I5(CLBLM_L_X10Y117_SLICE_X12Y117_DO6),
.O5(CLBLM_R_X11Y117_SLICE_X14Y117_CO5),
.O6(CLBLM_R_X11Y117_SLICE_X14Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3311333331313333)
  ) CLBLM_R_X11Y117_SLICE_X14Y117_BLUT (
.I0(CLBLM_L_X10Y116_SLICE_X13Y116_AQ),
.I1(CLBLM_L_X10Y117_SLICE_X12Y117_DO6),
.I2(CLBLM_L_X10Y117_SLICE_X13Y117_BO6),
.I3(CLBLM_L_X10Y117_SLICE_X13Y117_DO6),
.I4(CLBLM_R_X7Y118_SLICE_X9Y118_CO5),
.I5(CLBLM_R_X11Y117_SLICE_X15Y117_CQ),
.O5(CLBLM_R_X11Y117_SLICE_X14Y117_BO5),
.O6(CLBLM_R_X11Y117_SLICE_X14Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h2303330333333333)
  ) CLBLM_R_X11Y117_SLICE_X14Y117_ALUT (
.I0(CLBLM_R_X11Y117_SLICE_X14Y117_DO6),
.I1(CLBLM_L_X10Y117_SLICE_X12Y117_DO6),
.I2(CLBLM_R_X7Y118_SLICE_X9Y118_CO5),
.I3(CLBLM_L_X10Y119_SLICE_X12Y119_CO6),
.I4(CLBLM_R_X11Y116_SLICE_X14Y116_BQ),
.I5(CLBLM_L_X10Y116_SLICE_X12Y116_AQ),
.O5(CLBLM_R_X11Y117_SLICE_X14Y117_AO5),
.O6(CLBLM_R_X11Y117_SLICE_X14Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y117_SLICE_X15Y117_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y117_SLICE_X15Y117_AO6),
.Q(CLBLM_R_X11Y117_SLICE_X15Y117_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y117_SLICE_X15Y117_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y117_SLICE_X15Y117_CO6),
.Q(CLBLM_R_X11Y117_SLICE_X15Y117_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y117_SLICE_X15Y117_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y117_SLICE_X15Y117_DO6),
.Q(CLBLM_R_X11Y117_SLICE_X15Y117_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffecce33332002)
  ) CLBLM_R_X11Y117_SLICE_X15Y117_DLUT (
.I0(CLBLM_L_X10Y116_SLICE_X12Y116_DO5),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X11Y117_SLICE_X15Y117_DQ),
.I3(CLBLM_R_X11Y117_SLICE_X14Y117_BO6),
.I4(CLBLM_L_X10Y118_SLICE_X13Y118_CO6),
.I5(CLBLM_R_X11Y110_SLICE_X15Y110_A5Q),
.O5(CLBLM_R_X11Y117_SLICE_X15Y117_DO5),
.O6(CLBLM_R_X11Y117_SLICE_X15Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaf3aaf3aaf0aaf0)
  ) CLBLM_R_X11Y117_SLICE_X15Y117_CLUT (
.I0(CLBLM_R_X11Y116_SLICE_X15Y116_AQ),
.I1(CLBLM_R_X11Y117_SLICE_X14Y117_CO6),
.I2(CLBLM_L_X10Y118_SLICE_X13Y118_CO6),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLM_L_X10Y116_SLICE_X12Y116_DO5),
.O5(CLBLM_R_X11Y117_SLICE_X15Y117_CO5),
.O6(CLBLM_R_X11Y117_SLICE_X15Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaccaacc0000aaaa)
  ) CLBLM_R_X11Y117_SLICE_X15Y117_BLUT (
.I0(CLBLM_L_X10Y116_SLICE_X13Y116_AQ),
.I1(CLBLM_L_X10Y117_SLICE_X12Y117_A5Q),
.I2(1'b1),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y118_SLICE_X8Y118_DO6),
.I5(1'b1),
.O5(CLBLM_R_X11Y117_SLICE_X15Y117_BO5),
.O6(CLBLM_R_X11Y117_SLICE_X15Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff005e0000005e)
  ) CLBLM_R_X11Y117_SLICE_X15Y117_ALUT (
.I0(CLBLM_R_X11Y117_SLICE_X15Y117_BO5),
.I1(CLBLM_L_X10Y117_SLICE_X13Y117_AO6),
.I2(CLBLM_R_X11Y117_SLICE_X15Y117_AQ),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X12Y112_SLICE_X17Y112_A5Q),
.O5(CLBLM_R_X11Y117_SLICE_X15Y117_AO5),
.O6(CLBLM_R_X11Y117_SLICE_X15Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y118_SLICE_X14Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y118_SLICE_X14Y118_DO5),
.O6(CLBLM_R_X11Y118_SLICE_X14Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y118_SLICE_X14Y118_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y118_SLICE_X14Y118_CO5),
.O6(CLBLM_R_X11Y118_SLICE_X14Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y118_SLICE_X14Y118_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y118_SLICE_X14Y118_BO5),
.O6(CLBLM_R_X11Y118_SLICE_X14Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y118_SLICE_X14Y118_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y118_SLICE_X14Y118_AO5),
.O6(CLBLM_R_X11Y118_SLICE_X14Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y118_SLICE_X15Y118_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y118_SLICE_X15Y118_AO5),
.Q(CLBLM_R_X11Y118_SLICE_X15Y118_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y118_SLICE_X15Y118_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y118_SLICE_X15Y118_AO6),
.Q(CLBLM_R_X11Y118_SLICE_X15Y118_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y118_SLICE_X15Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y118_SLICE_X15Y118_DO5),
.O6(CLBLM_R_X11Y118_SLICE_X15Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y118_SLICE_X15Y118_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y118_SLICE_X15Y118_CO5),
.O6(CLBLM_R_X11Y118_SLICE_X15Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y118_SLICE_X15Y118_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y118_SLICE_X15Y118_BO5),
.O6(CLBLM_R_X11Y118_SLICE_X15Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdddd8888ff55aa00)
  ) CLBLM_R_X11Y118_SLICE_X15Y118_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLL_L_X4Y118_SLICE_X4Y118_AQ),
.I2(1'b1),
.I3(CLBLM_L_X12Y107_SLICE_X16Y107_BQ),
.I4(RIOB33_X105Y125_IOB_X1Y126_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y118_SLICE_X15Y118_AO5),
.O6(CLBLM_R_X11Y118_SLICE_X15Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y119_SLICE_X14Y119_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y119_SLICE_X14Y119_AO6),
.Q(CLBLM_R_X11Y119_SLICE_X14Y119_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y119_SLICE_X14Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y119_SLICE_X14Y119_DO5),
.O6(CLBLM_R_X11Y119_SLICE_X14Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y119_SLICE_X14Y119_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y119_SLICE_X14Y119_CO5),
.O6(CLBLM_R_X11Y119_SLICE_X14Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y119_SLICE_X14Y119_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y119_SLICE_X14Y119_BO5),
.O6(CLBLM_R_X11Y119_SLICE_X14Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccf0f0ccccfff0)
  ) CLBLM_R_X11Y119_SLICE_X14Y119_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y116_SLICE_X13Y116_BQ),
.I2(CLBLM_R_X11Y119_SLICE_X14Y119_AQ),
.I3(RIOB33_X105Y141_IOB_X1Y142_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y119_SLICE_X10Y119_AQ),
.O5(CLBLM_R_X11Y119_SLICE_X14Y119_AO5),
.O6(CLBLM_R_X11Y119_SLICE_X14Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y119_SLICE_X15Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y119_SLICE_X15Y119_DO5),
.O6(CLBLM_R_X11Y119_SLICE_X15Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y119_SLICE_X15Y119_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y119_SLICE_X15Y119_CO5),
.O6(CLBLM_R_X11Y119_SLICE_X15Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y119_SLICE_X15Y119_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y119_SLICE_X15Y119_BO5),
.O6(CLBLM_R_X11Y119_SLICE_X15Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y119_SLICE_X15Y119_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y119_SLICE_X15Y119_AO5),
.O6(CLBLM_R_X11Y119_SLICE_X15Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000011)
  ) CLBLM_R_X13Y106_SLICE_X18Y106_DLUT (
.I0(CLBLM_R_X13Y107_SLICE_X19Y107_AQ),
.I1(CLBLM_L_X12Y107_SLICE_X16Y107_AQ),
.I2(1'b1),
.I3(CLBLM_R_X13Y106_SLICE_X18Y106_CO6),
.I4(CLBLM_R_X13Y107_SLICE_X19Y107_BQ),
.I5(CLBLM_R_X13Y107_SLICE_X18Y107_AQ),
.O5(CLBLM_R_X13Y106_SLICE_X18Y106_DO5),
.O6(CLBLM_R_X13Y106_SLICE_X18Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffff1f)
  ) CLBLM_R_X13Y106_SLICE_X18Y106_CLUT (
.I0(CLBLM_R_X13Y109_SLICE_X19Y109_BQ),
.I1(CLBLM_L_X12Y107_SLICE_X17Y107_BQ),
.I2(CLBLM_R_X13Y113_SLICE_X18Y113_BQ),
.I3(CLBLM_L_X12Y107_SLICE_X16Y107_BQ),
.I4(CLBLM_R_X13Y108_SLICE_X19Y108_BQ),
.I5(CLBLM_L_X12Y108_SLICE_X16Y108_BQ),
.O5(CLBLM_R_X13Y106_SLICE_X18Y106_CO5),
.O6(CLBLM_R_X13Y106_SLICE_X18Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5ffd5ffffffffff)
  ) CLBLM_R_X13Y106_SLICE_X18Y106_BLUT (
.I0(CLBLM_R_X13Y108_SLICE_X19Y108_BQ),
.I1(CLBLM_R_X13Y109_SLICE_X19Y109_BQ),
.I2(CLBLM_R_X13Y113_SLICE_X18Y113_BQ),
.I3(CLBLM_L_X12Y108_SLICE_X16Y108_BQ),
.I4(CLBLM_L_X12Y107_SLICE_X17Y107_BQ),
.I5(CLBLM_L_X12Y107_SLICE_X16Y107_BQ),
.O5(CLBLM_R_X13Y106_SLICE_X18Y106_BO5),
.O6(CLBLM_R_X13Y106_SLICE_X18Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ffdf0000efcf)
  ) CLBLM_R_X13Y106_SLICE_X18Y106_ALUT (
.I0(CLBLM_R_X13Y107_SLICE_X19Y107_BQ),
.I1(CLBLM_L_X12Y105_SLICE_X17Y105_AO5),
.I2(CLBLM_L_X12Y107_SLICE_X16Y107_DQ),
.I3(CLBLM_R_X13Y106_SLICE_X18Y106_BO6),
.I4(CLBLM_L_X12Y105_SLICE_X17Y105_CO6),
.I5(CLBLM_R_X13Y106_SLICE_X18Y106_CO6),
.O5(CLBLM_R_X13Y106_SLICE_X18Y106_AO5),
.O6(CLBLM_R_X13Y106_SLICE_X18Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y106_SLICE_X19Y106_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y106_SLICE_X19Y106_DO5),
.O6(CLBLM_R_X13Y106_SLICE_X19Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y106_SLICE_X19Y106_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y106_SLICE_X19Y106_CO5),
.O6(CLBLM_R_X13Y106_SLICE_X19Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y106_SLICE_X19Y106_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y106_SLICE_X19Y106_BO5),
.O6(CLBLM_R_X13Y106_SLICE_X19Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y106_SLICE_X19Y106_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y106_SLICE_X19Y106_AO5),
.O6(CLBLM_R_X13Y106_SLICE_X19Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y107_SLICE_X18Y107_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y107_SLICE_X18Y107_AO6),
.Q(CLBLM_R_X13Y107_SLICE_X18Y107_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff7f7fffff)
  ) CLBLM_R_X13Y107_SLICE_X18Y107_DLUT (
.I0(CLBLM_R_X13Y107_SLICE_X19Y107_AQ),
.I1(CLBLM_R_X13Y107_SLICE_X18Y107_AQ),
.I2(CLBLM_L_X12Y107_SLICE_X16Y107_AQ),
.I3(1'b1),
.I4(CLBLM_R_X13Y107_SLICE_X19Y107_BQ),
.I5(CLBLM_R_X13Y106_SLICE_X18Y106_BO6),
.O5(CLBLM_R_X13Y107_SLICE_X18Y107_DO5),
.O6(CLBLM_R_X13Y107_SLICE_X18Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000080000000)
  ) CLBLM_R_X13Y107_SLICE_X18Y107_CLUT (
.I0(CLBLM_R_X13Y107_SLICE_X19Y107_AQ),
.I1(CLBLM_R_X13Y107_SLICE_X19Y107_BQ),
.I2(CLBLM_R_X13Y107_SLICE_X18Y107_AQ),
.I3(CLBLM_R_X13Y108_SLICE_X18Y108_AQ),
.I4(CLBLM_L_X12Y107_SLICE_X16Y107_AQ),
.I5(CLBLM_R_X13Y106_SLICE_X18Y106_BO6),
.O5(CLBLM_R_X13Y107_SLICE_X18Y107_CO5),
.O6(CLBLM_R_X13Y107_SLICE_X18Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000001)
  ) CLBLM_R_X13Y107_SLICE_X18Y107_BLUT (
.I0(CLBLM_L_X12Y107_SLICE_X16Y107_AQ),
.I1(CLBLM_R_X13Y106_SLICE_X18Y106_CO6),
.I2(CLBLM_R_X13Y107_SLICE_X18Y107_AQ),
.I3(CLBLM_R_X13Y107_SLICE_X19Y107_BQ),
.I4(CLBLM_R_X13Y107_SLICE_X19Y107_AQ),
.I5(CLBLM_R_X13Y108_SLICE_X18Y108_AQ),
.O5(CLBLM_R_X13Y107_SLICE_X18Y107_BO5),
.O6(CLBLM_R_X13Y107_SLICE_X18Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa3333aaaa0330)
  ) CLBLM_R_X13Y107_SLICE_X18Y107_ALUT (
.I0(CLBLM_R_X13Y112_SLICE_X18Y112_CQ),
.I1(CLBLM_L_X12Y108_SLICE_X17Y108_CO5),
.I2(CLBLM_R_X13Y107_SLICE_X18Y107_AQ),
.I3(CLBLM_L_X12Y106_SLICE_X17Y106_BO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X12Y107_SLICE_X17Y107_CO5),
.O5(CLBLM_R_X13Y107_SLICE_X18Y107_AO5),
.O6(CLBLM_R_X13Y107_SLICE_X18Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y107_SLICE_X19Y107_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y107_SLICE_X19Y107_AO6),
.Q(CLBLM_R_X13Y107_SLICE_X19Y107_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y107_SLICE_X19Y107_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y107_SLICE_X19Y107_BO6),
.Q(CLBLM_R_X13Y107_SLICE_X19Y107_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h04cc000000003200)
  ) CLBLM_R_X13Y107_SLICE_X19Y107_DLUT (
.I0(CLBLM_L_X12Y107_SLICE_X17Y107_BQ),
.I1(CLBLM_L_X12Y107_SLICE_X16Y107_BQ),
.I2(CLBLM_R_X13Y109_SLICE_X19Y109_BQ),
.I3(CLBLM_R_X13Y113_SLICE_X18Y113_BQ),
.I4(CLBLM_R_X13Y108_SLICE_X19Y108_BQ),
.I5(CLBLM_L_X12Y108_SLICE_X16Y108_BQ),
.O5(CLBLM_R_X13Y107_SLICE_X19Y107_DO5),
.O6(CLBLM_R_X13Y107_SLICE_X19Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff66566666)
  ) CLBLM_R_X13Y107_SLICE_X19Y107_CLUT (
.I0(CLBLM_R_X13Y107_SLICE_X19Y107_BQ),
.I1(CLBLM_L_X12Y105_SLICE_X17Y105_CO6),
.I2(CLBLM_L_X12Y108_SLICE_X16Y108_CQ),
.I3(CLBLM_L_X12Y105_SLICE_X17Y105_AO5),
.I4(CLBLM_R_X13Y107_SLICE_X19Y107_DO6),
.I5(CLBLM_L_X12Y107_SLICE_X17Y107_CO5),
.O5(CLBLM_R_X13Y107_SLICE_X19Y107_CO5),
.O6(CLBLM_R_X13Y107_SLICE_X19Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa00ffaaaa0000)
  ) CLBLM_R_X13Y107_SLICE_X19Y107_BLUT (
.I0(CLBLM_L_X10Y115_SLICE_X12Y115_CQ),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_L_X12Y108_SLICE_X17Y108_CO5),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X13Y107_SLICE_X19Y107_CO6),
.O5(CLBLM_R_X13Y107_SLICE_X19Y107_BO5),
.O6(CLBLM_R_X13Y107_SLICE_X19Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000feef5445)
  ) CLBLM_R_X13Y107_SLICE_X19Y107_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X12Y107_SLICE_X17Y107_CO5),
.I2(CLBLM_R_X13Y107_SLICE_X19Y107_AQ),
.I3(CLBLM_R_X13Y106_SLICE_X18Y106_AO6),
.I4(CLBLM_R_X7Y108_SLICE_X8Y108_BQ),
.I5(CLBLM_L_X12Y108_SLICE_X17Y108_CO5),
.O5(CLBLM_R_X13Y107_SLICE_X19Y107_AO5),
.O6(CLBLM_R_X13Y107_SLICE_X19Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y108_SLICE_X18Y108_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y108_SLICE_X18Y108_AO6),
.Q(CLBLM_R_X13Y108_SLICE_X18Y108_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ba00ffff45ff00)
  ) CLBLM_R_X13Y108_SLICE_X18Y108_DLUT (
.I0(CLBLM_L_X12Y105_SLICE_X17Y105_AO5),
.I1(CLBLM_R_X13Y106_SLICE_X18Y106_DO6),
.I2(CLBLM_R_X13Y107_SLICE_X18Y107_DO6),
.I3(CLBLM_L_X12Y105_SLICE_X17Y105_CO6),
.I4(CLBLM_L_X12Y108_SLICE_X17Y108_AQ),
.I5(CLBLM_R_X13Y108_SLICE_X18Y108_AQ),
.O5(CLBLM_R_X13Y108_SLICE_X18Y108_DO5),
.O6(CLBLM_R_X13Y108_SLICE_X18Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h333333339c9c9ccc)
  ) CLBLM_R_X13Y108_SLICE_X18Y108_CLUT (
.I0(CLBLM_L_X12Y105_SLICE_X17Y105_AO5),
.I1(CLBLM_R_X13Y108_SLICE_X19Y108_AQ),
.I2(CLBLM_R_X11Y108_SLICE_X14Y108_AQ),
.I3(CLBLM_R_X13Y107_SLICE_X18Y107_BO6),
.I4(CLBLM_R_X13Y107_SLICE_X18Y107_CO6),
.I5(CLBLM_L_X12Y105_SLICE_X17Y105_CO6),
.O5(CLBLM_R_X13Y108_SLICE_X18Y108_CO5),
.O6(CLBLM_R_X13Y108_SLICE_X18Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h2222330022223300)
  ) CLBLM_R_X13Y108_SLICE_X18Y108_BLUT (
.I0(CLBLM_R_X13Y107_SLICE_X18Y107_CO6),
.I1(CLBLM_L_X12Y105_SLICE_X17Y105_AO5),
.I2(1'b1),
.I3(CLBLM_R_X13Y107_SLICE_X18Y107_BO6),
.I4(CLBLM_R_X13Y108_SLICE_X19Y108_AQ),
.I5(1'b1),
.O5(CLBLM_R_X13Y108_SLICE_X18Y108_BO5),
.O6(CLBLM_R_X13Y108_SLICE_X18Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0f5e4f5e4)
  ) CLBLM_R_X13Y108_SLICE_X18Y108_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X13Y108_SLICE_X18Y108_DO6),
.I2(CLBLM_L_X12Y109_SLICE_X17Y109_DQ),
.I3(CLBLM_L_X12Y107_SLICE_X17Y107_CO5),
.I4(1'b1),
.I5(CLBLM_L_X12Y108_SLICE_X17Y108_CO5),
.O5(CLBLM_R_X13Y108_SLICE_X18Y108_AO5),
.O6(CLBLM_R_X13Y108_SLICE_X18Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y108_SLICE_X19Y108_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y108_SLICE_X19Y108_AO6),
.Q(CLBLM_R_X13Y108_SLICE_X19Y108_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y108_SLICE_X19Y108_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y108_SLICE_X19Y108_BO6),
.Q(CLBLM_R_X13Y108_SLICE_X19Y108_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y108_SLICE_X19Y108_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y108_SLICE_X19Y108_DO5),
.O6(CLBLM_R_X13Y108_SLICE_X19Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff0fb40fb4)
  ) CLBLM_R_X13Y108_SLICE_X19Y108_CLUT (
.I0(CLBLM_L_X12Y105_SLICE_X17Y105_AO5),
.I1(CLBLM_L_X12Y108_SLICE_X16Y108_DQ),
.I2(CLBLM_R_X13Y108_SLICE_X19Y108_BQ),
.I3(CLBLM_L_X12Y105_SLICE_X17Y105_CO6),
.I4(1'b1),
.I5(CLBLM_L_X12Y107_SLICE_X17Y107_CO5),
.O5(CLBLM_R_X13Y108_SLICE_X19Y108_CO5),
.O6(CLBLM_R_X13Y108_SLICE_X19Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbbb1111aaaa0000)
  ) CLBLM_R_X13Y108_SLICE_X19Y108_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X12Y108_SLICE_X17Y108_CO5),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_L_X10Y114_SLICE_X12Y114_CQ),
.I5(CLBLM_R_X13Y108_SLICE_X19Y108_CO6),
.O5(CLBLM_R_X13Y108_SLICE_X19Y108_BO5),
.O6(CLBLM_R_X13Y108_SLICE_X19Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbba1110bbba1110)
  ) CLBLM_R_X13Y108_SLICE_X19Y108_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X12Y108_SLICE_X17Y108_CO5),
.I2(CLBLM_R_X13Y108_SLICE_X18Y108_CO6),
.I3(CLBLM_L_X12Y107_SLICE_X17Y107_CO5),
.I4(CLBLM_L_X12Y107_SLICE_X17Y107_BQ),
.I5(1'b1),
.O5(CLBLM_R_X13Y108_SLICE_X19Y108_AO5),
.O6(CLBLM_R_X13Y108_SLICE_X19Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y109_SLICE_X18Y109_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y109_SLICE_X18Y109_AO6),
.Q(CLBLM_R_X13Y109_SLICE_X18Y109_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hc8ffc8888cff8ccc)
  ) CLBLM_R_X13Y109_SLICE_X18Y109_DLUT (
.I0(CLBLM_L_X12Y108_SLICE_X17Y108_DO6),
.I1(CLBLM_R_X13Y109_SLICE_X18Y109_AQ),
.I2(CLBLM_R_X11Y110_SLICE_X15Y110_A5Q),
.I3(CLBLM_L_X12Y107_SLICE_X17Y107_AQ),
.I4(CLBLM_R_X13Y109_SLICE_X18Y109_BO5),
.I5(CLBLM_R_X13Y109_SLICE_X18Y109_BO6),
.O5(CLBLM_R_X13Y109_SLICE_X18Y109_DO5),
.O6(CLBLM_R_X13Y109_SLICE_X18Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0ea3cbe00000000)
  ) CLBLM_R_X13Y109_SLICE_X18Y109_CLUT (
.I0(CLBLM_L_X12Y107_SLICE_X17Y107_DO5),
.I1(CLBLM_R_X13Y109_SLICE_X19Y109_BQ),
.I2(CLBLM_R_X13Y113_SLICE_X18Y113_BQ),
.I3(CLBLM_L_X12Y107_SLICE_X17Y107_AQ),
.I4(CLBLM_L_X12Y107_SLICE_X17Y107_BQ),
.I5(CLBLM_R_X13Y108_SLICE_X18Y108_BO6),
.O5(CLBLM_R_X13Y109_SLICE_X18Y109_CO5),
.O6(CLBLM_R_X13Y109_SLICE_X18Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0acaca00003300)
  ) CLBLM_R_X13Y109_SLICE_X18Y109_BLUT (
.I0(CLBLM_L_X12Y105_SLICE_X16Y105_AQ),
.I1(CLBLM_R_X13Y113_SLICE_X18Y113_BQ),
.I2(CLBLM_R_X11Y105_SLICE_X14Y105_DQ),
.I3(CLBLM_R_X13Y109_SLICE_X19Y109_BQ),
.I4(CLBLM_L_X12Y107_SLICE_X17Y107_BQ),
.I5(1'b1),
.O5(CLBLM_R_X13Y109_SLICE_X18Y109_BO5),
.O6(CLBLM_R_X13Y109_SLICE_X18Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000fa0afa0a)
  ) CLBLM_R_X13Y109_SLICE_X18Y109_ALUT (
.I0(CLBLM_R_X13Y109_SLICE_X18Y109_DO6),
.I1(1'b1),
.I2(CLBLM_L_X12Y105_SLICE_X16Y105_BO6),
.I3(CLBLM_R_X7Y116_SLICE_X9Y116_BO6),
.I4(CLBLM_R_X13Y108_SLICE_X19Y108_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X13Y109_SLICE_X18Y109_AO5),
.O6(CLBLM_R_X13Y109_SLICE_X18Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y109_SLICE_X19Y109_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y109_SLICE_X19Y109_AO6),
.Q(CLBLM_R_X13Y109_SLICE_X19Y109_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y109_SLICE_X19Y109_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y109_SLICE_X19Y109_BO6),
.Q(CLBLM_R_X13Y109_SLICE_X19Y109_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y109_SLICE_X19Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y109_SLICE_X19Y109_DO5),
.O6(CLBLM_R_X13Y109_SLICE_X19Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y109_SLICE_X19Y109_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y109_SLICE_X19Y109_CO5),
.O6(CLBLM_R_X13Y109_SLICE_X19Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc55cc00ccfacc00)
  ) CLBLM_R_X13Y109_SLICE_X19Y109_BLUT (
.I0(CLBLM_R_X13Y109_SLICE_X18Y109_CO6),
.I1(CLBLM_R_X13Y110_SLICE_X19Y110_AQ),
.I2(CLBLM_L_X12Y105_SLICE_X16Y105_BO6),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(CLBLM_R_X13Y109_SLICE_X19Y109_BQ),
.O5(CLBLM_R_X13Y109_SLICE_X19Y109_BO5),
.O6(CLBLM_R_X13Y109_SLICE_X19Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff4fff400f400f4)
  ) CLBLM_R_X13Y109_SLICE_X19Y109_ALUT (
.I0(CLBLM_L_X8Y119_SLICE_X10Y119_AQ),
.I1(RIOB33_X105Y141_IOB_X1Y142_I),
.I2(CLBLM_R_X13Y109_SLICE_X19Y109_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLM_R_X13Y112_SLICE_X18Y112_A5Q),
.O5(CLBLM_R_X13Y109_SLICE_X19Y109_AO5),
.O6(CLBLM_R_X13Y109_SLICE_X19Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y110_SLICE_X18Y110_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y110_SLICE_X18Y110_AO6),
.Q(CLBLM_R_X13Y110_SLICE_X18Y110_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y110_SLICE_X18Y110_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y110_SLICE_X18Y110_BO6),
.Q(CLBLM_R_X13Y110_SLICE_X18Y110_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y110_SLICE_X18Y110_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y110_SLICE_X18Y110_CO6),
.Q(CLBLM_R_X13Y110_SLICE_X18Y110_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000eeee0000fff0)
  ) CLBLM_R_X13Y110_SLICE_X18Y110_DLUT (
.I0(CLBLM_R_X13Y110_SLICE_X18Y110_CQ),
.I1(CLBLM_R_X11Y107_SLICE_X15Y107_CQ),
.I2(CLBLM_L_X12Y109_SLICE_X17Y109_DQ),
.I3(CLBLM_R_X13Y110_SLICE_X19Y110_CQ),
.I4(CLBLM_L_X10Y113_SLICE_X13Y113_CQ),
.I5(1'b1),
.O5(CLBLM_R_X13Y110_SLICE_X18Y110_DO5),
.O6(CLBLM_R_X13Y110_SLICE_X18Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaafcfcfc00)
  ) CLBLM_R_X13Y110_SLICE_X18Y110_CLUT (
.I0(CLBLL_L_X4Y110_SLICE_X4Y110_B5Q),
.I1(CLBLM_R_X13Y110_SLICE_X18Y110_CQ),
.I2(CLBLM_L_X10Y109_SLICE_X13Y109_CO6),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X13Y110_SLICE_X18Y110_CO5),
.O6(CLBLM_R_X13Y110_SLICE_X18Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0cfc0cfc0)
  ) CLBLM_R_X13Y110_SLICE_X18Y110_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X13Y108_SLICE_X19Y108_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X11Y111_SLICE_X15Y111_BQ),
.I4(1'b1),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X13Y110_SLICE_X18Y110_BO5),
.O6(CLBLM_R_X13Y110_SLICE_X18Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000ffa800a8)
  ) CLBLM_R_X13Y110_SLICE_X18Y110_ALUT (
.I0(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.I1(CLBLM_L_X12Y109_SLICE_X16Y109_BQ),
.I2(CLBLM_R_X13Y110_SLICE_X18Y110_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X13Y110_SLICE_X18Y110_CQ),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_R_X13Y110_SLICE_X18Y110_AO5),
.O6(CLBLM_R_X13Y110_SLICE_X18Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y110_SLICE_X19Y110_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y110_SLICE_X19Y110_AO6),
.Q(CLBLM_R_X13Y110_SLICE_X19Y110_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y110_SLICE_X19Y110_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y110_SLICE_X19Y110_BO6),
.Q(CLBLM_R_X13Y110_SLICE_X19Y110_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y110_SLICE_X19Y110_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y110_SLICE_X19Y110_CO6),
.Q(CLBLM_R_X13Y110_SLICE_X19Y110_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y110_SLICE_X19Y110_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y110_SLICE_X19Y110_DO5),
.O6(CLBLM_R_X13Y110_SLICE_X19Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffe4e4ffffe4a0)
  ) CLBLM_R_X13Y110_SLICE_X19Y110_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X13Y110_SLICE_X19Y110_CQ),
.I2(CLBLM_R_X11Y112_SLICE_X14Y112_C5Q),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_L_X10Y109_SLICE_X12Y109_DO6),
.I5(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.O5(CLBLM_R_X13Y110_SLICE_X19Y110_CO5),
.O6(CLBLM_R_X13Y110_SLICE_X19Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafafcfcfafafcf0)
  ) CLBLM_R_X13Y110_SLICE_X19Y110_BLUT (
.I0(CLBLM_L_X12Y110_SLICE_X16Y110_AQ),
.I1(CLBLM_R_X13Y110_SLICE_X19Y110_BQ),
.I2(CLBLM_L_X10Y109_SLICE_X12Y109_DO6),
.I3(CLBLM_L_X8Y116_SLICE_X10Y116_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_R_X13Y110_SLICE_X19Y110_BO5),
.O6(CLBLM_R_X13Y110_SLICE_X19Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff400040ff040004)
  ) CLBLM_R_X13Y110_SLICE_X19Y110_ALUT (
.I0(CLBLM_R_X7Y115_SLICE_X8Y115_DQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X13Y110_SLICE_X19Y110_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X13Y109_SLICE_X18Y109_AQ),
.I5(CLBLM_L_X12Y110_SLICE_X16Y110_DO6),
.O5(CLBLM_R_X13Y110_SLICE_X19Y110_AO5),
.O6(CLBLM_R_X13Y110_SLICE_X19Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y112_SLICE_X18Y112_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y112_SLICE_X18Y112_AO5),
.Q(CLBLM_R_X13Y112_SLICE_X18Y112_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y112_SLICE_X18Y112_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y112_SLICE_X18Y112_AO6),
.Q(CLBLM_R_X13Y112_SLICE_X18Y112_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y112_SLICE_X18Y112_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y112_SLICE_X18Y112_BO6),
.Q(CLBLM_R_X13Y112_SLICE_X18Y112_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y112_SLICE_X18Y112_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y112_SLICE_X18Y112_CO6),
.Q(CLBLM_R_X13Y112_SLICE_X18Y112_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h999999999c9c9c9c)
  ) CLBLM_R_X13Y112_SLICE_X18Y112_DLUT (
.I0(CLBLM_R_X13Y110_SLICE_X18Y110_BQ),
.I1(CLBLM_L_X12Y111_SLICE_X16Y111_DQ),
.I2(CLBLM_R_X13Y112_SLICE_X18Y112_BQ),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X10Y112_SLICE_X13Y112_AO6),
.O5(CLBLM_R_X13Y112_SLICE_X18Y112_DO5),
.O6(CLBLM_R_X13Y112_SLICE_X18Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hee44ee44aa00aa00)
  ) CLBLM_R_X13Y112_SLICE_X18Y112_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(1'b1),
.I3(CLBLM_L_X10Y114_SLICE_X13Y114_AQ),
.I4(1'b1),
.I5(CLBLM_L_X12Y109_SLICE_X17Y109_CQ),
.O5(CLBLM_R_X13Y112_SLICE_X18Y112_CO5),
.O6(CLBLM_R_X13Y112_SLICE_X18Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f10001f6f80608)
  ) CLBLM_R_X13Y112_SLICE_X18Y112_BLUT (
.I0(CLBLM_R_X13Y112_SLICE_X18Y112_DO6),
.I1(CLBLM_R_X13Y112_SLICE_X18Y112_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X12Y111_SLICE_X16Y111_CQ),
.I4(CLBLM_L_X12Y113_SLICE_X17Y113_B5Q),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X13Y112_SLICE_X18Y112_BO5),
.O6(CLBLM_R_X13Y112_SLICE_X18Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00f0f0ccccaaaa)
  ) CLBLM_R_X13Y112_SLICE_X18Y112_ALUT (
.I0(CLBLM_L_X12Y112_SLICE_X16Y112_A5Q),
.I1(CLBLM_R_X5Y112_SLICE_X6Y112_BQ),
.I2(RIOB33_X105Y103_IOB_X1Y104_I),
.I3(CLBLM_L_X12Y114_SLICE_X17Y114_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X13Y112_SLICE_X18Y112_AO5),
.O6(CLBLM_R_X13Y112_SLICE_X18Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y112_SLICE_X19Y112_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y112_SLICE_X19Y112_DO5),
.O6(CLBLM_R_X13Y112_SLICE_X19Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y112_SLICE_X19Y112_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y112_SLICE_X19Y112_CO5),
.O6(CLBLM_R_X13Y112_SLICE_X19Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y112_SLICE_X19Y112_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y112_SLICE_X19Y112_BO5),
.O6(CLBLM_R_X13Y112_SLICE_X19Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y112_SLICE_X19Y112_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y112_SLICE_X19Y112_AO5),
.O6(CLBLM_R_X13Y112_SLICE_X19Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y113_SLICE_X18Y113_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y113_SLICE_X18Y113_AO6),
.Q(CLBLM_R_X13Y113_SLICE_X18Y113_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y113_SLICE_X18Y113_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y113_SLICE_X18Y113_BO6),
.Q(CLBLM_R_X13Y113_SLICE_X18Y113_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y113_SLICE_X18Y113_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y113_SLICE_X18Y113_CO6),
.Q(CLBLM_R_X13Y113_SLICE_X18Y113_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_R_X13Y113_SLICE_X18Y113_DLUT (
.I0(RIOB33_X105Y133_IOB_X1Y133_I),
.I1(RIOB33_X105Y127_IOB_X1Y128_I),
.I2(RIOB33_X105Y129_IOB_X1Y130_I),
.I3(RIOB33_X105Y133_IOB_X1Y134_I),
.I4(RIOB33_X105Y137_IOB_X1Y137_I),
.I5(RIOB33_X105Y131_IOB_X1Y132_I),
.O5(CLBLM_R_X13Y113_SLICE_X18Y113_DO5),
.O6(CLBLM_R_X13Y113_SLICE_X18Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haafe0054aafe0054)
  ) CLBLM_R_X13Y113_SLICE_X18Y113_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X13Y113_SLICE_X18Y113_CQ),
.I2(CLBLM_L_X12Y114_SLICE_X17Y114_BQ),
.I3(CLBLM_R_X5Y115_SLICE_X7Y115_CO6),
.I4(CLBLM_L_X12Y112_SLICE_X16Y112_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X13Y113_SLICE_X18Y113_CO5),
.O6(CLBLM_R_X13Y113_SLICE_X18Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hae04ae04af05aa00)
  ) CLBLM_R_X13Y113_SLICE_X18Y113_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X13Y109_SLICE_X19Y109_BQ),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLM_R_X7Y115_SLICE_X8Y115_D5Q),
.I4(CLBLM_R_X13Y113_SLICE_X18Y113_BQ),
.I5(CLBLM_R_X13Y108_SLICE_X18Y108_BO6),
.O5(CLBLM_R_X13Y113_SLICE_X18Y113_BO5),
.O6(CLBLM_R_X13Y113_SLICE_X18Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f3f3e2f3f3f3f3)
  ) CLBLM_R_X13Y113_SLICE_X18Y113_ALUT (
.I0(CLBLM_R_X13Y113_SLICE_X18Y113_DO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X12Y115_SLICE_X16Y115_AQ),
.I3(RIOB33_X105Y135_IOB_X1Y136_I),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(RIOB33_X105Y135_IOB_X1Y135_I),
.O5(CLBLM_R_X13Y113_SLICE_X18Y113_AO5),
.O6(CLBLM_R_X13Y113_SLICE_X18Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y113_SLICE_X19Y113_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y113_SLICE_X19Y113_AO6),
.Q(CLBLM_R_X13Y113_SLICE_X19Y113_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y113_SLICE_X19Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y113_SLICE_X19Y113_DO5),
.O6(CLBLM_R_X13Y113_SLICE_X19Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y113_SLICE_X19Y113_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y113_SLICE_X19Y113_CO5),
.O6(CLBLM_R_X13Y113_SLICE_X19Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y113_SLICE_X19Y113_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y113_SLICE_X19Y113_BO5),
.O6(CLBLM_R_X13Y113_SLICE_X19Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000f3f0f3f0)
  ) CLBLM_R_X13Y113_SLICE_X19Y113_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y119_SLICE_X10Y119_AQ),
.I2(CLBLM_R_X13Y113_SLICE_X19Y113_AQ),
.I3(RIOB33_X105Y141_IOB_X1Y142_I),
.I4(CLBLM_R_X13Y108_SLICE_X18Y108_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X13Y113_SLICE_X19Y113_AO5),
.O6(CLBLM_R_X13Y113_SLICE_X19Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y117_SLICE_X18Y117_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y118_SLICE_X18Y118_AO5),
.Q(CLBLM_R_X13Y117_SLICE_X18Y117_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y117_SLICE_X18Y117_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y117_SLICE_X18Y117_AO6),
.Q(CLBLM_R_X13Y117_SLICE_X18Y117_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y117_SLICE_X18Y117_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y117_SLICE_X18Y117_DO5),
.O6(CLBLM_R_X13Y117_SLICE_X18Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y117_SLICE_X18Y117_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y117_SLICE_X18Y117_CO5),
.O6(CLBLM_R_X13Y117_SLICE_X18Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y117_SLICE_X18Y117_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y117_SLICE_X18Y117_BO5),
.O6(CLBLM_R_X13Y117_SLICE_X18Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000fc0cff55ff55)
  ) CLBLM_R_X13Y117_SLICE_X18Y117_ALUT (
.I0(RIOB33_X105Y143_IOB_X1Y143_I),
.I1(CLBLM_R_X7Y115_SLICE_X9Y115_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X12Y117_SLICE_X16Y117_AQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_R_X13Y117_SLICE_X18Y117_AO5),
.O6(CLBLM_R_X13Y117_SLICE_X18Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y117_SLICE_X19Y117_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y117_SLICE_X19Y117_DO5),
.O6(CLBLM_R_X13Y117_SLICE_X19Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y117_SLICE_X19Y117_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y117_SLICE_X19Y117_CO5),
.O6(CLBLM_R_X13Y117_SLICE_X19Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y117_SLICE_X19Y117_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y117_SLICE_X19Y117_BO5),
.O6(CLBLM_R_X13Y117_SLICE_X19Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y117_SLICE_X19Y117_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y117_SLICE_X19Y117_AO5),
.O6(CLBLM_R_X13Y117_SLICE_X19Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y118_SLICE_X18Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y118_SLICE_X18Y118_DO5),
.O6(CLBLM_R_X13Y118_SLICE_X18Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y118_SLICE_X18Y118_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y118_SLICE_X18Y118_CO5),
.O6(CLBLM_R_X13Y118_SLICE_X18Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y118_SLICE_X18Y118_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y118_SLICE_X18Y118_BO5),
.O6(CLBLM_R_X13Y118_SLICE_X18Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00fffffc0cfc0c)
  ) CLBLM_R_X13Y118_SLICE_X18Y118_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X12Y115_SLICE_X16Y115_AQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X12Y118_SLICE_X16Y118_AQ),
.I4(RIOB33_X105Y143_IOB_X1Y143_I),
.I5(1'b1),
.O5(CLBLM_R_X13Y118_SLICE_X18Y118_AO5),
.O6(CLBLM_R_X13Y118_SLICE_X18Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y118_SLICE_X19Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y118_SLICE_X19Y118_DO5),
.O6(CLBLM_R_X13Y118_SLICE_X19Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y118_SLICE_X19Y118_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y118_SLICE_X19Y118_CO5),
.O6(CLBLM_R_X13Y118_SLICE_X19Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y118_SLICE_X19Y118_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y118_SLICE_X19Y118_BO5),
.O6(CLBLM_R_X13Y118_SLICE_X19Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y118_SLICE_X19Y118_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y118_SLICE_X19Y118_AO5),
.O6(CLBLM_R_X13Y118_SLICE_X19Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X37Y117_SLICE_X56Y117_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X37Y117_SLICE_X56Y117_DO5),
.O6(CLBLM_R_X37Y117_SLICE_X56Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X37Y117_SLICE_X56Y117_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X37Y117_SLICE_X56Y117_CO5),
.O6(CLBLM_R_X37Y117_SLICE_X56Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X37Y117_SLICE_X56Y117_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X37Y117_SLICE_X56Y117_BO5),
.O6(CLBLM_R_X37Y117_SLICE_X56Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000050505050)
  ) CLBLM_R_X37Y117_SLICE_X56Y117_ALUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(1'b1),
.I2(RIOB33_X105Y119_IOB_X1Y119_I),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X8Y113_SLICE_X10Y113_DQ),
.O5(CLBLM_R_X37Y117_SLICE_X56Y117_AO5),
.O6(CLBLM_R_X37Y117_SLICE_X56Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X37Y117_SLICE_X57Y117_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X37Y117_SLICE_X57Y117_DO5),
.O6(CLBLM_R_X37Y117_SLICE_X57Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X37Y117_SLICE_X57Y117_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X37Y117_SLICE_X57Y117_CO5),
.O6(CLBLM_R_X37Y117_SLICE_X57Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X37Y117_SLICE_X57Y117_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X37Y117_SLICE_X57Y117_BO5),
.O6(CLBLM_R_X37Y117_SLICE_X57Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X37Y117_SLICE_X57Y117_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X37Y117_SLICE_X57Y117_AO5),
.O6(CLBLM_R_X37Y117_SLICE_X57Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y138_SLICE_X162Y138_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y138_SLICE_X162Y138_DO5),
.O6(CLBLM_R_X103Y138_SLICE_X162Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y138_SLICE_X162Y138_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y138_SLICE_X162Y138_CO5),
.O6(CLBLM_R_X103Y138_SLICE_X162Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y138_SLICE_X162Y138_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y138_SLICE_X162Y138_BO5),
.O6(CLBLM_R_X103Y138_SLICE_X162Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y138_SLICE_X162Y138_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y138_SLICE_X162Y138_AO5),
.O6(CLBLM_R_X103Y138_SLICE_X162Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y138_SLICE_X163Y138_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y138_SLICE_X163Y138_DO5),
.O6(CLBLM_R_X103Y138_SLICE_X163Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y138_SLICE_X163Y138_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y138_SLICE_X163Y138_CO5),
.O6(CLBLM_R_X103Y138_SLICE_X163Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y138_SLICE_X163Y138_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y138_SLICE_X163Y138_BO5),
.O6(CLBLM_R_X103Y138_SLICE_X163Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa0000000000)
  ) CLBLM_R_X103Y138_SLICE_X163Y138_ALUT (
.I0(RIOB33_X105Y139_IOB_X1Y139_I),
.I1(1'b1),
.I2(1'b1),
.I3(RIOB33_X105Y137_IOB_X1Y138_I),
.I4(1'b1),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X103Y138_SLICE_X163Y138_AO5),
.O6(CLBLM_R_X103Y138_SLICE_X163Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y169_SLICE_X162Y169_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y169_SLICE_X162Y169_DO5),
.O6(CLBLM_R_X103Y169_SLICE_X162Y169_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y169_SLICE_X162Y169_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y169_SLICE_X162Y169_CO5),
.O6(CLBLM_R_X103Y169_SLICE_X162Y169_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y169_SLICE_X162Y169_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y169_SLICE_X162Y169_BO5),
.O6(CLBLM_R_X103Y169_SLICE_X162Y169_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y169_SLICE_X162Y169_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y169_SLICE_X162Y169_AO5),
.O6(CLBLM_R_X103Y169_SLICE_X162Y169_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y169_SLICE_X163Y169_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y169_SLICE_X163Y169_DO5),
.O6(CLBLM_R_X103Y169_SLICE_X163Y169_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y169_SLICE_X163Y169_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y169_SLICE_X163Y169_CO5),
.O6(CLBLM_R_X103Y169_SLICE_X163Y169_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y169_SLICE_X163Y169_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y169_SLICE_X163Y169_BO5),
.O6(CLBLM_R_X103Y169_SLICE_X163Y169_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0fff0fff0fff0f)
  ) CLBLM_R_X103Y169_SLICE_X163Y169_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(RIOB33_X105Y143_IOB_X1Y143_I),
.I3(CLBLM_R_X11Y115_SLICE_X14Y115_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y169_SLICE_X163Y169_AO5),
.O6(CLBLM_R_X103Y169_SLICE_X163Y169_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y170_SLICE_X162Y170_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y170_SLICE_X162Y170_DO5),
.O6(CLBLM_R_X103Y170_SLICE_X162Y170_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y170_SLICE_X162Y170_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y170_SLICE_X162Y170_CO5),
.O6(CLBLM_R_X103Y170_SLICE_X162Y170_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y170_SLICE_X162Y170_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y170_SLICE_X162Y170_BO5),
.O6(CLBLM_R_X103Y170_SLICE_X162Y170_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y170_SLICE_X162Y170_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y170_SLICE_X162Y170_AO5),
.O6(CLBLM_R_X103Y170_SLICE_X162Y170_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y170_SLICE_X163Y170_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y170_SLICE_X163Y170_DO5),
.O6(CLBLM_R_X103Y170_SLICE_X163Y170_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y170_SLICE_X163Y170_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y170_SLICE_X163Y170_CO5),
.O6(CLBLM_R_X103Y170_SLICE_X163Y170_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y170_SLICE_X163Y170_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y170_SLICE_X163Y170_BO5),
.O6(CLBLM_R_X103Y170_SLICE_X163Y170_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ffffccccffff)
  ) CLBLM_R_X103Y170_SLICE_X163Y170_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y112_SLICE_X13Y112_AQ),
.I2(CLBLM_L_X12Y117_SLICE_X17Y117_AQ),
.I3(1'b1),
.I4(RIOB33_X105Y143_IOB_X1Y143_I),
.I5(1'b1),
.O5(CLBLM_R_X103Y170_SLICE_X163Y170_AO5),
.O6(CLBLM_R_X103Y170_SLICE_X163Y170_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y173_SLICE_X162Y173_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y173_SLICE_X162Y173_DO5),
.O6(CLBLM_R_X103Y173_SLICE_X162Y173_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y173_SLICE_X162Y173_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y173_SLICE_X162Y173_CO5),
.O6(CLBLM_R_X103Y173_SLICE_X162Y173_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y173_SLICE_X162Y173_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y173_SLICE_X162Y173_BO5),
.O6(CLBLM_R_X103Y173_SLICE_X162Y173_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y173_SLICE_X162Y173_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y173_SLICE_X162Y173_AO5),
.O6(CLBLM_R_X103Y173_SLICE_X162Y173_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y173_SLICE_X163Y173_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y173_SLICE_X163Y173_DO5),
.O6(CLBLM_R_X103Y173_SLICE_X163Y173_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y173_SLICE_X163Y173_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y173_SLICE_X163Y173_CO5),
.O6(CLBLM_R_X103Y173_SLICE_X163Y173_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y173_SLICE_X163Y173_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y173_SLICE_X163Y173_BO5),
.O6(CLBLM_R_X103Y173_SLICE_X163Y173_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff00fff0fff0ff)
  ) CLBLM_R_X103Y173_SLICE_X163Y173_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X11Y115_SLICE_X14Y115_AQ),
.I3(RIOB33_X105Y143_IOB_X1Y143_I),
.I4(CLBLM_R_X13Y113_SLICE_X19Y113_AQ),
.I5(1'b1),
.O5(CLBLM_R_X103Y173_SLICE_X163Y173_AO5),
.O6(CLBLM_R_X103Y173_SLICE_X163Y173_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y174_SLICE_X162Y174_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y174_SLICE_X162Y174_DO5),
.O6(CLBLM_R_X103Y174_SLICE_X162Y174_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y174_SLICE_X162Y174_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y174_SLICE_X162Y174_CO5),
.O6(CLBLM_R_X103Y174_SLICE_X162Y174_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y174_SLICE_X162Y174_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y174_SLICE_X162Y174_BO5),
.O6(CLBLM_R_X103Y174_SLICE_X162Y174_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y174_SLICE_X162Y174_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y174_SLICE_X162Y174_AO5),
.O6(CLBLM_R_X103Y174_SLICE_X162Y174_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y174_SLICE_X163Y174_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y174_SLICE_X163Y174_DO5),
.O6(CLBLM_R_X103Y174_SLICE_X163Y174_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y174_SLICE_X163Y174_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y174_SLICE_X163Y174_CO5),
.O6(CLBLM_R_X103Y174_SLICE_X163Y174_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y174_SLICE_X163Y174_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y174_SLICE_X163Y174_BO5),
.O6(CLBLM_R_X103Y174_SLICE_X163Y174_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00fffff0f0ffff)
  ) CLBLM_R_X103Y174_SLICE_X163Y174_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X11Y119_SLICE_X14Y119_AQ),
.I3(CLBLM_R_X13Y109_SLICE_X19Y109_AQ),
.I4(RIOB33_X105Y143_IOB_X1Y143_I),
.I5(1'b1),
.O5(CLBLM_R_X103Y174_SLICE_X163Y174_AO5),
.O6(CLBLM_R_X103Y174_SLICE_X163Y174_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y177_SLICE_X162Y177_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X162Y177_DO5),
.O6(CLBLM_R_X103Y177_SLICE_X162Y177_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y177_SLICE_X162Y177_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X162Y177_CO5),
.O6(CLBLM_R_X103Y177_SLICE_X162Y177_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y177_SLICE_X162Y177_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X162Y177_BO5),
.O6(CLBLM_R_X103Y177_SLICE_X162Y177_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y177_SLICE_X162Y177_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X162Y177_AO5),
.O6(CLBLM_R_X103Y177_SLICE_X162Y177_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y177_SLICE_X163Y177_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X163Y177_DO5),
.O6(CLBLM_R_X103Y177_SLICE_X163Y177_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y177_SLICE_X163Y177_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X163Y177_CO5),
.O6(CLBLM_R_X103Y177_SLICE_X163Y177_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y177_SLICE_X163Y177_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X163Y177_BO5),
.O6(CLBLM_R_X103Y177_SLICE_X163Y177_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ffffaaaaffff)
  ) CLBLM_R_X103Y177_SLICE_X163Y177_ALUT (
.I0(CLBLM_L_X12Y110_SLICE_X16Y110_AQ),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_L_X12Y111_SLICE_X16Y111_AQ),
.I4(RIOB33_X105Y143_IOB_X1Y143_I),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X163Y177_AO5),
.O6(CLBLM_R_X103Y177_SLICE_X163Y177_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFGCTRL" *)
  BUFGCTRL #(
    .INIT_OUT(0),
    .IS_CE0_INVERTED(0),
    .IS_CE1_INVERTED(1),
    .IS_IGNORE0_INVERTED(1),
    .IS_IGNORE1_INVERTED(0),
    .IS_S0_INVERTED(0),
    .IS_S1_INVERTED(1),
    .PRESELECT_I0("TRUE"),
    .PRESELECT_I1("FALSE")
  ) CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_BUFGCTRL (
.CE0(1'b1),
.CE1(1'b1),
.I0(LIOB33_X0Y77_IOB_X0Y78_I),
.I1(1'b1),
.IGNORE0(1'b1),
.IGNORE1(1'b1),
.O(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.S0(1'b1),
.S1(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFHCE" *)
  BUFHCE #(
    .CE_TYPE("SYNC"),
    .INIT_OUT(0),
    .IS_CE_INVERTED(0)
  ) CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_BUFHCE (
.CE(1'b1),
.I(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.O(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y51_IOB_X0Y51_IBUF (
.I(LIOB33_X0Y51_IOB_X0Y51_IPAD),
.O(LIOB33_X0Y51_IOB_X0Y51_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y51_IOB_X0Y52_IBUF (
.I(LIOB33_X0Y51_IOB_X0Y52_IPAD),
.O(LIOB33_X0Y51_IOB_X0Y52_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y53_IOB_X0Y53_IBUF (
.I(LIOB33_X0Y53_IOB_X0Y53_IPAD),
.O(LIOB33_X0Y53_IOB_X0Y53_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y53_IOB_X0Y54_IBUF (
.I(LIOB33_X0Y53_IOB_X0Y54_IPAD),
.O(LIOB33_X0Y53_IOB_X0Y54_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y55_IOB_X0Y55_IBUF (
.I(LIOB33_X0Y55_IOB_X0Y55_IPAD),
.O(LIOB33_X0Y55_IOB_X0Y55_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y55_IOB_X0Y56_IBUF (
.I(LIOB33_X0Y55_IOB_X0Y56_IPAD),
.O(LIOB33_X0Y55_IOB_X0Y56_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y57_IOB_X0Y57_IBUF (
.I(LIOB33_X0Y57_IOB_X0Y57_IPAD),
.O(LIOB33_X0Y57_IOB_X0Y57_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y57_IOB_X0Y58_IBUF (
.I(LIOB33_X0Y57_IOB_X0Y58_IPAD),
.O(LIOB33_X0Y57_IOB_X0Y58_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y59_IOB_X0Y59_IBUF (
.I(LIOB33_X0Y59_IOB_X0Y59_IPAD),
.O(LIOB33_X0Y59_IOB_X0Y59_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y59_IOB_X0Y60_IBUF (
.I(LIOB33_X0Y59_IOB_X0Y60_IPAD),
.O(LIOB33_X0Y59_IOB_X0Y60_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y61_IOB_X0Y61_IBUF (
.I(LIOB33_X0Y61_IOB_X0Y61_IPAD),
.O(LIOB33_X0Y61_IOB_X0Y61_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y61_IOB_X0Y62_IBUF (
.I(LIOB33_X0Y61_IOB_X0Y62_IPAD),
.O(LIOB33_X0Y61_IOB_X0Y62_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y63_IOB_X0Y63_IBUF (
.I(LIOB33_X0Y63_IOB_X0Y63_IPAD),
.O(LIOB33_X0Y63_IOB_X0Y63_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y63_IOB_X0Y64_IBUF (
.I(LIOB33_X0Y63_IOB_X0Y64_IPAD),
.O(LIOB33_X0Y63_IOB_X0Y64_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y65_IOB_X0Y65_IBUF (
.I(LIOB33_X0Y65_IOB_X0Y65_IPAD),
.O(LIOB33_X0Y65_IOB_X0Y65_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y65_IOB_X0Y66_IBUF (
.I(LIOB33_X0Y65_IOB_X0Y66_IPAD),
.O(LIOB33_X0Y65_IOB_X0Y66_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y67_IOB_X0Y67_IBUF (
.I(LIOB33_X0Y67_IOB_X0Y67_IPAD),
.O(LIOB33_X0Y67_IOB_X0Y67_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y67_IOB_X0Y68_IBUF (
.I(LIOB33_X0Y67_IOB_X0Y68_IPAD),
.O(LIOB33_X0Y67_IOB_X0Y68_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y69_IOB_X0Y69_IBUF (
.I(LIOB33_X0Y69_IOB_X0Y69_IPAD),
.O(LIOB33_X0Y69_IOB_X0Y69_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y69_IOB_X0Y70_IBUF (
.I(LIOB33_X0Y69_IOB_X0Y70_IPAD),
.O(LIOB33_X0Y69_IOB_X0Y70_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y71_IOB_X0Y71_IBUF (
.I(LIOB33_X0Y71_IOB_X0Y71_IPAD),
.O(LIOB33_X0Y71_IOB_X0Y71_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y71_IOB_X0Y72_IBUF (
.I(LIOB33_X0Y71_IOB_X0Y72_IPAD),
.O(LIOB33_X0Y71_IOB_X0Y72_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y73_IOB_X0Y73_IBUF (
.I(LIOB33_X0Y73_IOB_X0Y73_IPAD),
.O(LIOB33_X0Y73_IOB_X0Y73_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y73_IOB_X0Y74_IBUF (
.I(LIOB33_X0Y73_IOB_X0Y74_IPAD),
.O(LIOB33_X0Y73_IOB_X0Y74_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y75_IOB_X0Y75_IBUF (
.I(LIOB33_X0Y75_IOB_X0Y75_IPAD),
.O(LIOB33_X0Y75_IOB_X0Y75_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y75_IOB_X0Y76_IBUF (
.I(LIOB33_X0Y75_IOB_X0Y76_IPAD),
.O(LIOB33_X0Y75_IOB_X0Y76_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y77_IOB_X0Y77_IBUF (
.I(LIOB33_X0Y77_IOB_X0Y77_IPAD),
.O(LIOB33_X0Y77_IOB_X0Y77_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y77_IOB_X0Y78_IBUF (
.I(LIOB33_X0Y77_IOB_X0Y78_IPAD),
.O(LIOB33_X0Y77_IOB_X0Y78_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y79_IOB_X0Y79_IBUF (
.I(LIOB33_X0Y79_IOB_X0Y79_IPAD),
.O(LIOB33_X0Y79_IOB_X0Y79_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y79_IOB_X0Y80_OBUF (
.I(CLBLL_L_X2Y106_SLICE_X0Y106_AO6),
.O(LIOB33_X0Y79_IOB_X0Y80_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y101_IOB_X0Y101_OBUF (
.I(CLBLL_L_X2Y107_SLICE_X0Y107_AO6),
.O(LIOB33_X0Y101_IOB_X0Y101_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y101_IOB_X0Y102_OBUF (
.I(CLBLL_L_X2Y106_SLICE_X0Y106_BO5),
.O(LIOB33_X0Y101_IOB_X0Y102_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y103_IOB_X0Y103_OBUF (
.I(CLBLM_R_X3Y107_SLICE_X3Y107_BO6),
.O(LIOB33_X0Y103_IOB_X0Y103_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y103_IOB_X0Y104_OBUF (
.I(CLBLL_L_X2Y106_SLICE_X0Y106_CO6),
.O(LIOB33_X0Y103_IOB_X0Y104_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y105_IOB_X0Y105_OBUF (
.I(CLBLL_L_X2Y106_SLICE_X0Y106_CO5),
.O(LIOB33_X0Y105_IOB_X0Y105_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y105_IOB_X0Y106_OBUF (
.I(CLBLL_L_X2Y106_SLICE_X0Y106_AO5),
.O(LIOB33_X0Y105_IOB_X0Y106_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y107_IOB_X0Y107_OBUF (
.I(CLBLM_R_X3Y106_SLICE_X2Y106_BO6),
.O(LIOB33_X0Y107_IOB_X0Y107_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y107_IOB_X0Y108_OBUF (
.I(CLBLL_L_X2Y107_SLICE_X0Y107_AO5),
.O(LIOB33_X0Y107_IOB_X0Y108_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y109_IOB_X0Y109_OBUF (
.I(CLBLL_L_X2Y107_SLICE_X1Y107_AO5),
.O(LIOB33_X0Y109_IOB_X0Y109_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y109_IOB_X0Y110_OBUF (
.I(CLBLM_R_X3Y106_SLICE_X2Y106_AO6),
.O(LIOB33_X0Y109_IOB_X0Y110_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y111_IOB_X0Y111_OBUF (
.I(1'b0),
.O(LIOB33_X0Y111_IOB_X0Y111_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y111_IOB_X0Y112_OBUF (
.I(CLBLM_R_X11Y110_SLICE_X14Y110_D5Q),
.O(LIOB33_X0Y111_IOB_X0Y112_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y113_IOB_X0Y113_OBUF (
.I(RIOB33_X105Y121_IOB_X1Y121_I),
.O(LIOB33_X0Y113_IOB_X0Y113_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y113_IOB_X0Y114_OBUF (
.I(CLBLM_R_X7Y113_SLICE_X8Y113_CQ),
.O(LIOB33_X0Y113_IOB_X0Y114_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y115_IOB_X0Y115_OBUF (
.I(CLBLM_R_X11Y110_SLICE_X14Y110_DQ),
.O(LIOB33_X0Y115_IOB_X0Y115_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y115_IOB_X0Y116_OBUF (
.I(CLBLM_R_X11Y118_SLICE_X15Y118_AQ),
.O(LIOB33_X0Y115_IOB_X0Y116_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y117_IOB_X0Y117_OBUF (
.I(CLBLL_L_X4Y116_SLICE_X5Y116_BQ),
.O(LIOB33_X0Y117_IOB_X0Y117_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y117_IOB_X0Y118_OBUF (
.I(CLBLM_R_X5Y114_SLICE_X7Y114_CQ),
.O(LIOB33_X0Y117_IOB_X0Y118_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y119_IOB_X0Y119_OBUF (
.I(CLBLM_L_X10Y111_SLICE_X13Y111_CQ),
.O(LIOB33_X0Y119_IOB_X0Y119_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y119_IOB_X0Y120_OBUF (
.I(CLBLM_R_X13Y112_SLICE_X18Y112_AQ),
.O(LIOB33_X0Y119_IOB_X0Y120_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y121_IOB_X0Y121_OBUF (
.I(CLBLM_R_X11Y118_SLICE_X15Y118_A5Q),
.O(LIOB33_X0Y121_IOB_X0Y121_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y121_IOB_X0Y122_OBUF (
.I(CLBLM_R_X5Y116_SLICE_X7Y116_A5Q),
.O(LIOB33_X0Y121_IOB_X0Y122_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y123_IOB_X0Y123_OBUF (
.I(CLBLM_R_X7Y113_SLICE_X8Y113_C5Q),
.O(LIOB33_X0Y123_IOB_X0Y123_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y123_IOB_X0Y124_OBUF (
.I(CLBLM_R_X5Y114_SLICE_X7Y114_C5Q),
.O(LIOB33_X0Y123_IOB_X0Y124_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y125_IOB_X0Y125_OBUF (
.I(CLBLM_R_X11Y115_SLICE_X15Y115_B5Q),
.O(LIOB33_X0Y125_IOB_X0Y125_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y125_IOB_X0Y126_OBUF (
.I(CLBLL_L_X4Y117_SLICE_X4Y117_CQ),
.O(LIOB33_X0Y125_IOB_X0Y126_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y127_IOB_X0Y127_OBUF (
.I(CLBLL_L_X4Y113_SLICE_X4Y113_BQ),
.O(LIOB33_X0Y127_IOB_X0Y127_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y127_IOB_X0Y128_OBUF (
.I(CLBLM_R_X3Y115_SLICE_X2Y115_AQ),
.O(LIOB33_X0Y127_IOB_X0Y128_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y129_IOB_X0Y129_OBUF (
.I(CLBLM_R_X5Y109_SLICE_X6Y109_CQ),
.O(LIOB33_X0Y129_IOB_X0Y129_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y129_IOB_X0Y130_OBUF (
.I(CLBLL_L_X52Y126_SLICE_X78Y126_AO6),
.O(LIOB33_X0Y129_IOB_X0Y130_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y131_IOB_X0Y131_OBUF (
.I(CLBLM_L_X8Y119_SLICE_X10Y119_AO5),
.O(LIOB33_X0Y131_IOB_X0Y131_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y131_IOB_X0Y132_OBUF (
.I(CLBLM_L_X8Y119_SLICE_X10Y119_AQ),
.O(LIOB33_X0Y131_IOB_X0Y132_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y133_IOB_X0Y133_OBUF (
.I(CLBLL_L_X4Y118_SLICE_X4Y118_A5Q),
.O(LIOB33_X0Y133_IOB_X0Y133_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y133_IOB_X0Y134_OBUF (
.I(CLBLL_L_X4Y116_SLICE_X5Y116_AQ),
.O(LIOB33_X0Y133_IOB_X0Y134_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y135_IOB_X0Y135_OBUF (
.I(CLBLL_L_X4Y118_SLICE_X4Y118_AQ),
.O(LIOB33_X0Y135_IOB_X0Y135_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y135_IOB_X0Y136_OBUF (
.I(CLBLL_L_X4Y117_SLICE_X4Y117_DQ),
.O(LIOB33_X0Y135_IOB_X0Y136_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y137_IOB_X0Y137_OBUF (
.I(CLBLL_L_X4Y117_SLICE_X4Y117_AQ),
.O(LIOB33_X0Y137_IOB_X0Y137_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y137_IOB_X0Y138_OBUF (
.I(CLBLL_L_X4Y117_SLICE_X5Y117_AQ),
.O(LIOB33_X0Y137_IOB_X0Y138_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y139_IOB_X0Y139_OBUF (
.I(CLBLL_L_X4Y118_SLICE_X4Y118_BQ),
.O(LIOB33_X0Y139_IOB_X0Y139_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y139_IOB_X0Y140_OBUF (
.I(CLBLL_L_X4Y116_SLICE_X4Y116_AQ),
.O(LIOB33_X0Y139_IOB_X0Y140_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y141_IOB_X0Y141_OBUF (
.I(CLBLL_L_X4Y117_SLICE_X4Y117_BQ),
.O(LIOB33_X0Y141_IOB_X0Y141_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y141_IOB_X0Y142_OBUF (
.I(LIOB33_X0Y53_IOB_X0Y54_I),
.O(LIOB33_X0Y141_IOB_X0Y142_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y143_IOB_X0Y143_OBUF (
.I(LIOB33_X0Y55_IOB_X0Y55_I),
.O(LIOB33_X0Y143_IOB_X0Y143_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y145_IOB_X0Y145_OBUF (
.I(LIOB33_X0Y57_IOB_X0Y58_I),
.O(LIOB33_X0Y145_IOB_X0Y145_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y145_IOB_X0Y146_OBUF (
.I(LIOB33_X0Y59_IOB_X0Y59_I),
.O(LIOB33_X0Y145_IOB_X0Y146_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y147_IOB_X0Y147_OBUF (
.I(LIOB33_X0Y71_IOB_X0Y71_I),
.O(LIOB33_X0Y147_IOB_X0Y147_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y147_IOB_X0Y148_OBUF (
.I(LIOB33_X0Y61_IOB_X0Y61_I),
.O(LIOB33_X0Y147_IOB_X0Y148_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y151_IOB_X0Y151_OBUF (
.I(LIOB33_X0Y65_IOB_X0Y65_I),
.O(LIOB33_X0Y151_IOB_X0Y151_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y151_IOB_X0Y152_OBUF (
.I(LIOB33_X0Y65_IOB_X0Y66_I),
.O(LIOB33_X0Y151_IOB_X0Y152_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y153_IOB_X0Y153_OBUF (
.I(LIOB33_X0Y67_IOB_X0Y67_I),
.O(LIOB33_X0Y153_IOB_X0Y153_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y153_IOB_X0Y154_OBUF (
.I(LIOB33_X0Y67_IOB_X0Y68_I),
.O(LIOB33_X0Y153_IOB_X0Y154_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y155_IOB_X0Y155_OBUF (
.I(LIOB33_X0Y69_IOB_X0Y70_I),
.O(LIOB33_X0Y155_IOB_X0Y155_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y155_IOB_X0Y156_OBUF (
.I(RIOB33_X105Y105_IOB_X1Y106_I),
.O(LIOB33_X0Y155_IOB_X0Y156_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y157_IOB_X0Y157_OBUF (
.I(RIOB33_X105Y115_IOB_X1Y115_I),
.O(LIOB33_X0Y157_IOB_X0Y157_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y157_IOB_X0Y158_OBUF (
.I(RIOB33_X105Y115_IOB_X1Y116_I),
.O(LIOB33_X0Y157_IOB_X0Y158_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y159_IOB_X0Y159_OBUF (
.I(RIOB33_X105Y117_IOB_X1Y117_I),
.O(LIOB33_X0Y159_IOB_X0Y159_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y159_IOB_X0Y160_OBUF (
.I(RIOB33_X105Y107_IOB_X1Y107_I),
.O(LIOB33_X0Y159_IOB_X0Y160_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y161_IOB_X0Y161_OBUF (
.I(RIOB33_X105Y107_IOB_X1Y108_I),
.O(LIOB33_X0Y161_IOB_X0Y161_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y161_IOB_X0Y162_OBUF (
.I(RIOB33_X105Y109_IOB_X1Y109_I),
.O(LIOB33_X0Y161_IOB_X0Y162_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y163_IOB_X0Y163_OBUF (
.I(RIOB33_X105Y109_IOB_X1Y110_I),
.O(LIOB33_X0Y163_IOB_X0Y163_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y163_IOB_X0Y164_OBUF (
.I(RIOB33_X105Y111_IOB_X1Y111_I),
.O(LIOB33_X0Y163_IOB_X0Y164_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y165_IOB_X0Y165_OBUF (
.I(RIOB33_X105Y111_IOB_X1Y112_I),
.O(LIOB33_X0Y165_IOB_X0Y165_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y165_IOB_X0Y166_OBUF (
.I(RIOB33_X105Y113_IOB_X1Y113_I),
.O(LIOB33_X0Y165_IOB_X0Y166_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y167_IOB_X0Y167_OBUF (
.I(RIOB33_X105Y113_IOB_X1Y114_I),
.O(LIOB33_X0Y167_IOB_X0Y167_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y167_IOB_X0Y168_OBUF (
.I(RIOB33_X105Y123_IOB_X1Y123_I),
.O(LIOB33_X0Y167_IOB_X0Y168_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y169_IOB_X0Y169_OBUF (
.I(RIOB33_X105Y121_IOB_X1Y122_I),
.O(LIOB33_X0Y169_IOB_X0Y169_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y169_IOB_X0Y170_OBUF (
.I(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.O(LIOB33_X0Y169_IOB_X0Y170_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y171_IOB_X0Y171_OBUF (
.I(LIOB33_SING_X0Y50_IOB_X0Y50_I),
.O(LIOB33_X0Y171_IOB_X0Y171_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y171_IOB_X0Y172_OBUF (
.I(CLBLM_R_X103Y138_SLICE_X163Y138_AO6),
.O(LIOB33_X0Y171_IOB_X0Y172_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y173_IOB_X0Y173_OBUF (
.I(CLBLM_R_X7Y132_SLICE_X9Y132_AO5),
.O(LIOB33_X0Y173_IOB_X0Y173_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y173_IOB_X0Y174_OBUF (
.I(CLBLM_L_X10Y148_SLICE_X12Y148_AO6),
.O(LIOB33_X0Y173_IOB_X0Y174_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y175_IOB_X0Y175_OBUF (
.I(RIOB33_X105Y127_IOB_X1Y127_I),
.O(LIOB33_X0Y175_IOB_X0Y175_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y175_IOB_X0Y176_OBUF (
.I(RIOB33_X105Y127_IOB_X1Y128_I),
.O(LIOB33_X0Y175_IOB_X0Y176_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y177_IOB_X0Y177_OBUF (
.I(RIOB33_X105Y129_IOB_X1Y129_I),
.O(LIOB33_X0Y177_IOB_X0Y177_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y177_IOB_X0Y178_OBUF (
.I(RIOB33_X105Y129_IOB_X1Y130_I),
.O(LIOB33_X0Y177_IOB_X0Y178_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y179_IOB_X0Y179_OBUF (
.I(RIOB33_X105Y131_IOB_X1Y131_I),
.O(LIOB33_X0Y179_IOB_X0Y179_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y179_IOB_X0Y180_OBUF (
.I(RIOB33_X105Y131_IOB_X1Y132_I),
.O(LIOB33_X0Y179_IOB_X0Y180_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y181_IOB_X0Y181_OBUF (
.I(RIOB33_X105Y133_IOB_X1Y133_I),
.O(LIOB33_X0Y181_IOB_X0Y181_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y181_IOB_X0Y182_OBUF (
.I(RIOB33_X105Y133_IOB_X1Y134_I),
.O(LIOB33_X0Y181_IOB_X0Y182_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y183_IOB_X0Y183_OBUF (
.I(RIOB33_X105Y135_IOB_X1Y135_I),
.O(LIOB33_X0Y183_IOB_X0Y183_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y183_IOB_X0Y184_OBUF (
.I(RIOB33_X105Y135_IOB_X1Y136_I),
.O(LIOB33_X0Y183_IOB_X0Y184_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y185_IOB_X0Y185_OBUF (
.I(RIOB33_X105Y137_IOB_X1Y137_I),
.O(LIOB33_X0Y185_IOB_X0Y185_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y185_IOB_X0Y186_OBUF (
.I(RIOB33_X105Y143_IOB_X1Y143_I),
.O(LIOB33_X0Y185_IOB_X0Y186_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y187_IOB_X0Y187_OBUF (
.I(RIOB33_X105Y143_IOB_X1Y144_I),
.O(LIOB33_X0Y187_IOB_X0Y187_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y187_IOB_X0Y188_OBUF (
.I(RIOB33_X105Y145_IOB_X1Y145_I),
.O(LIOB33_X0Y187_IOB_X0Y188_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y189_IOB_X0Y189_OBUF (
.I(RIOB33_X105Y145_IOB_X1Y146_I),
.O(LIOB33_X0Y189_IOB_X0Y189_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y189_IOB_X0Y190_OBUF (
.I(RIOB33_X105Y147_IOB_X1Y147_I),
.O(LIOB33_X0Y189_IOB_X0Y190_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y191_IOB_X0Y191_OBUF (
.I(RIOB33_X105Y147_IOB_X1Y148_I),
.O(LIOB33_X0Y191_IOB_X0Y191_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y191_IOB_X0Y192_OBUF (
.I(LIOB33_X0Y51_IOB_X0Y52_I),
.O(LIOB33_X0Y191_IOB_X0Y192_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y193_IOB_X0Y193_OBUF (
.I(LIOB33_X0Y55_IOB_X0Y56_I),
.O(LIOB33_X0Y193_IOB_X0Y193_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y193_IOB_X0Y194_OBUF (
.I(LIOB33_X0Y59_IOB_X0Y60_I),
.O(LIOB33_X0Y193_IOB_X0Y194_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y195_IOB_X0Y195_OBUF (
.I(LIOB33_X0Y63_IOB_X0Y64_I),
.O(LIOB33_X0Y195_IOB_X0Y195_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y195_IOB_X0Y196_OBUF (
.I(LIOB33_X0Y69_IOB_X0Y69_I),
.O(LIOB33_X0Y195_IOB_X0Y196_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y197_IOB_X0Y197_OBUF (
.I(LIOB33_X0Y71_IOB_X0Y72_I),
.O(LIOB33_X0Y197_IOB_X0Y197_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y197_IOB_X0Y198_OBUF (
.I(LIOB33_X0Y73_IOB_X0Y73_I),
.O(LIOB33_X0Y197_IOB_X0Y198_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_SING_X0Y50_IOB_X0Y50_IBUF (
.I(LIOB33_SING_X0Y50_IOB_X0Y50_IPAD),
.O(LIOB33_SING_X0Y50_IOB_X0Y50_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y100_IOB_X0Y100_OBUF (
.I(CLBLL_L_X2Y106_SLICE_X0Y106_BO6),
.O(LIOB33_SING_X0Y100_IOB_X0Y100_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y149_IOB_X0Y149_OBUF (
.I(LIOB33_X0Y61_IOB_X0Y62_I),
.O(LIOB33_SING_X0Y149_IOB_X0Y149_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y150_IOB_X0Y150_OBUF (
.I(LIOB33_X0Y63_IOB_X0Y63_I),
.O(LIOB33_SING_X0Y150_IOB_X0Y150_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y199_IOB_X0Y199_OBUF (
.I(LIOB33_X0Y73_IOB_X0Y74_I),
.O(LIOB33_SING_X0Y199_IOB_X0Y199_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y101_IOB_X1Y101_IBUF (
.I(RIOB33_X105Y101_IOB_X1Y101_IPAD),
.O(RIOB33_X105Y101_IOB_X1Y101_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y101_IOB_X1Y102_IBUF (
.I(RIOB33_X105Y101_IOB_X1Y102_IPAD),
.O(RIOB33_X105Y101_IOB_X1Y102_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y103_IOB_X1Y103_IBUF (
.I(RIOB33_X105Y103_IOB_X1Y103_IPAD),
.O(RIOB33_X105Y103_IOB_X1Y103_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y103_IOB_X1Y104_IBUF (
.I(RIOB33_X105Y103_IOB_X1Y104_IPAD),
.O(RIOB33_X105Y103_IOB_X1Y104_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y105_IOB_X1Y105_IBUF (
.I(RIOB33_X105Y105_IOB_X1Y105_IPAD),
.O(RIOB33_X105Y105_IOB_X1Y105_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y105_IOB_X1Y106_IBUF (
.I(RIOB33_X105Y105_IOB_X1Y106_IPAD),
.O(RIOB33_X105Y105_IOB_X1Y106_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y107_IOB_X1Y107_IBUF (
.I(RIOB33_X105Y107_IOB_X1Y107_IPAD),
.O(RIOB33_X105Y107_IOB_X1Y107_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y107_IOB_X1Y108_IBUF (
.I(RIOB33_X105Y107_IOB_X1Y108_IPAD),
.O(RIOB33_X105Y107_IOB_X1Y108_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y109_IOB_X1Y109_IBUF (
.I(RIOB33_X105Y109_IOB_X1Y109_IPAD),
.O(RIOB33_X105Y109_IOB_X1Y109_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y109_IOB_X1Y110_IBUF (
.I(RIOB33_X105Y109_IOB_X1Y110_IPAD),
.O(RIOB33_X105Y109_IOB_X1Y110_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y111_IOB_X1Y111_IBUF (
.I(RIOB33_X105Y111_IOB_X1Y111_IPAD),
.O(RIOB33_X105Y111_IOB_X1Y111_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y111_IOB_X1Y112_IBUF (
.I(RIOB33_X105Y111_IOB_X1Y112_IPAD),
.O(RIOB33_X105Y111_IOB_X1Y112_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y113_IOB_X1Y113_IBUF (
.I(RIOB33_X105Y113_IOB_X1Y113_IPAD),
.O(RIOB33_X105Y113_IOB_X1Y113_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y113_IOB_X1Y114_IBUF (
.I(RIOB33_X105Y113_IOB_X1Y114_IPAD),
.O(RIOB33_X105Y113_IOB_X1Y114_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y115_IOB_X1Y115_IBUF (
.I(RIOB33_X105Y115_IOB_X1Y115_IPAD),
.O(RIOB33_X105Y115_IOB_X1Y115_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y115_IOB_X1Y116_IBUF (
.I(RIOB33_X105Y115_IOB_X1Y116_IPAD),
.O(RIOB33_X105Y115_IOB_X1Y116_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y117_IOB_X1Y117_IBUF (
.I(RIOB33_X105Y117_IOB_X1Y117_IPAD),
.O(RIOB33_X105Y117_IOB_X1Y117_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y117_IOB_X1Y118_IBUF (
.I(RIOB33_X105Y117_IOB_X1Y118_IPAD),
.O(RIOB33_X105Y117_IOB_X1Y118_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y119_IOB_X1Y119_IBUF (
.I(RIOB33_X105Y119_IOB_X1Y119_IPAD),
.O(RIOB33_X105Y119_IOB_X1Y119_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y119_IOB_X1Y120_IBUF (
.I(RIOB33_X105Y119_IOB_X1Y120_IPAD),
.O(RIOB33_X105Y119_IOB_X1Y120_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y121_IOB_X1Y121_IBUF (
.I(RIOB33_X105Y121_IOB_X1Y121_IPAD),
.O(RIOB33_X105Y121_IOB_X1Y121_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y121_IOB_X1Y122_IBUF (
.I(RIOB33_X105Y121_IOB_X1Y122_IPAD),
.O(RIOB33_X105Y121_IOB_X1Y122_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y123_IOB_X1Y123_IBUF (
.I(RIOB33_X105Y123_IOB_X1Y123_IPAD),
.O(RIOB33_X105Y123_IOB_X1Y123_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y123_IOB_X1Y124_IBUF (
.I(RIOB33_X105Y123_IOB_X1Y124_IPAD),
.O(RIOB33_X105Y123_IOB_X1Y124_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y125_IOB_X1Y125_IBUF (
.I(RIOB33_X105Y125_IOB_X1Y125_IPAD),
.O(RIOB33_X105Y125_IOB_X1Y125_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y125_IOB_X1Y126_IBUF (
.I(RIOB33_X105Y125_IOB_X1Y126_IPAD),
.O(RIOB33_X105Y125_IOB_X1Y126_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y127_IOB_X1Y127_IBUF (
.I(RIOB33_X105Y127_IOB_X1Y127_IPAD),
.O(RIOB33_X105Y127_IOB_X1Y127_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y127_IOB_X1Y128_IBUF (
.I(RIOB33_X105Y127_IOB_X1Y128_IPAD),
.O(RIOB33_X105Y127_IOB_X1Y128_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y129_IOB_X1Y129_IBUF (
.I(RIOB33_X105Y129_IOB_X1Y129_IPAD),
.O(RIOB33_X105Y129_IOB_X1Y129_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y129_IOB_X1Y130_IBUF (
.I(RIOB33_X105Y129_IOB_X1Y130_IPAD),
.O(RIOB33_X105Y129_IOB_X1Y130_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y131_IOB_X1Y131_IBUF (
.I(RIOB33_X105Y131_IOB_X1Y131_IPAD),
.O(RIOB33_X105Y131_IOB_X1Y131_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y131_IOB_X1Y132_IBUF (
.I(RIOB33_X105Y131_IOB_X1Y132_IPAD),
.O(RIOB33_X105Y131_IOB_X1Y132_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y133_IOB_X1Y133_IBUF (
.I(RIOB33_X105Y133_IOB_X1Y133_IPAD),
.O(RIOB33_X105Y133_IOB_X1Y133_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y133_IOB_X1Y134_IBUF (
.I(RIOB33_X105Y133_IOB_X1Y134_IPAD),
.O(RIOB33_X105Y133_IOB_X1Y134_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y135_IOB_X1Y135_IBUF (
.I(RIOB33_X105Y135_IOB_X1Y135_IPAD),
.O(RIOB33_X105Y135_IOB_X1Y135_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y135_IOB_X1Y136_IBUF (
.I(RIOB33_X105Y135_IOB_X1Y136_IPAD),
.O(RIOB33_X105Y135_IOB_X1Y136_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y137_IOB_X1Y137_IBUF (
.I(RIOB33_X105Y137_IOB_X1Y137_IPAD),
.O(RIOB33_X105Y137_IOB_X1Y137_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y137_IOB_X1Y138_IBUF (
.I(RIOB33_X105Y137_IOB_X1Y138_IPAD),
.O(RIOB33_X105Y137_IOB_X1Y138_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y139_IOB_X1Y139_IBUF (
.I(RIOB33_X105Y139_IOB_X1Y139_IPAD),
.O(RIOB33_X105Y139_IOB_X1Y139_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y139_IOB_X1Y140_IBUF (
.I(RIOB33_X105Y139_IOB_X1Y140_IPAD),
.O(RIOB33_X105Y139_IOB_X1Y140_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y141_IOB_X1Y141_IBUF (
.I(RIOB33_X105Y141_IOB_X1Y141_IPAD),
.O(RIOB33_X105Y141_IOB_X1Y141_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y141_IOB_X1Y142_IBUF (
.I(RIOB33_X105Y141_IOB_X1Y142_IPAD),
.O(RIOB33_X105Y141_IOB_X1Y142_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y143_IOB_X1Y143_IBUF (
.I(RIOB33_X105Y143_IOB_X1Y143_IPAD),
.O(RIOB33_X105Y143_IOB_X1Y143_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y143_IOB_X1Y144_IBUF (
.I(RIOB33_X105Y143_IOB_X1Y144_IPAD),
.O(RIOB33_X105Y143_IOB_X1Y144_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y145_IOB_X1Y145_IBUF (
.I(RIOB33_X105Y145_IOB_X1Y145_IPAD),
.O(RIOB33_X105Y145_IOB_X1Y145_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y145_IOB_X1Y146_IBUF (
.I(RIOB33_X105Y145_IOB_X1Y146_IPAD),
.O(RIOB33_X105Y145_IOB_X1Y146_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y147_IOB_X1Y147_IBUF (
.I(RIOB33_X105Y147_IOB_X1Y147_IPAD),
.O(RIOB33_X105Y147_IOB_X1Y147_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y147_IOB_X1Y148_IBUF (
.I(RIOB33_X105Y147_IOB_X1Y148_IPAD),
.O(RIOB33_X105Y147_IOB_X1Y148_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y151_IOB_X1Y151_OBUF (
.I(LIOB33_X0Y75_IOB_X0Y76_I),
.O(RIOB33_X105Y151_IOB_X1Y151_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y151_IOB_X1Y152_OBUF (
.I(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.O(RIOB33_X105Y151_IOB_X1Y152_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y153_IOB_X1Y153_OBUF (
.I(RIOB33_X105Y101_IOB_X1Y101_I),
.O(RIOB33_X105Y153_IOB_X1Y153_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y153_IOB_X1Y154_OBUF (
.I(RIOB33_X105Y101_IOB_X1Y102_I),
.O(RIOB33_X105Y153_IOB_X1Y154_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y155_IOB_X1Y155_OBUF (
.I(RIOB33_X105Y103_IOB_X1Y103_I),
.O(RIOB33_X105Y155_IOB_X1Y155_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y155_IOB_X1Y156_OBUF (
.I(RIOB33_X105Y103_IOB_X1Y104_I),
.O(RIOB33_X105Y155_IOB_X1Y156_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y157_IOB_X1Y157_OBUF (
.I(RIOB33_X105Y125_IOB_X1Y126_I),
.O(RIOB33_X105Y157_IOB_X1Y157_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y157_IOB_X1Y158_OBUF (
.I(CLBLM_R_X37Y117_SLICE_X56Y117_AO6),
.O(RIOB33_X105Y157_IOB_X1Y158_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y159_IOB_X1Y159_OBUF (
.I(CLBLM_R_X13Y110_SLICE_X18Y110_DO6),
.O(RIOB33_X105Y159_IOB_X1Y159_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y159_IOB_X1Y160_OBUF (
.I(CLBLM_R_X13Y110_SLICE_X18Y110_DO5),
.O(RIOB33_X105Y159_IOB_X1Y160_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y161_IOB_X1Y161_OBUF (
.I(CLBLM_L_X12Y114_SLICE_X16Y114_DO6),
.O(RIOB33_X105Y161_IOB_X1Y161_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y161_IOB_X1Y162_OBUF (
.I(CLBLM_L_X12Y114_SLICE_X16Y114_DO5),
.O(RIOB33_X105Y161_IOB_X1Y162_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y163_IOB_X1Y163_OBUF (
.I(CLBLM_L_X8Y110_SLICE_X10Y110_CO6),
.O(RIOB33_X105Y163_IOB_X1Y163_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y163_IOB_X1Y164_OBUF (
.I(CLBLM_L_X8Y110_SLICE_X10Y110_CO5),
.O(RIOB33_X105Y163_IOB_X1Y164_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y165_IOB_X1Y165_OBUF (
.I(RIOB33_X105Y125_IOB_X1Y125_I),
.O(RIOB33_X105Y165_IOB_X1Y165_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y165_IOB_X1Y166_OBUF (
.I(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.O(RIOB33_X105Y165_IOB_X1Y166_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y167_IOB_X1Y167_OBUF (
.I(LIOB33_SING_X0Y50_IOB_X0Y50_I),
.O(RIOB33_X105Y167_IOB_X1Y167_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y167_IOB_X1Y168_OBUF (
.I(CLBLM_L_X10Y148_SLICE_X12Y148_AO6),
.O(RIOB33_X105Y167_IOB_X1Y168_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y169_IOB_X1Y169_OBUF (
.I(CLBLM_R_X103Y169_SLICE_X163Y169_AO6),
.O(RIOB33_X105Y169_IOB_X1Y169_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y169_IOB_X1Y170_OBUF (
.I(CLBLM_R_X103Y170_SLICE_X163Y170_AO6),
.O(RIOB33_X105Y169_IOB_X1Y170_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y171_IOB_X1Y171_OBUF (
.I(CLBLM_R_X103Y170_SLICE_X163Y170_AO5),
.O(RIOB33_X105Y171_IOB_X1Y171_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y171_IOB_X1Y172_OBUF (
.I(CLBLM_R_X103Y173_SLICE_X163Y173_AO6),
.O(RIOB33_X105Y171_IOB_X1Y172_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y173_IOB_X1Y173_OBUF (
.I(CLBLM_R_X103Y173_SLICE_X163Y173_AO5),
.O(RIOB33_X105Y173_IOB_X1Y173_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y173_IOB_X1Y174_OBUF (
.I(CLBLM_R_X103Y174_SLICE_X163Y174_AO6),
.O(RIOB33_X105Y173_IOB_X1Y174_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y175_IOB_X1Y175_OBUF (
.I(CLBLM_R_X13Y118_SLICE_X18Y118_AO6),
.O(RIOB33_X105Y175_IOB_X1Y175_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y175_IOB_X1Y176_OBUF (
.I(CLBLM_R_X103Y174_SLICE_X163Y174_AO5),
.O(RIOB33_X105Y175_IOB_X1Y176_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y177_IOB_X1Y177_OBUF (
.I(CLBLM_R_X103Y177_SLICE_X163Y177_AO6),
.O(RIOB33_X105Y177_IOB_X1Y177_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y177_IOB_X1Y178_OBUF (
.I(CLBLM_R_X103Y177_SLICE_X163Y177_AO5),
.O(RIOB33_X105Y177_IOB_X1Y178_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y179_IOB_X1Y179_OBUF (
.I(CLBLM_R_X13Y117_SLICE_X18Y117_AO5),
.O(RIOB33_X105Y179_IOB_X1Y179_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y179_IOB_X1Y180_OBUF (
.I(CLBLM_R_X13Y110_SLICE_X18Y110_DO6),
.O(RIOB33_X105Y179_IOB_X1Y180_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y181_IOB_X1Y181_OBUF (
.I(CLBLM_R_X13Y110_SLICE_X18Y110_DO5),
.O(RIOB33_X105Y181_IOB_X1Y181_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y181_IOB_X1Y182_OBUF (
.I(CLBLM_L_X12Y114_SLICE_X16Y114_DO6),
.O(RIOB33_X105Y181_IOB_X1Y182_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y183_IOB_X1Y183_OBUF (
.I(CLBLM_L_X12Y114_SLICE_X16Y114_DO5),
.O(RIOB33_X105Y183_IOB_X1Y183_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y183_IOB_X1Y184_OBUF (
.I(CLBLM_L_X8Y110_SLICE_X10Y110_CO6),
.O(RIOB33_X105Y183_IOB_X1Y184_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y185_IOB_X1Y185_OBUF (
.I(CLBLM_L_X8Y110_SLICE_X10Y110_CO5),
.O(RIOB33_X105Y185_IOB_X1Y185_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y185_IOB_X1Y186_OBUF (
.I(CLBLM_L_X12Y111_SLICE_X16Y111_AQ),
.O(RIOB33_X105Y185_IOB_X1Y186_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y187_IOB_X1Y187_OBUF (
.I(CLBLM_R_X11Y115_SLICE_X14Y115_BQ),
.O(RIOB33_X105Y187_IOB_X1Y187_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y187_IOB_X1Y188_OBUF (
.I(CLBLM_L_X12Y117_SLICE_X17Y117_AQ),
.O(RIOB33_X105Y187_IOB_X1Y188_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y189_IOB_X1Y189_OBUF (
.I(CLBLM_L_X10Y112_SLICE_X13Y112_AQ),
.O(RIOB33_X105Y189_IOB_X1Y189_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y189_IOB_X1Y190_OBUF (
.I(CLBLM_R_X13Y113_SLICE_X19Y113_AQ),
.O(RIOB33_X105Y189_IOB_X1Y190_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y191_IOB_X1Y191_OBUF (
.I(CLBLM_R_X11Y115_SLICE_X14Y115_AQ),
.O(RIOB33_X105Y191_IOB_X1Y191_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y191_IOB_X1Y192_OBUF (
.I(CLBLM_R_X13Y109_SLICE_X19Y109_AQ),
.O(RIOB33_X105Y191_IOB_X1Y192_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y193_IOB_X1Y193_OBUF (
.I(CLBLM_L_X12Y118_SLICE_X16Y118_AQ),
.O(RIOB33_X105Y193_IOB_X1Y193_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y193_IOB_X1Y194_OBUF (
.I(CLBLM_R_X11Y119_SLICE_X14Y119_AQ),
.O(RIOB33_X105Y193_IOB_X1Y194_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y195_IOB_X1Y195_OBUF (
.I(CLBLM_L_X12Y110_SLICE_X16Y110_AQ),
.O(RIOB33_X105Y195_IOB_X1Y195_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y195_IOB_X1Y196_OBUF (
.I(CLBLM_L_X12Y117_SLICE_X16Y117_AQ),
.O(RIOB33_X105Y195_IOB_X1Y196_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y197_IOB_X1Y197_OBUF (
.I(CLBLL_L_X26Y136_SLICE_X38Y136_AO5),
.O(RIOB33_X105Y197_IOB_X1Y197_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y197_IOB_X1Y198_OBUF (
.I(CLBLL_L_X26Y136_SLICE_X38Y136_AO5),
.O(RIOB33_X105Y197_IOB_X1Y198_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_SING_X105Y100_IOB_X1Y100_IBUF (
.I(RIOB33_SING_X105Y100_IOB_X1Y100_IPAD),
.O(RIOB33_SING_X105Y100_IOB_X1Y100_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_SING_X105Y149_IOB_X1Y149_IBUF (
.I(RIOB33_SING_X105Y149_IOB_X1Y149_IPAD),
.O(RIOB33_SING_X105Y149_IOB_X1Y149_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_SING_X105Y150_IOB_X1Y150_OBUF (
.I(LIOB33_X0Y75_IOB_X0Y75_I),
.O(RIOB33_SING_X105Y150_IOB_X1Y150_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_SING_X105Y199_IOB_X1Y199_OBUF (
.I(CLBLM_R_X11Y119_SLICE_X14Y119_AQ),
.O(RIOB33_SING_X105Y199_IOB_X1Y199_OPAD)
  );
  assign CLBLL_L_X2Y106_SLICE_X0Y106_A = CLBLL_L_X2Y106_SLICE_X0Y106_AO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_B = CLBLL_L_X2Y106_SLICE_X0Y106_BO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_C = CLBLL_L_X2Y106_SLICE_X0Y106_CO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_D = CLBLL_L_X2Y106_SLICE_X0Y106_DO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_AMUX = CLBLL_L_X2Y106_SLICE_X0Y106_AO5;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_BMUX = CLBLL_L_X2Y106_SLICE_X0Y106_BO5;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_CMUX = CLBLL_L_X2Y106_SLICE_X0Y106_CO5;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_A = CLBLL_L_X2Y106_SLICE_X1Y106_AO6;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_B = CLBLL_L_X2Y106_SLICE_X1Y106_BO6;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_C = CLBLL_L_X2Y106_SLICE_X1Y106_CO6;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_D = CLBLL_L_X2Y106_SLICE_X1Y106_DO6;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_A = CLBLL_L_X2Y107_SLICE_X0Y107_AO6;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_B = CLBLL_L_X2Y107_SLICE_X0Y107_BO6;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_C = CLBLL_L_X2Y107_SLICE_X0Y107_CO6;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_D = CLBLL_L_X2Y107_SLICE_X0Y107_DO6;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_AMUX = CLBLL_L_X2Y107_SLICE_X0Y107_AO5;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_A = CLBLL_L_X2Y107_SLICE_X1Y107_AO6;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_B = CLBLL_L_X2Y107_SLICE_X1Y107_BO6;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_C = CLBLL_L_X2Y107_SLICE_X1Y107_CO6;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_D = CLBLL_L_X2Y107_SLICE_X1Y107_DO6;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_AMUX = CLBLL_L_X2Y107_SLICE_X1Y107_AO5;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_A = CLBLL_L_X2Y108_SLICE_X0Y108_AO6;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_B = CLBLL_L_X2Y108_SLICE_X0Y108_BO6;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_C = CLBLL_L_X2Y108_SLICE_X0Y108_CO6;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_D = CLBLL_L_X2Y108_SLICE_X0Y108_DO6;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_A = CLBLL_L_X2Y108_SLICE_X1Y108_AO6;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_B = CLBLL_L_X2Y108_SLICE_X1Y108_BO6;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_C = CLBLL_L_X2Y108_SLICE_X1Y108_CO6;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_D = CLBLL_L_X2Y108_SLICE_X1Y108_DO6;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_AMUX = CLBLL_L_X2Y108_SLICE_X1Y108_AO5;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_BMUX = CLBLL_L_X2Y108_SLICE_X1Y108_BO5;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_CMUX = CLBLL_L_X2Y108_SLICE_X1Y108_CO6;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_A = CLBLL_L_X2Y109_SLICE_X0Y109_AO6;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_B = CLBLL_L_X2Y109_SLICE_X0Y109_BO6;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_C = CLBLL_L_X2Y109_SLICE_X0Y109_CO6;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_D = CLBLL_L_X2Y109_SLICE_X0Y109_DO6;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_AMUX = CLBLL_L_X2Y109_SLICE_X0Y109_AO5;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_BMUX = CLBLL_L_X2Y109_SLICE_X0Y109_BO5;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_CMUX = CLBLL_L_X2Y109_SLICE_X0Y109_CO6;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_A = CLBLL_L_X2Y109_SLICE_X1Y109_AO6;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_B = CLBLL_L_X2Y109_SLICE_X1Y109_BO6;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_C = CLBLL_L_X2Y109_SLICE_X1Y109_CO6;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_D = CLBLL_L_X2Y109_SLICE_X1Y109_DO6;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_BMUX = CLBLL_L_X2Y109_SLICE_X1Y109_BO6;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_DMUX = CLBLL_L_X2Y109_SLICE_X1Y109_DO6;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_A = CLBLL_L_X2Y110_SLICE_X0Y110_AO6;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_B = CLBLL_L_X2Y110_SLICE_X0Y110_BO6;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_C = CLBLL_L_X2Y110_SLICE_X0Y110_CO6;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_D = CLBLL_L_X2Y110_SLICE_X0Y110_DO6;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_AMUX = CLBLL_L_X2Y110_SLICE_X0Y110_AO5;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_BMUX = CLBLL_L_X2Y110_SLICE_X0Y110_BO5;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_CMUX = CLBLL_L_X2Y110_SLICE_X0Y110_CO5;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_A = CLBLL_L_X2Y110_SLICE_X1Y110_AO6;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_B = CLBLL_L_X2Y110_SLICE_X1Y110_BO6;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_C = CLBLL_L_X2Y110_SLICE_X1Y110_CO6;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_D = CLBLL_L_X2Y110_SLICE_X1Y110_DO6;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_AMUX = CLBLL_L_X2Y110_SLICE_X1Y110_AO5;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_CMUX = CLBLL_L_X2Y110_SLICE_X1Y110_CO6;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_A = CLBLL_L_X2Y111_SLICE_X0Y111_AO6;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_B = CLBLL_L_X2Y111_SLICE_X0Y111_BO6;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_C = CLBLL_L_X2Y111_SLICE_X0Y111_CO6;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_D = CLBLL_L_X2Y111_SLICE_X0Y111_DO6;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_BMUX = CLBLL_L_X2Y111_SLICE_X0Y111_BO6;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_A = CLBLL_L_X2Y111_SLICE_X1Y111_AO6;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_B = CLBLL_L_X2Y111_SLICE_X1Y111_BO6;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_C = CLBLL_L_X2Y111_SLICE_X1Y111_CO6;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_D = CLBLL_L_X2Y111_SLICE_X1Y111_DO6;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_AMUX = CLBLL_L_X2Y111_SLICE_X1Y111_AO5;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_BMUX = CLBLL_L_X2Y111_SLICE_X1Y111_BO5;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_A = CLBLL_L_X2Y112_SLICE_X0Y112_AO6;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_B = CLBLL_L_X2Y112_SLICE_X0Y112_BO6;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_C = CLBLL_L_X2Y112_SLICE_X0Y112_CO6;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_D = CLBLL_L_X2Y112_SLICE_X0Y112_DO6;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_AMUX = CLBLL_L_X2Y112_SLICE_X0Y112_AO5;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_A = CLBLL_L_X2Y112_SLICE_X1Y112_AO6;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_B = CLBLL_L_X2Y112_SLICE_X1Y112_BO6;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_C = CLBLL_L_X2Y112_SLICE_X1Y112_CO6;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_D = CLBLL_L_X2Y112_SLICE_X1Y112_DO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_A = CLBLL_L_X2Y113_SLICE_X0Y113_AO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_B = CLBLL_L_X2Y113_SLICE_X0Y113_BO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_C = CLBLL_L_X2Y113_SLICE_X0Y113_CO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_D = CLBLL_L_X2Y113_SLICE_X0Y113_DO6;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_A = CLBLL_L_X2Y113_SLICE_X1Y113_AO6;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_B = CLBLL_L_X2Y113_SLICE_X1Y113_BO6;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_C = CLBLL_L_X2Y113_SLICE_X1Y113_CO6;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_D = CLBLL_L_X2Y113_SLICE_X1Y113_DO6;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_AMUX = CLBLL_L_X2Y113_SLICE_X1Y113_AO5;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_CMUX = CLBLL_L_X2Y113_SLICE_X1Y113_CO6;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_A = CLBLL_L_X2Y114_SLICE_X0Y114_AO6;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_B = CLBLL_L_X2Y114_SLICE_X0Y114_BO6;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_C = CLBLL_L_X2Y114_SLICE_X0Y114_CO6;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_D = CLBLL_L_X2Y114_SLICE_X0Y114_DO6;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_AMUX = CLBLL_L_X2Y114_SLICE_X0Y114_AO5;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_A = CLBLL_L_X2Y114_SLICE_X1Y114_AO6;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_B = CLBLL_L_X2Y114_SLICE_X1Y114_BO6;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_C = CLBLL_L_X2Y114_SLICE_X1Y114_CO6;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_D = CLBLL_L_X2Y114_SLICE_X1Y114_DO6;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_AMUX = CLBLL_L_X2Y114_SLICE_X1Y114_AO5;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_A = CLBLL_L_X4Y106_SLICE_X4Y106_AO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_B = CLBLL_L_X4Y106_SLICE_X4Y106_BO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_C = CLBLL_L_X4Y106_SLICE_X4Y106_CO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_D = CLBLL_L_X4Y106_SLICE_X4Y106_DO6;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_A = CLBLL_L_X4Y106_SLICE_X5Y106_AO6;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_B = CLBLL_L_X4Y106_SLICE_X5Y106_BO6;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_C = CLBLL_L_X4Y106_SLICE_X5Y106_CO6;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_D = CLBLL_L_X4Y106_SLICE_X5Y106_DO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_A = CLBLL_L_X4Y107_SLICE_X4Y107_AO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_B = CLBLL_L_X4Y107_SLICE_X4Y107_BO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_C = CLBLL_L_X4Y107_SLICE_X4Y107_CO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_D = CLBLL_L_X4Y107_SLICE_X4Y107_DO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_AMUX = CLBLL_L_X4Y107_SLICE_X4Y107_A5Q;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_BMUX = CLBLL_L_X4Y107_SLICE_X4Y107_BO5;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_A = CLBLL_L_X4Y107_SLICE_X5Y107_AO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_B = CLBLL_L_X4Y107_SLICE_X5Y107_BO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_C = CLBLL_L_X4Y107_SLICE_X5Y107_CO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_D = CLBLL_L_X4Y107_SLICE_X5Y107_DO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_BMUX = CLBLL_L_X4Y107_SLICE_X5Y107_BO5;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_A = CLBLL_L_X4Y108_SLICE_X4Y108_AO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_B = CLBLL_L_X4Y108_SLICE_X4Y108_BO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_C = CLBLL_L_X4Y108_SLICE_X4Y108_CO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_D = CLBLL_L_X4Y108_SLICE_X4Y108_DO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_A = CLBLL_L_X4Y108_SLICE_X5Y108_AO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_B = CLBLL_L_X4Y108_SLICE_X5Y108_BO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_C = CLBLL_L_X4Y108_SLICE_X5Y108_CO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_D = CLBLL_L_X4Y108_SLICE_X5Y108_DO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_AMUX = CLBLL_L_X4Y108_SLICE_X5Y108_AO5;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A = CLBLL_L_X4Y109_SLICE_X4Y109_AO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B = CLBLL_L_X4Y109_SLICE_X4Y109_BO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C = CLBLL_L_X4Y109_SLICE_X4Y109_CO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D = CLBLL_L_X4Y109_SLICE_X4Y109_DO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A = CLBLL_L_X4Y109_SLICE_X5Y109_AO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B = CLBLL_L_X4Y109_SLICE_X5Y109_BO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C = CLBLL_L_X4Y109_SLICE_X5Y109_CO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D = CLBLL_L_X4Y109_SLICE_X5Y109_DO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_BMUX = CLBLL_L_X4Y109_SLICE_X5Y109_BO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_A = CLBLL_L_X4Y110_SLICE_X4Y110_AO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_B = CLBLL_L_X4Y110_SLICE_X4Y110_BO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_C = CLBLL_L_X4Y110_SLICE_X4Y110_CO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_D = CLBLL_L_X4Y110_SLICE_X4Y110_DO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_BMUX = CLBLL_L_X4Y110_SLICE_X4Y110_B5Q;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_CMUX = CLBLL_L_X4Y110_SLICE_X4Y110_C5Q;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_A = CLBLL_L_X4Y110_SLICE_X5Y110_AO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_B = CLBLL_L_X4Y110_SLICE_X5Y110_BO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_C = CLBLL_L_X4Y110_SLICE_X5Y110_CO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_D = CLBLL_L_X4Y110_SLICE_X5Y110_DO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_CMUX = CLBLL_L_X4Y110_SLICE_X5Y110_CO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_DMUX = CLBLL_L_X4Y110_SLICE_X5Y110_DO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_A = CLBLL_L_X4Y111_SLICE_X4Y111_AO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_B = CLBLL_L_X4Y111_SLICE_X4Y111_BO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_C = CLBLL_L_X4Y111_SLICE_X4Y111_CO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_D = CLBLL_L_X4Y111_SLICE_X4Y111_DO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_A = CLBLL_L_X4Y111_SLICE_X5Y111_AO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_B = CLBLL_L_X4Y111_SLICE_X5Y111_BO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_C = CLBLL_L_X4Y111_SLICE_X5Y111_CO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_D = CLBLL_L_X4Y111_SLICE_X5Y111_DO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_A = CLBLL_L_X4Y112_SLICE_X4Y112_AO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_B = CLBLL_L_X4Y112_SLICE_X4Y112_BO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_C = CLBLL_L_X4Y112_SLICE_X4Y112_CO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_D = CLBLL_L_X4Y112_SLICE_X4Y112_DO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_CMUX = CLBLL_L_X4Y112_SLICE_X4Y112_CO5;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_A = CLBLL_L_X4Y112_SLICE_X5Y112_AO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_B = CLBLL_L_X4Y112_SLICE_X5Y112_BO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_C = CLBLL_L_X4Y112_SLICE_X5Y112_CO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_D = CLBLL_L_X4Y112_SLICE_X5Y112_DO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_BMUX = CLBLL_L_X4Y112_SLICE_X5Y112_BO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A = CLBLL_L_X4Y113_SLICE_X4Y113_AO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B = CLBLL_L_X4Y113_SLICE_X4Y113_BO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C = CLBLL_L_X4Y113_SLICE_X4Y113_CO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D = CLBLL_L_X4Y113_SLICE_X4Y113_DO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_CMUX = CLBLL_L_X4Y113_SLICE_X4Y113_CO5;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A = CLBLL_L_X4Y113_SLICE_X5Y113_AO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B = CLBLL_L_X4Y113_SLICE_X5Y113_BO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C = CLBLL_L_X4Y113_SLICE_X5Y113_CO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D = CLBLL_L_X4Y113_SLICE_X5Y113_DO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_BMUX = CLBLL_L_X4Y113_SLICE_X5Y113_B5Q;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_A = CLBLL_L_X4Y114_SLICE_X4Y114_AO6;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_B = CLBLL_L_X4Y114_SLICE_X4Y114_BO6;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_C = CLBLL_L_X4Y114_SLICE_X4Y114_CO6;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_D = CLBLL_L_X4Y114_SLICE_X4Y114_DO6;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_A = CLBLL_L_X4Y114_SLICE_X5Y114_AO6;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_B = CLBLL_L_X4Y114_SLICE_X5Y114_BO6;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_C = CLBLL_L_X4Y114_SLICE_X5Y114_CO6;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_D = CLBLL_L_X4Y114_SLICE_X5Y114_DO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_A = CLBLL_L_X4Y115_SLICE_X4Y115_AO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_B = CLBLL_L_X4Y115_SLICE_X4Y115_BO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_C = CLBLL_L_X4Y115_SLICE_X4Y115_CO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_D = CLBLL_L_X4Y115_SLICE_X4Y115_DO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_A = CLBLL_L_X4Y115_SLICE_X5Y115_AO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_B = CLBLL_L_X4Y115_SLICE_X5Y115_BO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_C = CLBLL_L_X4Y115_SLICE_X5Y115_CO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_D = CLBLL_L_X4Y115_SLICE_X5Y115_DO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_AMUX = CLBLL_L_X4Y115_SLICE_X5Y115_A5Q;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_A = CLBLL_L_X4Y116_SLICE_X4Y116_AO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_B = CLBLL_L_X4Y116_SLICE_X4Y116_BO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_C = CLBLL_L_X4Y116_SLICE_X4Y116_CO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_D = CLBLL_L_X4Y116_SLICE_X4Y116_DO6;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_AMUX = CLBLL_L_X4Y116_SLICE_X4Y116_A5Q;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_BMUX = CLBLL_L_X4Y116_SLICE_X4Y116_BO5;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_A = CLBLL_L_X4Y116_SLICE_X5Y116_AO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_B = CLBLL_L_X4Y116_SLICE_X5Y116_BO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_C = CLBLL_L_X4Y116_SLICE_X5Y116_CO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_D = CLBLL_L_X4Y116_SLICE_X5Y116_DO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_AMUX = CLBLL_L_X4Y116_SLICE_X5Y116_A5Q;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_BMUX = CLBLL_L_X4Y116_SLICE_X5Y116_B5Q;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_A = CLBLL_L_X4Y117_SLICE_X4Y117_AO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_B = CLBLL_L_X4Y117_SLICE_X4Y117_BO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_C = CLBLL_L_X4Y117_SLICE_X4Y117_CO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_D = CLBLL_L_X4Y117_SLICE_X4Y117_DO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_A = CLBLL_L_X4Y117_SLICE_X5Y117_AO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_B = CLBLL_L_X4Y117_SLICE_X5Y117_BO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_C = CLBLL_L_X4Y117_SLICE_X5Y117_CO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_D = CLBLL_L_X4Y117_SLICE_X5Y117_DO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_BMUX = CLBLL_L_X4Y117_SLICE_X5Y117_BO5;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_A = CLBLL_L_X4Y118_SLICE_X4Y118_AO6;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_B = CLBLL_L_X4Y118_SLICE_X4Y118_BO6;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_C = CLBLL_L_X4Y118_SLICE_X4Y118_CO6;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_D = CLBLL_L_X4Y118_SLICE_X4Y118_DO6;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_AMUX = CLBLL_L_X4Y118_SLICE_X4Y118_A5Q;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_CMUX = CLBLL_L_X4Y118_SLICE_X4Y118_CO5;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_DMUX = CLBLL_L_X4Y118_SLICE_X4Y118_DO5;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_A = CLBLL_L_X4Y118_SLICE_X5Y118_AO6;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_B = CLBLL_L_X4Y118_SLICE_X5Y118_BO6;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_C = CLBLL_L_X4Y118_SLICE_X5Y118_CO6;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_D = CLBLL_L_X4Y118_SLICE_X5Y118_DO6;
  assign CLBLL_L_X26Y136_SLICE_X38Y136_A = CLBLL_L_X26Y136_SLICE_X38Y136_AO6;
  assign CLBLL_L_X26Y136_SLICE_X38Y136_B = CLBLL_L_X26Y136_SLICE_X38Y136_BO6;
  assign CLBLL_L_X26Y136_SLICE_X38Y136_C = CLBLL_L_X26Y136_SLICE_X38Y136_CO6;
  assign CLBLL_L_X26Y136_SLICE_X38Y136_D = CLBLL_L_X26Y136_SLICE_X38Y136_DO6;
  assign CLBLL_L_X26Y136_SLICE_X38Y136_AMUX = CLBLL_L_X26Y136_SLICE_X38Y136_AO5;
  assign CLBLL_L_X26Y136_SLICE_X39Y136_A = CLBLL_L_X26Y136_SLICE_X39Y136_AO6;
  assign CLBLL_L_X26Y136_SLICE_X39Y136_B = CLBLL_L_X26Y136_SLICE_X39Y136_BO6;
  assign CLBLL_L_X26Y136_SLICE_X39Y136_C = CLBLL_L_X26Y136_SLICE_X39Y136_CO6;
  assign CLBLL_L_X26Y136_SLICE_X39Y136_D = CLBLL_L_X26Y136_SLICE_X39Y136_DO6;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_A = CLBLL_L_X52Y126_SLICE_X78Y126_AO6;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_B = CLBLL_L_X52Y126_SLICE_X78Y126_BO6;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_C = CLBLL_L_X52Y126_SLICE_X78Y126_CO6;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_D = CLBLL_L_X52Y126_SLICE_X78Y126_DO6;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_A = CLBLL_L_X52Y126_SLICE_X79Y126_AO6;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_B = CLBLL_L_X52Y126_SLICE_X79Y126_BO6;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_C = CLBLL_L_X52Y126_SLICE_X79Y126_CO6;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_D = CLBLL_L_X52Y126_SLICE_X79Y126_DO6;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_A = CLBLM_L_X8Y104_SLICE_X10Y104_AO6;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_B = CLBLM_L_X8Y104_SLICE_X10Y104_BO6;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_C = CLBLM_L_X8Y104_SLICE_X10Y104_CO6;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_D = CLBLM_L_X8Y104_SLICE_X10Y104_DO6;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_A = CLBLM_L_X8Y104_SLICE_X11Y104_AO6;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_B = CLBLM_L_X8Y104_SLICE_X11Y104_BO6;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_C = CLBLM_L_X8Y104_SLICE_X11Y104_CO6;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_D = CLBLM_L_X8Y104_SLICE_X11Y104_DO6;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_AMUX = CLBLM_L_X8Y104_SLICE_X11Y104_AO5;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_A = CLBLM_L_X8Y105_SLICE_X10Y105_AO6;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_B = CLBLM_L_X8Y105_SLICE_X10Y105_BO6;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_C = CLBLM_L_X8Y105_SLICE_X10Y105_CO6;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_D = CLBLM_L_X8Y105_SLICE_X10Y105_DO6;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_A = CLBLM_L_X8Y105_SLICE_X11Y105_AO6;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_B = CLBLM_L_X8Y105_SLICE_X11Y105_BO6;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_C = CLBLM_L_X8Y105_SLICE_X11Y105_CO6;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_D = CLBLM_L_X8Y105_SLICE_X11Y105_DO6;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_CMUX = CLBLM_L_X8Y105_SLICE_X11Y105_CO6;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_A = CLBLM_L_X8Y106_SLICE_X10Y106_AO6;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_B = CLBLM_L_X8Y106_SLICE_X10Y106_BO6;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_C = CLBLM_L_X8Y106_SLICE_X10Y106_CO6;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_D = CLBLM_L_X8Y106_SLICE_X10Y106_DO6;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_DMUX = CLBLM_L_X8Y106_SLICE_X10Y106_DO6;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_A = CLBLM_L_X8Y106_SLICE_X11Y106_AO6;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_B = CLBLM_L_X8Y106_SLICE_X11Y106_BO6;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_C = CLBLM_L_X8Y106_SLICE_X11Y106_CO6;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_D = CLBLM_L_X8Y106_SLICE_X11Y106_DO6;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_AMUX = CLBLM_L_X8Y106_SLICE_X11Y106_A5Q;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_CMUX = CLBLM_L_X8Y106_SLICE_X11Y106_CO5;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_A = CLBLM_L_X8Y107_SLICE_X10Y107_AO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_B = CLBLM_L_X8Y107_SLICE_X10Y107_BO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_C = CLBLM_L_X8Y107_SLICE_X10Y107_CO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_D = CLBLM_L_X8Y107_SLICE_X10Y107_DO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_A = CLBLM_L_X8Y107_SLICE_X11Y107_AO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_B = CLBLM_L_X8Y107_SLICE_X11Y107_BO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_C = CLBLM_L_X8Y107_SLICE_X11Y107_CO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_D = CLBLM_L_X8Y107_SLICE_X11Y107_DO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_AMUX = CLBLM_L_X8Y107_SLICE_X11Y107_A5Q;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_BMUX = CLBLM_L_X8Y107_SLICE_X11Y107_B5Q;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_DMUX = CLBLM_L_X8Y107_SLICE_X11Y107_DO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_A = CLBLM_L_X8Y108_SLICE_X10Y108_AO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_B = CLBLM_L_X8Y108_SLICE_X10Y108_BO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_C = CLBLM_L_X8Y108_SLICE_X10Y108_CO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_D = CLBLM_L_X8Y108_SLICE_X10Y108_DO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_AMUX = CLBLM_L_X8Y108_SLICE_X10Y108_AO5;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_A = CLBLM_L_X8Y108_SLICE_X11Y108_AO6;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_B = CLBLM_L_X8Y108_SLICE_X11Y108_BO6;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_C = CLBLM_L_X8Y108_SLICE_X11Y108_CO6;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_D = CLBLM_L_X8Y108_SLICE_X11Y108_DO6;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_A = CLBLM_L_X8Y109_SLICE_X10Y109_AO6;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_B = CLBLM_L_X8Y109_SLICE_X10Y109_BO6;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_C = CLBLM_L_X8Y109_SLICE_X10Y109_CO6;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_D = CLBLM_L_X8Y109_SLICE_X10Y109_DO6;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_CMUX = CLBLM_L_X8Y109_SLICE_X10Y109_C5Q;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_A = CLBLM_L_X8Y109_SLICE_X11Y109_AO6;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_B = CLBLM_L_X8Y109_SLICE_X11Y109_BO6;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_C = CLBLM_L_X8Y109_SLICE_X11Y109_CO6;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_D = CLBLM_L_X8Y109_SLICE_X11Y109_DO6;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_AMUX = CLBLM_L_X8Y109_SLICE_X11Y109_A5Q;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_A = CLBLM_L_X8Y110_SLICE_X10Y110_AO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_B = CLBLM_L_X8Y110_SLICE_X10Y110_BO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_C = CLBLM_L_X8Y110_SLICE_X10Y110_CO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_D = CLBLM_L_X8Y110_SLICE_X10Y110_DO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_CMUX = CLBLM_L_X8Y110_SLICE_X10Y110_CO5;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_A = CLBLM_L_X8Y110_SLICE_X11Y110_AO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_B = CLBLM_L_X8Y110_SLICE_X11Y110_BO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_C = CLBLM_L_X8Y110_SLICE_X11Y110_CO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_D = CLBLM_L_X8Y110_SLICE_X11Y110_DO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_AMUX = CLBLM_L_X8Y110_SLICE_X11Y110_A5Q;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_BMUX = CLBLM_L_X8Y110_SLICE_X11Y110_BO5;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_A = CLBLM_L_X8Y111_SLICE_X10Y111_AO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_B = CLBLM_L_X8Y111_SLICE_X10Y111_BO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_C = CLBLM_L_X8Y111_SLICE_X10Y111_CO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_D = CLBLM_L_X8Y111_SLICE_X10Y111_DO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_AMUX = CLBLM_L_X8Y111_SLICE_X10Y111_A5Q;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_BMUX = CLBLM_L_X8Y111_SLICE_X10Y111_BO5;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_CMUX = CLBLM_L_X8Y111_SLICE_X10Y111_CO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_DMUX = CLBLM_L_X8Y111_SLICE_X10Y111_DO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_A = CLBLM_L_X8Y111_SLICE_X11Y111_AO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_B = CLBLM_L_X8Y111_SLICE_X11Y111_BO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_C = CLBLM_L_X8Y111_SLICE_X11Y111_CO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_D = CLBLM_L_X8Y111_SLICE_X11Y111_DO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_DMUX = CLBLM_L_X8Y111_SLICE_X11Y111_DO5;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_A = CLBLM_L_X8Y112_SLICE_X10Y112_AO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_B = CLBLM_L_X8Y112_SLICE_X10Y112_BO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_C = CLBLM_L_X8Y112_SLICE_X10Y112_CO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_D = CLBLM_L_X8Y112_SLICE_X10Y112_DO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_AMUX = CLBLM_L_X8Y112_SLICE_X10Y112_A5Q;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_A = CLBLM_L_X8Y112_SLICE_X11Y112_AO6;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_B = CLBLM_L_X8Y112_SLICE_X11Y112_BO6;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_C = CLBLM_L_X8Y112_SLICE_X11Y112_CO6;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_D = CLBLM_L_X8Y112_SLICE_X11Y112_DO6;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_AMUX = CLBLM_L_X8Y112_SLICE_X11Y112_AO5;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_DMUX = CLBLM_L_X8Y112_SLICE_X11Y112_DO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_A = CLBLM_L_X8Y113_SLICE_X10Y113_AO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_B = CLBLM_L_X8Y113_SLICE_X10Y113_BO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_C = CLBLM_L_X8Y113_SLICE_X10Y113_CO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_D = CLBLM_L_X8Y113_SLICE_X10Y113_DO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_DMUX = CLBLM_L_X8Y113_SLICE_X10Y113_D5Q;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_A = CLBLM_L_X8Y113_SLICE_X11Y113_AO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_B = CLBLM_L_X8Y113_SLICE_X11Y113_BO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_C = CLBLM_L_X8Y113_SLICE_X11Y113_CO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_D = CLBLM_L_X8Y113_SLICE_X11Y113_DO6;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_A = CLBLM_L_X8Y114_SLICE_X10Y114_AO6;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_B = CLBLM_L_X8Y114_SLICE_X10Y114_BO6;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_C = CLBLM_L_X8Y114_SLICE_X10Y114_CO6;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_D = CLBLM_L_X8Y114_SLICE_X10Y114_DO6;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_A = CLBLM_L_X8Y114_SLICE_X11Y114_AO6;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_B = CLBLM_L_X8Y114_SLICE_X11Y114_BO6;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_C = CLBLM_L_X8Y114_SLICE_X11Y114_CO6;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_D = CLBLM_L_X8Y114_SLICE_X11Y114_DO6;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_BMUX = CLBLM_L_X8Y114_SLICE_X11Y114_B5Q;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_A = CLBLM_L_X8Y115_SLICE_X10Y115_AO6;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_B = CLBLM_L_X8Y115_SLICE_X10Y115_BO6;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_C = CLBLM_L_X8Y115_SLICE_X10Y115_CO6;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_D = CLBLM_L_X8Y115_SLICE_X10Y115_DO6;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_AMUX = CLBLM_L_X8Y115_SLICE_X10Y115_A5Q;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_A = CLBLM_L_X8Y115_SLICE_X11Y115_AO6;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_B = CLBLM_L_X8Y115_SLICE_X11Y115_BO6;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_C = CLBLM_L_X8Y115_SLICE_X11Y115_CO6;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_D = CLBLM_L_X8Y115_SLICE_X11Y115_DO6;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_A = CLBLM_L_X8Y116_SLICE_X10Y116_AO6;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_B = CLBLM_L_X8Y116_SLICE_X10Y116_BO6;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_C = CLBLM_L_X8Y116_SLICE_X10Y116_CO6;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_D = CLBLM_L_X8Y116_SLICE_X10Y116_DO6;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_A = CLBLM_L_X8Y116_SLICE_X11Y116_AO6;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_B = CLBLM_L_X8Y116_SLICE_X11Y116_BO6;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_C = CLBLM_L_X8Y116_SLICE_X11Y116_CO6;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_D = CLBLM_L_X8Y116_SLICE_X11Y116_DO6;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_A = CLBLM_L_X8Y117_SLICE_X10Y117_AO6;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_B = CLBLM_L_X8Y117_SLICE_X10Y117_BO6;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_C = CLBLM_L_X8Y117_SLICE_X10Y117_CO6;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_D = CLBLM_L_X8Y117_SLICE_X10Y117_DO6;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_A = CLBLM_L_X8Y117_SLICE_X11Y117_AO6;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_B = CLBLM_L_X8Y117_SLICE_X11Y117_BO6;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_C = CLBLM_L_X8Y117_SLICE_X11Y117_CO6;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_D = CLBLM_L_X8Y117_SLICE_X11Y117_DO6;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_A = CLBLM_L_X8Y118_SLICE_X10Y118_AO6;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_B = CLBLM_L_X8Y118_SLICE_X10Y118_BO6;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_C = CLBLM_L_X8Y118_SLICE_X10Y118_CO6;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_D = CLBLM_L_X8Y118_SLICE_X10Y118_DO6;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_CMUX = CLBLM_L_X8Y118_SLICE_X10Y118_CO5;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_DMUX = CLBLM_L_X8Y118_SLICE_X10Y118_DO5;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_A = CLBLM_L_X8Y118_SLICE_X11Y118_AO6;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_B = CLBLM_L_X8Y118_SLICE_X11Y118_BO6;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_C = CLBLM_L_X8Y118_SLICE_X11Y118_CO6;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_D = CLBLM_L_X8Y118_SLICE_X11Y118_DO6;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_A = CLBLM_L_X8Y119_SLICE_X10Y119_AO6;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_B = CLBLM_L_X8Y119_SLICE_X10Y119_BO6;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_C = CLBLM_L_X8Y119_SLICE_X10Y119_CO6;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_D = CLBLM_L_X8Y119_SLICE_X10Y119_DO6;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_AMUX = CLBLM_L_X8Y119_SLICE_X10Y119_AO5;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_A = CLBLM_L_X8Y119_SLICE_X11Y119_AO6;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_B = CLBLM_L_X8Y119_SLICE_X11Y119_BO6;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_C = CLBLM_L_X8Y119_SLICE_X11Y119_CO6;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_D = CLBLM_L_X8Y119_SLICE_X11Y119_DO6;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_A = CLBLM_L_X10Y104_SLICE_X12Y104_AO6;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_B = CLBLM_L_X10Y104_SLICE_X12Y104_BO6;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_C = CLBLM_L_X10Y104_SLICE_X12Y104_CO6;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_D = CLBLM_L_X10Y104_SLICE_X12Y104_DO6;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_A = CLBLM_L_X10Y104_SLICE_X13Y104_AO6;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_B = CLBLM_L_X10Y104_SLICE_X13Y104_BO6;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_C = CLBLM_L_X10Y104_SLICE_X13Y104_CO6;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_D = CLBLM_L_X10Y104_SLICE_X13Y104_DO6;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_A = CLBLM_L_X10Y105_SLICE_X12Y105_AO6;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_B = CLBLM_L_X10Y105_SLICE_X12Y105_BO6;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_C = CLBLM_L_X10Y105_SLICE_X12Y105_CO6;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_D = CLBLM_L_X10Y105_SLICE_X12Y105_DO6;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_CMUX = CLBLM_L_X10Y105_SLICE_X12Y105_CO5;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_A = CLBLM_L_X10Y105_SLICE_X13Y105_AO6;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_B = CLBLM_L_X10Y105_SLICE_X13Y105_BO6;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_C = CLBLM_L_X10Y105_SLICE_X13Y105_CO6;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_D = CLBLM_L_X10Y105_SLICE_X13Y105_DO6;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_A = CLBLM_L_X10Y106_SLICE_X12Y106_AO6;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_B = CLBLM_L_X10Y106_SLICE_X12Y106_BO6;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_C = CLBLM_L_X10Y106_SLICE_X12Y106_CO6;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_D = CLBLM_L_X10Y106_SLICE_X12Y106_DO6;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_BMUX = CLBLM_L_X10Y106_SLICE_X12Y106_BO5;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_A = CLBLM_L_X10Y106_SLICE_X13Y106_AO6;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_B = CLBLM_L_X10Y106_SLICE_X13Y106_BO6;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_C = CLBLM_L_X10Y106_SLICE_X13Y106_CO6;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_D = CLBLM_L_X10Y106_SLICE_X13Y106_DO6;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_A = CLBLM_L_X10Y107_SLICE_X12Y107_AO6;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_B = CLBLM_L_X10Y107_SLICE_X12Y107_BO6;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_C = CLBLM_L_X10Y107_SLICE_X12Y107_CO6;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_D = CLBLM_L_X10Y107_SLICE_X12Y107_DO6;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_DMUX = CLBLM_L_X10Y107_SLICE_X12Y107_DO6;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_A = CLBLM_L_X10Y107_SLICE_X13Y107_AO6;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_B = CLBLM_L_X10Y107_SLICE_X13Y107_BO6;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_C = CLBLM_L_X10Y107_SLICE_X13Y107_CO6;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_D = CLBLM_L_X10Y107_SLICE_X13Y107_DO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_A = CLBLM_L_X10Y108_SLICE_X12Y108_AO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_B = CLBLM_L_X10Y108_SLICE_X12Y108_BO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_C = CLBLM_L_X10Y108_SLICE_X12Y108_CO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_D = CLBLM_L_X10Y108_SLICE_X12Y108_DO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_AMUX = CLBLM_L_X10Y108_SLICE_X12Y108_AO5;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_A = CLBLM_L_X10Y108_SLICE_X13Y108_AO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_B = CLBLM_L_X10Y108_SLICE_X13Y108_BO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_C = CLBLM_L_X10Y108_SLICE_X13Y108_CO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_D = CLBLM_L_X10Y108_SLICE_X13Y108_DO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_A = CLBLM_L_X10Y109_SLICE_X12Y109_AO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_B = CLBLM_L_X10Y109_SLICE_X12Y109_BO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_C = CLBLM_L_X10Y109_SLICE_X12Y109_CO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_D = CLBLM_L_X10Y109_SLICE_X12Y109_DO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_CMUX = CLBLM_L_X10Y109_SLICE_X12Y109_CO5;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_A = CLBLM_L_X10Y109_SLICE_X13Y109_AO6;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_B = CLBLM_L_X10Y109_SLICE_X13Y109_BO6;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_C = CLBLM_L_X10Y109_SLICE_X13Y109_CO6;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_D = CLBLM_L_X10Y109_SLICE_X13Y109_DO6;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_AMUX = CLBLM_L_X10Y109_SLICE_X13Y109_AO5;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_BMUX = CLBLM_L_X10Y109_SLICE_X13Y109_BO5;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_DMUX = CLBLM_L_X10Y109_SLICE_X13Y109_DO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_A = CLBLM_L_X10Y110_SLICE_X12Y110_AO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_B = CLBLM_L_X10Y110_SLICE_X12Y110_BO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_C = CLBLM_L_X10Y110_SLICE_X12Y110_CO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_D = CLBLM_L_X10Y110_SLICE_X12Y110_DO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_BMUX = CLBLM_L_X10Y110_SLICE_X12Y110_B5Q;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_CMUX = CLBLM_L_X10Y110_SLICE_X12Y110_CO5;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_A = CLBLM_L_X10Y110_SLICE_X13Y110_AO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_B = CLBLM_L_X10Y110_SLICE_X13Y110_BO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_C = CLBLM_L_X10Y110_SLICE_X13Y110_CO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_D = CLBLM_L_X10Y110_SLICE_X13Y110_DO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_A = CLBLM_L_X10Y111_SLICE_X12Y111_AO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_B = CLBLM_L_X10Y111_SLICE_X12Y111_BO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_C = CLBLM_L_X10Y111_SLICE_X12Y111_CO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_D = CLBLM_L_X10Y111_SLICE_X12Y111_DO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_AMUX = CLBLM_L_X10Y111_SLICE_X12Y111_A5Q;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_CMUX = CLBLM_L_X10Y111_SLICE_X12Y111_C5Q;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_A = CLBLM_L_X10Y111_SLICE_X13Y111_AO6;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_B = CLBLM_L_X10Y111_SLICE_X13Y111_BO6;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_C = CLBLM_L_X10Y111_SLICE_X13Y111_CO6;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_D = CLBLM_L_X10Y111_SLICE_X13Y111_DO6;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_CMUX = CLBLM_L_X10Y111_SLICE_X13Y111_C5Q;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_A = CLBLM_L_X10Y112_SLICE_X12Y112_AO6;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_B = CLBLM_L_X10Y112_SLICE_X12Y112_BO6;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_C = CLBLM_L_X10Y112_SLICE_X12Y112_CO6;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_D = CLBLM_L_X10Y112_SLICE_X12Y112_DO6;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_CMUX = CLBLM_L_X10Y112_SLICE_X12Y112_C5Q;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_A = CLBLM_L_X10Y112_SLICE_X13Y112_AO6;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_B = CLBLM_L_X10Y112_SLICE_X13Y112_BO6;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_C = CLBLM_L_X10Y112_SLICE_X13Y112_CO6;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_D = CLBLM_L_X10Y112_SLICE_X13Y112_DO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_A = CLBLM_L_X10Y113_SLICE_X12Y113_AO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_B = CLBLM_L_X10Y113_SLICE_X12Y113_BO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_C = CLBLM_L_X10Y113_SLICE_X12Y113_CO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_D = CLBLM_L_X10Y113_SLICE_X12Y113_DO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_DMUX = CLBLM_L_X10Y113_SLICE_X12Y113_DO5;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_A = CLBLM_L_X10Y113_SLICE_X13Y113_AO6;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_B = CLBLM_L_X10Y113_SLICE_X13Y113_BO6;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_C = CLBLM_L_X10Y113_SLICE_X13Y113_CO6;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_D = CLBLM_L_X10Y113_SLICE_X13Y113_DO6;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_CMUX = CLBLM_L_X10Y113_SLICE_X13Y113_C5Q;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_A = CLBLM_L_X10Y114_SLICE_X12Y114_AO6;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_B = CLBLM_L_X10Y114_SLICE_X12Y114_BO6;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_C = CLBLM_L_X10Y114_SLICE_X12Y114_CO6;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_D = CLBLM_L_X10Y114_SLICE_X12Y114_DO6;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_A = CLBLM_L_X10Y114_SLICE_X13Y114_AO6;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_B = CLBLM_L_X10Y114_SLICE_X13Y114_BO6;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_C = CLBLM_L_X10Y114_SLICE_X13Y114_CO6;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_D = CLBLM_L_X10Y114_SLICE_X13Y114_DO6;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_A = CLBLM_L_X10Y115_SLICE_X12Y115_AO6;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_B = CLBLM_L_X10Y115_SLICE_X12Y115_BO6;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_C = CLBLM_L_X10Y115_SLICE_X12Y115_CO6;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_D = CLBLM_L_X10Y115_SLICE_X12Y115_DO6;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_A = CLBLM_L_X10Y115_SLICE_X13Y115_AO6;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_B = CLBLM_L_X10Y115_SLICE_X13Y115_BO6;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_C = CLBLM_L_X10Y115_SLICE_X13Y115_CO6;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_D = CLBLM_L_X10Y115_SLICE_X13Y115_DO6;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_DMUX = CLBLM_L_X10Y115_SLICE_X13Y115_DO5;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_A = CLBLM_L_X10Y116_SLICE_X12Y116_AO6;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_B = CLBLM_L_X10Y116_SLICE_X12Y116_BO6;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_C = CLBLM_L_X10Y116_SLICE_X12Y116_CO6;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_D = CLBLM_L_X10Y116_SLICE_X12Y116_DO6;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_DMUX = CLBLM_L_X10Y116_SLICE_X12Y116_DO5;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_A = CLBLM_L_X10Y116_SLICE_X13Y116_AO6;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_B = CLBLM_L_X10Y116_SLICE_X13Y116_BO6;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_C = CLBLM_L_X10Y116_SLICE_X13Y116_CO6;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_D = CLBLM_L_X10Y116_SLICE_X13Y116_DO6;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_A = CLBLM_L_X10Y117_SLICE_X12Y117_AO6;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_B = CLBLM_L_X10Y117_SLICE_X12Y117_BO6;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_C = CLBLM_L_X10Y117_SLICE_X12Y117_CO6;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_D = CLBLM_L_X10Y117_SLICE_X12Y117_DO6;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_AMUX = CLBLM_L_X10Y117_SLICE_X12Y117_A5Q;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_A = CLBLM_L_X10Y117_SLICE_X13Y117_AO6;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_B = CLBLM_L_X10Y117_SLICE_X13Y117_BO6;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_C = CLBLM_L_X10Y117_SLICE_X13Y117_CO6;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_D = CLBLM_L_X10Y117_SLICE_X13Y117_DO6;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_AMUX = CLBLM_L_X10Y117_SLICE_X13Y117_AO5;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_BMUX = CLBLM_L_X10Y117_SLICE_X13Y117_BO5;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_A = CLBLM_L_X10Y118_SLICE_X12Y118_AO6;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_B = CLBLM_L_X10Y118_SLICE_X12Y118_BO6;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_C = CLBLM_L_X10Y118_SLICE_X12Y118_CO6;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_D = CLBLM_L_X10Y118_SLICE_X12Y118_DO6;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_A = CLBLM_L_X10Y118_SLICE_X13Y118_AO6;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_B = CLBLM_L_X10Y118_SLICE_X13Y118_BO6;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_C = CLBLM_L_X10Y118_SLICE_X13Y118_CO6;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_D = CLBLM_L_X10Y118_SLICE_X13Y118_DO6;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_CMUX = CLBLM_L_X10Y118_SLICE_X13Y118_CO6;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_A = CLBLM_L_X10Y119_SLICE_X12Y119_AO6;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_B = CLBLM_L_X10Y119_SLICE_X12Y119_BO6;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_C = CLBLM_L_X10Y119_SLICE_X12Y119_CO6;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_D = CLBLM_L_X10Y119_SLICE_X12Y119_DO6;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_CMUX = CLBLM_L_X10Y119_SLICE_X12Y119_CO6;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_A = CLBLM_L_X10Y119_SLICE_X13Y119_AO6;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_B = CLBLM_L_X10Y119_SLICE_X13Y119_BO6;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_C = CLBLM_L_X10Y119_SLICE_X13Y119_CO6;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_D = CLBLM_L_X10Y119_SLICE_X13Y119_DO6;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_A = CLBLM_L_X10Y148_SLICE_X12Y148_AO6;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_B = CLBLM_L_X10Y148_SLICE_X12Y148_BO6;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_C = CLBLM_L_X10Y148_SLICE_X12Y148_CO6;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_D = CLBLM_L_X10Y148_SLICE_X12Y148_DO6;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_A = CLBLM_L_X10Y148_SLICE_X13Y148_AO6;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_B = CLBLM_L_X10Y148_SLICE_X13Y148_BO6;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_C = CLBLM_L_X10Y148_SLICE_X13Y148_CO6;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_D = CLBLM_L_X10Y148_SLICE_X13Y148_DO6;
  assign CLBLM_L_X12Y105_SLICE_X16Y105_A = CLBLM_L_X12Y105_SLICE_X16Y105_AO6;
  assign CLBLM_L_X12Y105_SLICE_X16Y105_B = CLBLM_L_X12Y105_SLICE_X16Y105_BO6;
  assign CLBLM_L_X12Y105_SLICE_X16Y105_C = CLBLM_L_X12Y105_SLICE_X16Y105_CO6;
  assign CLBLM_L_X12Y105_SLICE_X16Y105_D = CLBLM_L_X12Y105_SLICE_X16Y105_DO6;
  assign CLBLM_L_X12Y105_SLICE_X16Y105_BMUX = CLBLM_L_X12Y105_SLICE_X16Y105_BO5;
  assign CLBLM_L_X12Y105_SLICE_X16Y105_CMUX = CLBLM_L_X12Y105_SLICE_X16Y105_CO5;
  assign CLBLM_L_X12Y105_SLICE_X17Y105_A = CLBLM_L_X12Y105_SLICE_X17Y105_AO6;
  assign CLBLM_L_X12Y105_SLICE_X17Y105_B = CLBLM_L_X12Y105_SLICE_X17Y105_BO6;
  assign CLBLM_L_X12Y105_SLICE_X17Y105_C = CLBLM_L_X12Y105_SLICE_X17Y105_CO6;
  assign CLBLM_L_X12Y105_SLICE_X17Y105_D = CLBLM_L_X12Y105_SLICE_X17Y105_DO6;
  assign CLBLM_L_X12Y105_SLICE_X17Y105_AMUX = CLBLM_L_X12Y105_SLICE_X17Y105_AO5;
  assign CLBLM_L_X12Y105_SLICE_X17Y105_BMUX = CLBLM_L_X12Y105_SLICE_X17Y105_BO5;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_A = CLBLM_L_X12Y106_SLICE_X16Y106_AO6;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_B = CLBLM_L_X12Y106_SLICE_X16Y106_BO6;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_C = CLBLM_L_X12Y106_SLICE_X16Y106_CO6;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_D = CLBLM_L_X12Y106_SLICE_X16Y106_DO6;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_A = CLBLM_L_X12Y106_SLICE_X17Y106_AO6;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_B = CLBLM_L_X12Y106_SLICE_X17Y106_BO6;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_C = CLBLM_L_X12Y106_SLICE_X17Y106_CO6;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_D = CLBLM_L_X12Y106_SLICE_X17Y106_DO6;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_A = CLBLM_L_X12Y107_SLICE_X16Y107_AO6;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_B = CLBLM_L_X12Y107_SLICE_X16Y107_BO6;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_C = CLBLM_L_X12Y107_SLICE_X16Y107_CO6;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_D = CLBLM_L_X12Y107_SLICE_X16Y107_DO6;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_A = CLBLM_L_X12Y107_SLICE_X17Y107_AO6;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_B = CLBLM_L_X12Y107_SLICE_X17Y107_BO6;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_C = CLBLM_L_X12Y107_SLICE_X17Y107_CO6;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_D = CLBLM_L_X12Y107_SLICE_X17Y107_DO6;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_CMUX = CLBLM_L_X12Y107_SLICE_X17Y107_CO5;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_DMUX = CLBLM_L_X12Y107_SLICE_X17Y107_DO5;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_A = CLBLM_L_X12Y108_SLICE_X16Y108_AO6;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_B = CLBLM_L_X12Y108_SLICE_X16Y108_BO6;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_C = CLBLM_L_X12Y108_SLICE_X16Y108_CO6;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_D = CLBLM_L_X12Y108_SLICE_X16Y108_DO6;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_AMUX = CLBLM_L_X12Y108_SLICE_X16Y108_AO5;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_A = CLBLM_L_X12Y108_SLICE_X17Y108_AO6;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_B = CLBLM_L_X12Y108_SLICE_X17Y108_BO6;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_C = CLBLM_L_X12Y108_SLICE_X17Y108_CO6;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_D = CLBLM_L_X12Y108_SLICE_X17Y108_DO6;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_CMUX = CLBLM_L_X12Y108_SLICE_X17Y108_CO5;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_A = CLBLM_L_X12Y109_SLICE_X16Y109_AO6;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_B = CLBLM_L_X12Y109_SLICE_X16Y109_BO6;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_C = CLBLM_L_X12Y109_SLICE_X16Y109_CO6;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_D = CLBLM_L_X12Y109_SLICE_X16Y109_DO6;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_DMUX = CLBLM_L_X12Y109_SLICE_X16Y109_D5Q;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_A = CLBLM_L_X12Y109_SLICE_X17Y109_AO6;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_B = CLBLM_L_X12Y109_SLICE_X17Y109_BO6;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_C = CLBLM_L_X12Y109_SLICE_X17Y109_CO6;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_D = CLBLM_L_X12Y109_SLICE_X17Y109_DO6;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_A = CLBLM_L_X12Y110_SLICE_X16Y110_AO6;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_B = CLBLM_L_X12Y110_SLICE_X16Y110_BO6;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_C = CLBLM_L_X12Y110_SLICE_X16Y110_CO6;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_D = CLBLM_L_X12Y110_SLICE_X16Y110_DO6;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_AMUX = CLBLM_L_X12Y110_SLICE_X16Y110_AO5;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_BMUX = CLBLM_L_X12Y110_SLICE_X16Y110_BO5;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_CMUX = CLBLM_L_X12Y110_SLICE_X16Y110_CO5;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_DMUX = CLBLM_L_X12Y110_SLICE_X16Y110_DO5;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_A = CLBLM_L_X12Y110_SLICE_X17Y110_AO6;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_B = CLBLM_L_X12Y110_SLICE_X17Y110_BO6;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_C = CLBLM_L_X12Y110_SLICE_X17Y110_CO6;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_D = CLBLM_L_X12Y110_SLICE_X17Y110_DO6;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_A = CLBLM_L_X12Y111_SLICE_X16Y111_AO6;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_B = CLBLM_L_X12Y111_SLICE_X16Y111_BO6;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_C = CLBLM_L_X12Y111_SLICE_X16Y111_CO6;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_D = CLBLM_L_X12Y111_SLICE_X16Y111_DO6;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_A = CLBLM_L_X12Y111_SLICE_X17Y111_AO6;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_B = CLBLM_L_X12Y111_SLICE_X17Y111_BO6;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_C = CLBLM_L_X12Y111_SLICE_X17Y111_CO6;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_D = CLBLM_L_X12Y111_SLICE_X17Y111_DO6;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_A = CLBLM_L_X12Y112_SLICE_X16Y112_AO6;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_B = CLBLM_L_X12Y112_SLICE_X16Y112_BO6;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_C = CLBLM_L_X12Y112_SLICE_X16Y112_CO6;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_D = CLBLM_L_X12Y112_SLICE_X16Y112_DO6;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_AMUX = CLBLM_L_X12Y112_SLICE_X16Y112_A5Q;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_BMUX = CLBLM_L_X12Y112_SLICE_X16Y112_B5Q;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_A = CLBLM_L_X12Y112_SLICE_X17Y112_AO6;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_B = CLBLM_L_X12Y112_SLICE_X17Y112_BO6;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_C = CLBLM_L_X12Y112_SLICE_X17Y112_CO6;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_D = CLBLM_L_X12Y112_SLICE_X17Y112_DO6;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_AMUX = CLBLM_L_X12Y112_SLICE_X17Y112_A5Q;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_BMUX = CLBLM_L_X12Y112_SLICE_X17Y112_B5Q;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_CMUX = CLBLM_L_X12Y112_SLICE_X17Y112_CO5;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_A = CLBLM_L_X12Y113_SLICE_X16Y113_AO6;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_B = CLBLM_L_X12Y113_SLICE_X16Y113_BO6;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_C = CLBLM_L_X12Y113_SLICE_X16Y113_CO6;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_D = CLBLM_L_X12Y113_SLICE_X16Y113_DO6;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_A = CLBLM_L_X12Y113_SLICE_X17Y113_AO6;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_B = CLBLM_L_X12Y113_SLICE_X17Y113_BO6;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_C = CLBLM_L_X12Y113_SLICE_X17Y113_CO6;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_D = CLBLM_L_X12Y113_SLICE_X17Y113_DO6;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_BMUX = CLBLM_L_X12Y113_SLICE_X17Y113_B5Q;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_A = CLBLM_L_X12Y114_SLICE_X16Y114_AO6;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_B = CLBLM_L_X12Y114_SLICE_X16Y114_BO6;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_C = CLBLM_L_X12Y114_SLICE_X16Y114_CO6;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_D = CLBLM_L_X12Y114_SLICE_X16Y114_DO6;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_DMUX = CLBLM_L_X12Y114_SLICE_X16Y114_DO5;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_A = CLBLM_L_X12Y114_SLICE_X17Y114_AO6;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_B = CLBLM_L_X12Y114_SLICE_X17Y114_BO6;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_C = CLBLM_L_X12Y114_SLICE_X17Y114_CO6;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_D = CLBLM_L_X12Y114_SLICE_X17Y114_DO6;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_A = CLBLM_L_X12Y115_SLICE_X16Y115_AO6;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_B = CLBLM_L_X12Y115_SLICE_X16Y115_BO6;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_C = CLBLM_L_X12Y115_SLICE_X16Y115_CO6;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_D = CLBLM_L_X12Y115_SLICE_X16Y115_DO6;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_A = CLBLM_L_X12Y115_SLICE_X17Y115_AO6;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_B = CLBLM_L_X12Y115_SLICE_X17Y115_BO6;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_C = CLBLM_L_X12Y115_SLICE_X17Y115_CO6;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_D = CLBLM_L_X12Y115_SLICE_X17Y115_DO6;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_A = CLBLM_L_X12Y117_SLICE_X16Y117_AO6;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_B = CLBLM_L_X12Y117_SLICE_X16Y117_BO6;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_C = CLBLM_L_X12Y117_SLICE_X16Y117_CO6;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_D = CLBLM_L_X12Y117_SLICE_X16Y117_DO6;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_AMUX = CLBLM_L_X12Y117_SLICE_X16Y117_AO6;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_A = CLBLM_L_X12Y117_SLICE_X17Y117_AO6;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_B = CLBLM_L_X12Y117_SLICE_X17Y117_BO6;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_C = CLBLM_L_X12Y117_SLICE_X17Y117_CO6;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_D = CLBLM_L_X12Y117_SLICE_X17Y117_DO6;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_A = CLBLM_L_X12Y118_SLICE_X16Y118_AO6;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_B = CLBLM_L_X12Y118_SLICE_X16Y118_BO6;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_C = CLBLM_L_X12Y118_SLICE_X16Y118_CO6;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_D = CLBLM_L_X12Y118_SLICE_X16Y118_DO6;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_A = CLBLM_L_X12Y118_SLICE_X17Y118_AO6;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_B = CLBLM_L_X12Y118_SLICE_X17Y118_BO6;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_C = CLBLM_L_X12Y118_SLICE_X17Y118_CO6;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_D = CLBLM_L_X12Y118_SLICE_X17Y118_DO6;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_A = CLBLM_R_X3Y106_SLICE_X2Y106_AO6;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_B = CLBLM_R_X3Y106_SLICE_X2Y106_BO6;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_C = CLBLM_R_X3Y106_SLICE_X2Y106_CO6;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_D = CLBLM_R_X3Y106_SLICE_X2Y106_DO6;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_A = CLBLM_R_X3Y106_SLICE_X3Y106_AO6;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_B = CLBLM_R_X3Y106_SLICE_X3Y106_BO6;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_C = CLBLM_R_X3Y106_SLICE_X3Y106_CO6;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_D = CLBLM_R_X3Y106_SLICE_X3Y106_DO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_A = CLBLM_R_X3Y107_SLICE_X2Y107_AO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_B = CLBLM_R_X3Y107_SLICE_X2Y107_BO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_C = CLBLM_R_X3Y107_SLICE_X2Y107_CO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_D = CLBLM_R_X3Y107_SLICE_X2Y107_DO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_A = CLBLM_R_X3Y107_SLICE_X3Y107_AO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_B = CLBLM_R_X3Y107_SLICE_X3Y107_BO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_C = CLBLM_R_X3Y107_SLICE_X3Y107_CO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_D = CLBLM_R_X3Y107_SLICE_X3Y107_DO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_BMUX = CLBLM_R_X3Y107_SLICE_X3Y107_BO5;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_A = CLBLM_R_X3Y108_SLICE_X2Y108_AO6;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_B = CLBLM_R_X3Y108_SLICE_X2Y108_BO6;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_C = CLBLM_R_X3Y108_SLICE_X2Y108_CO6;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_D = CLBLM_R_X3Y108_SLICE_X2Y108_DO6;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_CMUX = CLBLM_R_X3Y108_SLICE_X2Y108_CO6;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_DMUX = CLBLM_R_X3Y108_SLICE_X2Y108_DO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_A = CLBLM_R_X3Y108_SLICE_X3Y108_AO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_B = CLBLM_R_X3Y108_SLICE_X3Y108_BO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_C = CLBLM_R_X3Y108_SLICE_X3Y108_CO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_D = CLBLM_R_X3Y108_SLICE_X3Y108_DO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_DMUX = CLBLM_R_X3Y108_SLICE_X3Y108_DO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_A = CLBLM_R_X3Y109_SLICE_X2Y109_AO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_B = CLBLM_R_X3Y109_SLICE_X2Y109_BO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_C = CLBLM_R_X3Y109_SLICE_X2Y109_CO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_D = CLBLM_R_X3Y109_SLICE_X2Y109_DO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_AMUX = CLBLM_R_X3Y109_SLICE_X2Y109_A5Q;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_CMUX = CLBLM_R_X3Y109_SLICE_X2Y109_CO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_DMUX = CLBLM_R_X3Y109_SLICE_X2Y109_DO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_A = CLBLM_R_X3Y109_SLICE_X3Y109_AO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_B = CLBLM_R_X3Y109_SLICE_X3Y109_BO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_C = CLBLM_R_X3Y109_SLICE_X3Y109_CO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_D = CLBLM_R_X3Y109_SLICE_X3Y109_DO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_A = CLBLM_R_X3Y110_SLICE_X2Y110_AO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_B = CLBLM_R_X3Y110_SLICE_X2Y110_BO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_C = CLBLM_R_X3Y110_SLICE_X2Y110_CO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_D = CLBLM_R_X3Y110_SLICE_X2Y110_DO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_AMUX = CLBLM_R_X3Y110_SLICE_X2Y110_AO5;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_DMUX = CLBLM_R_X3Y110_SLICE_X2Y110_DO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_A = CLBLM_R_X3Y110_SLICE_X3Y110_AO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_B = CLBLM_R_X3Y110_SLICE_X3Y110_BO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_C = CLBLM_R_X3Y110_SLICE_X3Y110_CO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_D = CLBLM_R_X3Y110_SLICE_X3Y110_DO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_A = CLBLM_R_X3Y111_SLICE_X2Y111_AO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_B = CLBLM_R_X3Y111_SLICE_X2Y111_BO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_C = CLBLM_R_X3Y111_SLICE_X2Y111_CO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_D = CLBLM_R_X3Y111_SLICE_X2Y111_DO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_DMUX = CLBLM_R_X3Y111_SLICE_X2Y111_DO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_A = CLBLM_R_X3Y111_SLICE_X3Y111_AO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_B = CLBLM_R_X3Y111_SLICE_X3Y111_BO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_C = CLBLM_R_X3Y111_SLICE_X3Y111_CO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_D = CLBLM_R_X3Y111_SLICE_X3Y111_DO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_A = CLBLM_R_X3Y112_SLICE_X2Y112_AO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_B = CLBLM_R_X3Y112_SLICE_X2Y112_BO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_C = CLBLM_R_X3Y112_SLICE_X2Y112_CO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_D = CLBLM_R_X3Y112_SLICE_X2Y112_DO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_AMUX = CLBLM_R_X3Y112_SLICE_X2Y112_AO5;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_A = CLBLM_R_X3Y112_SLICE_X3Y112_AO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_B = CLBLM_R_X3Y112_SLICE_X3Y112_BO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_C = CLBLM_R_X3Y112_SLICE_X3Y112_CO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_D = CLBLM_R_X3Y112_SLICE_X3Y112_DO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_BMUX = CLBLM_R_X3Y112_SLICE_X3Y112_BO5;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_A = CLBLM_R_X3Y113_SLICE_X2Y113_AO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_B = CLBLM_R_X3Y113_SLICE_X2Y113_BO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_C = CLBLM_R_X3Y113_SLICE_X2Y113_CO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_D = CLBLM_R_X3Y113_SLICE_X2Y113_DO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_A = CLBLM_R_X3Y113_SLICE_X3Y113_AO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_B = CLBLM_R_X3Y113_SLICE_X3Y113_BO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_C = CLBLM_R_X3Y113_SLICE_X3Y113_CO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_D = CLBLM_R_X3Y113_SLICE_X3Y113_DO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_A = CLBLM_R_X3Y114_SLICE_X2Y114_AO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_B = CLBLM_R_X3Y114_SLICE_X2Y114_BO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_C = CLBLM_R_X3Y114_SLICE_X2Y114_CO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_D = CLBLM_R_X3Y114_SLICE_X2Y114_DO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_CMUX = CLBLM_R_X3Y114_SLICE_X2Y114_CO5;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_A = CLBLM_R_X3Y114_SLICE_X3Y114_AO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_B = CLBLM_R_X3Y114_SLICE_X3Y114_BO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_C = CLBLM_R_X3Y114_SLICE_X3Y114_CO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_D = CLBLM_R_X3Y114_SLICE_X3Y114_DO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_CMUX = CLBLM_R_X3Y114_SLICE_X3Y114_CO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_A = CLBLM_R_X3Y115_SLICE_X2Y115_AO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_B = CLBLM_R_X3Y115_SLICE_X2Y115_BO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_C = CLBLM_R_X3Y115_SLICE_X2Y115_CO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_D = CLBLM_R_X3Y115_SLICE_X2Y115_DO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_AMUX = CLBLM_R_X3Y115_SLICE_X2Y115_AO5;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_CMUX = CLBLM_R_X3Y115_SLICE_X2Y115_CO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_A = CLBLM_R_X3Y115_SLICE_X3Y115_AO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_B = CLBLM_R_X3Y115_SLICE_X3Y115_BO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_C = CLBLM_R_X3Y115_SLICE_X3Y115_CO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_D = CLBLM_R_X3Y115_SLICE_X3Y115_DO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_AMUX = CLBLM_R_X3Y115_SLICE_X3Y115_AO5;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_BMUX = CLBLM_R_X3Y115_SLICE_X3Y115_BO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_CMUX = CLBLM_R_X3Y115_SLICE_X3Y115_CO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_DMUX = CLBLM_R_X3Y115_SLICE_X3Y115_DO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_A = CLBLM_R_X3Y116_SLICE_X2Y116_AO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_B = CLBLM_R_X3Y116_SLICE_X2Y116_BO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_C = CLBLM_R_X3Y116_SLICE_X2Y116_CO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_D = CLBLM_R_X3Y116_SLICE_X2Y116_DO6;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_AMUX = CLBLM_R_X3Y116_SLICE_X2Y116_AO6;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_A = CLBLM_R_X3Y116_SLICE_X3Y116_AO6;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_B = CLBLM_R_X3Y116_SLICE_X3Y116_BO6;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_C = CLBLM_R_X3Y116_SLICE_X3Y116_CO6;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_D = CLBLM_R_X3Y116_SLICE_X3Y116_DO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_A = CLBLM_R_X3Y118_SLICE_X2Y118_AO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_B = CLBLM_R_X3Y118_SLICE_X2Y118_BO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_C = CLBLM_R_X3Y118_SLICE_X2Y118_CO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_D = CLBLM_R_X3Y118_SLICE_X2Y118_DO6;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_A = CLBLM_R_X3Y118_SLICE_X3Y118_AO6;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_B = CLBLM_R_X3Y118_SLICE_X3Y118_BO6;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_C = CLBLM_R_X3Y118_SLICE_X3Y118_CO6;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_D = CLBLM_R_X3Y118_SLICE_X3Y118_DO6;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_A = CLBLM_R_X5Y105_SLICE_X6Y105_AO6;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_B = CLBLM_R_X5Y105_SLICE_X6Y105_BO6;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_C = CLBLM_R_X5Y105_SLICE_X6Y105_CO6;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_D = CLBLM_R_X5Y105_SLICE_X6Y105_DO6;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_A = CLBLM_R_X5Y105_SLICE_X7Y105_AO6;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_B = CLBLM_R_X5Y105_SLICE_X7Y105_BO6;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_C = CLBLM_R_X5Y105_SLICE_X7Y105_CO6;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_D = CLBLM_R_X5Y105_SLICE_X7Y105_DO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_A = CLBLM_R_X5Y106_SLICE_X6Y106_AO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_B = CLBLM_R_X5Y106_SLICE_X6Y106_BO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_C = CLBLM_R_X5Y106_SLICE_X6Y106_CO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_D = CLBLM_R_X5Y106_SLICE_X6Y106_DO6;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_A = CLBLM_R_X5Y106_SLICE_X7Y106_AO6;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_B = CLBLM_R_X5Y106_SLICE_X7Y106_BO6;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_C = CLBLM_R_X5Y106_SLICE_X7Y106_CO6;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_D = CLBLM_R_X5Y106_SLICE_X7Y106_DO6;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_BMUX = CLBLM_R_X5Y106_SLICE_X7Y106_BO5;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_A = CLBLM_R_X5Y107_SLICE_X6Y107_AO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_B = CLBLM_R_X5Y107_SLICE_X6Y107_BO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_C = CLBLM_R_X5Y107_SLICE_X6Y107_CO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_D = CLBLM_R_X5Y107_SLICE_X6Y107_DO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_A = CLBLM_R_X5Y107_SLICE_X7Y107_AO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_B = CLBLM_R_X5Y107_SLICE_X7Y107_BO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_C = CLBLM_R_X5Y107_SLICE_X7Y107_CO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_D = CLBLM_R_X5Y107_SLICE_X7Y107_DO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_BMUX = CLBLM_R_X5Y107_SLICE_X7Y107_B5Q;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_CMUX = CLBLM_R_X5Y107_SLICE_X7Y107_CO5;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_DMUX = CLBLM_R_X5Y107_SLICE_X7Y107_DO5;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_A = CLBLM_R_X5Y108_SLICE_X6Y108_AO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_B = CLBLM_R_X5Y108_SLICE_X6Y108_BO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_C = CLBLM_R_X5Y108_SLICE_X6Y108_CO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_D = CLBLM_R_X5Y108_SLICE_X6Y108_DO6;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_A = CLBLM_R_X5Y108_SLICE_X7Y108_AO6;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_B = CLBLM_R_X5Y108_SLICE_X7Y108_BO6;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_C = CLBLM_R_X5Y108_SLICE_X7Y108_CO6;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_D = CLBLM_R_X5Y108_SLICE_X7Y108_DO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_A = CLBLM_R_X5Y109_SLICE_X6Y109_AO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_B = CLBLM_R_X5Y109_SLICE_X6Y109_BO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_C = CLBLM_R_X5Y109_SLICE_X6Y109_CO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_D = CLBLM_R_X5Y109_SLICE_X6Y109_DO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_A = CLBLM_R_X5Y109_SLICE_X7Y109_AO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_B = CLBLM_R_X5Y109_SLICE_X7Y109_BO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_C = CLBLM_R_X5Y109_SLICE_X7Y109_CO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_D = CLBLM_R_X5Y109_SLICE_X7Y109_DO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_AMUX = CLBLM_R_X5Y109_SLICE_X7Y109_A5Q;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_BMUX = CLBLM_R_X5Y109_SLICE_X7Y109_B5Q;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_CMUX = CLBLM_R_X5Y109_SLICE_X7Y109_CO5;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_A = CLBLM_R_X5Y110_SLICE_X6Y110_AO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_B = CLBLM_R_X5Y110_SLICE_X6Y110_BO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_C = CLBLM_R_X5Y110_SLICE_X6Y110_CO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_D = CLBLM_R_X5Y110_SLICE_X6Y110_DO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_BMUX = CLBLM_R_X5Y110_SLICE_X6Y110_B5Q;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_A = CLBLM_R_X5Y110_SLICE_X7Y110_AO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_B = CLBLM_R_X5Y110_SLICE_X7Y110_BO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_C = CLBLM_R_X5Y110_SLICE_X7Y110_CO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_D = CLBLM_R_X5Y110_SLICE_X7Y110_DO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_BMUX = CLBLM_R_X5Y110_SLICE_X7Y110_B5Q;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_CMUX = CLBLM_R_X5Y110_SLICE_X7Y110_CO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_A = CLBLM_R_X5Y111_SLICE_X6Y111_AO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_B = CLBLM_R_X5Y111_SLICE_X6Y111_BO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_C = CLBLM_R_X5Y111_SLICE_X6Y111_CO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_D = CLBLM_R_X5Y111_SLICE_X6Y111_DO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_A = CLBLM_R_X5Y111_SLICE_X7Y111_AO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_B = CLBLM_R_X5Y111_SLICE_X7Y111_BO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_C = CLBLM_R_X5Y111_SLICE_X7Y111_CO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_D = CLBLM_R_X5Y111_SLICE_X7Y111_DO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_A = CLBLM_R_X5Y112_SLICE_X6Y112_AO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_B = CLBLM_R_X5Y112_SLICE_X6Y112_BO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_C = CLBLM_R_X5Y112_SLICE_X6Y112_CO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_D = CLBLM_R_X5Y112_SLICE_X6Y112_DO6;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_A = CLBLM_R_X5Y112_SLICE_X7Y112_AO6;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_B = CLBLM_R_X5Y112_SLICE_X7Y112_BO6;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_C = CLBLM_R_X5Y112_SLICE_X7Y112_CO6;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_D = CLBLM_R_X5Y112_SLICE_X7Y112_DO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_A = CLBLM_R_X5Y113_SLICE_X6Y113_AO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_B = CLBLM_R_X5Y113_SLICE_X6Y113_BO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_C = CLBLM_R_X5Y113_SLICE_X6Y113_CO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_D = CLBLM_R_X5Y113_SLICE_X6Y113_DO6;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_A = CLBLM_R_X5Y113_SLICE_X7Y113_AO6;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_B = CLBLM_R_X5Y113_SLICE_X7Y113_BO6;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_C = CLBLM_R_X5Y113_SLICE_X7Y113_CO6;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_D = CLBLM_R_X5Y113_SLICE_X7Y113_DO6;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_A = CLBLM_R_X5Y114_SLICE_X6Y114_AO6;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_B = CLBLM_R_X5Y114_SLICE_X6Y114_BO6;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_C = CLBLM_R_X5Y114_SLICE_X6Y114_CO6;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_D = CLBLM_R_X5Y114_SLICE_X6Y114_DO6;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_A = CLBLM_R_X5Y114_SLICE_X7Y114_AO6;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_B = CLBLM_R_X5Y114_SLICE_X7Y114_BO6;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_C = CLBLM_R_X5Y114_SLICE_X7Y114_CO6;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_D = CLBLM_R_X5Y114_SLICE_X7Y114_DO6;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_BMUX = CLBLM_R_X5Y114_SLICE_X7Y114_B5Q;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_CMUX = CLBLM_R_X5Y114_SLICE_X7Y114_C5Q;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_A = CLBLM_R_X5Y115_SLICE_X6Y115_AO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_B = CLBLM_R_X5Y115_SLICE_X6Y115_BO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_C = CLBLM_R_X5Y115_SLICE_X6Y115_CO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_D = CLBLM_R_X5Y115_SLICE_X6Y115_DO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_DMUX = CLBLM_R_X5Y115_SLICE_X6Y115_DO5;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_A = CLBLM_R_X5Y115_SLICE_X7Y115_AO6;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_B = CLBLM_R_X5Y115_SLICE_X7Y115_BO6;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_C = CLBLM_R_X5Y115_SLICE_X7Y115_CO6;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_D = CLBLM_R_X5Y115_SLICE_X7Y115_DO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_A = CLBLM_R_X5Y116_SLICE_X6Y116_AO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_B = CLBLM_R_X5Y116_SLICE_X6Y116_BO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_C = CLBLM_R_X5Y116_SLICE_X6Y116_CO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_D = CLBLM_R_X5Y116_SLICE_X6Y116_DO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_AMUX = CLBLM_R_X5Y116_SLICE_X6Y116_AO5;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_DMUX = CLBLM_R_X5Y116_SLICE_X6Y116_D5Q;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_A = CLBLM_R_X5Y116_SLICE_X7Y116_AO6;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_B = CLBLM_R_X5Y116_SLICE_X7Y116_BO6;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_C = CLBLM_R_X5Y116_SLICE_X7Y116_CO6;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_D = CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_AMUX = CLBLM_R_X5Y116_SLICE_X7Y116_A5Q;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_CMUX = CLBLM_R_X5Y116_SLICE_X7Y116_CO5;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_A = CLBLM_R_X5Y117_SLICE_X6Y117_AO6;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_B = CLBLM_R_X5Y117_SLICE_X6Y117_BO6;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_C = CLBLM_R_X5Y117_SLICE_X6Y117_CO6;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_D = CLBLM_R_X5Y117_SLICE_X6Y117_DO6;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_A = CLBLM_R_X5Y117_SLICE_X7Y117_AO6;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_B = CLBLM_R_X5Y117_SLICE_X7Y117_BO6;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_C = CLBLM_R_X5Y117_SLICE_X7Y117_CO6;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_D = CLBLM_R_X5Y117_SLICE_X7Y117_DO6;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_A = CLBLM_R_X7Y105_SLICE_X8Y105_AO6;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_B = CLBLM_R_X7Y105_SLICE_X8Y105_BO6;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_C = CLBLM_R_X7Y105_SLICE_X8Y105_CO6;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_D = CLBLM_R_X7Y105_SLICE_X8Y105_DO6;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_AMUX = CLBLM_R_X7Y105_SLICE_X8Y105_A5Q;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_BMUX = CLBLM_R_X7Y105_SLICE_X8Y105_BO5;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_A = CLBLM_R_X7Y105_SLICE_X9Y105_AO6;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_B = CLBLM_R_X7Y105_SLICE_X9Y105_BO6;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_C = CLBLM_R_X7Y105_SLICE_X9Y105_CO6;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_D = CLBLM_R_X7Y105_SLICE_X9Y105_DO6;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_AMUX = CLBLM_R_X7Y105_SLICE_X9Y105_AO5;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_A = CLBLM_R_X7Y106_SLICE_X8Y106_AO6;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_B = CLBLM_R_X7Y106_SLICE_X8Y106_BO6;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_C = CLBLM_R_X7Y106_SLICE_X8Y106_CO6;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_D = CLBLM_R_X7Y106_SLICE_X8Y106_DO6;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_A = CLBLM_R_X7Y106_SLICE_X9Y106_AO6;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_B = CLBLM_R_X7Y106_SLICE_X9Y106_BO6;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_C = CLBLM_R_X7Y106_SLICE_X9Y106_CO6;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_D = CLBLM_R_X7Y106_SLICE_X9Y106_DO6;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_DMUX = CLBLM_R_X7Y106_SLICE_X9Y106_DO5;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_A = CLBLM_R_X7Y107_SLICE_X8Y107_AO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_B = CLBLM_R_X7Y107_SLICE_X8Y107_BO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_C = CLBLM_R_X7Y107_SLICE_X8Y107_CO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_D = CLBLM_R_X7Y107_SLICE_X8Y107_DO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_A = CLBLM_R_X7Y107_SLICE_X9Y107_AO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_B = CLBLM_R_X7Y107_SLICE_X9Y107_BO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_C = CLBLM_R_X7Y107_SLICE_X9Y107_CO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_D = CLBLM_R_X7Y107_SLICE_X9Y107_DO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_CMUX = CLBLM_R_X7Y107_SLICE_X9Y107_C5Q;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_A = CLBLM_R_X7Y108_SLICE_X8Y108_AO6;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_B = CLBLM_R_X7Y108_SLICE_X8Y108_BO6;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_C = CLBLM_R_X7Y108_SLICE_X8Y108_CO6;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_D = CLBLM_R_X7Y108_SLICE_X8Y108_DO6;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_DMUX = CLBLM_R_X7Y108_SLICE_X8Y108_DO5;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_A = CLBLM_R_X7Y108_SLICE_X9Y108_AO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_B = CLBLM_R_X7Y108_SLICE_X9Y108_BO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_C = CLBLM_R_X7Y108_SLICE_X9Y108_CO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_D = CLBLM_R_X7Y108_SLICE_X9Y108_DO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_BMUX = CLBLM_R_X7Y108_SLICE_X9Y108_BO5;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_A = CLBLM_R_X7Y109_SLICE_X8Y109_AO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_B = CLBLM_R_X7Y109_SLICE_X8Y109_BO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_C = CLBLM_R_X7Y109_SLICE_X8Y109_CO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_D = CLBLM_R_X7Y109_SLICE_X8Y109_DO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_CMUX = CLBLM_R_X7Y109_SLICE_X8Y109_CO5;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_DMUX = CLBLM_R_X7Y109_SLICE_X8Y109_DO5;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_A = CLBLM_R_X7Y109_SLICE_X9Y109_AO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_B = CLBLM_R_X7Y109_SLICE_X9Y109_BO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_C = CLBLM_R_X7Y109_SLICE_X9Y109_CO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_D = CLBLM_R_X7Y109_SLICE_X9Y109_DO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_A = CLBLM_R_X7Y110_SLICE_X8Y110_AO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_B = CLBLM_R_X7Y110_SLICE_X8Y110_BO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_C = CLBLM_R_X7Y110_SLICE_X8Y110_CO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_D = CLBLM_R_X7Y110_SLICE_X8Y110_DO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_DMUX = CLBLM_R_X7Y110_SLICE_X8Y110_DO5;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_A = CLBLM_R_X7Y110_SLICE_X9Y110_AO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_B = CLBLM_R_X7Y110_SLICE_X9Y110_BO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_C = CLBLM_R_X7Y110_SLICE_X9Y110_CO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_D = CLBLM_R_X7Y110_SLICE_X9Y110_DO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_A = CLBLM_R_X7Y111_SLICE_X8Y111_AO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_B = CLBLM_R_X7Y111_SLICE_X8Y111_BO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_C = CLBLM_R_X7Y111_SLICE_X8Y111_CO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_D = CLBLM_R_X7Y111_SLICE_X8Y111_DO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_A = CLBLM_R_X7Y111_SLICE_X9Y111_AO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_B = CLBLM_R_X7Y111_SLICE_X9Y111_BO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_C = CLBLM_R_X7Y111_SLICE_X9Y111_CO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_D = CLBLM_R_X7Y111_SLICE_X9Y111_DO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_DMUX = CLBLM_R_X7Y111_SLICE_X9Y111_DO5;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_A = CLBLM_R_X7Y112_SLICE_X8Y112_AO6;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_B = CLBLM_R_X7Y112_SLICE_X8Y112_BO6;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_C = CLBLM_R_X7Y112_SLICE_X8Y112_CO6;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_D = CLBLM_R_X7Y112_SLICE_X8Y112_DO6;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_CMUX = CLBLM_R_X7Y112_SLICE_X8Y112_C5Q;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_A = CLBLM_R_X7Y112_SLICE_X9Y112_AO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_B = CLBLM_R_X7Y112_SLICE_X9Y112_BO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_C = CLBLM_R_X7Y112_SLICE_X9Y112_CO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_D = CLBLM_R_X7Y112_SLICE_X9Y112_DO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_A = CLBLM_R_X7Y113_SLICE_X8Y113_AO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_B = CLBLM_R_X7Y113_SLICE_X8Y113_BO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_C = CLBLM_R_X7Y113_SLICE_X8Y113_CO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_D = CLBLM_R_X7Y113_SLICE_X8Y113_DO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_CMUX = CLBLM_R_X7Y113_SLICE_X8Y113_C5Q;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_A = CLBLM_R_X7Y113_SLICE_X9Y113_AO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_B = CLBLM_R_X7Y113_SLICE_X9Y113_BO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_C = CLBLM_R_X7Y113_SLICE_X9Y113_CO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_D = CLBLM_R_X7Y113_SLICE_X9Y113_DO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_AMUX = CLBLM_R_X7Y113_SLICE_X9Y113_A5Q;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_BMUX = CLBLM_R_X7Y113_SLICE_X9Y113_BO5;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_A = CLBLM_R_X7Y114_SLICE_X8Y114_AO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_B = CLBLM_R_X7Y114_SLICE_X8Y114_BO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_C = CLBLM_R_X7Y114_SLICE_X8Y114_CO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_D = CLBLM_R_X7Y114_SLICE_X8Y114_DO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_AMUX = CLBLM_R_X7Y114_SLICE_X8Y114_A5Q;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_A = CLBLM_R_X7Y114_SLICE_X9Y114_AO6;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_B = CLBLM_R_X7Y114_SLICE_X9Y114_BO6;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_C = CLBLM_R_X7Y114_SLICE_X9Y114_CO6;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_D = CLBLM_R_X7Y114_SLICE_X9Y114_DO6;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_AMUX = CLBLM_R_X7Y114_SLICE_X9Y114_AO5;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_A = CLBLM_R_X7Y115_SLICE_X8Y115_AO6;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_B = CLBLM_R_X7Y115_SLICE_X8Y115_BO6;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_C = CLBLM_R_X7Y115_SLICE_X8Y115_CO6;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_D = CLBLM_R_X7Y115_SLICE_X8Y115_DO6;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_BMUX = CLBLM_R_X7Y115_SLICE_X8Y115_B5Q;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_DMUX = CLBLM_R_X7Y115_SLICE_X8Y115_D5Q;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_A = CLBLM_R_X7Y115_SLICE_X9Y115_AO6;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_B = CLBLM_R_X7Y115_SLICE_X9Y115_BO6;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_C = CLBLM_R_X7Y115_SLICE_X9Y115_CO6;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_D = CLBLM_R_X7Y115_SLICE_X9Y115_DO6;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_AMUX = CLBLM_R_X7Y115_SLICE_X9Y115_A5Q;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_BMUX = CLBLM_R_X7Y115_SLICE_X9Y115_B5Q;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_CMUX = CLBLM_R_X7Y115_SLICE_X9Y115_CO5;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_A = CLBLM_R_X7Y116_SLICE_X8Y116_AO6;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_B = CLBLM_R_X7Y116_SLICE_X8Y116_BO6;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_C = CLBLM_R_X7Y116_SLICE_X8Y116_CO6;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_D = CLBLM_R_X7Y116_SLICE_X8Y116_DO6;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_A = CLBLM_R_X7Y116_SLICE_X9Y116_AO6;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_B = CLBLM_R_X7Y116_SLICE_X9Y116_BO6;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_C = CLBLM_R_X7Y116_SLICE_X9Y116_CO6;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_D = CLBLM_R_X7Y116_SLICE_X9Y116_DO6;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_BMUX = CLBLM_R_X7Y116_SLICE_X9Y116_BO5;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_A = CLBLM_R_X7Y117_SLICE_X8Y117_AO6;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_B = CLBLM_R_X7Y117_SLICE_X8Y117_BO6;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_C = CLBLM_R_X7Y117_SLICE_X8Y117_CO6;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_D = CLBLM_R_X7Y117_SLICE_X8Y117_DO6;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_A = CLBLM_R_X7Y117_SLICE_X9Y117_AO6;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_B = CLBLM_R_X7Y117_SLICE_X9Y117_BO6;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_C = CLBLM_R_X7Y117_SLICE_X9Y117_CO6;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_D = CLBLM_R_X7Y117_SLICE_X9Y117_DO6;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_AMUX = CLBLM_R_X7Y117_SLICE_X9Y117_A5Q;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_CMUX = CLBLM_R_X7Y117_SLICE_X9Y117_CO5;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_A = CLBLM_R_X7Y118_SLICE_X8Y118_AO6;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_B = CLBLM_R_X7Y118_SLICE_X8Y118_BO6;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_C = CLBLM_R_X7Y118_SLICE_X8Y118_CO6;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_D = CLBLM_R_X7Y118_SLICE_X8Y118_DO6;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_A = CLBLM_R_X7Y118_SLICE_X9Y118_AO6;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_B = CLBLM_R_X7Y118_SLICE_X9Y118_BO6;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_C = CLBLM_R_X7Y118_SLICE_X9Y118_CO6;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_D = CLBLM_R_X7Y118_SLICE_X9Y118_DO6;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_BMUX = CLBLM_R_X7Y118_SLICE_X9Y118_BO5;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_CMUX = CLBLM_R_X7Y118_SLICE_X9Y118_CO5;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_A = CLBLM_R_X7Y132_SLICE_X8Y132_AO6;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_B = CLBLM_R_X7Y132_SLICE_X8Y132_BO6;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_C = CLBLM_R_X7Y132_SLICE_X8Y132_CO6;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_D = CLBLM_R_X7Y132_SLICE_X8Y132_DO6;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_A = CLBLM_R_X7Y132_SLICE_X9Y132_AO6;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_B = CLBLM_R_X7Y132_SLICE_X9Y132_BO6;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_C = CLBLM_R_X7Y132_SLICE_X9Y132_CO6;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_D = CLBLM_R_X7Y132_SLICE_X9Y132_DO6;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_AMUX = CLBLM_R_X7Y132_SLICE_X9Y132_AO5;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_A = CLBLM_R_X11Y105_SLICE_X14Y105_AO6;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_B = CLBLM_R_X11Y105_SLICE_X14Y105_BO6;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_C = CLBLM_R_X11Y105_SLICE_X14Y105_CO6;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_D = CLBLM_R_X11Y105_SLICE_X14Y105_DO6;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_CMUX = CLBLM_R_X11Y105_SLICE_X14Y105_C5Q;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_A = CLBLM_R_X11Y105_SLICE_X15Y105_AO6;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_B = CLBLM_R_X11Y105_SLICE_X15Y105_BO6;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_C = CLBLM_R_X11Y105_SLICE_X15Y105_CO6;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_D = CLBLM_R_X11Y105_SLICE_X15Y105_DO6;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_AMUX = CLBLM_R_X11Y105_SLICE_X15Y105_A5Q;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_DMUX = CLBLM_R_X11Y105_SLICE_X15Y105_DO5;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_A = CLBLM_R_X11Y106_SLICE_X14Y106_AO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_B = CLBLM_R_X11Y106_SLICE_X14Y106_BO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_C = CLBLM_R_X11Y106_SLICE_X14Y106_CO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_D = CLBLM_R_X11Y106_SLICE_X14Y106_DO6;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_A = CLBLM_R_X11Y106_SLICE_X15Y106_AO6;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_B = CLBLM_R_X11Y106_SLICE_X15Y106_BO6;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_C = CLBLM_R_X11Y106_SLICE_X15Y106_CO6;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_D = CLBLM_R_X11Y106_SLICE_X15Y106_DO6;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_BMUX = CLBLM_R_X11Y106_SLICE_X15Y106_BO5;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_CMUX = CLBLM_R_X11Y106_SLICE_X15Y106_CO5;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_DMUX = CLBLM_R_X11Y106_SLICE_X15Y106_DO5;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_A = CLBLM_R_X11Y107_SLICE_X14Y107_AO6;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_B = CLBLM_R_X11Y107_SLICE_X14Y107_BO6;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_C = CLBLM_R_X11Y107_SLICE_X14Y107_CO6;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_D = CLBLM_R_X11Y107_SLICE_X14Y107_DO6;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_AMUX = CLBLM_R_X11Y107_SLICE_X14Y107_AO5;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_A = CLBLM_R_X11Y107_SLICE_X15Y107_AO6;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_B = CLBLM_R_X11Y107_SLICE_X15Y107_BO6;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_C = CLBLM_R_X11Y107_SLICE_X15Y107_CO6;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_D = CLBLM_R_X11Y107_SLICE_X15Y107_DO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_A = CLBLM_R_X11Y108_SLICE_X14Y108_AO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_B = CLBLM_R_X11Y108_SLICE_X14Y108_BO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_C = CLBLM_R_X11Y108_SLICE_X14Y108_CO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_D = CLBLM_R_X11Y108_SLICE_X14Y108_DO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_BMUX = CLBLM_R_X11Y108_SLICE_X14Y108_BO6;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_A = CLBLM_R_X11Y108_SLICE_X15Y108_AO6;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_B = CLBLM_R_X11Y108_SLICE_X15Y108_BO6;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_C = CLBLM_R_X11Y108_SLICE_X15Y108_CO6;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_D = CLBLM_R_X11Y108_SLICE_X15Y108_DO6;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_AMUX = CLBLM_R_X11Y108_SLICE_X15Y108_AO5;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_BMUX = CLBLM_R_X11Y108_SLICE_X15Y108_BO5;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_CMUX = CLBLM_R_X11Y108_SLICE_X15Y108_CO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_A = CLBLM_R_X11Y109_SLICE_X14Y109_AO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_B = CLBLM_R_X11Y109_SLICE_X14Y109_BO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_C = CLBLM_R_X11Y109_SLICE_X14Y109_CO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_D = CLBLM_R_X11Y109_SLICE_X14Y109_DO6;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_A = CLBLM_R_X11Y109_SLICE_X15Y109_AO6;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_B = CLBLM_R_X11Y109_SLICE_X15Y109_BO6;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_C = CLBLM_R_X11Y109_SLICE_X15Y109_CO6;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_D = CLBLM_R_X11Y109_SLICE_X15Y109_DO6;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_AMUX = CLBLM_R_X11Y109_SLICE_X15Y109_AO5;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_CMUX = CLBLM_R_X11Y109_SLICE_X15Y109_CO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_A = CLBLM_R_X11Y110_SLICE_X14Y110_AO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_B = CLBLM_R_X11Y110_SLICE_X14Y110_BO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_C = CLBLM_R_X11Y110_SLICE_X14Y110_CO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_D = CLBLM_R_X11Y110_SLICE_X14Y110_DO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_AMUX = CLBLM_R_X11Y110_SLICE_X14Y110_A5Q;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_BMUX = CLBLM_R_X11Y110_SLICE_X14Y110_BO5;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_DMUX = CLBLM_R_X11Y110_SLICE_X14Y110_D5Q;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_A = CLBLM_R_X11Y110_SLICE_X15Y110_AO6;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_B = CLBLM_R_X11Y110_SLICE_X15Y110_BO6;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_C = CLBLM_R_X11Y110_SLICE_X15Y110_CO6;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_D = CLBLM_R_X11Y110_SLICE_X15Y110_DO6;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_AMUX = CLBLM_R_X11Y110_SLICE_X15Y110_A5Q;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_A = CLBLM_R_X11Y111_SLICE_X14Y111_AO6;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_B = CLBLM_R_X11Y111_SLICE_X14Y111_BO6;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_C = CLBLM_R_X11Y111_SLICE_X14Y111_CO6;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_D = CLBLM_R_X11Y111_SLICE_X14Y111_DO6;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_AMUX = CLBLM_R_X11Y111_SLICE_X14Y111_AO6;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_A = CLBLM_R_X11Y111_SLICE_X15Y111_AO6;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_B = CLBLM_R_X11Y111_SLICE_X15Y111_BO6;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_C = CLBLM_R_X11Y111_SLICE_X15Y111_CO6;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_D = CLBLM_R_X11Y111_SLICE_X15Y111_DO6;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_CMUX = CLBLM_R_X11Y111_SLICE_X15Y111_C5Q;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_A = CLBLM_R_X11Y112_SLICE_X14Y112_AO6;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_B = CLBLM_R_X11Y112_SLICE_X14Y112_BO6;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_C = CLBLM_R_X11Y112_SLICE_X14Y112_CO6;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_D = CLBLM_R_X11Y112_SLICE_X14Y112_DO6;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_AMUX = CLBLM_R_X11Y112_SLICE_X14Y112_AO5;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_BMUX = CLBLM_R_X11Y112_SLICE_X14Y112_B5Q;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_CMUX = CLBLM_R_X11Y112_SLICE_X14Y112_C5Q;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_A = CLBLM_R_X11Y112_SLICE_X15Y112_AO6;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_B = CLBLM_R_X11Y112_SLICE_X15Y112_BO6;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_C = CLBLM_R_X11Y112_SLICE_X15Y112_CO6;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_D = CLBLM_R_X11Y112_SLICE_X15Y112_DO6;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_A = CLBLM_R_X11Y113_SLICE_X14Y113_AO6;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_B = CLBLM_R_X11Y113_SLICE_X14Y113_BO6;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_C = CLBLM_R_X11Y113_SLICE_X14Y113_CO6;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_D = CLBLM_R_X11Y113_SLICE_X14Y113_DO6;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_A = CLBLM_R_X11Y113_SLICE_X15Y113_AO6;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_B = CLBLM_R_X11Y113_SLICE_X15Y113_BO6;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_C = CLBLM_R_X11Y113_SLICE_X15Y113_CO6;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_D = CLBLM_R_X11Y113_SLICE_X15Y113_DO6;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_A = CLBLM_R_X11Y114_SLICE_X14Y114_AO6;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_B = CLBLM_R_X11Y114_SLICE_X14Y114_BO6;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_C = CLBLM_R_X11Y114_SLICE_X14Y114_CO6;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_D = CLBLM_R_X11Y114_SLICE_X14Y114_DO6;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_A = CLBLM_R_X11Y114_SLICE_X15Y114_AO6;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_B = CLBLM_R_X11Y114_SLICE_X15Y114_BO6;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_C = CLBLM_R_X11Y114_SLICE_X15Y114_CO6;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_D = CLBLM_R_X11Y114_SLICE_X15Y114_DO6;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_A = CLBLM_R_X11Y115_SLICE_X14Y115_AO6;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_B = CLBLM_R_X11Y115_SLICE_X14Y115_BO6;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_C = CLBLM_R_X11Y115_SLICE_X14Y115_CO6;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_D = CLBLM_R_X11Y115_SLICE_X14Y115_DO6;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_AMUX = CLBLM_R_X11Y115_SLICE_X14Y115_AO5;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_BMUX = CLBLM_R_X11Y115_SLICE_X14Y115_BO5;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_A = CLBLM_R_X11Y115_SLICE_X15Y115_AO6;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_B = CLBLM_R_X11Y115_SLICE_X15Y115_BO6;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_C = CLBLM_R_X11Y115_SLICE_X15Y115_CO6;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_D = CLBLM_R_X11Y115_SLICE_X15Y115_DO6;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_BMUX = CLBLM_R_X11Y115_SLICE_X15Y115_B5Q;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_DMUX = CLBLM_R_X11Y115_SLICE_X15Y115_DO6;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_A = CLBLM_R_X11Y116_SLICE_X14Y116_AO6;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_B = CLBLM_R_X11Y116_SLICE_X14Y116_BO6;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_C = CLBLM_R_X11Y116_SLICE_X14Y116_CO6;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_D = CLBLM_R_X11Y116_SLICE_X14Y116_DO6;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_AMUX = CLBLM_R_X11Y116_SLICE_X14Y116_A5Q;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_A = CLBLM_R_X11Y116_SLICE_X15Y116_AO6;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_B = CLBLM_R_X11Y116_SLICE_X15Y116_BO6;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_C = CLBLM_R_X11Y116_SLICE_X15Y116_CO6;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_D = CLBLM_R_X11Y116_SLICE_X15Y116_DO6;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_A = CLBLM_R_X11Y117_SLICE_X14Y117_AO6;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_B = CLBLM_R_X11Y117_SLICE_X14Y117_BO6;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_C = CLBLM_R_X11Y117_SLICE_X14Y117_CO6;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_D = CLBLM_R_X11Y117_SLICE_X14Y117_DO6;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_A = CLBLM_R_X11Y117_SLICE_X15Y117_AO6;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_B = CLBLM_R_X11Y117_SLICE_X15Y117_BO6;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_C = CLBLM_R_X11Y117_SLICE_X15Y117_CO6;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_D = CLBLM_R_X11Y117_SLICE_X15Y117_DO6;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_BMUX = CLBLM_R_X11Y117_SLICE_X15Y117_BO5;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_A = CLBLM_R_X11Y118_SLICE_X14Y118_AO6;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_B = CLBLM_R_X11Y118_SLICE_X14Y118_BO6;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_C = CLBLM_R_X11Y118_SLICE_X14Y118_CO6;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_D = CLBLM_R_X11Y118_SLICE_X14Y118_DO6;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_A = CLBLM_R_X11Y118_SLICE_X15Y118_AO6;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_B = CLBLM_R_X11Y118_SLICE_X15Y118_BO6;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_C = CLBLM_R_X11Y118_SLICE_X15Y118_CO6;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_D = CLBLM_R_X11Y118_SLICE_X15Y118_DO6;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_AMUX = CLBLM_R_X11Y118_SLICE_X15Y118_A5Q;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_A = CLBLM_R_X11Y119_SLICE_X14Y119_AO6;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_B = CLBLM_R_X11Y119_SLICE_X14Y119_BO6;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_C = CLBLM_R_X11Y119_SLICE_X14Y119_CO6;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_D = CLBLM_R_X11Y119_SLICE_X14Y119_DO6;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_A = CLBLM_R_X11Y119_SLICE_X15Y119_AO6;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_B = CLBLM_R_X11Y119_SLICE_X15Y119_BO6;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_C = CLBLM_R_X11Y119_SLICE_X15Y119_CO6;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_D = CLBLM_R_X11Y119_SLICE_X15Y119_DO6;
  assign CLBLM_R_X13Y106_SLICE_X18Y106_A = CLBLM_R_X13Y106_SLICE_X18Y106_AO6;
  assign CLBLM_R_X13Y106_SLICE_X18Y106_B = CLBLM_R_X13Y106_SLICE_X18Y106_BO6;
  assign CLBLM_R_X13Y106_SLICE_X18Y106_C = CLBLM_R_X13Y106_SLICE_X18Y106_CO6;
  assign CLBLM_R_X13Y106_SLICE_X18Y106_D = CLBLM_R_X13Y106_SLICE_X18Y106_DO6;
  assign CLBLM_R_X13Y106_SLICE_X19Y106_A = CLBLM_R_X13Y106_SLICE_X19Y106_AO6;
  assign CLBLM_R_X13Y106_SLICE_X19Y106_B = CLBLM_R_X13Y106_SLICE_X19Y106_BO6;
  assign CLBLM_R_X13Y106_SLICE_X19Y106_C = CLBLM_R_X13Y106_SLICE_X19Y106_CO6;
  assign CLBLM_R_X13Y106_SLICE_X19Y106_D = CLBLM_R_X13Y106_SLICE_X19Y106_DO6;
  assign CLBLM_R_X13Y107_SLICE_X18Y107_A = CLBLM_R_X13Y107_SLICE_X18Y107_AO6;
  assign CLBLM_R_X13Y107_SLICE_X18Y107_B = CLBLM_R_X13Y107_SLICE_X18Y107_BO6;
  assign CLBLM_R_X13Y107_SLICE_X18Y107_C = CLBLM_R_X13Y107_SLICE_X18Y107_CO6;
  assign CLBLM_R_X13Y107_SLICE_X18Y107_D = CLBLM_R_X13Y107_SLICE_X18Y107_DO6;
  assign CLBLM_R_X13Y107_SLICE_X18Y107_BMUX = CLBLM_R_X13Y107_SLICE_X18Y107_BO6;
  assign CLBLM_R_X13Y107_SLICE_X19Y107_A = CLBLM_R_X13Y107_SLICE_X19Y107_AO6;
  assign CLBLM_R_X13Y107_SLICE_X19Y107_B = CLBLM_R_X13Y107_SLICE_X19Y107_BO6;
  assign CLBLM_R_X13Y107_SLICE_X19Y107_C = CLBLM_R_X13Y107_SLICE_X19Y107_CO6;
  assign CLBLM_R_X13Y107_SLICE_X19Y107_D = CLBLM_R_X13Y107_SLICE_X19Y107_DO6;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_A = CLBLM_R_X13Y108_SLICE_X18Y108_AO6;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_B = CLBLM_R_X13Y108_SLICE_X18Y108_BO6;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_C = CLBLM_R_X13Y108_SLICE_X18Y108_CO6;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_D = CLBLM_R_X13Y108_SLICE_X18Y108_DO6;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_BMUX = CLBLM_R_X13Y108_SLICE_X18Y108_BO5;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_CMUX = CLBLM_R_X13Y108_SLICE_X18Y108_CO6;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_A = CLBLM_R_X13Y108_SLICE_X19Y108_AO6;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_B = CLBLM_R_X13Y108_SLICE_X19Y108_BO6;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_C = CLBLM_R_X13Y108_SLICE_X19Y108_CO6;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_D = CLBLM_R_X13Y108_SLICE_X19Y108_DO6;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_A = CLBLM_R_X13Y109_SLICE_X18Y109_AO6;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_B = CLBLM_R_X13Y109_SLICE_X18Y109_BO6;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_C = CLBLM_R_X13Y109_SLICE_X18Y109_CO6;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_D = CLBLM_R_X13Y109_SLICE_X18Y109_DO6;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_BMUX = CLBLM_R_X13Y109_SLICE_X18Y109_BO5;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_A = CLBLM_R_X13Y109_SLICE_X19Y109_AO6;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_B = CLBLM_R_X13Y109_SLICE_X19Y109_BO6;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_C = CLBLM_R_X13Y109_SLICE_X19Y109_CO6;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_D = CLBLM_R_X13Y109_SLICE_X19Y109_DO6;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_A = CLBLM_R_X13Y110_SLICE_X18Y110_AO6;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_B = CLBLM_R_X13Y110_SLICE_X18Y110_BO6;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_C = CLBLM_R_X13Y110_SLICE_X18Y110_CO6;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_D = CLBLM_R_X13Y110_SLICE_X18Y110_DO6;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_DMUX = CLBLM_R_X13Y110_SLICE_X18Y110_DO5;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_A = CLBLM_R_X13Y110_SLICE_X19Y110_AO6;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_B = CLBLM_R_X13Y110_SLICE_X19Y110_BO6;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_C = CLBLM_R_X13Y110_SLICE_X19Y110_CO6;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_D = CLBLM_R_X13Y110_SLICE_X19Y110_DO6;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_A = CLBLM_R_X13Y112_SLICE_X18Y112_AO6;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_B = CLBLM_R_X13Y112_SLICE_X18Y112_BO6;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_C = CLBLM_R_X13Y112_SLICE_X18Y112_CO6;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_D = CLBLM_R_X13Y112_SLICE_X18Y112_DO6;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_AMUX = CLBLM_R_X13Y112_SLICE_X18Y112_A5Q;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_A = CLBLM_R_X13Y112_SLICE_X19Y112_AO6;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_B = CLBLM_R_X13Y112_SLICE_X19Y112_BO6;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_C = CLBLM_R_X13Y112_SLICE_X19Y112_CO6;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_D = CLBLM_R_X13Y112_SLICE_X19Y112_DO6;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_A = CLBLM_R_X13Y113_SLICE_X18Y113_AO6;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_B = CLBLM_R_X13Y113_SLICE_X18Y113_BO6;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_C = CLBLM_R_X13Y113_SLICE_X18Y113_CO6;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_D = CLBLM_R_X13Y113_SLICE_X18Y113_DO6;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_A = CLBLM_R_X13Y113_SLICE_X19Y113_AO6;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_B = CLBLM_R_X13Y113_SLICE_X19Y113_BO6;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_C = CLBLM_R_X13Y113_SLICE_X19Y113_CO6;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_D = CLBLM_R_X13Y113_SLICE_X19Y113_DO6;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_A = CLBLM_R_X13Y117_SLICE_X18Y117_AO6;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_B = CLBLM_R_X13Y117_SLICE_X18Y117_BO6;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_C = CLBLM_R_X13Y117_SLICE_X18Y117_CO6;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_D = CLBLM_R_X13Y117_SLICE_X18Y117_DO6;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_AMUX = CLBLM_R_X13Y117_SLICE_X18Y117_AO5;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_A = CLBLM_R_X13Y117_SLICE_X19Y117_AO6;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_B = CLBLM_R_X13Y117_SLICE_X19Y117_BO6;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_C = CLBLM_R_X13Y117_SLICE_X19Y117_CO6;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_D = CLBLM_R_X13Y117_SLICE_X19Y117_DO6;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_A = CLBLM_R_X13Y118_SLICE_X18Y118_AO6;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_B = CLBLM_R_X13Y118_SLICE_X18Y118_BO6;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_C = CLBLM_R_X13Y118_SLICE_X18Y118_CO6;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_D = CLBLM_R_X13Y118_SLICE_X18Y118_DO6;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_AMUX = CLBLM_R_X13Y118_SLICE_X18Y118_AO5;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_A = CLBLM_R_X13Y118_SLICE_X19Y118_AO6;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_B = CLBLM_R_X13Y118_SLICE_X19Y118_BO6;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_C = CLBLM_R_X13Y118_SLICE_X19Y118_CO6;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_D = CLBLM_R_X13Y118_SLICE_X19Y118_DO6;
  assign CLBLM_R_X37Y117_SLICE_X56Y117_A = CLBLM_R_X37Y117_SLICE_X56Y117_AO6;
  assign CLBLM_R_X37Y117_SLICE_X56Y117_B = CLBLM_R_X37Y117_SLICE_X56Y117_BO6;
  assign CLBLM_R_X37Y117_SLICE_X56Y117_C = CLBLM_R_X37Y117_SLICE_X56Y117_CO6;
  assign CLBLM_R_X37Y117_SLICE_X56Y117_D = CLBLM_R_X37Y117_SLICE_X56Y117_DO6;
  assign CLBLM_R_X37Y117_SLICE_X57Y117_A = CLBLM_R_X37Y117_SLICE_X57Y117_AO6;
  assign CLBLM_R_X37Y117_SLICE_X57Y117_B = CLBLM_R_X37Y117_SLICE_X57Y117_BO6;
  assign CLBLM_R_X37Y117_SLICE_X57Y117_C = CLBLM_R_X37Y117_SLICE_X57Y117_CO6;
  assign CLBLM_R_X37Y117_SLICE_X57Y117_D = CLBLM_R_X37Y117_SLICE_X57Y117_DO6;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_A = CLBLM_R_X103Y138_SLICE_X162Y138_AO6;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_B = CLBLM_R_X103Y138_SLICE_X162Y138_BO6;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_C = CLBLM_R_X103Y138_SLICE_X162Y138_CO6;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_D = CLBLM_R_X103Y138_SLICE_X162Y138_DO6;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_A = CLBLM_R_X103Y138_SLICE_X163Y138_AO6;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_B = CLBLM_R_X103Y138_SLICE_X163Y138_BO6;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_C = CLBLM_R_X103Y138_SLICE_X163Y138_CO6;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_D = CLBLM_R_X103Y138_SLICE_X163Y138_DO6;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_A = CLBLM_R_X103Y169_SLICE_X162Y169_AO6;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_B = CLBLM_R_X103Y169_SLICE_X162Y169_BO6;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_C = CLBLM_R_X103Y169_SLICE_X162Y169_CO6;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_D = CLBLM_R_X103Y169_SLICE_X162Y169_DO6;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_A = CLBLM_R_X103Y169_SLICE_X163Y169_AO6;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_B = CLBLM_R_X103Y169_SLICE_X163Y169_BO6;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_C = CLBLM_R_X103Y169_SLICE_X163Y169_CO6;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_D = CLBLM_R_X103Y169_SLICE_X163Y169_DO6;
  assign CLBLM_R_X103Y170_SLICE_X162Y170_A = CLBLM_R_X103Y170_SLICE_X162Y170_AO6;
  assign CLBLM_R_X103Y170_SLICE_X162Y170_B = CLBLM_R_X103Y170_SLICE_X162Y170_BO6;
  assign CLBLM_R_X103Y170_SLICE_X162Y170_C = CLBLM_R_X103Y170_SLICE_X162Y170_CO6;
  assign CLBLM_R_X103Y170_SLICE_X162Y170_D = CLBLM_R_X103Y170_SLICE_X162Y170_DO6;
  assign CLBLM_R_X103Y170_SLICE_X163Y170_A = CLBLM_R_X103Y170_SLICE_X163Y170_AO6;
  assign CLBLM_R_X103Y170_SLICE_X163Y170_B = CLBLM_R_X103Y170_SLICE_X163Y170_BO6;
  assign CLBLM_R_X103Y170_SLICE_X163Y170_C = CLBLM_R_X103Y170_SLICE_X163Y170_CO6;
  assign CLBLM_R_X103Y170_SLICE_X163Y170_D = CLBLM_R_X103Y170_SLICE_X163Y170_DO6;
  assign CLBLM_R_X103Y170_SLICE_X163Y170_AMUX = CLBLM_R_X103Y170_SLICE_X163Y170_AO5;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_A = CLBLM_R_X103Y173_SLICE_X162Y173_AO6;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_B = CLBLM_R_X103Y173_SLICE_X162Y173_BO6;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_C = CLBLM_R_X103Y173_SLICE_X162Y173_CO6;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_D = CLBLM_R_X103Y173_SLICE_X162Y173_DO6;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_A = CLBLM_R_X103Y173_SLICE_X163Y173_AO6;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_B = CLBLM_R_X103Y173_SLICE_X163Y173_BO6;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_C = CLBLM_R_X103Y173_SLICE_X163Y173_CO6;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_D = CLBLM_R_X103Y173_SLICE_X163Y173_DO6;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_AMUX = CLBLM_R_X103Y173_SLICE_X163Y173_AO5;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_A = CLBLM_R_X103Y174_SLICE_X162Y174_AO6;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_B = CLBLM_R_X103Y174_SLICE_X162Y174_BO6;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_C = CLBLM_R_X103Y174_SLICE_X162Y174_CO6;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_D = CLBLM_R_X103Y174_SLICE_X162Y174_DO6;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_A = CLBLM_R_X103Y174_SLICE_X163Y174_AO6;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_B = CLBLM_R_X103Y174_SLICE_X163Y174_BO6;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_C = CLBLM_R_X103Y174_SLICE_X163Y174_CO6;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_D = CLBLM_R_X103Y174_SLICE_X163Y174_DO6;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_AMUX = CLBLM_R_X103Y174_SLICE_X163Y174_AO5;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_A = CLBLM_R_X103Y177_SLICE_X162Y177_AO6;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_B = CLBLM_R_X103Y177_SLICE_X162Y177_BO6;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_C = CLBLM_R_X103Y177_SLICE_X162Y177_CO6;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_D = CLBLM_R_X103Y177_SLICE_X162Y177_DO6;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_A = CLBLM_R_X103Y177_SLICE_X163Y177_AO6;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_B = CLBLM_R_X103Y177_SLICE_X163Y177_BO6;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_C = CLBLM_R_X103Y177_SLICE_X163Y177_CO6;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_D = CLBLM_R_X103Y177_SLICE_X163Y177_DO6;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_AMUX = CLBLM_R_X103Y177_SLICE_X163Y177_AO5;
  assign LIOI3_X0Y51_ILOGIC_X0Y52_O = LIOB33_X0Y51_IOB_X0Y52_I;
  assign LIOI3_X0Y51_ILOGIC_X0Y51_O = LIOB33_X0Y51_IOB_X0Y51_I;
  assign LIOI3_X0Y53_ILOGIC_X0Y54_O = LIOB33_X0Y53_IOB_X0Y54_I;
  assign LIOI3_X0Y53_ILOGIC_X0Y53_O = LIOB33_X0Y53_IOB_X0Y53_I;
  assign LIOI3_X0Y55_ILOGIC_X0Y56_O = LIOB33_X0Y55_IOB_X0Y56_I;
  assign LIOI3_X0Y55_ILOGIC_X0Y55_O = LIOB33_X0Y55_IOB_X0Y55_I;
  assign LIOI3_X0Y59_ILOGIC_X0Y60_O = LIOB33_X0Y59_IOB_X0Y60_I;
  assign LIOI3_X0Y59_ILOGIC_X0Y59_O = LIOB33_X0Y59_IOB_X0Y59_I;
  assign LIOI3_X0Y61_ILOGIC_X0Y62_O = LIOB33_X0Y61_IOB_X0Y62_I;
  assign LIOI3_X0Y61_ILOGIC_X0Y61_O = LIOB33_X0Y61_IOB_X0Y61_I;
  assign LIOI3_X0Y65_ILOGIC_X0Y66_O = LIOB33_X0Y65_IOB_X0Y66_I;
  assign LIOI3_X0Y65_ILOGIC_X0Y65_O = LIOB33_X0Y65_IOB_X0Y65_I;
  assign LIOI3_X0Y67_ILOGIC_X0Y68_O = LIOB33_X0Y67_IOB_X0Y68_I;
  assign LIOI3_X0Y67_ILOGIC_X0Y67_O = LIOB33_X0Y67_IOB_X0Y67_I;
  assign LIOI3_X0Y71_ILOGIC_X0Y72_O = LIOB33_X0Y71_IOB_X0Y72_I;
  assign LIOI3_X0Y71_ILOGIC_X0Y71_O = LIOB33_X0Y71_IOB_X0Y71_I;
  assign LIOI3_X0Y73_ILOGIC_X0Y74_O = LIOB33_X0Y73_IOB_X0Y74_I;
  assign LIOI3_X0Y73_ILOGIC_X0Y73_O = LIOB33_X0Y73_IOB_X0Y73_I;
  assign LIOI3_X0Y75_ILOGIC_X0Y76_O = LIOB33_X0Y75_IOB_X0Y76_I;
  assign LIOI3_X0Y75_ILOGIC_X0Y75_O = LIOB33_X0Y75_IOB_X0Y75_I;
  assign LIOI3_X0Y77_ILOGIC_X0Y78_O = LIOB33_X0Y77_IOB_X0Y78_I;
  assign LIOI3_X0Y77_ILOGIC_X0Y77_O = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOI3_X0Y79_ILOGIC_X0Y79_O = LIOB33_X0Y79_IOB_X0Y79_I;
  assign LIOI3_X0Y79_OLOGIC_X0Y80_OQ = CLBLL_L_X2Y106_SLICE_X0Y106_AO6;
  assign LIOI3_X0Y79_OLOGIC_X0Y80_TQ = 1'b1;
  assign LIOI3_X0Y101_OLOGIC_X0Y102_OQ = CLBLL_L_X2Y106_SLICE_X0Y106_BO5;
  assign LIOI3_X0Y101_OLOGIC_X0Y102_TQ = 1'b1;
  assign LIOI3_X0Y101_OLOGIC_X0Y101_OQ = CLBLL_L_X2Y107_SLICE_X0Y107_AO6;
  assign LIOI3_X0Y101_OLOGIC_X0Y101_TQ = 1'b1;
  assign LIOI3_X0Y103_OLOGIC_X0Y104_OQ = CLBLL_L_X2Y106_SLICE_X0Y106_CO6;
  assign LIOI3_X0Y103_OLOGIC_X0Y104_TQ = 1'b1;
  assign LIOI3_X0Y103_OLOGIC_X0Y103_OQ = CLBLM_R_X3Y107_SLICE_X3Y107_BO6;
  assign LIOI3_X0Y103_OLOGIC_X0Y103_TQ = 1'b1;
  assign LIOI3_X0Y105_OLOGIC_X0Y106_OQ = CLBLL_L_X2Y106_SLICE_X0Y106_AO5;
  assign LIOI3_X0Y105_OLOGIC_X0Y106_TQ = 1'b1;
  assign LIOI3_X0Y105_OLOGIC_X0Y105_OQ = CLBLL_L_X2Y106_SLICE_X0Y106_CO5;
  assign LIOI3_X0Y105_OLOGIC_X0Y105_TQ = 1'b1;
  assign LIOI3_X0Y109_OLOGIC_X0Y110_OQ = CLBLM_R_X3Y106_SLICE_X2Y106_AO6;
  assign LIOI3_X0Y109_OLOGIC_X0Y110_TQ = 1'b1;
  assign LIOI3_X0Y109_OLOGIC_X0Y109_OQ = CLBLL_L_X2Y107_SLICE_X1Y107_AO5;
  assign LIOI3_X0Y109_OLOGIC_X0Y109_TQ = 1'b1;
  assign LIOI3_X0Y111_OLOGIC_X0Y112_OQ = CLBLM_R_X11Y110_SLICE_X14Y110_D5Q;
  assign LIOI3_X0Y111_OLOGIC_X0Y112_TQ = 1'b1;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_OQ = 1'b0;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_TQ = 1'b1;
  assign LIOI3_X0Y115_OLOGIC_X0Y116_OQ = CLBLM_R_X11Y118_SLICE_X15Y118_AQ;
  assign LIOI3_X0Y115_OLOGIC_X0Y116_TQ = 1'b1;
  assign LIOI3_X0Y115_OLOGIC_X0Y115_OQ = CLBLM_R_X11Y110_SLICE_X14Y110_DQ;
  assign LIOI3_X0Y115_OLOGIC_X0Y115_TQ = 1'b1;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_OQ = CLBLM_R_X5Y114_SLICE_X7Y114_CQ;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_TQ = 1'b1;
  assign LIOI3_X0Y117_OLOGIC_X0Y117_OQ = CLBLL_L_X4Y116_SLICE_X5Y116_BQ;
  assign LIOI3_X0Y117_OLOGIC_X0Y117_TQ = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_OQ = CLBLM_R_X5Y116_SLICE_X7Y116_A5Q;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_TQ = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_OQ = CLBLM_R_X11Y118_SLICE_X15Y118_A5Q;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_TQ = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_OQ = CLBLM_R_X5Y114_SLICE_X7Y114_C5Q;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_TQ = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_OQ = CLBLM_R_X7Y113_SLICE_X8Y113_C5Q;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_TQ = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_OQ = CLBLL_L_X4Y117_SLICE_X4Y117_CQ;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_TQ = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_OQ = CLBLM_R_X11Y115_SLICE_X15Y115_B5Q;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_TQ = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_OQ = CLBLM_R_X3Y115_SLICE_X2Y115_AQ;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_TQ = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_OQ = CLBLL_L_X4Y113_SLICE_X4Y113_BQ;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_TQ = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_OQ = CLBLL_L_X52Y126_SLICE_X78Y126_AO6;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_TQ = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_OQ = CLBLM_R_X5Y109_SLICE_X6Y109_CQ;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_TQ = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_OQ = CLBLL_L_X4Y116_SLICE_X5Y116_AQ;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_TQ = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_OQ = CLBLL_L_X4Y118_SLICE_X4Y118_A5Q;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_TQ = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_OQ = CLBLL_L_X4Y117_SLICE_X4Y117_DQ;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_TQ = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_OQ = CLBLL_L_X4Y118_SLICE_X4Y118_AQ;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_TQ = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_OQ = CLBLL_L_X4Y116_SLICE_X4Y116_AQ;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_TQ = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_OQ = CLBLL_L_X4Y118_SLICE_X4Y118_BQ;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_TQ = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_OQ = LIOB33_X0Y53_IOB_X0Y54_I;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_TQ = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_OQ = CLBLL_L_X4Y117_SLICE_X4Y117_BQ;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_TQ = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_OQ = LIOB33_X0Y59_IOB_X0Y59_I;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_TQ = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_OQ = LIOB33_X0Y57_IOB_X0Y58_I;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_TQ = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_OQ = LIOB33_X0Y61_IOB_X0Y61_I;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_TQ = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_OQ = LIOB33_X0Y71_IOB_X0Y71_I;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_TQ = 1'b1;
  assign LIOI3_X0Y151_OLOGIC_X0Y152_OQ = LIOB33_X0Y65_IOB_X0Y66_I;
  assign LIOI3_X0Y151_OLOGIC_X0Y152_TQ = 1'b1;
  assign LIOI3_X0Y151_OLOGIC_X0Y151_OQ = LIOB33_X0Y65_IOB_X0Y65_I;
  assign LIOI3_X0Y151_OLOGIC_X0Y151_TQ = 1'b1;
  assign LIOI3_X0Y153_OLOGIC_X0Y154_OQ = LIOB33_X0Y67_IOB_X0Y68_I;
  assign LIOI3_X0Y153_OLOGIC_X0Y154_TQ = 1'b1;
  assign LIOI3_X0Y153_OLOGIC_X0Y153_OQ = LIOB33_X0Y67_IOB_X0Y67_I;
  assign LIOI3_X0Y153_OLOGIC_X0Y153_TQ = 1'b1;
  assign LIOI3_X0Y155_OLOGIC_X0Y156_OQ = RIOB33_X105Y105_IOB_X1Y106_I;
  assign LIOI3_X0Y155_OLOGIC_X0Y156_TQ = 1'b1;
  assign LIOI3_X0Y155_OLOGIC_X0Y155_OQ = LIOB33_X0Y69_IOB_X0Y70_I;
  assign LIOI3_X0Y155_OLOGIC_X0Y155_TQ = 1'b1;
  assign LIOI3_X0Y159_OLOGIC_X0Y160_OQ = RIOB33_X105Y107_IOB_X1Y107_I;
  assign LIOI3_X0Y159_OLOGIC_X0Y160_TQ = 1'b1;
  assign LIOI3_X0Y159_OLOGIC_X0Y159_OQ = RIOB33_X105Y117_IOB_X1Y117_I;
  assign LIOI3_X0Y159_OLOGIC_X0Y159_TQ = 1'b1;
  assign LIOI3_X0Y161_OLOGIC_X0Y162_OQ = RIOB33_X105Y109_IOB_X1Y109_I;
  assign LIOI3_X0Y161_OLOGIC_X0Y162_TQ = 1'b1;
  assign LIOI3_X0Y161_OLOGIC_X0Y161_OQ = RIOB33_X105Y107_IOB_X1Y108_I;
  assign LIOI3_X0Y161_OLOGIC_X0Y161_TQ = 1'b1;
  assign LIOI3_X0Y165_OLOGIC_X0Y166_OQ = RIOB33_X105Y113_IOB_X1Y113_I;
  assign LIOI3_X0Y165_OLOGIC_X0Y166_TQ = 1'b1;
  assign LIOI3_X0Y165_OLOGIC_X0Y165_OQ = RIOB33_X105Y111_IOB_X1Y112_I;
  assign LIOI3_X0Y165_OLOGIC_X0Y165_TQ = 1'b1;
  assign LIOI3_X0Y167_OLOGIC_X0Y168_OQ = RIOB33_X105Y123_IOB_X1Y123_I;
  assign LIOI3_X0Y167_OLOGIC_X0Y168_TQ = 1'b1;
  assign LIOI3_X0Y167_OLOGIC_X0Y167_OQ = RIOB33_X105Y113_IOB_X1Y114_I;
  assign LIOI3_X0Y167_OLOGIC_X0Y167_TQ = 1'b1;
  assign LIOI3_X0Y171_OLOGIC_X0Y172_OQ = CLBLM_R_X103Y138_SLICE_X163Y138_AO6;
  assign LIOI3_X0Y171_OLOGIC_X0Y172_TQ = 1'b1;
  assign LIOI3_X0Y171_OLOGIC_X0Y171_OQ = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign LIOI3_X0Y171_OLOGIC_X0Y171_TQ = 1'b1;
  assign LIOI3_X0Y173_OLOGIC_X0Y174_OQ = CLBLM_L_X10Y148_SLICE_X12Y148_AO6;
  assign LIOI3_X0Y173_OLOGIC_X0Y174_TQ = 1'b1;
  assign LIOI3_X0Y173_OLOGIC_X0Y173_OQ = CLBLM_R_X7Y132_SLICE_X9Y132_AO5;
  assign LIOI3_X0Y173_OLOGIC_X0Y173_TQ = 1'b1;
  assign LIOI3_X0Y175_OLOGIC_X0Y176_OQ = RIOB33_X105Y127_IOB_X1Y128_I;
  assign LIOI3_X0Y175_OLOGIC_X0Y176_TQ = 1'b1;
  assign LIOI3_X0Y175_OLOGIC_X0Y175_OQ = RIOB33_X105Y127_IOB_X1Y127_I;
  assign LIOI3_X0Y175_OLOGIC_X0Y175_TQ = 1'b1;
  assign LIOI3_X0Y177_OLOGIC_X0Y178_OQ = RIOB33_X105Y129_IOB_X1Y130_I;
  assign LIOI3_X0Y177_OLOGIC_X0Y178_TQ = 1'b1;
  assign LIOI3_X0Y177_OLOGIC_X0Y177_OQ = RIOB33_X105Y129_IOB_X1Y129_I;
  assign LIOI3_X0Y177_OLOGIC_X0Y177_TQ = 1'b1;
  assign LIOI3_X0Y179_OLOGIC_X0Y180_OQ = RIOB33_X105Y131_IOB_X1Y132_I;
  assign LIOI3_X0Y179_OLOGIC_X0Y180_TQ = 1'b1;
  assign LIOI3_X0Y179_OLOGIC_X0Y179_OQ = RIOB33_X105Y131_IOB_X1Y131_I;
  assign LIOI3_X0Y179_OLOGIC_X0Y179_TQ = 1'b1;
  assign LIOI3_X0Y183_OLOGIC_X0Y184_OQ = RIOB33_X105Y135_IOB_X1Y136_I;
  assign LIOI3_X0Y183_OLOGIC_X0Y184_TQ = 1'b1;
  assign LIOI3_X0Y183_OLOGIC_X0Y183_OQ = RIOB33_X105Y135_IOB_X1Y135_I;
  assign LIOI3_X0Y183_OLOGIC_X0Y183_TQ = 1'b1;
  assign LIOI3_X0Y185_OLOGIC_X0Y186_OQ = RIOB33_X105Y143_IOB_X1Y143_I;
  assign LIOI3_X0Y185_OLOGIC_X0Y186_TQ = 1'b1;
  assign LIOI3_X0Y185_OLOGIC_X0Y185_OQ = RIOB33_X105Y137_IOB_X1Y137_I;
  assign LIOI3_X0Y185_OLOGIC_X0Y185_TQ = 1'b1;
  assign LIOI3_X0Y189_OLOGIC_X0Y190_OQ = RIOB33_X105Y147_IOB_X1Y147_I;
  assign LIOI3_X0Y189_OLOGIC_X0Y190_TQ = 1'b1;
  assign LIOI3_X0Y189_OLOGIC_X0Y189_OQ = RIOB33_X105Y145_IOB_X1Y146_I;
  assign LIOI3_X0Y189_OLOGIC_X0Y189_TQ = 1'b1;
  assign LIOI3_X0Y191_OLOGIC_X0Y192_OQ = LIOB33_X0Y51_IOB_X0Y52_I;
  assign LIOI3_X0Y191_OLOGIC_X0Y192_TQ = 1'b1;
  assign LIOI3_X0Y191_OLOGIC_X0Y191_OQ = RIOB33_X105Y147_IOB_X1Y148_I;
  assign LIOI3_X0Y191_OLOGIC_X0Y191_TQ = 1'b1;
  assign LIOI3_X0Y195_OLOGIC_X0Y196_OQ = LIOB33_X0Y69_IOB_X0Y69_I;
  assign LIOI3_X0Y195_OLOGIC_X0Y196_TQ = 1'b1;
  assign LIOI3_X0Y195_OLOGIC_X0Y195_OQ = LIOB33_X0Y63_IOB_X0Y64_I;
  assign LIOI3_X0Y195_OLOGIC_X0Y195_TQ = 1'b1;
  assign LIOI3_X0Y197_OLOGIC_X0Y198_OQ = LIOB33_X0Y73_IOB_X0Y73_I;
  assign LIOI3_X0Y197_OLOGIC_X0Y198_TQ = 1'b1;
  assign LIOI3_X0Y197_OLOGIC_X0Y197_OQ = LIOB33_X0Y71_IOB_X0Y72_I;
  assign LIOI3_X0Y197_OLOGIC_X0Y197_TQ = 1'b1;
  assign LIOI3_SING_X0Y50_ILOGIC_X0Y50_O = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign LIOI3_SING_X0Y100_OLOGIC_X0Y100_OQ = CLBLL_L_X2Y106_SLICE_X0Y106_BO6;
  assign LIOI3_SING_X0Y100_OLOGIC_X0Y100_TQ = 1'b1;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_OQ = LIOB33_X0Y61_IOB_X0Y62_I;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_TQ = 1'b1;
  assign LIOI3_SING_X0Y150_OLOGIC_X0Y150_OQ = LIOB33_X0Y63_IOB_X0Y63_I;
  assign LIOI3_SING_X0Y150_OLOGIC_X0Y150_TQ = 1'b1;
  assign LIOI3_SING_X0Y199_OLOGIC_X0Y199_OQ = LIOB33_X0Y73_IOB_X0Y74_I;
  assign LIOI3_SING_X0Y199_OLOGIC_X0Y199_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y58_O = LIOB33_X0Y57_IOB_X0Y58_I;
  assign LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y57_O = LIOB33_X0Y57_IOB_X0Y57_I;
  assign LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y70_O = LIOB33_X0Y69_IOB_X0Y70_I;
  assign LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y69_O = LIOB33_X0Y69_IOB_X0Y69_I;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_OQ = CLBLL_L_X2Y107_SLICE_X0Y107_AO5;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_OQ = CLBLM_R_X3Y106_SLICE_X2Y106_BO6;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_OQ = CLBLM_R_X13Y112_SLICE_X18Y112_AQ;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_OQ = CLBLM_L_X10Y111_SLICE_X13Y111_CQ;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_OQ = CLBLM_L_X8Y119_SLICE_X10Y119_AQ;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_OQ = CLBLM_L_X8Y119_SLICE_X10Y119_AO5;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_OQ = LIOB33_X0Y57_IOB_X0Y57_I;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_OQ = LIOB33_X0Y55_IOB_X0Y55_I;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_OQ = RIOB33_X105Y115_IOB_X1Y116_I;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_OQ = RIOB33_X105Y115_IOB_X1Y115_I;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_OQ = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_OQ = RIOB33_X105Y121_IOB_X1Y122_I;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_OQ = RIOB33_X105Y133_IOB_X1Y134_I;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_OQ = RIOB33_X105Y133_IOB_X1Y133_I;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_OQ = LIOB33_X0Y59_IOB_X0Y60_I;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_OQ = LIOB33_X0Y55_IOB_X0Y56_I;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y64_O = LIOB33_X0Y63_IOB_X0Y64_I;
  assign LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y63_O = LIOB33_X0Y63_IOB_X0Y63_I;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_OQ = CLBLM_R_X7Y113_SLICE_X8Y113_CQ;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_OQ = RIOB33_X105Y121_IOB_X1Y121_I;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_OQ = CLBLL_L_X4Y117_SLICE_X5Y117_AQ;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_OQ = CLBLL_L_X4Y117_SLICE_X4Y117_AQ;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_OQ = RIOB33_X105Y111_IOB_X1Y111_I;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_OQ = RIOB33_X105Y109_IOB_X1Y110_I;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_OQ = RIOB33_X105Y145_IOB_X1Y145_I;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_OQ = RIOB33_X105Y143_IOB_X1Y144_I;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_TQ = 1'b1;
  assign RIOI3_X105Y101_ILOGIC_X1Y102_O = RIOB33_X105Y101_IOB_X1Y102_I;
  assign RIOI3_X105Y101_ILOGIC_X1Y101_O = RIOB33_X105Y101_IOB_X1Y101_I;
  assign RIOI3_X105Y103_ILOGIC_X1Y104_O = RIOB33_X105Y103_IOB_X1Y104_I;
  assign RIOI3_X105Y103_ILOGIC_X1Y103_O = RIOB33_X105Y103_IOB_X1Y103_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y106_O = RIOB33_X105Y105_IOB_X1Y106_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y105_O = RIOB33_X105Y105_IOB_X1Y105_I;
  assign RIOI3_X105Y109_ILOGIC_X1Y110_O = RIOB33_X105Y109_IOB_X1Y110_I;
  assign RIOI3_X105Y109_ILOGIC_X1Y109_O = RIOB33_X105Y109_IOB_X1Y109_I;
  assign RIOI3_X105Y111_ILOGIC_X1Y112_O = RIOB33_X105Y111_IOB_X1Y112_I;
  assign RIOI3_X105Y111_ILOGIC_X1Y111_O = RIOB33_X105Y111_IOB_X1Y111_I;
  assign RIOI3_X105Y115_ILOGIC_X1Y116_O = RIOB33_X105Y115_IOB_X1Y116_I;
  assign RIOI3_X105Y115_ILOGIC_X1Y115_O = RIOB33_X105Y115_IOB_X1Y115_I;
  assign RIOI3_X105Y117_ILOGIC_X1Y118_O = RIOB33_X105Y117_IOB_X1Y118_I;
  assign RIOI3_X105Y117_ILOGIC_X1Y117_O = RIOB33_X105Y117_IOB_X1Y117_I;
  assign RIOI3_X105Y121_ILOGIC_X1Y122_O = RIOB33_X105Y121_IOB_X1Y122_I;
  assign RIOI3_X105Y121_ILOGIC_X1Y121_O = RIOB33_X105Y121_IOB_X1Y121_I;
  assign RIOI3_X105Y123_ILOGIC_X1Y124_O = RIOB33_X105Y123_IOB_X1Y124_I;
  assign RIOI3_X105Y123_ILOGIC_X1Y123_O = RIOB33_X105Y123_IOB_X1Y123_I;
  assign RIOI3_X105Y125_ILOGIC_X1Y126_O = RIOB33_X105Y125_IOB_X1Y126_I;
  assign RIOI3_X105Y125_ILOGIC_X1Y125_O = RIOB33_X105Y125_IOB_X1Y125_I;
  assign RIOI3_X105Y127_ILOGIC_X1Y128_O = RIOB33_X105Y127_IOB_X1Y128_I;
  assign RIOI3_X105Y127_ILOGIC_X1Y127_O = RIOB33_X105Y127_IOB_X1Y127_I;
  assign RIOI3_X105Y129_ILOGIC_X1Y130_O = RIOB33_X105Y129_IOB_X1Y130_I;
  assign RIOI3_X105Y129_ILOGIC_X1Y129_O = RIOB33_X105Y129_IOB_X1Y129_I;
  assign RIOI3_X105Y133_ILOGIC_X1Y134_O = RIOB33_X105Y133_IOB_X1Y134_I;
  assign RIOI3_X105Y133_ILOGIC_X1Y133_O = RIOB33_X105Y133_IOB_X1Y133_I;
  assign RIOI3_X105Y135_ILOGIC_X1Y136_O = RIOB33_X105Y135_IOB_X1Y136_I;
  assign RIOI3_X105Y135_ILOGIC_X1Y135_O = RIOB33_X105Y135_IOB_X1Y135_I;
  assign RIOI3_X105Y139_ILOGIC_X1Y140_O = RIOB33_X105Y139_IOB_X1Y140_I;
  assign RIOI3_X105Y139_ILOGIC_X1Y139_O = RIOB33_X105Y139_IOB_X1Y139_I;
  assign RIOI3_X105Y141_ILOGIC_X1Y142_O = RIOB33_X105Y141_IOB_X1Y142_I;
  assign RIOI3_X105Y141_ILOGIC_X1Y141_O = RIOB33_X105Y141_IOB_X1Y141_I;
  assign RIOI3_X105Y145_ILOGIC_X1Y146_O = RIOB33_X105Y145_IOB_X1Y146_I;
  assign RIOI3_X105Y145_ILOGIC_X1Y145_O = RIOB33_X105Y145_IOB_X1Y145_I;
  assign RIOI3_X105Y147_ILOGIC_X1Y148_O = RIOB33_X105Y147_IOB_X1Y148_I;
  assign RIOI3_X105Y147_ILOGIC_X1Y147_O = RIOB33_X105Y147_IOB_X1Y147_I;
  assign RIOI3_X105Y151_OLOGIC_X1Y152_OQ = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign RIOI3_X105Y151_OLOGIC_X1Y152_TQ = 1'b1;
  assign RIOI3_X105Y151_OLOGIC_X1Y151_OQ = LIOB33_X0Y75_IOB_X0Y76_I;
  assign RIOI3_X105Y151_OLOGIC_X1Y151_TQ = 1'b1;
  assign RIOI3_X105Y153_OLOGIC_X1Y154_OQ = RIOB33_X105Y101_IOB_X1Y102_I;
  assign RIOI3_X105Y153_OLOGIC_X1Y154_TQ = 1'b1;
  assign RIOI3_X105Y153_OLOGIC_X1Y153_OQ = RIOB33_X105Y101_IOB_X1Y101_I;
  assign RIOI3_X105Y153_OLOGIC_X1Y153_TQ = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y156_OQ = RIOB33_X105Y103_IOB_X1Y104_I;
  assign RIOI3_X105Y155_OLOGIC_X1Y156_TQ = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y155_OQ = RIOB33_X105Y103_IOB_X1Y103_I;
  assign RIOI3_X105Y155_OLOGIC_X1Y155_TQ = 1'b1;
  assign RIOI3_X105Y159_OLOGIC_X1Y160_OQ = CLBLM_R_X13Y110_SLICE_X18Y110_DO5;
  assign RIOI3_X105Y159_OLOGIC_X1Y160_TQ = 1'b1;
  assign RIOI3_X105Y159_OLOGIC_X1Y159_OQ = CLBLM_R_X13Y110_SLICE_X18Y110_DO6;
  assign RIOI3_X105Y159_OLOGIC_X1Y159_TQ = 1'b1;
  assign RIOI3_X105Y161_OLOGIC_X1Y162_OQ = CLBLM_L_X12Y114_SLICE_X16Y114_DO5;
  assign RIOI3_X105Y161_OLOGIC_X1Y162_TQ = 1'b1;
  assign RIOI3_X105Y161_OLOGIC_X1Y161_OQ = CLBLM_L_X12Y114_SLICE_X16Y114_DO6;
  assign RIOI3_X105Y161_OLOGIC_X1Y161_TQ = 1'b1;
  assign RIOI3_X105Y165_OLOGIC_X1Y166_OQ = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign RIOI3_X105Y165_OLOGIC_X1Y166_TQ = 1'b1;
  assign RIOI3_X105Y165_OLOGIC_X1Y165_OQ = RIOB33_X105Y125_IOB_X1Y125_I;
  assign RIOI3_X105Y165_OLOGIC_X1Y165_TQ = 1'b1;
  assign RIOI3_X105Y167_OLOGIC_X1Y168_OQ = CLBLM_L_X10Y148_SLICE_X12Y148_AO6;
  assign RIOI3_X105Y167_OLOGIC_X1Y168_TQ = 1'b1;
  assign RIOI3_X105Y167_OLOGIC_X1Y167_OQ = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign RIOI3_X105Y167_OLOGIC_X1Y167_TQ = 1'b1;
  assign RIOI3_X105Y171_OLOGIC_X1Y172_OQ = CLBLM_R_X103Y173_SLICE_X163Y173_AO6;
  assign RIOI3_X105Y171_OLOGIC_X1Y172_TQ = 1'b1;
  assign RIOI3_X105Y171_OLOGIC_X1Y171_OQ = CLBLM_R_X103Y170_SLICE_X163Y170_AO5;
  assign RIOI3_X105Y171_OLOGIC_X1Y171_TQ = 1'b1;
  assign RIOI3_X105Y173_OLOGIC_X1Y174_OQ = CLBLM_R_X103Y174_SLICE_X163Y174_AO6;
  assign RIOI3_X105Y173_OLOGIC_X1Y174_TQ = 1'b1;
  assign RIOI3_X105Y173_OLOGIC_X1Y173_OQ = CLBLM_R_X103Y173_SLICE_X163Y173_AO5;
  assign RIOI3_X105Y173_OLOGIC_X1Y173_TQ = 1'b1;
  assign RIOI3_X105Y175_OLOGIC_X1Y176_OQ = CLBLM_R_X103Y174_SLICE_X163Y174_AO5;
  assign RIOI3_X105Y175_OLOGIC_X1Y176_TQ = 1'b1;
  assign RIOI3_X105Y175_OLOGIC_X1Y175_OQ = CLBLM_R_X13Y118_SLICE_X18Y118_AO6;
  assign RIOI3_X105Y175_OLOGIC_X1Y175_TQ = 1'b1;
  assign RIOI3_X105Y177_OLOGIC_X1Y178_OQ = CLBLM_R_X103Y177_SLICE_X163Y177_AO5;
  assign RIOI3_X105Y177_OLOGIC_X1Y178_TQ = 1'b1;
  assign RIOI3_X105Y177_OLOGIC_X1Y177_OQ = CLBLM_R_X103Y177_SLICE_X163Y177_AO6;
  assign RIOI3_X105Y177_OLOGIC_X1Y177_TQ = 1'b1;
  assign RIOI3_X105Y179_OLOGIC_X1Y180_OQ = CLBLM_R_X13Y110_SLICE_X18Y110_DO6;
  assign RIOI3_X105Y179_OLOGIC_X1Y180_TQ = 1'b1;
  assign RIOI3_X105Y179_OLOGIC_X1Y179_OQ = CLBLM_R_X13Y117_SLICE_X18Y117_AO5;
  assign RIOI3_X105Y179_OLOGIC_X1Y179_TQ = 1'b1;
  assign RIOI3_X105Y183_OLOGIC_X1Y184_OQ = CLBLM_L_X8Y110_SLICE_X10Y110_CO6;
  assign RIOI3_X105Y183_OLOGIC_X1Y184_TQ = 1'b1;
  assign RIOI3_X105Y183_OLOGIC_X1Y183_OQ = CLBLM_L_X12Y114_SLICE_X16Y114_DO5;
  assign RIOI3_X105Y183_OLOGIC_X1Y183_TQ = 1'b1;
  assign RIOI3_X105Y185_OLOGIC_X1Y186_OQ = CLBLM_L_X12Y111_SLICE_X16Y111_AQ;
  assign RIOI3_X105Y185_OLOGIC_X1Y186_TQ = 1'b1;
  assign RIOI3_X105Y185_OLOGIC_X1Y185_OQ = CLBLM_L_X8Y110_SLICE_X10Y110_CO5;
  assign RIOI3_X105Y185_OLOGIC_X1Y185_TQ = 1'b1;
  assign RIOI3_X105Y189_OLOGIC_X1Y190_OQ = CLBLM_R_X13Y113_SLICE_X19Y113_AQ;
  assign RIOI3_X105Y189_OLOGIC_X1Y190_TQ = 1'b1;
  assign RIOI3_X105Y189_OLOGIC_X1Y189_OQ = CLBLM_L_X10Y112_SLICE_X13Y112_AQ;
  assign RIOI3_X105Y189_OLOGIC_X1Y189_TQ = 1'b1;
  assign RIOI3_X105Y191_OLOGIC_X1Y192_OQ = CLBLM_R_X13Y109_SLICE_X19Y109_AQ;
  assign RIOI3_X105Y191_OLOGIC_X1Y192_TQ = 1'b1;
  assign RIOI3_X105Y191_OLOGIC_X1Y191_OQ = CLBLM_R_X11Y115_SLICE_X14Y115_AQ;
  assign RIOI3_X105Y191_OLOGIC_X1Y191_TQ = 1'b1;
  assign RIOI3_X105Y195_OLOGIC_X1Y196_OQ = CLBLM_L_X12Y117_SLICE_X16Y117_AQ;
  assign RIOI3_X105Y195_OLOGIC_X1Y196_TQ = 1'b1;
  assign RIOI3_X105Y195_OLOGIC_X1Y195_OQ = CLBLM_L_X12Y110_SLICE_X16Y110_AQ;
  assign RIOI3_X105Y195_OLOGIC_X1Y195_TQ = 1'b1;
  assign RIOI3_X105Y197_OLOGIC_X1Y198_OQ = CLBLL_L_X26Y136_SLICE_X38Y136_AO5;
  assign RIOI3_X105Y197_OLOGIC_X1Y198_TQ = 1'b1;
  assign RIOI3_X105Y197_OLOGIC_X1Y197_OQ = CLBLL_L_X26Y136_SLICE_X38Y136_AO5;
  assign RIOI3_X105Y197_OLOGIC_X1Y197_TQ = 1'b1;
  assign RIOI3_SING_X105Y100_ILOGIC_X1Y100_O = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign RIOI3_SING_X105Y149_ILOGIC_X1Y149_O = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign RIOI3_SING_X105Y150_OLOGIC_X1Y150_OQ = LIOB33_X0Y75_IOB_X0Y75_I;
  assign RIOI3_SING_X105Y150_OLOGIC_X1Y150_TQ = 1'b1;
  assign RIOI3_SING_X105Y199_OLOGIC_X1Y199_OQ = CLBLM_R_X11Y119_SLICE_X14Y119_AQ;
  assign RIOI3_SING_X105Y199_OLOGIC_X1Y199_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_O = RIOB33_X105Y107_IOB_X1Y108_I;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_O = RIOB33_X105Y107_IOB_X1Y107_I;
  assign RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_O = RIOB33_X105Y119_IOB_X1Y119_I;
  assign RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y132_O = RIOB33_X105Y131_IOB_X1Y132_I;
  assign RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y131_O = RIOB33_X105Y131_IOB_X1Y131_I;
  assign RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y144_O = RIOB33_X105Y143_IOB_X1Y144_I;
  assign RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y143_O = RIOB33_X105Y143_IOB_X1Y143_I;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_OQ = CLBLM_R_X37Y117_SLICE_X56Y117_AO6;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_OQ = RIOB33_X105Y125_IOB_X1Y126_I;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_OQ = CLBLM_R_X103Y170_SLICE_X163Y170_AO6;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_OQ = CLBLM_R_X103Y169_SLICE_X163Y169_AO6;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_OQ = CLBLM_L_X12Y114_SLICE_X16Y114_DO6;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_OQ = CLBLM_R_X13Y110_SLICE_X18Y110_DO5;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_OQ = CLBLM_R_X11Y119_SLICE_X14Y119_AQ;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_OQ = CLBLM_L_X12Y118_SLICE_X16Y118_AQ;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y114_O = RIOB33_X105Y113_IOB_X1Y114_I;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_O = RIOB33_X105Y113_IOB_X1Y113_I;
  assign RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y138_O = RIOB33_X105Y137_IOB_X1Y138_I;
  assign RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y137_O = RIOB33_X105Y137_IOB_X1Y137_I;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_OQ = CLBLM_L_X8Y110_SLICE_X10Y110_CO5;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_OQ = CLBLM_L_X8Y110_SLICE_X10Y110_CO6;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_OQ = CLBLM_L_X12Y117_SLICE_X17Y117_AQ;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_OQ = CLBLM_R_X11Y115_SLICE_X14Y115_BQ;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_TQ = 1'b1;
  assign CLBLM_R_X37Y117_SLICE_X56Y117_C1 = 1'b1;
  assign CLBLM_R_X37Y117_SLICE_X56Y117_C2 = 1'b1;
  assign CLBLM_R_X37Y117_SLICE_X56Y117_C3 = 1'b1;
  assign CLBLM_R_X37Y117_SLICE_X56Y117_C4 = 1'b1;
  assign CLBLM_R_X37Y117_SLICE_X56Y117_C5 = 1'b1;
  assign CLBLM_R_X37Y117_SLICE_X56Y117_C6 = 1'b1;
  assign LIOI3_SING_X0Y199_OLOGIC_X0Y199_T1 = 1'b1;
  assign LIOB33_X0Y79_IOB_X0Y80_O = CLBLL_L_X2Y106_SLICE_X0Y106_AO6;
  assign LIOB33_X0Y147_IOB_X0Y147_O = LIOB33_X0Y71_IOB_X0Y71_I;
  assign LIOB33_X0Y147_IOB_X0Y148_O = LIOB33_X0Y61_IOB_X0Y61_I;
  assign CLBLM_R_X37Y117_SLICE_X56Y117_D1 = 1'b1;
  assign CLBLM_R_X37Y117_SLICE_X56Y117_D2 = 1'b1;
  assign CLBLM_R_X37Y117_SLICE_X56Y117_D3 = 1'b1;
  assign CLBLM_R_X37Y117_SLICE_X56Y117_D4 = 1'b1;
  assign CLBLM_R_X37Y117_SLICE_X56Y117_D5 = 1'b1;
  assign CLBLM_R_X37Y117_SLICE_X56Y117_D6 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_B1 = CLBLL_L_X4Y112_SLICE_X4Y112_CO5;
  assign CLBLM_R_X13Y107_SLICE_X19Y107_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_B2 = CLBLM_R_X7Y109_SLICE_X9Y109_BQ;
  assign CLBLM_R_X13Y107_SLICE_X19Y107_A2 = CLBLM_L_X12Y107_SLICE_X17Y107_CO5;
  assign CLBLM_R_X13Y107_SLICE_X19Y107_A3 = CLBLM_R_X13Y107_SLICE_X19Y107_AQ;
  assign CLBLM_R_X13Y107_SLICE_X19Y107_A4 = CLBLM_R_X13Y106_SLICE_X18Y106_AO6;
  assign CLBLM_R_X13Y107_SLICE_X19Y107_A5 = CLBLM_R_X7Y108_SLICE_X8Y108_BQ;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y107_SLICE_X19Y107_A6 = CLBLM_L_X12Y108_SLICE_X17Y108_CO5;
  assign CLBLM_R_X13Y107_SLICE_X19Y107_B1 = CLBLM_L_X10Y115_SLICE_X12Y115_CQ;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_B4 = CLBLM_L_X10Y108_SLICE_X12Y108_CQ;
  assign CLBLM_R_X13Y107_SLICE_X19Y107_B2 = 1'b1;
  assign CLBLM_R_X13Y107_SLICE_X19Y107_B3 = 1'b1;
  assign CLBLM_R_X13Y107_SLICE_X19Y107_B4 = CLBLM_L_X12Y108_SLICE_X17Y108_CO5;
  assign CLBLM_R_X13Y107_SLICE_X19Y107_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_B5 = CLBLM_L_X12Y108_SLICE_X16Y108_AQ;
  assign CLBLM_R_X13Y107_SLICE_X19Y107_B6 = CLBLM_R_X13Y107_SLICE_X19Y107_CO6;
  assign CLBLM_R_X13Y107_SLICE_X19Y107_C1 = CLBLM_R_X13Y107_SLICE_X19Y107_BQ;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_B6 = 1'b1;
  assign CLBLM_R_X13Y107_SLICE_X19Y107_C2 = CLBLM_L_X12Y105_SLICE_X17Y105_CO6;
  assign CLBLM_R_X13Y107_SLICE_X19Y107_C3 = CLBLM_L_X12Y108_SLICE_X16Y108_CQ;
  assign CLBLM_R_X13Y107_SLICE_X19Y107_C4 = CLBLM_L_X12Y105_SLICE_X17Y105_AO5;
  assign CLBLM_R_X13Y107_SLICE_X19Y107_C5 = CLBLM_R_X13Y107_SLICE_X19Y107_DO6;
  assign CLBLM_R_X13Y107_SLICE_X19Y107_C6 = CLBLM_L_X12Y107_SLICE_X17Y107_CO5;
  assign CLBLM_R_X13Y107_SLICE_X19Y107_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y155_OLOGIC_X0Y156_D1 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X13Y107_SLICE_X19Y107_D1 = CLBLM_L_X12Y107_SLICE_X17Y107_BQ;
  assign CLBLM_R_X13Y107_SLICE_X19Y107_D2 = CLBLM_L_X12Y107_SLICE_X16Y107_BQ;
  assign CLBLM_R_X13Y107_SLICE_X19Y107_D3 = CLBLM_R_X13Y109_SLICE_X19Y109_BQ;
  assign CLBLM_R_X13Y107_SLICE_X19Y107_D4 = CLBLM_R_X13Y113_SLICE_X18Y113_BQ;
  assign CLBLM_R_X13Y107_SLICE_X19Y107_D5 = CLBLM_R_X13Y108_SLICE_X19Y108_BQ;
  assign CLBLM_R_X13Y107_SLICE_X19Y107_D6 = CLBLM_L_X12Y108_SLICE_X16Y108_BQ;
  assign LIOI3_X0Y155_OLOGIC_X0Y156_T1 = 1'b1;
  assign CLBLM_R_X13Y107_SLICE_X18Y107_A1 = CLBLM_R_X13Y112_SLICE_X18Y112_CQ;
  assign CLBLM_R_X13Y107_SLICE_X18Y107_A2 = CLBLM_L_X12Y108_SLICE_X17Y108_CO5;
  assign CLBLM_R_X13Y107_SLICE_X18Y107_A3 = CLBLM_R_X13Y107_SLICE_X18Y107_AQ;
  assign CLBLM_R_X13Y107_SLICE_X18Y107_A4 = CLBLM_L_X12Y106_SLICE_X17Y106_BO6;
  assign CLBLM_R_X13Y107_SLICE_X18Y107_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y107_SLICE_X18Y107_A6 = CLBLM_L_X12Y107_SLICE_X17Y107_CO5;
  assign LIOI3_X0Y155_OLOGIC_X0Y155_D1 = LIOB33_X0Y69_IOB_X0Y70_I;
  assign CLBLM_R_X13Y107_SLICE_X18Y107_B1 = CLBLM_L_X12Y107_SLICE_X16Y107_AQ;
  assign CLBLM_R_X13Y107_SLICE_X18Y107_B2 = CLBLM_R_X13Y106_SLICE_X18Y106_CO6;
  assign CLBLM_R_X13Y107_SLICE_X18Y107_B3 = CLBLM_R_X13Y107_SLICE_X18Y107_AQ;
  assign CLBLM_R_X13Y107_SLICE_X18Y107_B4 = CLBLM_R_X13Y107_SLICE_X19Y107_BQ;
  assign CLBLM_R_X13Y107_SLICE_X18Y107_B5 = CLBLM_R_X13Y107_SLICE_X19Y107_AQ;
  assign CLBLM_R_X13Y107_SLICE_X18Y107_B6 = CLBLM_R_X13Y108_SLICE_X18Y108_AQ;
  assign LIOI3_X0Y155_OLOGIC_X0Y155_T1 = 1'b1;
  assign CLBLM_R_X13Y107_SLICE_X18Y107_C1 = CLBLM_R_X13Y107_SLICE_X19Y107_AQ;
  assign CLBLM_R_X13Y107_SLICE_X18Y107_C2 = CLBLM_R_X13Y107_SLICE_X19Y107_BQ;
  assign CLBLM_R_X13Y107_SLICE_X18Y107_C3 = CLBLM_R_X13Y107_SLICE_X18Y107_AQ;
  assign CLBLM_R_X13Y107_SLICE_X18Y107_C4 = CLBLM_R_X13Y108_SLICE_X18Y108_AQ;
  assign CLBLM_R_X13Y107_SLICE_X18Y107_C5 = CLBLM_L_X12Y107_SLICE_X16Y107_AQ;
  assign CLBLM_R_X13Y107_SLICE_X18Y107_C6 = CLBLM_R_X13Y106_SLICE_X18Y106_BO6;
  assign CLBLM_R_X13Y107_SLICE_X18Y107_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y107_SLICE_X18Y107_D1 = CLBLM_R_X13Y107_SLICE_X19Y107_AQ;
  assign CLBLM_R_X13Y107_SLICE_X18Y107_D2 = CLBLM_R_X13Y107_SLICE_X18Y107_AQ;
  assign CLBLM_R_X13Y107_SLICE_X18Y107_D3 = CLBLM_L_X12Y107_SLICE_X16Y107_AQ;
  assign CLBLM_R_X13Y107_SLICE_X18Y107_D4 = 1'b1;
  assign CLBLM_R_X13Y107_SLICE_X18Y107_D5 = CLBLM_R_X13Y107_SLICE_X19Y107_BQ;
  assign CLBLM_R_X13Y107_SLICE_X18Y107_D6 = CLBLM_R_X13Y106_SLICE_X18Y106_BO6;
  assign RIOB33_SING_X105Y150_IOB_X1Y150_O = LIOB33_X0Y75_IOB_X0Y75_I;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_D1 = CLBLM_L_X12Y114_SLICE_X16Y114_DO6;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_D1 = CLBLM_R_X13Y110_SLICE_X18Y110_DO5;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_T1 = 1'b1;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_A1 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_A2 = CLBLM_R_X5Y115_SLICE_X7Y115_CO6;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_A3 = CLBLM_L_X12Y114_SLICE_X17Y114_AQ;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_A5 = 1'b1;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_A6 = CLBLM_L_X12Y111_SLICE_X16Y111_BQ;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_B1 = CLBLM_R_X11Y115_SLICE_X15Y115_AQ;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_B2 = CLBLM_L_X12Y114_SLICE_X17Y114_BQ;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_B3 = CLBLM_L_X12Y114_SLICE_X17Y114_AQ;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_B5 = 1'b1;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_B6 = CLBLM_R_X5Y115_SLICE_X7Y115_CO6;
  assign RIOB33_X105Y157_IOB_X1Y158_O = CLBLM_R_X37Y117_SLICE_X56Y117_AO6;
  assign RIOB33_X105Y157_IOB_X1Y157_O = RIOB33_X105Y125_IOB_X1Y126_I;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_A1 = 1'b1;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_A2 = 1'b1;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_A3 = 1'b1;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_A4 = 1'b1;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_A5 = 1'b1;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_A6 = 1'b1;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_C1 = CLBLM_L_X12Y112_SLICE_X16Y112_DQ;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_C2 = CLBLM_L_X12Y114_SLICE_X17Y114_AQ;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_C3 = 1'b1;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_B1 = 1'b1;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_B2 = 1'b1;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_B3 = 1'b1;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_B4 = 1'b1;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_B5 = 1'b1;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_B6 = 1'b1;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_D2 = 1'b1;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_D3 = 1'b1;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_D4 = 1'b1;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_C1 = 1'b1;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_C2 = 1'b1;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_C3 = 1'b1;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_C4 = 1'b1;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_C5 = 1'b1;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_C6 = 1'b1;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_D5 = 1'b1;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_D6 = 1'b1;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_A1 = 1'b1;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_A3 = CLBLM_R_X11Y111_SLICE_X15Y111_CQ;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_A4 = CLBLM_L_X12Y114_SLICE_X16Y114_AQ;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_A5 = CLBLM_R_X7Y115_SLICE_X9Y115_DO6;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_A6 = CLBLM_L_X8Y114_SLICE_X10Y114_BQ;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_D1 = 1'b1;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_D2 = 1'b1;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_D3 = 1'b1;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_D4 = 1'b1;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_D5 = 1'b1;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_D6 = 1'b1;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_B1 = CLBLM_R_X11Y115_SLICE_X15Y115_CQ;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_B6 = CLBLM_R_X11Y114_SLICE_X14Y114_DQ;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_B2 = CLBLM_L_X12Y114_SLICE_X16Y114_BQ;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_B3 = CLBLM_R_X5Y115_SLICE_X7Y115_CO6;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_B5 = 1'b1;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_A2 = CLBLM_L_X10Y106_SLICE_X13Y106_BQ;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_A3 = CLBLM_L_X10Y104_SLICE_X12Y104_AQ;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_A4 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_A5 = 1'b1;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_A6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_C1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_C2 = CLBLM_L_X12Y114_SLICE_X16Y114_CQ;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_C3 = CLBLM_L_X12Y117_SLICE_X17Y117_BQ;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_B1 = CLBLM_L_X10Y105_SLICE_X13Y105_CO6;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_B2 = CLBLM_L_X8Y104_SLICE_X11Y104_BO6;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_B3 = CLBLM_L_X10Y105_SLICE_X12Y105_DO6;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_B4 = CLBLM_L_X12Y110_SLICE_X16Y110_DO5;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_B5 = CLBLM_R_X3Y108_SLICE_X3Y108_CO6;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_B6 = CLBLM_L_X10Y106_SLICE_X12Y106_BO6;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_D1 = CLBLM_L_X10Y113_SLICE_X13Y113_CQ;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_C1 = CLBLM_R_X3Y108_SLICE_X3Y108_CO6;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_C2 = 1'b1;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_C3 = CLBLM_L_X10Y105_SLICE_X12Y105_DO6;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_C4 = CLBLM_L_X12Y110_SLICE_X16Y110_DO5;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_C5 = CLBLM_L_X10Y105_SLICE_X13Y105_CO6;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_C6 = CLBLM_L_X8Y104_SLICE_X11Y104_BO6;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_D2 = CLBLM_L_X12Y114_SLICE_X16Y114_CQ;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_D3 = CLBLM_L_X10Y110_SLICE_X13Y110_DQ;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_D4 = CLBLM_L_X8Y115_SLICE_X11Y115_AQ;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_D6 = 1'b1;
  assign RIOI3_X105Y139_ILOGIC_X1Y140_D = RIOB33_X105Y139_IOB_X1Y140_I;
  assign RIOI3_X105Y139_ILOGIC_X1Y139_D = RIOB33_X105Y139_IOB_X1Y139_I;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_D1 = 1'b1;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_D2 = 1'b1;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_D3 = 1'b1;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_D4 = 1'b1;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_D5 = 1'b1;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_D6 = 1'b1;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_A2 = CLBLM_L_X12Y108_SLICE_X17Y108_CO5;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_A3 = CLBLM_R_X13Y108_SLICE_X18Y108_CO6;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_A4 = CLBLM_L_X12Y107_SLICE_X17Y107_CO5;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_A5 = CLBLM_L_X12Y107_SLICE_X17Y107_BQ;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_A6 = 1'b1;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_B2 = CLBLM_L_X12Y108_SLICE_X17Y108_CO5;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_B3 = 1'b1;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_B4 = 1'b1;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_B5 = CLBLM_L_X10Y114_SLICE_X12Y114_CQ;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_B6 = CLBLM_R_X13Y108_SLICE_X19Y108_CO6;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_C1 = CLBLM_L_X12Y105_SLICE_X17Y105_AO5;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_C2 = CLBLM_L_X12Y108_SLICE_X16Y108_DQ;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_C3 = CLBLM_R_X13Y108_SLICE_X19Y108_BQ;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_C4 = CLBLM_L_X12Y105_SLICE_X17Y105_CO6;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_C5 = 1'b1;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_C6 = CLBLM_L_X12Y107_SLICE_X17Y107_CO5;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_D1 = 1'b1;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_D2 = 1'b1;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_D3 = 1'b1;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_D4 = 1'b1;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_D5 = 1'b1;
  assign CLBLM_R_X13Y108_SLICE_X19Y108_D6 = 1'b1;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_A2 = CLBLM_R_X13Y108_SLICE_X18Y108_DO6;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_A3 = CLBLM_L_X12Y109_SLICE_X17Y109_DQ;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_A4 = CLBLM_L_X12Y107_SLICE_X17Y107_CO5;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_A5 = 1'b1;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_A6 = CLBLM_L_X12Y108_SLICE_X17Y108_CO5;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_B1 = CLBLM_R_X13Y107_SLICE_X18Y107_CO6;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_B2 = CLBLM_L_X12Y105_SLICE_X17Y105_AO5;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_B3 = 1'b1;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_B4 = CLBLM_R_X13Y107_SLICE_X18Y107_BO6;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_B5 = CLBLM_R_X13Y108_SLICE_X19Y108_AQ;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_B6 = 1'b1;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_C1 = CLBLM_L_X12Y105_SLICE_X17Y105_AO5;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_C2 = CLBLM_R_X13Y108_SLICE_X19Y108_AQ;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_C3 = CLBLM_R_X11Y108_SLICE_X14Y108_AQ;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_C4 = CLBLM_R_X13Y107_SLICE_X18Y107_BO6;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_C5 = CLBLM_R_X13Y107_SLICE_X18Y107_CO6;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_C6 = CLBLM_L_X12Y105_SLICE_X17Y105_CO6;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_D1 = CLBLM_L_X12Y105_SLICE_X17Y105_AO5;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_D2 = CLBLM_R_X13Y106_SLICE_X18Y106_DO6;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_D3 = CLBLM_R_X13Y107_SLICE_X18Y107_DO6;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_D4 = CLBLM_L_X12Y105_SLICE_X17Y105_CO6;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_D5 = CLBLM_L_X12Y108_SLICE_X17Y108_AQ;
  assign CLBLM_R_X13Y108_SLICE_X18Y108_D6 = CLBLM_R_X13Y108_SLICE_X18Y108_AQ;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_A1 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_A2 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_A3 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_A4 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_A5 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_A6 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_B1 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_B2 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_B3 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_B4 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_B5 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_B6 = 1'b1;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_A1 = CLBLM_R_X7Y106_SLICE_X9Y106_DO6;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_A2 = CLBLM_R_X11Y105_SLICE_X14Y105_CQ;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_A3 = CLBLM_L_X10Y106_SLICE_X12Y106_AQ;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_A4 = CLBLM_R_X11Y105_SLICE_X14Y105_C5Q;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_A5 = CLBLM_L_X10Y105_SLICE_X12Y105_AQ;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_A6 = CLBLM_R_X5Y115_SLICE_X7Y115_CO6;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_C1 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_C2 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_C3 = 1'b1;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_B1 = CLBLM_R_X7Y106_SLICE_X9Y106_DO6;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_B2 = CLBLM_R_X11Y105_SLICE_X14Y105_CQ;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_B3 = CLBLM_L_X10Y106_SLICE_X12Y106_AQ;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_B4 = CLBLM_R_X11Y105_SLICE_X14Y105_C5Q;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_B5 = CLBLM_L_X10Y105_SLICE_X12Y105_AQ;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_B6 = CLBLM_R_X5Y115_SLICE_X7Y115_CO6;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_D1 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_D2 = 1'b1;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_C1 = CLBLM_R_X11Y105_SLICE_X14Y105_BQ;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_C2 = CLBLM_L_X10Y111_SLICE_X13Y111_BQ;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_C3 = CLBLM_L_X10Y106_SLICE_X12Y106_DO6;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_C4 = 1'b1;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_C5 = CLBLM_L_X10Y105_SLICE_X13Y105_DO6;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_C6 = CLBLM_L_X8Y105_SLICE_X10Y105_DO6;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_D3 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_D4 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_A1 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_A2 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_A3 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_A4 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_A5 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_A6 = 1'b1;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_D1 = CLBLM_L_X10Y107_SLICE_X12Y107_AQ;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_D2 = CLBLM_R_X11Y105_SLICE_X14Y105_AQ;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_D3 = 1'b1;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_D4 = CLBLM_L_X8Y105_SLICE_X11Y105_BQ;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_D5 = 1'b1;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_D6 = CLBLM_L_X10Y105_SLICE_X12Y105_BQ;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_AX = CLBLM_R_X11Y115_SLICE_X14Y115_BO6;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_B1 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_B2 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_B3 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_B4 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_B6 = 1'b1;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_A1 = CLBLM_R_X7Y106_SLICE_X9Y106_DO6;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_A2 = CLBLM_R_X5Y115_SLICE_X7Y115_CO6;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_A3 = CLBLM_L_X10Y105_SLICE_X12Y105_AQ;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_A5 = CLBLM_L_X10Y105_SLICE_X12Y105_CO5;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_C4 = 1'b1;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_A6 = CLBLM_L_X8Y107_SLICE_X10Y107_CQ;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_C1 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_C2 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_C3 = 1'b1;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_B1 = CLBLM_L_X10Y106_SLICE_X12Y106_BO6;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_B2 = CLBLM_L_X10Y105_SLICE_X12Y105_BQ;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_B3 = CLBLM_L_X8Y105_SLICE_X10Y105_AQ;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_C5 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_C6 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_D1 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_D2 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_D3 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_D4 = 1'b1;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_C2 = CLBLM_L_X10Y105_SLICE_X12Y105_AQ;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_C3 = CLBLM_R_X11Y105_SLICE_X14Y105_CQ;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_C4 = CLBLM_R_X5Y115_SLICE_X7Y115_CO6;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_D5 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_D6 = 1'b1;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_C1 = CLBLM_L_X10Y106_SLICE_X12Y106_AQ;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_C5 = CLBLM_R_X11Y105_SLICE_X14Y105_C5Q;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_C6 = 1'b1;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_D1 = CLBLM_L_X8Y106_SLICE_X11Y106_BQ;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_D2 = CLBLM_L_X10Y108_SLICE_X12Y108_BQ;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_D3 = CLBLM_L_X8Y107_SLICE_X10Y107_BQ;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_D4 = CLBLM_L_X8Y106_SLICE_X11Y106_DO6;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_D5 = CLBLM_R_X11Y106_SLICE_X14Y106_AQ;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_D6 = 1'b1;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_A1 = CLBLM_L_X8Y119_SLICE_X10Y119_AQ;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_A2 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_A3 = CLBLM_R_X13Y109_SLICE_X19Y109_AQ;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_A5 = 1'b1;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_A6 = CLBLM_R_X13Y112_SLICE_X18Y112_A5Q;
  assign RIOI3_X105Y195_OLOGIC_X1Y196_D1 = CLBLM_L_X12Y117_SLICE_X16Y117_AQ;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_B1 = CLBLM_R_X13Y109_SLICE_X18Y109_CO6;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_B2 = CLBLM_R_X13Y110_SLICE_X19Y110_AQ;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_B3 = CLBLM_L_X12Y105_SLICE_X16Y105_BO6;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_B5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_B6 = CLBLM_R_X13Y109_SLICE_X19Y109_BQ;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_C1 = 1'b1;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_C2 = 1'b1;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_C3 = 1'b1;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_C4 = 1'b1;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_C5 = 1'b1;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_C6 = 1'b1;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_D1 = 1'b1;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_D2 = 1'b1;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_D3 = 1'b1;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_D4 = 1'b1;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_D5 = 1'b1;
  assign CLBLM_R_X13Y109_SLICE_X19Y109_D6 = 1'b1;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_A1 = CLBLM_R_X13Y109_SLICE_X18Y109_DO6;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_A2 = 1'b1;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_A3 = CLBLM_L_X12Y105_SLICE_X16Y105_BO6;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_A4 = CLBLM_R_X7Y116_SLICE_X9Y116_BO6;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_A5 = CLBLM_R_X13Y108_SLICE_X19Y108_AQ;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_B1 = CLBLM_L_X12Y105_SLICE_X16Y105_AQ;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_B2 = CLBLM_R_X13Y113_SLICE_X18Y113_BQ;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_B3 = CLBLM_R_X11Y105_SLICE_X14Y105_DQ;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_B4 = CLBLM_R_X13Y109_SLICE_X19Y109_BQ;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_B5 = CLBLM_L_X12Y107_SLICE_X17Y107_BQ;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_B6 = 1'b1;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_C1 = CLBLM_L_X12Y107_SLICE_X17Y107_DO5;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_C2 = CLBLM_R_X13Y109_SLICE_X19Y109_BQ;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_C3 = CLBLM_R_X13Y113_SLICE_X18Y113_BQ;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_C4 = CLBLM_L_X12Y107_SLICE_X17Y107_AQ;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_C5 = CLBLM_L_X12Y107_SLICE_X17Y107_BQ;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_C6 = CLBLM_R_X13Y108_SLICE_X18Y108_BO6;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_D1 = CLBLM_L_X12Y108_SLICE_X17Y108_DO6;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_D2 = CLBLM_R_X13Y109_SLICE_X18Y109_AQ;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_D3 = CLBLM_R_X11Y110_SLICE_X15Y110_A5Q;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_D4 = CLBLM_L_X12Y107_SLICE_X17Y107_AQ;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_D5 = CLBLM_R_X13Y109_SLICE_X18Y109_BO5;
  assign CLBLM_R_X13Y109_SLICE_X18Y109_D6 = CLBLM_R_X13Y109_SLICE_X18Y109_BO6;
  assign LIOI3_X0Y159_OLOGIC_X0Y160_D1 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign LIOI3_X0Y159_OLOGIC_X0Y160_T1 = 1'b1;
  assign LIOI3_X0Y159_OLOGIC_X0Y159_D1 = RIOB33_X105Y117_IOB_X1Y117_I;
  assign LIOI3_X0Y159_OLOGIC_X0Y159_T1 = 1'b1;
  assign LIOB33_X0Y155_IOB_X0Y156_O = RIOB33_X105Y105_IOB_X1Y106_I;
  assign LIOB33_X0Y155_IOB_X0Y155_O = LIOB33_X0Y69_IOB_X0Y70_I;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_A1 = CLBLM_R_X11Y106_SLICE_X14Y106_CQ;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_A2 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_A3 = CLBLM_L_X10Y106_SLICE_X13Y106_AQ;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_A5 = CLBLM_L_X10Y107_SLICE_X13Y107_AQ;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_A6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign LIOB33_X0Y153_IOB_X0Y153_O = LIOB33_X0Y67_IOB_X0Y67_I;
  assign LIOB33_X0Y153_IOB_X0Y154_O = LIOB33_X0Y67_IOB_X0Y68_I;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_B1 = CLBLM_R_X7Y107_SLICE_X9Y107_C5Q;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_B2 = CLBLM_L_X10Y106_SLICE_X13Y106_BQ;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_B3 = 1'b1;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_B4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_B5 = 1'b1;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_C1 = CLBLM_L_X10Y106_SLICE_X12Y106_BO6;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_C2 = CLBLM_L_X10Y106_SLICE_X12Y106_CO6;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_C3 = CLBLM_R_X13Y109_SLICE_X19Y109_AQ;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_C5 = CLBLM_L_X10Y106_SLICE_X13Y106_CQ;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_C6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_D1 = CLBLM_L_X12Y105_SLICE_X17Y105_AO6;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_D2 = CLBLL_L_X4Y107_SLICE_X4Y107_BO5;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_D3 = CLBLM_R_X11Y105_SLICE_X15Y105_BQ;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_D4 = CLBLM_L_X12Y107_SLICE_X17Y107_BQ;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_D5 = CLBLM_L_X8Y106_SLICE_X10Y106_BQ;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_D6 = CLBLM_R_X5Y107_SLICE_X6Y107_BQ;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_D1 = CLBLM_R_X11Y119_SLICE_X14Y119_AQ;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_T1 = 1'b1;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_A2 = CLBLM_L_X10Y105_SLICE_X12Y105_CO6;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_A3 = CLBLM_L_X10Y106_SLICE_X12Y106_AQ;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_A5 = CLBLM_L_X8Y115_SLICE_X10Y115_AQ;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_A6 = CLBLM_L_X10Y111_SLICE_X12Y111_CQ;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_A6 = 1'b1;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_B1 = CLBLM_L_X10Y107_SLICE_X12Y107_BQ;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_B2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_B3 = CLBLM_L_X10Y113_SLICE_X13Y113_AQ;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_B4 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_B5 = CLBLM_R_X7Y105_SLICE_X8Y105_AQ;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_B6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_D1 = CLBLM_L_X12Y118_SLICE_X16Y118_AQ;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_C1 = CLBLM_R_X11Y110_SLICE_X14Y110_AQ;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_C2 = CLBLM_R_X3Y108_SLICE_X2Y108_DO6;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_C3 = CLBLM_R_X5Y107_SLICE_X7Y107_AQ;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_C4 = CLBLM_L_X10Y105_SLICE_X13Y105_CO6;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_C5 = CLBLM_L_X10Y112_SLICE_X12Y112_DO6;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_C6 = CLBLM_L_X12Y110_SLICE_X16Y110_DO5;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_T1 = 1'b1;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_D1 = CLBLM_L_X10Y110_SLICE_X13Y110_AQ;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_D2 = CLBLM_L_X10Y110_SLICE_X13Y110_BQ;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_D3 = CLBLM_L_X8Y106_SLICE_X11Y106_BQ;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_D4 = CLBLM_L_X10Y106_SLICE_X13Y106_CQ;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_D5 = CLBLM_L_X10Y107_SLICE_X12Y107_BQ;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_D6 = CLBLM_L_X8Y107_SLICE_X10Y107_BQ;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_C1 = 1'b1;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_C2 = 1'b1;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_C3 = 1'b1;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_C4 = 1'b1;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_C5 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_A1 = CLBLM_R_X7Y115_SLICE_X8Y115_DQ;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_C6 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_A3 = CLBLM_R_X13Y110_SLICE_X19Y110_AQ;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_A5 = CLBLM_R_X13Y109_SLICE_X18Y109_AQ;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_A6 = CLBLM_L_X12Y110_SLICE_X16Y110_DO6;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_B1 = CLBLM_L_X12Y110_SLICE_X16Y110_AQ;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_B2 = CLBLM_R_X13Y110_SLICE_X19Y110_BQ;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_B3 = CLBLM_L_X10Y109_SLICE_X12Y109_DO6;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_B4 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_B6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_C2 = CLBLM_R_X13Y110_SLICE_X19Y110_CQ;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_C3 = CLBLM_R_X11Y112_SLICE_X14Y112_C5Q;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_C4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_C5 = CLBLM_L_X10Y109_SLICE_X12Y109_DO6;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_C6 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_D1 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_D2 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_D3 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_D4 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_D5 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X19Y110_D6 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_A1 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_A2 = CLBLM_L_X12Y109_SLICE_X16Y109_BQ;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_A3 = CLBLM_R_X13Y110_SLICE_X18Y110_AQ;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_D1 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_A5 = CLBLM_R_X13Y110_SLICE_X18Y110_CQ;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_A6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_D2 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_B1 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_B2 = CLBLM_R_X13Y108_SLICE_X19Y108_BQ;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_D3 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_B4 = CLBLM_R_X11Y111_SLICE_X15Y111_BQ;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_B5 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign RIOI3_X105Y141_ILOGIC_X1Y142_D = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_D4 = 1'b1;
  assign RIOI3_X105Y141_ILOGIC_X1Y141_D = RIOB33_X105Y141_IOB_X1Y141_I;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_C1 = CLBLL_L_X4Y110_SLICE_X4Y110_B5Q;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_C2 = CLBLM_R_X13Y110_SLICE_X18Y110_CQ;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_D5 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_C3 = CLBLM_L_X10Y109_SLICE_X13Y109_CO6;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_C4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_C5 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_D6 = 1'b1;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_D1 = CLBLM_R_X13Y110_SLICE_X18Y110_CQ;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_D2 = CLBLM_R_X11Y107_SLICE_X15Y107_CQ;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_D3 = CLBLM_L_X12Y109_SLICE_X17Y109_DQ;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_D4 = CLBLM_R_X13Y110_SLICE_X19Y110_CQ;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_D5 = CLBLM_L_X10Y113_SLICE_X13Y113_CQ;
  assign CLBLM_R_X13Y110_SLICE_X18Y110_D6 = 1'b1;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_A1 = 1'b1;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_A2 = 1'b1;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_C4 = CLBLM_R_X7Y117_SLICE_X9Y117_A5Q;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_A3 = 1'b1;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_A4 = 1'b1;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_A5 = 1'b1;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_A6 = 1'b1;
  assign LIOB33_X0Y157_IOB_X0Y158_O = RIOB33_X105Y115_IOB_X1Y116_I;
  assign LIOB33_X0Y157_IOB_X0Y157_O = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_A1 = 1'b1;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_A2 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_A3 = CLBLM_L_X12Y117_SLICE_X17Y117_AQ;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_A4 = CLBLM_R_X11Y117_SLICE_X15Y117_CQ;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_A5 = CLBLM_L_X8Y119_SLICE_X10Y119_AQ;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_B1 = 1'b1;
  assign RIOI3_X105Y159_OLOGIC_X1Y160_D1 = CLBLM_R_X13Y110_SLICE_X18Y110_DO5;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_B2 = 1'b1;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_B1 = CLBLM_L_X12Y107_SLICE_X17Y107_AQ;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_B2 = CLBLM_L_X12Y117_SLICE_X17Y117_BQ;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_B3 = CLBLM_L_X10Y116_SLICE_X12Y116_DO5;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_B4 = CLBLM_L_X10Y118_SLICE_X13Y118_BO6;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_B5 = CLBLM_L_X10Y118_SLICE_X13Y118_CO6;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_B3 = 1'b1;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_B4 = 1'b1;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_A1 = 1'b1;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_A2 = CLBLM_L_X8Y119_SLICE_X10Y119_AQ;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_A3 = CLBLM_R_X7Y106_SLICE_X8Y106_AQ;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_A5 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_A6 = CLBLM_L_X10Y108_SLICE_X13Y108_BO6;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_C1 = 1'b1;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_C2 = 1'b1;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_B1 = CLBLM_L_X10Y106_SLICE_X12Y106_BO5;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_B2 = CLBLM_L_X8Y107_SLICE_X11Y107_BQ;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_B3 = CLBLM_R_X11Y105_SLICE_X15Y105_BQ;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_B4 = CLBLM_L_X12Y110_SLICE_X17Y110_BQ;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_B5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_B6 = CLBLM_R_X11Y107_SLICE_X14Y107_BO6;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_D3 = 1'b1;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_D4 = 1'b1;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_C1 = CLBLM_L_X10Y105_SLICE_X12Y105_CO5;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_C2 = CLBLM_L_X8Y115_SLICE_X11Y115_BQ;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_C3 = CLBLM_L_X10Y105_SLICE_X12Y105_AQ;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_C4 = CLBLM_R_X5Y115_SLICE_X7Y115_DO6;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_C5 = CLBLM_L_X10Y107_SLICE_X13Y107_DO6;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_C6 = CLBLM_R_X3Y107_SLICE_X3Y107_CO6;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_D5 = 1'b1;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_D6 = 1'b1;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_A1 = 1'b1;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_A2 = CLBLM_L_X8Y119_SLICE_X10Y119_AQ;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_A3 = 1'b1;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_A4 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_A5 = 1'b1;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_D1 = CLBLL_L_X2Y108_SLICE_X1Y108_AO6;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_D2 = CLBLM_R_X11Y106_SLICE_X14Y106_CQ;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_D3 = CLBLM_L_X12Y105_SLICE_X17Y105_CO6;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_D4 = CLBLM_R_X7Y114_SLICE_X9Y114_CO6;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_D5 = CLBLM_R_X11Y106_SLICE_X15Y106_CO5;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_D6 = CLBLM_L_X10Y107_SLICE_X13Y107_BO6;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_AX = CLBLM_R_X13Y109_SLICE_X19Y109_BQ;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_B1 = 1'b1;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_B2 = 1'b1;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_B3 = 1'b1;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_B4 = 1'b1;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_A1 = CLBLM_L_X8Y108_SLICE_X10Y108_CQ;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_A2 = CLBLM_L_X10Y107_SLICE_X12Y107_BQ;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_A3 = CLBLM_L_X10Y107_SLICE_X12Y107_AQ;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_A6 = CLBLM_L_X10Y106_SLICE_X12Y106_BO6;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_C1 = 1'b1;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_C2 = 1'b1;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_C3 = 1'b1;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_B2 = CLBLM_L_X8Y105_SLICE_X11Y105_BQ;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_B3 = CLBLM_L_X10Y107_SLICE_X12Y107_BQ;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_B4 = CLBLM_L_X10Y106_SLICE_X12Y106_BO6;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_B6 = CLBLM_R_X11Y116_SLICE_X14Y116_BQ;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_CE = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_D1 = 1'b1;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_C1 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_C2 = CLBLM_R_X5Y115_SLICE_X7Y115_CO6;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_C3 = CLBLM_L_X10Y112_SLICE_X12Y112_DO6;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_C4 = CLBLM_R_X3Y108_SLICE_X2Y108_DO6;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_C5 = CLBLM_R_X11Y108_SLICE_X15Y108_DO6;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_C6 = CLBLM_L_X8Y119_SLICE_X10Y119_AQ;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_D6 = 1'b1;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_SR = CLBLM_L_X12Y117_SLICE_X16Y117_AO6;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X37Y117_SLICE_X57Y117_B5 = 1'b1;
  assign CLBLM_R_X37Y117_SLICE_X57Y117_B6 = 1'b1;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_D1 = CLBLM_L_X10Y104_SLICE_X12Y104_AQ;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_D2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_D3 = CLBLM_L_X10Y110_SLICE_X12Y110_CO6;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_D4 = CLBLM_R_X3Y108_SLICE_X2Y108_DO6;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_D5 = 1'b1;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_D6 = CLBLM_R_X7Y116_SLICE_X8Y116_CQ;
  assign RIOI3_X105Y159_OLOGIC_X1Y159_D1 = CLBLM_R_X13Y110_SLICE_X18Y110_DO6;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_T1 = 1'b1;
  assign CLBLM_R_X37Y117_SLICE_X57Y117_C3 = 1'b1;
  assign CLBLM_R_X37Y117_SLICE_X57Y117_C5 = 1'b1;
  assign CLBLM_R_X37Y117_SLICE_X57Y117_C6 = 1'b1;
  assign RIOI3_X105Y159_OLOGIC_X1Y159_T1 = 1'b1;
  assign CLBLM_R_X37Y117_SLICE_X57Y117_D4 = 1'b1;
  assign CLBLM_R_X37Y117_SLICE_X57Y117_D5 = 1'b1;
  assign CLBLM_R_X37Y117_SLICE_X57Y117_D6 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_B6 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_D1 = CLBLM_R_X11Y115_SLICE_X14Y115_BQ;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_A4 = CLBLM_R_X11Y105_SLICE_X14Y105_CQ;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_A5 = CLBLM_L_X12Y110_SLICE_X17Y110_AQ;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_A6 = 1'b1;
  assign LIOB33_X0Y159_IOB_X0Y159_O = RIOB33_X105Y117_IOB_X1Y117_I;
  assign LIOB33_X0Y159_IOB_X0Y160_O = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_A2 = CLBLM_R_X7Y115_SLICE_X9Y115_BQ;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_A1 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_A2 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_A3 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_A4 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_A5 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_A6 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_B1 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_B2 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_B3 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_B4 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_B5 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_B6 = 1'b1;
  assign CLBLM_R_X37Y117_SLICE_X56Y117_B2 = 1'b1;
  assign CLBLM_R_X37Y117_SLICE_X56Y117_B3 = 1'b1;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_A1 = 1'b1;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_A2 = CLBLM_R_X13Y110_SLICE_X19Y110_CQ;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_A4 = CLBLM_L_X8Y119_SLICE_X10Y119_AQ;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_A5 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_A6 = CLBLM_L_X10Y108_SLICE_X13Y108_CO6;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_C1 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_C2 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_C3 = 1'b1;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_B1 = CLBLM_R_X5Y115_SLICE_X7Y115_CO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_B2 = CLBLM_R_X11Y108_SLICE_X15Y108_AQ;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_B3 = CLBLM_L_X10Y107_SLICE_X13Y107_AQ;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_B4 = CLBLM_L_X10Y109_SLICE_X13Y109_AO5;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_B5 = CLBLM_L_X12Y110_SLICE_X17Y110_AQ;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_B6 = CLBLM_R_X11Y105_SLICE_X14Y105_CQ;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_D1 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_D2 = 1'b1;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_C1 = CLBLM_R_X5Y115_SLICE_X7Y115_CO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_C2 = CLBLM_L_X8Y115_SLICE_X11Y115_BQ;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_C3 = CLBLM_L_X10Y109_SLICE_X13Y109_AO5;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_C4 = CLBLM_R_X11Y105_SLICE_X14Y105_CQ;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_C5 = CLBLM_L_X10Y108_SLICE_X13Y108_AQ;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_C6 = CLBLM_R_X13Y112_SLICE_X18Y112_A5Q;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_D4 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_D5 = 1'b1;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_A1 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_A2 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_A3 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_A4 = 1'b1;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_D3 = CLBLM_R_X13Y113_SLICE_X18Y113_DO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_D1 = CLBLM_R_X3Y110_SLICE_X2Y110_BO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_D2 = CLBLL_L_X4Y107_SLICE_X5Y107_BO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_D3 = CLBLM_R_X5Y115_SLICE_X7Y115_DO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_D4 = CLBLM_R_X7Y107_SLICE_X9Y107_C5Q;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_D5 = CLBLM_L_X10Y109_SLICE_X13Y109_BO5;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_D6 = CLBLM_L_X8Y109_SLICE_X11Y109_CQ;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_B3 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_B2 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_B4 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_AX = CLBLM_R_X11Y117_SLICE_X15Y117_AQ;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_B5 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_B6 = 1'b1;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_A1 = CLBLM_L_X10Y105_SLICE_X12Y105_AQ;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_A2 = CLBLM_R_X11Y105_SLICE_X14Y105_C5Q;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_A3 = CLBLM_L_X10Y106_SLICE_X12Y106_AQ;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_A4 = CLBLM_R_X11Y105_SLICE_X14Y105_CQ;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_A5 = CLBLM_L_X8Y115_SLICE_X10Y115_AQ;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_A6 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_C1 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_CE = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_C2 = 1'b1;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_B1 = CLBLM_R_X5Y112_SLICE_X6Y112_CQ;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_B2 = CLBLM_L_X10Y108_SLICE_X12Y108_BQ;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_B3 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_B4 = CLBLM_R_X11Y108_SLICE_X14Y108_AQ;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_B6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_D1 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_D4 = 1'b1;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_C1 = CLBLM_L_X10Y110_SLICE_X12Y110_CO5;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_C2 = 1'b1;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_C3 = CLBLM_R_X5Y108_SLICE_X7Y108_AQ;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_C4 = CLBLM_R_X11Y105_SLICE_X15Y105_A5Q;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_C6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_D6 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_SR = CLBLM_L_X12Y117_SLICE_X16Y117_AO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y161_OLOGIC_X0Y162_T1 = 1'b1;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_D1 = CLBLM_L_X10Y110_SLICE_X12Y110_AQ;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_D2 = CLBLM_L_X8Y112_SLICE_X10Y112_AQ;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_D3 = CLBLM_R_X11Y108_SLICE_X15Y108_AO5;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_D4 = CLBLM_L_X10Y108_SLICE_X12Y108_AO5;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_D5 = CLBLM_R_X5Y115_SLICE_X7Y115_CO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_D6 = CLBLM_L_X8Y108_SLICE_X10Y108_CQ;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOI3_X0Y101_OLOGIC_X0Y102_D1 = CLBLL_L_X2Y106_SLICE_X0Y106_BO5;
  assign LIOI3_X0Y161_OLOGIC_X0Y161_D1 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign LIOI3_X0Y101_OLOGIC_X0Y102_T1 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_A5 = CLBLM_R_X11Y110_SLICE_X14Y110_AQ;
  assign LIOI3_X0Y161_OLOGIC_X0Y161_T1 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_A6 = CLBLM_L_X8Y112_SLICE_X10Y112_BO6;
  assign LIOI3_X0Y101_OLOGIC_X0Y101_D1 = CLBLL_L_X2Y107_SLICE_X0Y107_AO6;
  assign LIOI3_X0Y101_OLOGIC_X0Y101_T1 = 1'b1;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_A1 = 1'b1;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_A2 = 1'b1;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_A3 = 1'b1;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_A4 = 1'b1;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_A5 = 1'b1;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_A6 = 1'b1;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_B1 = 1'b1;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_B2 = 1'b1;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_B3 = 1'b1;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_B4 = 1'b1;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_B5 = 1'b1;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_B6 = 1'b1;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_C1 = 1'b1;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_C2 = 1'b1;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_C3 = 1'b1;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_C4 = 1'b1;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_C5 = 1'b1;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_C6 = 1'b1;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_D1 = 1'b1;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_D2 = 1'b1;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_D3 = 1'b1;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_D4 = 1'b1;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_D5 = 1'b1;
  assign CLBLM_R_X13Y112_SLICE_X19Y112_D6 = 1'b1;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_A1 = CLBLM_L_X12Y112_SLICE_X16Y112_A5Q;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_A2 = CLBLM_R_X5Y112_SLICE_X6Y112_BQ;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_A3 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_A4 = CLBLM_L_X12Y114_SLICE_X17Y114_BQ;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_A6 = 1'b1;
  assign CLBLM_R_X13Y106_SLICE_X18Y106_D4 = CLBLM_R_X13Y106_SLICE_X18Y106_CO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X13Y106_SLICE_X18Y106_D5 = CLBLM_R_X13Y107_SLICE_X19Y107_BQ;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_B1 = CLBLM_R_X13Y112_SLICE_X18Y112_DO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_C2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_B2 = CLBLM_R_X13Y112_SLICE_X18Y112_BQ;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y106_SLICE_X18Y106_D6 = CLBLM_R_X13Y107_SLICE_X18Y107_AQ;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_B4 = CLBLM_L_X12Y111_SLICE_X16Y111_CQ;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_C3 = CLBLM_R_X7Y116_SLICE_X8Y116_CQ;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_B5 = CLBLM_L_X12Y113_SLICE_X17Y113_B5Q;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_C2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_C3 = 1'b1;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_C4 = CLBLM_L_X10Y114_SLICE_X13Y114_AQ;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_C5 = 1'b1;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_C6 = CLBLM_L_X12Y109_SLICE_X17Y109_CQ;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_C5 = CLBLM_R_X3Y110_SLICE_X3Y110_DO6;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_D1 = CLBLM_R_X13Y110_SLICE_X18Y110_BQ;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_D2 = CLBLM_L_X12Y111_SLICE_X16Y111_DQ;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_D3 = CLBLM_R_X13Y112_SLICE_X18Y112_BQ;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_D4 = 1'b1;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_D5 = 1'b1;
  assign CLBLM_R_X13Y112_SLICE_X18Y112_D6 = CLBLM_L_X10Y112_SLICE_X13Y112_AO6;
  assign LIOB33_X0Y161_IOB_X0Y161_O = RIOB33_X105Y107_IOB_X1Y108_I;
  assign LIOB33_X0Y161_IOB_X0Y162_O = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_B4 = 1'b1;
  assign RIOI3_X105Y145_ILOGIC_X1Y146_D = RIOB33_X105Y145_IOB_X1Y146_I;
  assign RIOI3_X105Y145_ILOGIC_X1Y145_D = RIOB33_X105Y145_IOB_X1Y145_I;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_A1 = CLBLM_L_X10Y105_SLICE_X12Y105_AQ;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_A2 = CLBLM_R_X11Y105_SLICE_X14Y105_C5Q;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_A3 = CLBLM_L_X10Y106_SLICE_X12Y106_AQ;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_A4 = CLBLM_R_X11Y105_SLICE_X14Y105_CQ;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_A5 = CLBLM_L_X10Y115_SLICE_X13Y115_BQ;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_A6 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_B5 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y64_D = LIOB33_X0Y63_IOB_X0Y64_I;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_B1 = CLBLM_L_X10Y105_SLICE_X12Y105_AQ;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_B2 = CLBLM_R_X11Y105_SLICE_X14Y105_C5Q;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_B3 = CLBLM_L_X10Y106_SLICE_X12Y106_AQ;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_B4 = CLBLM_R_X7Y110_SLICE_X8Y110_CQ;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_B5 = CLBLM_R_X11Y105_SLICE_X14Y105_CQ;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_B6 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y63_D = LIOB33_X0Y63_IOB_X0Y63_I;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_C1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_C2 = CLBLM_R_X11Y111_SLICE_X15Y111_BQ;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_C3 = CLBLM_L_X8Y109_SLICE_X11Y109_AQ;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_C4 = CLBLL_L_X2Y110_SLICE_X1Y110_DO6;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_C5 = CLBLM_R_X7Y109_SLICE_X8Y109_DO5;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_C6 = CLBLM_L_X10Y109_SLICE_X12Y109_CO5;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_B6 = 1'b1;
  assign LIOI3_X0Y179_OLOGIC_X0Y180_D1 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_D1 = CLBLM_R_X11Y111_SLICE_X15Y111_C5Q;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_D2 = CLBLM_R_X3Y107_SLICE_X3Y107_CO6;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_D3 = CLBLM_R_X5Y115_SLICE_X7Y115_DO6;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_D4 = CLBLM_R_X11Y115_SLICE_X15Y115_BQ;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_D5 = CLBLM_L_X10Y109_SLICE_X13Y109_AO6;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_D6 = CLBLM_L_X10Y109_SLICE_X13Y109_BO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_A1 = 1'b1;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_A2 = CLBLM_R_X7Y116_SLICE_X8Y116_CQ;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_A3 = CLBLM_L_X10Y109_SLICE_X12Y109_AQ;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_A4 = CLBLM_R_X5Y115_SLICE_X7Y115_CO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_A6 = CLBLM_L_X10Y114_SLICE_X12Y114_CQ;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_B2 = CLBLM_L_X10Y109_SLICE_X12Y109_BQ;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_B4 = CLBLM_R_X5Y108_SLICE_X7Y108_AQ;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_B5 = 1'b1;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_B6 = 1'b1;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_C1 = CLBLM_L_X10Y104_SLICE_X12Y104_AQ;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_C2 = CLBLM_R_X7Y116_SLICE_X8Y116_CQ;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_C3 = CLBLM_L_X8Y109_SLICE_X11Y109_DO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_C5 = CLBLM_R_X3Y111_SLICE_X2Y111_CO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_C6 = 1'b1;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_D1 = CLBLM_L_X10Y104_SLICE_X12Y104_AQ;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_D2 = CLBLM_L_X10Y110_SLICE_X12Y110_CO5;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_D3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_D4 = CLBLM_L_X8Y104_SLICE_X11Y104_AO5;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_D5 = CLBLM_R_X3Y111_SLICE_X2Y111_CO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_D6 = CLBLM_R_X7Y116_SLICE_X8Y116_CQ;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_D1 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_A1 = RIOB33_X105Y139_IOB_X1Y139_I;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_A2 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_A3 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_A4 = RIOB33_X105Y137_IOB_X1Y138_I;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_A5 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_A6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_B1 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_B2 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_B3 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_B4 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_B5 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_B6 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_C1 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_C2 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_C3 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_C4 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_C5 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_C6 = 1'b1;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_A1 = 1'b1;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_A2 = CLBLM_L_X8Y119_SLICE_X10Y119_AQ;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_A3 = CLBLM_R_X13Y113_SLICE_X19Y113_AQ;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_A4 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_A5 = CLBLM_R_X13Y108_SLICE_X18Y108_AQ;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_D1 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_D2 = 1'b1;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_B1 = 1'b1;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_B2 = 1'b1;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_B3 = 1'b1;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_B4 = 1'b1;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_B5 = 1'b1;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_B6 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_A1 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_A2 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_A3 = 1'b1;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_C1 = 1'b1;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_C2 = 1'b1;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_C3 = 1'b1;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_C4 = 1'b1;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_C5 = 1'b1;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_C6 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_A4 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_A5 = 1'b1;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_A6 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_B1 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_B2 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_B3 = 1'b1;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_D1 = 1'b1;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_D2 = 1'b1;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_D3 = 1'b1;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_D4 = 1'b1;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_D5 = 1'b1;
  assign CLBLM_R_X13Y113_SLICE_X19Y113_D6 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_C1 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_C2 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_C3 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_C4 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_C5 = 1'b1;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_A1 = CLBLM_R_X13Y113_SLICE_X18Y113_DO6;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_A3 = CLBLM_L_X12Y115_SLICE_X16Y115_AQ;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_A4 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_A5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_A6 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_D1 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_D2 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_D3 = 1'b1;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_B2 = CLBLM_R_X13Y109_SLICE_X19Y109_BQ;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_B3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_B4 = CLBLM_R_X7Y115_SLICE_X8Y115_D5Q;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_B5 = CLBLM_R_X13Y113_SLICE_X18Y113_BQ;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_B6 = CLBLM_R_X13Y108_SLICE_X18Y108_BO6;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_D4 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_D5 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_D6 = 1'b1;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_C2 = CLBLM_R_X13Y113_SLICE_X18Y113_CQ;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_C3 = CLBLM_L_X12Y114_SLICE_X17Y114_BQ;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_C4 = CLBLM_R_X5Y115_SLICE_X7Y115_CO6;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_C5 = CLBLM_L_X12Y112_SLICE_X16Y112_A5Q;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_C6 = 1'b1;
  assign LIOI3_X0Y59_ILOGIC_X0Y60_D = LIOB33_X0Y59_IOB_X0Y60_I;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_T1 = 1'b1;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_D1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_D2 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_D3 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_D4 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_D5 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X13Y113_SLICE_X18Y113_D6 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign LIOI3_X0Y59_ILOGIC_X0Y59_D = LIOB33_X0Y59_IOB_X0Y59_I;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_C4 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_D1 = CLBLL_L_X4Y117_SLICE_X4Y117_AQ;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_B3 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_B4 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_B5 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_C6 = 1'b1;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_A1 = CLBLM_R_X7Y111_SLICE_X8Y111_AQ;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_A4 = CLBLM_L_X10Y106_SLICE_X12Y106_BO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_A5 = CLBLM_R_X11Y105_SLICE_X14Y105_AQ;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_A6 = CLBLM_L_X10Y110_SLICE_X13Y110_AQ;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_B1 = CLBLM_L_X10Y118_SLICE_X12Y118_BQ;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_B2 = CLBLM_L_X10Y110_SLICE_X13Y110_BQ;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_B3 = CLBLM_L_X10Y107_SLICE_X12Y107_AQ;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_B4 = CLBLM_L_X10Y106_SLICE_X12Y106_BO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_C2 = CLBLM_L_X10Y110_SLICE_X13Y110_CQ;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_C3 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_C4 = CLBLM_L_X10Y109_SLICE_X12Y109_CO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_C5 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_C6 = CLBLM_L_X10Y112_SLICE_X12Y112_BQ;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_D2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_D3 = CLBLM_L_X10Y110_SLICE_X13Y110_DQ;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_D4 = CLBLM_L_X10Y109_SLICE_X12Y109_CO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_D5 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_D6 = CLBLM_L_X8Y111_SLICE_X11Y111_AQ;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_A1 = CLBLM_R_X7Y115_SLICE_X9Y115_DO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_A2 = 1'b1;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_A3 = CLBLM_L_X10Y110_SLICE_X12Y110_AQ;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_A4 = CLBLM_R_X7Y110_SLICE_X8Y110_CQ;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_A5 = CLBLM_L_X8Y108_SLICE_X10Y108_AQ;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_B2 = CLBLM_L_X10Y110_SLICE_X12Y110_BQ;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_B4 = CLBLM_R_X5Y110_SLICE_X6Y110_AQ;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_B5 = CLBLM_L_X10Y107_SLICE_X12Y107_AQ;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_B6 = 1'b1;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_C1 = CLBLM_L_X10Y113_SLICE_X12Y113_BQ;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_C2 = CLBLM_R_X13Y112_SLICE_X18Y112_CQ;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_C3 = CLBLM_L_X10Y112_SLICE_X12Y112_CQ;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_C4 = CLBLM_L_X8Y110_SLICE_X11Y110_CQ;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_C5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_C6 = 1'b1;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_A1 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_A2 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_A3 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_A4 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_A5 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_A6 = 1'b1;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_D1 = 1'b1;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_D2 = CLBLM_L_X10Y106_SLICE_X13Y106_BQ;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_B1 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_B2 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_B3 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_B4 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_B5 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_B6 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_C1 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_C2 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_C3 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_C4 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_C5 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_C6 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_D1 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_D2 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_D3 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_D4 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_D5 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_D6 = 1'b1;
  assign LIOB33_X0Y165_IOB_X0Y166_O = RIOB33_X105Y113_IOB_X1Y113_I;
  assign LIOB33_X0Y165_IOB_X0Y165_O = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_A1 = CLBLM_R_X5Y107_SLICE_X6Y107_CQ;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_A2 = CLBLM_R_X3Y110_SLICE_X2Y110_DO6;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_A3 = CLBLL_L_X4Y106_SLICE_X5Y106_AQ;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_A6 = CLBLM_R_X7Y105_SLICE_X8Y105_BO5;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_B2 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_B3 = CLBLL_L_X4Y106_SLICE_X5Y106_AQ;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_B4 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_B6 = CLBLM_R_X7Y108_SLICE_X8Y108_CQ;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_C1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_C2 = CLBLM_R_X3Y116_SLICE_X3Y116_AO6;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_C3 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_C4 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_C5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_C6 = CLBLM_R_X5Y106_SLICE_X6Y106_AQ;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y165_OLOGIC_X0Y166_D1 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_D1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_D2 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_D3 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_D4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_D5 = CLBLM_L_X12Y106_SLICE_X16Y106_AQ;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_D6 = CLBLM_R_X3Y116_SLICE_X3Y116_AO6;
  assign LIOI3_X0Y165_OLOGIC_X0Y166_T1 = 1'b1;
  assign LIOI3_X0Y103_OLOGIC_X0Y104_D1 = CLBLL_L_X2Y106_SLICE_X0Y106_CO6;
  assign LIOI3_X0Y165_OLOGIC_X0Y165_D1 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign LIOI3_X0Y103_OLOGIC_X0Y104_T1 = 1'b1;
  assign LIOI3_X0Y165_OLOGIC_X0Y165_T1 = 1'b1;
  assign LIOI3_X0Y103_OLOGIC_X0Y103_D1 = CLBLM_R_X3Y107_SLICE_X3Y107_BO6;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_B6 = 1'b1;
  assign LIOI3_X0Y103_OLOGIC_X0Y103_T1 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_C1 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_C2 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_C3 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_C4 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_C5 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_C6 = 1'b1;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_A2 = CLBLM_R_X11Y115_SLICE_X15Y115_AQ;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_A3 = CLBLM_L_X10Y111_SLICE_X13Y111_AQ;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_A4 = CLBLM_R_X11Y106_SLICE_X14Y106_BQ;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_A5 = CLBLL_L_X4Y116_SLICE_X4Y116_BO6;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_A6 = 1'b1;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_B1 = CLBLM_L_X10Y110_SLICE_X13Y110_AQ;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_B2 = CLBLM_L_X10Y111_SLICE_X13Y111_BQ;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_B3 = CLBLM_L_X10Y106_SLICE_X12Y106_BO6;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_B4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_B6 = CLBLM_L_X8Y114_SLICE_X11Y114_AQ;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_D1 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_D2 = 1'b1;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_C2 = CLBLM_L_X8Y106_SLICE_X10Y106_BQ;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_C3 = CLBLM_R_X11Y111_SLICE_X15Y111_AQ;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_C4 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_C5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_C6 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_D3 = 1'b1;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_D4 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_D5 = 1'b1;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_D1 = CLBLM_L_X10Y111_SLICE_X13Y111_C5Q;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_D2 = CLBLL_L_X2Y110_SLICE_X1Y110_DO6;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_D3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_D4 = CLBLM_R_X7Y109_SLICE_X8Y109_DO5;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_D5 = CLBLM_L_X10Y109_SLICE_X12Y109_CO5;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_D6 = CLBLM_L_X8Y111_SLICE_X11Y111_BQ;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_D6 = 1'b1;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_A1 = CLBLM_L_X10Y114_SLICE_X12Y114_DQ;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_A2 = CLBLM_L_X10Y110_SLICE_X12Y110_CO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_A5 = 1'b1;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_A6 = CLBLM_R_X5Y109_SLICE_X7Y109_AQ;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_AX = CLBLM_L_X10Y113_SLICE_X12Y113_DO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_B1 = 1'b1;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_B2 = CLBLM_L_X10Y111_SLICE_X12Y111_BQ;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_B4 = CLBLM_L_X8Y113_SLICE_X11Y113_BQ;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_B5 = 1'b1;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_C2 = CLBLM_R_X11Y109_SLICE_X14Y109_BQ;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_C3 = CLBLM_R_X11Y110_SLICE_X15Y110_BQ;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_C4 = CLBLM_R_X13Y113_SLICE_X18Y113_AQ;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_C5 = CLBLM_L_X8Y117_SLICE_X10Y117_BQ;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_C6 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_A1 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_A1 = CLBLM_L_X10Y108_SLICE_X13Y108_AQ;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_A3 = LIOB33_X0Y53_IOB_X0Y53_I;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_A4 = CLBLL_L_X4Y113_SLICE_X4Y113_BQ;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_A6 = CLBLM_R_X3Y109_SLICE_X2Y109_AQ;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_AX = CLBLL_L_X4Y107_SLICE_X4Y107_BO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_D2 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_B2 = CLBLM_R_X7Y105_SLICE_X8Y105_CQ;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_B3 = CLBLL_L_X4Y109_SLICE_X4Y109_AQ;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_B4 = CLBLL_L_X4Y110_SLICE_X4Y110_AQ;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_B6 = 1'b1;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_D3 = CLBLM_L_X10Y108_SLICE_X12Y108_BQ;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_D4 = CLBLM_L_X8Y112_SLICE_X10Y112_A5Q;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_D6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_C1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_C2 = CLBLL_L_X4Y107_SLICE_X4Y107_CQ;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_C4 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_C5 = CLBLL_L_X4Y110_SLICE_X4Y110_CQ;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_C6 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_A6 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_X105Y147_ILOGIC_X1Y148_D = RIOB33_X105Y147_IOB_X1Y148_I;
  assign RIOI3_X105Y147_ILOGIC_X1Y147_D = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_C1 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_D1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_D2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_D3 = CLBLL_L_X4Y107_SLICE_X4Y107_DQ;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_D4 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_D5 = CLBLM_L_X10Y108_SLICE_X13Y108_AQ;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_D6 = CLBLM_R_X3Y109_SLICE_X2Y109_A5Q;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_C2 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_C3 = 1'b1;
  assign LIOB33_X0Y167_IOB_X0Y167_O = RIOB33_X105Y113_IOB_X1Y114_I;
  assign LIOB33_X0Y167_IOB_X0Y168_O = RIOB33_X105Y123_IOB_X1Y123_I;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_C4 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_C5 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_C6 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_B2 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_B3 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_A1 = CLBLM_R_X11Y106_SLICE_X15Y106_DO5;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_A2 = CLBLM_R_X11Y115_SLICE_X14Y115_BQ;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_A3 = CLBLM_R_X11Y105_SLICE_X15Y105_AQ;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_A4 = CLBLM_R_X11Y105_SLICE_X15Y105_DO5;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_A1 = CLBLM_R_X5Y107_SLICE_X6Y107_CQ;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_A2 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_A3 = CLBLL_L_X4Y107_SLICE_X5Y107_AQ;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_A5 = CLBLL_L_X4Y112_SLICE_X4Y112_CO5;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_A6 = CLBLM_R_X5Y107_SLICE_X6Y107_DQ;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_B3 = CLBLL_L_X4Y107_SLICE_X4Y107_A5Q;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_A6 = CLBLM_L_X12Y105_SLICE_X16Y105_BO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_B1 = CLBLM_R_X3Y109_SLICE_X2Y109_CO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_B2 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_B3 = CLBLM_R_X3Y110_SLICE_X2Y110_DO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_B4 = CLBLM_R_X3Y110_SLICE_X3Y110_AO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_B5 = CLBLM_R_X3Y111_SLICE_X2Y111_CO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_B6 = 1'b1;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_B3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_B6 = CLBLM_R_X11Y106_SLICE_X15Y106_CO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_C1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_C2 = CLBLM_R_X7Y109_SLICE_X8Y109_AQ;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_C3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_C4 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_C5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_C6 = CLBLM_R_X3Y116_SLICE_X3Y116_AO6;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_C3 = CLBLM_L_X12Y105_SLICE_X16Y105_CO5;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_C4 = CLBLM_L_X12Y105_SLICE_X16Y105_BO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_C6 = CLBLM_L_X12Y108_SLICE_X17Y108_BQ;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_D2 = CLBLM_L_X12Y105_SLICE_X16Y105_BO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_D1 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_D2 = CLBLM_R_X3Y108_SLICE_X2Y108_DO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_D3 = CLBLL_L_X2Y111_SLICE_X1Y111_DO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_D4 = CLBLM_R_X3Y110_SLICE_X3Y110_DO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_D5 = CLBLL_L_X4Y107_SLICE_X5Y107_BO5;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_D6 = CLBLL_L_X2Y110_SLICE_X1Y110_DO6;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_D3 = CLBLM_L_X12Y112_SLICE_X16Y112_CQ;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_D4 = CLBLM_R_X11Y105_SLICE_X15Y105_A5Q;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_A1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_A3 = CLBLM_R_X11Y105_SLICE_X14Y105_AQ;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_A4 = CLBLM_L_X10Y106_SLICE_X12Y106_BO6;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_A5 = CLBLM_L_X10Y105_SLICE_X12Y105_BQ;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_A6 = CLBLM_R_X11Y105_SLICE_X15Y105_CQ;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_D2 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_D3 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_D4 = 1'b1;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_B2 = CLBLM_R_X11Y105_SLICE_X14Y105_BQ;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_B3 = CLBLM_L_X10Y111_SLICE_X13Y111_BQ;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_B4 = CLBLM_L_X10Y106_SLICE_X12Y106_BO6;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_B6 = CLBLM_R_X13Y112_SLICE_X18Y112_BQ;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_C4 = CLBLL_L_X2Y111_SLICE_X1Y111_DO6;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_D5 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_D6 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_C5 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_C5 = CLBLM_R_X3Y108_SLICE_X2Y108_DO6;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_C2 = CLBLL_L_X4Y112_SLICE_X4Y112_BQ;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_C3 = CLBLM_L_X10Y105_SLICE_X13Y105_AO6;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_C4 = CLBLM_L_X10Y105_SLICE_X13Y105_BO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_C6 = 1'b1;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_C5 = CLBLM_R_X13Y107_SLICE_X19Y107_AQ;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_C6 = 1'b1;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_D2 = CLBLM_R_X11Y106_SLICE_X15Y106_DO5;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_D3 = CLBLM_R_X11Y105_SLICE_X14Y105_DQ;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_D4 = CLBLM_L_X12Y105_SLICE_X16Y105_BO6;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_D5 = CLBLM_L_X12Y105_SLICE_X17Y105_AO6;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_D6 = CLBLL_L_X4Y107_SLICE_X4Y107_AQ;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_A1 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_A2 = CLBLM_L_X10Y116_SLICE_X13Y116_BQ;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_A3 = CLBLM_R_X11Y119_SLICE_X14Y119_AQ;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_A4 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_D1 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_D2 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_A6 = CLBLM_L_X8Y119_SLICE_X10Y119_AQ;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_D5 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_D6 = CLBLM_L_X10Y114_SLICE_X13Y114_BQ;
  assign RIOB33_X105Y165_IOB_X1Y166_O = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_B2 = 1'b1;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_A1 = CLBLM_R_X11Y112_SLICE_X14Y112_CQ;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_A2 = CLBLM_R_X13Y112_SLICE_X18Y112_CQ;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_A3 = CLBLM_R_X5Y109_SLICE_X6Y109_DQ;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_A4 = CLBLM_L_X10Y112_SLICE_X13Y112_BO6;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_A5 = CLBLM_R_X7Y112_SLICE_X8Y112_C5Q;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_A6 = CLBLM_L_X10Y112_SLICE_X13Y112_CO6;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_B3 = 1'b1;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_AX = CLBLM_R_X7Y115_SLICE_X9Y115_A5Q;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_B4 = 1'b1;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_B1 = CLBLM_L_X10Y112_SLICE_X13Y112_DO6;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_B2 = CLBLM_R_X7Y110_SLICE_X8Y110_BQ;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_B3 = CLBLM_L_X12Y112_SLICE_X17Y112_DO6;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_B4 = CLBLM_R_X11Y112_SLICE_X14Y112_DO6;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_B5 = CLBLM_R_X5Y114_SLICE_X7Y114_BQ;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_B6 = CLBLM_R_X11Y112_SLICE_X15Y112_BQ;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_B5 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_B6 = 1'b1;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_C1 = 1'b1;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_C2 = CLBLM_L_X10Y111_SLICE_X12Y111_DQ;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_C3 = CLBLM_L_X10Y112_SLICE_X12Y112_CQ;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_C4 = CLBLM_L_X8Y112_SLICE_X10Y112_A5Q;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_C5 = CLBLM_R_X11Y111_SLICE_X15Y111_AQ;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_C6 = 1'b1;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_CE = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_D1 = CLBLM_R_X11Y112_SLICE_X14Y112_BQ;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_D2 = CLBLM_R_X7Y112_SLICE_X9Y112_BQ;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_D3 = CLBLM_L_X10Y111_SLICE_X13Y111_C5Q;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_D4 = 1'b1;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_D5 = 1'b1;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_D6 = CLBLM_L_X12Y111_SLICE_X16Y111_DQ;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_SR = CLBLM_L_X12Y117_SLICE_X16Y117_AO6;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_A1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_A2 = CLBLM_R_X13Y113_SLICE_X18Y113_DO6;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_A3 = CLBLM_L_X8Y110_SLICE_X11Y110_A5Q;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_A4 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_A6 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_C1 = 1'b1;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_B1 = 1'b1;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_B2 = CLBLM_L_X10Y112_SLICE_X12Y112_BQ;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_B4 = CLBLM_R_X7Y112_SLICE_X8Y112_CQ;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_B5 = CLBLM_L_X12Y112_SLICE_X16Y112_BQ;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_C2 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_C3 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_C4 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_C5 = 1'b1;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_C2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_C3 = CLBLM_R_X7Y118_SLICE_X8Y118_CQ;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_C4 = CLBLM_L_X10Y111_SLICE_X12Y111_DQ;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_C5 = CLBLM_L_X12Y112_SLICE_X16Y112_B5Q;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_C6 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_A2 = CLBLL_L_X4Y110_SLICE_X4Y110_AQ;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_A3 = CLBLL_L_X4Y108_SLICE_X4Y108_AQ;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_A4 = CLBLM_R_X7Y106_SLICE_X9Y106_AQ;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_A5 = CLBLM_R_X7Y105_SLICE_X8Y105_CQ;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_A6 = CLBLL_L_X4Y108_SLICE_X4Y108_BQ;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_C6 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_B1 = CLBLL_L_X4Y112_SLICE_X4Y112_CO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_B3 = CLBLM_R_X7Y107_SLICE_X9Y107_CQ;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_D4 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_D5 = 1'b1;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_D6 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_B4 = CLBLM_R_X5Y114_SLICE_X7Y114_CQ;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_B5 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_B6 = CLBLL_L_X4Y108_SLICE_X4Y108_BQ;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_D1 = 1'b1;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_D2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_C1 = LIOB33_X0Y53_IOB_X0Y53_I;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_C2 = CLBLM_R_X3Y109_SLICE_X2Y109_AQ;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_C3 = CLBLM_R_X5Y110_SLICE_X6Y110_B5Q;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_C4 = CLBLL_L_X4Y113_SLICE_X4Y113_BQ;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_C6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_D1 = CLBLL_L_X2Y110_SLICE_X0Y110_AO5;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_D2 = CLBLL_L_X4Y107_SLICE_X5Y107_AQ;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_D3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_D4 = CLBLL_L_X4Y108_SLICE_X4Y108_BQ;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_D5 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_D6 = CLBLM_R_X3Y116_SLICE_X3Y116_AO6;
  assign RIOI3_X105Y185_OLOGIC_X1Y185_D1 = CLBLM_L_X8Y110_SLICE_X10Y110_CO5;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_A1 = CLBLL_L_X2Y111_SLICE_X1Y111_DO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_A3 = CLBLM_R_X3Y110_SLICE_X3Y110_DO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_A4 = CLBLM_R_X3Y109_SLICE_X2Y109_CO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_A5 = CLBLM_R_X3Y108_SLICE_X2Y108_DO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_A6 = 1'b1;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_A1 = CLBLM_R_X11Y106_SLICE_X15Y106_BO5;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_A2 = CLBLM_L_X12Y105_SLICE_X16Y105_BO6;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_A3 = CLBLM_R_X11Y106_SLICE_X15Y106_AQ;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_B1 = CLBLL_L_X4Y112_SLICE_X5Y112_CO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_B2 = CLBLL_L_X2Y110_SLICE_X0Y110_BO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_B3 = CLBLM_R_X7Y106_SLICE_X8Y106_CQ;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_B4 = CLBLM_R_X5Y111_SLICE_X6Y111_BQ;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_B5 = CLBLL_L_X4Y107_SLICE_X5Y107_CO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_B6 = CLBLL_L_X2Y108_SLICE_X1Y108_AO5;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_B1 = CLBLM_L_X10Y111_SLICE_X12Y111_A5Q;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_B2 = CLBLM_R_X11Y105_SLICE_X15Y105_AQ;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_C1 = CLBLL_L_X2Y112_SLICE_X0Y112_AO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_C2 = CLBLM_R_X3Y116_SLICE_X3Y116_AO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_C3 = CLBLM_R_X5Y109_SLICE_X7Y109_BQ;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_C4 = CLBLL_L_X2Y114_SLICE_X0Y114_AO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_C5 = CLBLM_R_X5Y105_SLICE_X7Y105_AQ;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_C6 = CLBLL_L_X2Y108_SLICE_X1Y108_BO6;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_C1 = CLBLM_L_X12Y105_SLICE_X16Y105_BO6;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_C2 = CLBLM_L_X12Y108_SLICE_X17Y108_BQ;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_C3 = CLBLM_R_X11Y105_SLICE_X15Y105_CQ;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_C4 = CLBLM_R_X11Y108_SLICE_X14Y108_AQ;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_C5 = CLBLM_L_X12Y105_SLICE_X16Y105_CO5;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_C6 = 1'b1;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_D1 = CLBLM_R_X7Y108_SLICE_X8Y108_BQ;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_D2 = CLBLL_L_X2Y114_SLICE_X0Y114_AO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_D3 = CLBLM_R_X5Y107_SLICE_X7Y107_B5Q;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_D4 = CLBLM_R_X3Y116_SLICE_X3Y116_AO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_D5 = CLBLL_L_X2Y109_SLICE_X0Y109_AO5;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_D6 = CLBLL_L_X2Y108_SLICE_X1Y108_BO6;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_D4 = CLBLM_L_X12Y112_SLICE_X16Y112_CQ;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_D5 = CLBLM_R_X11Y106_SLICE_X15Y106_AQ;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_D6 = 1'b1;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_D3 = CLBLM_R_X11Y106_SLICE_X14Y106_BQ;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_A1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_A2 = CLBLM_R_X11Y106_SLICE_X14Y106_DQ;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_A3 = CLBLM_R_X11Y106_SLICE_X14Y106_AQ;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_A4 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_A5 = CLBLM_L_X12Y111_SLICE_X16Y111_AQ;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign RIOI3_X105Y103_ILOGIC_X1Y104_D = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_B1 = 1'b1;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_B2 = CLBLM_R_X11Y106_SLICE_X14Y106_BQ;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_B3 = CLBLM_L_X12Y105_SLICE_X16Y105_BO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_B4 = CLBLM_R_X7Y106_SLICE_X8Y106_BQ;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_B6 = CLBLM_R_X11Y106_SLICE_X15Y106_DO6;
  assign LIOB33_X0Y131_IOB_X0Y131_O = CLBLM_L_X8Y119_SLICE_X10Y119_AO5;
  assign LIOB33_X0Y131_IOB_X0Y132_O = CLBLM_L_X8Y119_SLICE_X10Y119_AQ;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_C1 = CLBLM_L_X12Y105_SLICE_X16Y105_CO5;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_C2 = CLBLM_R_X11Y106_SLICE_X14Y106_CQ;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_C4 = CLBLM_R_X3Y113_SLICE_X3Y113_AQ;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_C5 = CLBLM_L_X12Y107_SLICE_X16Y107_DQ;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_C6 = CLBLM_L_X12Y105_SLICE_X16Y105_BO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_D1 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_D2 = CLBLM_R_X11Y109_SLICE_X14Y109_AQ;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_D3 = CLBLM_R_X11Y106_SLICE_X14Y106_DQ;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_D4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_D5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_D6 = CLBLM_R_X11Y105_SLICE_X14Y105_BQ;
  assign LIOI3_X0Y109_OLOGIC_X0Y109_T1 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_B4 = CLBLM_R_X11Y107_SLICE_X15Y107_BQ;
  assign LIOI3_X0Y167_OLOGIC_X0Y168_D1 = RIOB33_X105Y123_IOB_X1Y123_I;
  assign RIOI3_X105Y103_ILOGIC_X1Y103_D = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_B5 = CLBLM_R_X11Y109_SLICE_X15Y109_AO6;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_B6 = CLBLM_R_X11Y111_SLICE_X15Y111_CQ;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y167_OLOGIC_X0Y168_T1 = 1'b1;
  assign LIOI3_X0Y105_OLOGIC_X0Y106_D1 = CLBLL_L_X2Y106_SLICE_X0Y106_AO5;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_A1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_A2 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_A3 = CLBLM_L_X10Y113_SLICE_X13Y113_AQ;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_A5 = CLBLM_L_X10Y113_SLICE_X13Y113_C5Q;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_A6 = CLBLM_L_X10Y113_SLICE_X12Y113_CQ;
  assign LIOI3_X0Y167_OLOGIC_X0Y167_D1 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_B1 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_B2 = CLBLM_L_X10Y113_SLICE_X13Y113_BQ;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_B3 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_B5 = CLBLM_L_X10Y113_SLICE_X13Y113_C5Q;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_B6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign LIOI3_X0Y105_OLOGIC_X0Y106_T1 = 1'b1;
  assign RIOI3_X105Y151_OLOGIC_X1Y152_D1 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign LIOI3_X0Y167_OLOGIC_X0Y167_T1 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_C2 = CLBLM_L_X10Y113_SLICE_X13Y113_CQ;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_C3 = CLBLM_L_X8Y113_SLICE_X10Y113_DQ;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_C4 = RIOB33_X105Y119_IOB_X1Y119_I;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_C5 = CLBLM_R_X5Y109_SLICE_X7Y109_BQ;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_C6 = 1'b1;
  assign LIOI3_X0Y105_OLOGIC_X0Y105_D1 = CLBLL_L_X2Y106_SLICE_X0Y106_CO5;
  assign RIOI3_X105Y151_OLOGIC_X1Y152_T1 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_D1 = CLBLM_R_X7Y113_SLICE_X8Y113_CQ;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_D2 = CLBLM_L_X8Y114_SLICE_X11Y114_B5Q;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_D3 = CLBLM_L_X10Y113_SLICE_X13Y113_DQ;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_D4 = CLBLM_R_X7Y108_SLICE_X9Y108_AQ;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_D5 = CLBLM_R_X13Y113_SLICE_X18Y113_CQ;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_D6 = CLBLM_L_X10Y104_SLICE_X12Y104_BO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_D3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign LIOI3_X0Y105_OLOGIC_X0Y105_T1 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_D4 = CLBLM_L_X8Y107_SLICE_X10Y107_BQ;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_T1 = 1'b1;
  assign RIOI3_X105Y151_OLOGIC_X1Y151_D1 = LIOB33_X0Y75_IOB_X0Y76_I;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_A1 = CLBLM_L_X10Y110_SLICE_X13Y110_AQ;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_A3 = CLBLM_L_X10Y113_SLICE_X12Y113_AQ;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_A4 = CLBLM_R_X11Y110_SLICE_X15Y110_BQ;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_A5 = CLBLL_L_X4Y116_SLICE_X4Y116_BO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_A6 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_D6 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_D1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign RIOI3_X105Y151_OLOGIC_X1Y151_T1 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_B2 = CLBLM_L_X10Y113_SLICE_X12Y113_BQ;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_B3 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_B4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_B5 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_B6 = CLBLM_L_X8Y112_SLICE_X11Y112_CO6;
  assign LIOB33_X0Y171_IOB_X0Y171_O = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign LIOB33_X0Y171_IOB_X0Y172_O = CLBLM_R_X103Y138_SLICE_X163Y138_AO6;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_T1 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_C1 = CLBLM_L_X10Y111_SLICE_X12Y111_AQ;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A1 = CLBLL_L_X4Y112_SLICE_X4Y112_CO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A2 = CLBLL_L_X4Y110_SLICE_X4Y110_BQ;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A3 = CLBLL_L_X4Y109_SLICE_X4Y109_AQ;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_C5 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A4 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A5 = CLBLM_R_X5Y111_SLICE_X7Y111_AQ;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_C2 = CLBLM_L_X10Y113_SLICE_X12Y113_CQ;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_C3 = CLBLM_R_X11Y109_SLICE_X14Y109_BQ;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_C4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B1 = CLBLM_R_X7Y105_SLICE_X8Y105_BO5;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B2 = CLBLL_L_X4Y109_SLICE_X4Y109_BQ;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B3 = CLBLM_L_X12Y110_SLICE_X17Y110_BQ;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_D2 = CLBLM_L_X12Y113_SLICE_X17Y113_CQ;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B6 = CLBLL_L_X2Y110_SLICE_X1Y110_DO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_D5 = CLBLM_R_X5Y114_SLICE_X7Y114_BQ;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C1 = CLBLL_L_X2Y108_SLICE_X1Y108_AO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C2 = CLBLM_R_X7Y109_SLICE_X9Y109_BQ;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C3 = CLBLL_L_X2Y110_SLICE_X0Y110_BO5;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C4 = CLBLL_L_X2Y111_SLICE_X1Y111_AO5;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C5 = CLBLM_L_X12Y112_SLICE_X16Y112_AQ;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C6 = CLBLM_R_X7Y107_SLICE_X8Y107_AQ;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D1 = CLBLL_L_X2Y108_SLICE_X1Y108_AO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D2 = CLBLM_R_X3Y112_SLICE_X3Y112_BO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D3 = CLBLM_R_X11Y114_SLICE_X14Y114_AQ;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D4 = CLBLL_L_X4Y108_SLICE_X4Y108_DO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D5 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D6 = CLBLM_R_X7Y108_SLICE_X8Y108_AQ;
  assign RIOI3_X105Y185_OLOGIC_X1Y185_T1 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_A1 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_A2 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_A3 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_C2 = CLBLM_L_X8Y116_SLICE_X11Y116_BQ;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_A4 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_A5 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_A6 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_B1 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_B2 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_B3 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_B4 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X19Y117_B5 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A1 = CLBLM_R_X5Y109_SLICE_X7Y109_DQ;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A3 = CLBLL_L_X4Y109_SLICE_X5Y109_AQ;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A5 = CLBLM_R_X7Y113_SLICE_X9Y113_DO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A6 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_A1 = CLBLM_R_X11Y107_SLICE_X15Y107_DO6;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_A2 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_A3 = CLBLM_L_X8Y114_SLICE_X11Y114_B5Q;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B1 = CLBLM_R_X3Y112_SLICE_X2Y112_AO5;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B2 = CLBLL_L_X4Y106_SLICE_X5Y106_DO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B3 = CLBLL_L_X4Y106_SLICE_X5Y106_AQ;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B4 = CLBLL_L_X2Y110_SLICE_X0Y110_BO5;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B5 = CLBLL_L_X4Y113_SLICE_X5Y113_AQ;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B6 = CLBLL_L_X4Y109_SLICE_X5Y109_CO6;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_A4 = 1'b1;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_A6 = CLBLM_L_X8Y119_SLICE_X10Y119_AQ;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C2 = CLBLM_L_X12Y109_SLICE_X16Y109_D5Q;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C4 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C5 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C6 = CLBLM_R_X3Y116_SLICE_X3Y116_AO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_B5 = CLBLL_L_X4Y112_SLICE_X4Y112_CO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_B6 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_B6 = CLBLM_L_X8Y119_SLICE_X10Y119_AQ;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_C2 = CLBLM_R_X11Y107_SLICE_X15Y107_CQ;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_C3 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D1 = CLBLL_L_X4Y109_SLICE_X4Y109_AQ;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D2 = CLBLM_R_X7Y115_SLICE_X8Y115_AQ;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D3 = CLBLM_R_X3Y112_SLICE_X2Y112_AO5;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D4 = CLBLL_L_X2Y110_SLICE_X0Y110_BO5;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D5 = CLBLL_L_X2Y111_SLICE_X1Y111_AO5;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D6 = CLBLM_R_X5Y107_SLICE_X6Y107_AQ;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_D1 = CLBLM_L_X8Y109_SLICE_X10Y109_C5Q;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_D2 = CLBLM_R_X11Y108_SLICE_X15Y108_AO5;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_D3 = CLBLM_R_X5Y115_SLICE_X7Y115_CO6;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_D4 = CLBLM_R_X11Y107_SLICE_X15Y107_AQ;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_D5 = CLBLM_R_X11Y110_SLICE_X14Y110_CQ;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_D6 = CLBLM_R_X11Y107_SLICE_X14Y107_AO6;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_AX = CLBLM_R_X13Y118_SLICE_X18Y118_AO5;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_B1 = 1'b1;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_A1 = CLBLM_R_X11Y105_SLICE_X14Y105_CQ;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_A2 = CLBLM_L_X10Y105_SLICE_X12Y105_AQ;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_A3 = CLBLM_L_X10Y106_SLICE_X12Y106_AQ;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_A4 = CLBLM_L_X8Y115_SLICE_X11Y115_BQ;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_A5 = CLBLM_R_X11Y105_SLICE_X14Y105_C5Q;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_A6 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_BX = CLBLM_R_X13Y117_SLICE_X18Y117_AO6;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_C1 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_C2 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_C3 = 1'b1;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_B1 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_B2 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_B3 = CLBLM_L_X8Y107_SLICE_X11Y107_BQ;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_B4 = CLBLM_L_X12Y109_SLICE_X16Y109_AQ;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_B5 = CLBLM_L_X10Y116_SLICE_X13Y116_AQ;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_B6 = CLBLM_L_X8Y107_SLICE_X11Y107_B5Q;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_D5 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_D3 = CLBLM_L_X10Y115_SLICE_X12Y115_CQ;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_C1 = CLBLM_R_X11Y105_SLICE_X14Y105_C5Q;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_C2 = CLBLM_R_X11Y105_SLICE_X14Y105_CQ;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_C3 = CLBLM_L_X10Y106_SLICE_X12Y106_AQ;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_D4 = CLBLM_L_X10Y115_SLICE_X13Y115_DO5;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_C4 = 1'b1;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_C5 = CLBLM_R_X11Y110_SLICE_X14Y110_CQ;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_C6 = CLBLM_L_X10Y105_SLICE_X12Y105_AQ;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_D3 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_D4 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_D5 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_D6 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_D1 = CLBLM_L_X8Y109_SLICE_X10Y109_C5Q;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_D2 = CLBLM_R_X5Y115_SLICE_X7Y115_DO6;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_D3 = 1'b1;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_D4 = CLBLM_R_X11Y107_SLICE_X14Y107_CO6;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_D5 = CLBLM_R_X3Y110_SLICE_X2Y110_BO6;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_D6 = CLBLL_L_X4Y107_SLICE_X5Y107_BO6;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_A1 = CLBLM_L_X10Y114_SLICE_X13Y114_DO6;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_A3 = CLBLM_L_X10Y114_SLICE_X13Y114_AQ;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_A4 = CLBLM_L_X8Y115_SLICE_X11Y115_CO6;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_A5 = CLBLM_L_X12Y114_SLICE_X16Y114_AQ;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_A6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_B1 = CLBLL_L_X4Y116_SLICE_X4Y116_BO6;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_B2 = CLBLM_R_X11Y115_SLICE_X15Y115_BQ;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_B4 = CLBLM_L_X12Y112_SLICE_X17Y112_BQ;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_B5 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_B6 = CLBLM_L_X10Y114_SLICE_X13Y114_BQ;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_A1 = CLBLM_L_X10Y110_SLICE_X13Y110_CQ;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_A2 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_A3 = CLBLM_L_X8Y105_SLICE_X11Y105_CO6;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_A4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_A6 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_C2 = CLBLM_L_X10Y114_SLICE_X13Y114_CQ;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_C3 = CLBLM_L_X10Y114_SLICE_X13Y114_BQ;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_B1 = CLBLM_L_X8Y105_SLICE_X11Y105_DO6;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_B2 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_B3 = CLBLM_R_X5Y105_SLICE_X6Y105_AQ;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_B4 = CLBLM_L_X8Y105_SLICE_X11Y105_BQ;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_B5 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_B6 = CLBLM_L_X8Y105_SLICE_X10Y105_CO6;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_D1 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_C1 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_C2 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_C3 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_C4 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_C5 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_C6 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_D3 = CLBLM_L_X10Y115_SLICE_X13Y115_DO6;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_D4 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_A1 = CLBLM_R_X7Y115_SLICE_X8Y115_B5Q;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_A2 = CLBLM_L_X12Y114_SLICE_X16Y114_AQ;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_A3 = CLBLM_L_X10Y114_SLICE_X12Y114_AQ;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_A5 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_D1 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_D2 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_D3 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_D4 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_D5 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_D6 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_A6 = CLBLM_R_X7Y115_SLICE_X9Y115_DO6;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_B1 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_B2 = CLBLM_L_X8Y108_SLICE_X10Y108_BQ;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_A1 = CLBLL_L_X4Y110_SLICE_X4Y110_B5Q;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_A2 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_A3 = CLBLM_R_X7Y105_SLICE_X8Y105_CQ;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_A3 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_A5 = CLBLL_L_X4Y110_SLICE_X4Y110_C5Q;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_A4 = CLBLM_L_X10Y106_SLICE_X12Y106_BO6;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_A5 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_A6 = CLBLM_L_X12Y110_SLICE_X16Y110_DO5;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_A6 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_A1 = CLBLM_L_X8Y114_SLICE_X11Y114_B5Q;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_A2 = CLBLM_L_X10Y104_SLICE_X12Y104_CO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_B4 = CLBLM_R_X5Y109_SLICE_X7Y109_A5Q;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_B5 = CLBLL_L_X4Y110_SLICE_X5Y110_AQ;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_B6 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_B1 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_B2 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_C1 = CLBLM_R_X5Y110_SLICE_X6Y110_AQ;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_D2 = CLBLM_L_X10Y114_SLICE_X12Y114_AQ;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_D3 = CLBLM_L_X10Y114_SLICE_X12Y114_DQ;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_D4 = CLBLM_R_X7Y115_SLICE_X9Y115_DO6;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_D5 = CLBLM_L_X8Y108_SLICE_X10Y108_DQ;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_D6 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_C2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_B6 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_C3 = CLBLL_L_X4Y107_SLICE_X4Y107_A5Q;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_C1 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_C2 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_C3 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_C4 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_C5 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_C6 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_D1 = CLBLL_L_X2Y110_SLICE_X0Y110_CO5;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_D2 = CLBLM_R_X3Y112_SLICE_X3Y112_BO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_D3 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_D4 = CLBLM_L_X10Y111_SLICE_X13Y111_AQ;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_D1 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_D2 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_D3 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_D4 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_D5 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_D6 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_A1 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_A2 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_A3 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_A4 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_A5 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_A6 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_A1 = CLBLM_R_X5Y110_SLICE_X7Y110_B5Q;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_A2 = CLBLM_L_X8Y110_SLICE_X11Y110_BO5;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_A3 = CLBLM_R_X5Y115_SLICE_X7Y115_CO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_A4 = CLBLM_R_X5Y111_SLICE_X7Y111_AQ;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_A5 = CLBLM_R_X5Y110_SLICE_X7Y110_BQ;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_A6 = CLBLL_L_X4Y113_SLICE_X5Y113_BQ;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_B1 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_B2 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_AX = CLBLM_R_X7Y110_SLICE_X8Y110_DO6;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_B3 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_B1 = CLBLM_R_X3Y112_SLICE_X2Y112_AO5;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_B2 = CLBLM_R_X5Y112_SLICE_X7Y112_AQ;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_B3 = CLBLL_L_X2Y111_SLICE_X1Y111_AO5;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_B4 = CLBLM_R_X7Y112_SLICE_X8Y112_AQ;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_B5 = CLBLM_L_X8Y116_SLICE_X10Y116_DQ;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_B6 = CLBLM_R_X3Y112_SLICE_X3Y112_BO5;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_A1 = CLBLM_L_X10Y105_SLICE_X12Y105_AQ;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_A2 = CLBLM_L_X10Y106_SLICE_X12Y106_AQ;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_A3 = CLBLM_R_X11Y105_SLICE_X14Y105_C5Q;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_C1 = CLBLL_L_X2Y108_SLICE_X1Y108_AO5;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_C2 = CLBLM_R_X5Y109_SLICE_X7Y109_DQ;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_C3 = CLBLM_R_X5Y112_SLICE_X6Y112_DO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_C4 = CLBLL_L_X4Y106_SLICE_X5Y106_CO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_C5 = CLBLM_L_X8Y113_SLICE_X10Y113_AQ;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_C6 = CLBLL_L_X2Y110_SLICE_X0Y110_BO5;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_AX = CLBLM_R_X11Y106_SLICE_X15Y106_BO6;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_B1 = CLBLM_L_X10Y105_SLICE_X12Y105_AQ;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_B2 = CLBLM_L_X10Y106_SLICE_X12Y106_AQ;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_B3 = CLBLM_R_X11Y105_SLICE_X14Y105_C5Q;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_B4 = CLBLM_L_X10Y110_SLICE_X12Y110_AQ;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_B5 = CLBLM_R_X11Y105_SLICE_X14Y105_CQ;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_B6 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_D1 = CLBLL_L_X2Y110_SLICE_X0Y110_CO5;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_D2 = CLBLM_R_X3Y112_SLICE_X3Y112_BO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_D3 = CLBLM_R_X5Y114_SLICE_X6Y114_CO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_D4 = CLBLM_L_X8Y111_SLICE_X11Y111_AQ;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_D5 = CLBLL_L_X4Y108_SLICE_X5Y108_DO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_D6 = CLBLL_L_X4Y111_SLICE_X4Y111_AQ;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_C3 = CLBLM_R_X11Y109_SLICE_X15Y109_AO5;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_C4 = CLBLM_R_X11Y108_SLICE_X15Y108_AQ;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_C6 = CLBLM_R_X3Y107_SLICE_X3Y107_CO6;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_D1 = CLBLM_R_X11Y105_SLICE_X14Y105_CQ;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_D2 = CLBLM_L_X12Y109_SLICE_X16Y109_DQ;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_D3 = CLBLM_R_X11Y105_SLICE_X14Y105_C5Q;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_D4 = CLBLM_L_X10Y105_SLICE_X12Y105_AQ;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_D5 = CLBLM_L_X12Y113_SLICE_X17Y113_DO6;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_D6 = CLBLM_L_X10Y106_SLICE_X12Y106_AQ;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_B1 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_B2 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_B3 = 1'b1;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_A2 = CLBLM_L_X12Y108_SLICE_X17Y108_AQ;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_A3 = CLBLM_R_X11Y108_SLICE_X14Y108_AQ;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_A4 = CLBLM_L_X12Y105_SLICE_X16Y105_BO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_A5 = CLBLM_L_X12Y105_SLICE_X16Y105_CO5;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_A6 = CLBLM_L_X8Y116_SLICE_X10Y116_BQ;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_C1 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_C2 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_C3 = 1'b1;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_B1 = CLBLM_R_X11Y108_SLICE_X14Y108_DO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_B2 = CLBLM_L_X10Y109_SLICE_X13Y109_DO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_B3 = CLBLM_R_X11Y108_SLICE_X15Y108_CO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_B4 = CLBLM_R_X11Y107_SLICE_X14Y107_DO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_B5 = CLBLM_L_X10Y108_SLICE_X13Y108_DO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_B6 = CLBLM_R_X11Y108_SLICE_X14Y108_CO6;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_D1 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_D2 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_D3 = 1'b1;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_C1 = CLBLM_R_X5Y115_SLICE_X7Y115_DO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_C2 = CLBLM_R_X13Y112_SLICE_X18Y112_A5Q;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_C3 = CLBLM_R_X11Y108_SLICE_X15Y108_BO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_C4 = CLBLM_R_X11Y107_SLICE_X14Y107_AO5;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_C5 = CLBLM_L_X8Y112_SLICE_X10Y112_AQ;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_C6 = CLBLM_R_X3Y107_SLICE_X3Y107_CO6;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_D4 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_D5 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_D6 = 1'b1;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_D1 = CLBLM_R_X5Y115_SLICE_X7Y115_DO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_D2 = CLBLM_R_X3Y110_SLICE_X2Y110_BO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_D3 = CLBLL_L_X4Y107_SLICE_X5Y107_BO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_D4 = 1'b1;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_D5 = CLBLM_R_X13Y117_SLICE_X18Y117_AQ;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_D6 = CLBLM_L_X10Y108_SLICE_X12Y108_AO6;
  assign LIOB33_X0Y175_IOB_X0Y176_O = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_A1 = CLBLM_R_X7Y112_SLICE_X9Y112_DO6;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_A2 = CLBLM_R_X5Y114_SLICE_X7Y114_BQ;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_A3 = CLBLM_L_X10Y115_SLICE_X13Y115_AQ;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_A5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_A6 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign LIOB33_X0Y175_IOB_X0Y175_O = RIOB33_X105Y127_IOB_X1Y127_I;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_B1 = CLBLM_L_X12Y113_SLICE_X17Y113_DO6;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_B2 = CLBLM_L_X10Y115_SLICE_X13Y115_BQ;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_B4 = 1'b1;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_B5 = CLBLM_R_X7Y117_SLICE_X9Y117_A5Q;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_B6 = CLBLM_R_X7Y115_SLICE_X9Y115_DO6;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_A1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_A2 = CLBLM_L_X8Y107_SLICE_X10Y107_BQ;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_A3 = CLBLM_L_X8Y105_SLICE_X11Y105_AQ;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_C4 = CLBLM_L_X10Y113_SLICE_X13Y113_CQ;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_C5 = CLBLM_R_X5Y108_SLICE_X6Y108_BO6;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_C6 = CLBLM_L_X10Y114_SLICE_X13Y114_CQ;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_A5 = CLBLM_L_X10Y106_SLICE_X12Y106_BO6;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_A6 = CLBLM_L_X12Y107_SLICE_X16Y107_AQ;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_C2 = CLBLM_L_X10Y117_SLICE_X13Y117_AO5;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_B2 = CLBLM_L_X8Y105_SLICE_X11Y105_BQ;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_B3 = CLBLM_R_X5Y105_SLICE_X6Y105_BQ;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_D2 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_B5 = CLBLM_L_X10Y106_SLICE_X12Y106_BO6;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_B6 = CLBLM_L_X8Y106_SLICE_X11Y106_BQ;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_D1 = CLBLM_R_X11Y110_SLICE_X15Y110_BQ;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_C1 = CLBLM_L_X8Y104_SLICE_X11Y104_AQ;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_C2 = CLBLM_R_X3Y108_SLICE_X2Y108_DO6;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_C3 = CLBLM_R_X11Y106_SLICE_X14Y106_AQ;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_C4 = CLBLM_L_X10Y112_SLICE_X12Y112_DO6;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_C5 = CLBLM_L_X10Y108_SLICE_X12Y108_BQ;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_C6 = CLBLM_L_X8Y106_SLICE_X10Y106_DO6;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_A1 = CLBLM_R_X11Y116_SLICE_X14Y116_AQ;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_A2 = 1'b1;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_A4 = CLBLM_R_X7Y115_SLICE_X9Y115_A5Q;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_A5 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_D1 = CLBLM_L_X8Y106_SLICE_X11Y106_AQ;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_D2 = CLBLM_L_X8Y105_SLICE_X11Y105_AQ;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_D3 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_D4 = CLBLM_L_X8Y107_SLICE_X10Y107_AQ;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_D5 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_D6 = CLBLM_L_X10Y107_SLICE_X12Y107_AQ;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_A1 = CLBLM_R_X5Y112_SLICE_X7Y112_CQ;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_A3 = CLBLL_L_X4Y111_SLICE_X4Y111_AQ;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_A4 = CLBLL_L_X4Y116_SLICE_X4Y116_BO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_A5 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_A6 = CLBLM_R_X5Y109_SLICE_X7Y109_B5Q;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_A1 = CLBLM_R_X7Y117_SLICE_X9Y117_DQ;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_A2 = CLBLM_L_X10Y106_SLICE_X12Y106_BO6;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_A3 = CLBLM_L_X8Y105_SLICE_X10Y105_AQ;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_A5 = CLBLM_R_X7Y105_SLICE_X9Y105_BQ;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_B1 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_B2 = CLBLM_R_X5Y109_SLICE_X6Y109_BQ;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_B3 = CLBLL_L_X4Y112_SLICE_X4Y112_CO5;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_B1 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_B2 = CLBLM_L_X8Y107_SLICE_X10Y107_AQ;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_B3 = CLBLM_R_X7Y107_SLICE_X8Y107_BQ;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_C2 = CLBLL_L_X4Y111_SLICE_X4Y111_CQ;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_C3 = CLBLM_R_X7Y105_SLICE_X8Y105_BO5;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_B4 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_C5 = CLBLM_R_X3Y111_SLICE_X2Y111_CO6;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_B5 = CLBLM_L_X8Y106_SLICE_X11Y106_AQ;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_B6 = CLBLM_R_X5Y105_SLICE_X6Y105_AQ;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_C1 = CLBLM_R_X7Y105_SLICE_X9Y105_BQ;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_C2 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_C3 = CLBLM_R_X7Y107_SLICE_X8Y107_BQ;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_C4 = CLBLM_L_X8Y106_SLICE_X10Y106_AQ;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_C5 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_C6 = CLBLM_L_X10Y110_SLICE_X13Y110_BQ;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_D1 = CLBLL_L_X2Y108_SLICE_X1Y108_AO6;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_D2 = CLBLL_L_X4Y114_SLICE_X4Y114_BQ;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_D3 = CLBLM_R_X5Y111_SLICE_X6Y111_AQ;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_D4 = CLBLL_L_X2Y111_SLICE_X1Y111_AO5;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_D5 = CLBLM_R_X7Y114_SLICE_X8Y114_BQ;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_D6 = CLBLL_L_X2Y110_SLICE_X0Y110_BO5;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_D1 = CLBLM_R_X7Y105_SLICE_X9Y105_BQ;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_D2 = CLBLM_L_X8Y105_SLICE_X10Y105_AQ;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_D3 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_D4 = CLBLM_L_X8Y105_SLICE_X11Y105_AQ;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_D5 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_D6 = 1'b1;
  assign LIOI3_X0Y109_OLOGIC_X0Y110_D1 = CLBLM_R_X3Y106_SLICE_X2Y106_AO6;
  assign LIOI3_X0Y171_OLOGIC_X0Y172_T1 = 1'b1;
  assign LIOI3_X0Y171_OLOGIC_X0Y171_D1 = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign LIOI3_X0Y109_OLOGIC_X0Y110_T1 = 1'b1;
  assign RIOI3_X105Y153_OLOGIC_X1Y154_D1 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_A1 = CLBLL_L_X4Y110_SLICE_X4Y110_AQ;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_A2 = CLBLM_R_X5Y105_SLICE_X7Y105_BQ;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_A3 = CLBLL_L_X4Y111_SLICE_X5Y111_AQ;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_A5 = CLBLM_R_X7Y105_SLICE_X8Y105_CQ;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_A6 = CLBLM_R_X5Y110_SLICE_X7Y110_BQ;
  assign LIOI3_X0Y109_OLOGIC_X0Y109_D1 = CLBLL_L_X2Y107_SLICE_X1Y107_AO5;
  assign LIOI3_X0Y171_OLOGIC_X0Y171_T1 = 1'b1;
  assign RIOI3_X105Y153_OLOGIC_X1Y154_T1 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_B1 = CLBLM_R_X5Y110_SLICE_X7Y110_B5Q;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_B2 = CLBLM_R_X11Y112_SLICE_X15Y112_CO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_B3 = CLBLM_R_X5Y111_SLICE_X7Y111_AQ;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_B4 = CLBLL_L_X4Y113_SLICE_X5Y113_BQ;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_B5 = CLBLM_R_X5Y115_SLICE_X7Y115_CO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_B6 = CLBLM_R_X5Y110_SLICE_X7Y110_BQ;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_A1 = CLBLM_L_X10Y105_SLICE_X12Y105_AQ;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_A2 = CLBLM_R_X11Y105_SLICE_X14Y105_CQ;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_A3 = CLBLM_R_X11Y105_SLICE_X14Y105_C5Q;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_C1 = CLBLM_L_X8Y110_SLICE_X11Y110_BO5;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_C2 = CLBLL_L_X4Y113_SLICE_X5Y113_BQ;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_C3 = CLBLM_R_X5Y110_SLICE_X7Y110_B5Q;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_C4 = CLBLM_R_X5Y110_SLICE_X7Y110_BQ;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_C5 = CLBLM_R_X5Y111_SLICE_X7Y111_AQ;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_C6 = CLBLM_R_X5Y115_SLICE_X7Y115_CO6;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_A4 = CLBLM_R_X11Y113_SLICE_X15Y113_AQ;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_A5 = CLBLM_L_X10Y106_SLICE_X12Y106_AQ;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_A6 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_B1 = CLBLM_R_X5Y115_SLICE_X7Y115_CO6;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_B2 = CLBLM_R_X11Y113_SLICE_X15Y113_AQ;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_B3 = CLBLM_R_X11Y105_SLICE_X14Y105_CQ;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_D1 = CLBLL_L_X4Y108_SLICE_X5Y108_CO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_D2 = CLBLL_L_X2Y111_SLICE_X1Y111_AO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_D3 = CLBLL_L_X4Y114_SLICE_X5Y114_DO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_D4 = CLBLM_R_X5Y113_SLICE_X7Y113_CO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_D5 = CLBLM_R_X7Y111_SLICE_X9Y111_BQ;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_D6 = CLBLL_L_X4Y113_SLICE_X5Y113_CO6;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_C1 = CLBLM_R_X5Y115_SLICE_X7Y115_CO6;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_C2 = CLBLM_R_X11Y105_SLICE_X14Y105_C5Q;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_C3 = CLBLM_L_X12Y113_SLICE_X17Y113_DO6;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_C4 = CLBLM_L_X12Y109_SLICE_X16Y109_DQ;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_C5 = CLBLM_L_X10Y106_SLICE_X12Y106_AQ;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_C6 = CLBLM_R_X11Y108_SLICE_X15Y108_AO5;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_D1 = CLBLM_R_X11Y113_SLICE_X15Y113_AQ;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_D2 = CLBLM_L_X10Y110_SLICE_X12Y110_AQ;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_D3 = CLBLM_R_X11Y110_SLICE_X14Y110_CQ;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_D4 = CLBLM_L_X8Y109_SLICE_X11Y109_CQ;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_D5 = CLBLM_L_X12Y110_SLICE_X17Y110_AQ;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_D6 = CLBLM_R_X7Y110_SLICE_X8Y110_CQ;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_T1 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_A1 = CLBLM_R_X11Y109_SLICE_X14Y109_DO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_A2 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_A3 = CLBLM_L_X8Y119_SLICE_X10Y119_AQ;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_A4 = CLBLM_R_X7Y108_SLICE_X8Y108_AQ;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_A6 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_B2 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_B3 = CLBLM_L_X8Y119_SLICE_X10Y119_AQ;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_B4 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_B5 = CLBLM_L_X10Y109_SLICE_X12Y109_BQ;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_B6 = CLBLM_R_X11Y109_SLICE_X14Y109_CO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_C1 = CLBLM_R_X11Y109_SLICE_X14Y109_BQ;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_C2 = CLBLM_L_X10Y105_SLICE_X12Y105_AQ;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_C3 = CLBLM_R_X5Y115_SLICE_X7Y115_CO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_C4 = CLBLM_R_X11Y108_SLICE_X15Y108_BO5;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_C5 = CLBLM_L_X10Y115_SLICE_X13Y115_BQ;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_C6 = CLBLM_R_X11Y111_SLICE_X15Y111_C5Q;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_T1 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_B4 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_D1 = CLBLM_L_X8Y115_SLICE_X10Y115_AQ;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_D2 = CLBLM_R_X11Y109_SLICE_X14Y109_AQ;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_D3 = CLBLM_L_X10Y105_SLICE_X12Y105_AQ;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_D4 = CLBLM_R_X5Y115_SLICE_X7Y115_CO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_D5 = CLBLM_R_X13Y117_SLICE_X18Y117_AQ;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_A5 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_D6 = CLBLM_R_X11Y108_SLICE_X15Y108_BO5;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_B5 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_B6 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_A6 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_C1 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_C2 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_C3 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_C4 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_B3 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_C5 = 1'b1;
  assign LIOB33_X0Y177_IOB_X0Y177_O = RIOB33_X105Y129_IOB_X1Y129_I;
  assign LIOB33_X0Y177_IOB_X0Y178_O = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_B4 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_C6 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_B5 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_B6 = 1'b1;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_A1 = CLBLM_R_X7Y118_SLICE_X8Y118_DO6;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_A3 = CLBLM_L_X10Y116_SLICE_X13Y116_AQ;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_A4 = CLBLM_L_X10Y116_SLICE_X12Y116_BQ;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_A5 = CLBLM_L_X10Y117_SLICE_X13Y117_AO5;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_A6 = CLBLM_L_X10Y111_SLICE_X13Y111_CQ;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_B1 = CLBLM_R_X7Y118_SLICE_X8Y118_DO6;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_B2 = CLBLM_L_X10Y116_SLICE_X13Y116_BQ;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_B3 = CLBLM_L_X10Y116_SLICE_X13Y116_AQ;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_B5 = CLBLL_L_X4Y114_SLICE_X4Y114_BQ;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_B6 = CLBLM_L_X10Y117_SLICE_X13Y117_AO5;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_A1 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_A3 = CLBLM_L_X8Y106_SLICE_X11Y106_AQ;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_A4 = CLBLM_L_X10Y106_SLICE_X13Y106_AQ;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_A5 = CLBLM_L_X8Y109_SLICE_X10Y109_DQ;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_A6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_C1 = CLBLM_R_X11Y117_SLICE_X14Y117_AO6;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_C2 = CLBLM_L_X10Y116_SLICE_X13Y116_CQ;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_AX = CLBLM_L_X8Y106_SLICE_X11Y106_CO6;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_C3 = CLBLM_L_X10Y116_SLICE_X12Y116_DO5;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_B2 = CLBLM_L_X8Y106_SLICE_X11Y106_BQ;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_B3 = CLBLM_L_X10Y106_SLICE_X12Y106_BO6;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_B4 = CLBLM_L_X8Y109_SLICE_X11Y109_AQ;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_B6 = CLBLM_L_X10Y106_SLICE_X13Y106_CQ;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_D1 = CLBLM_L_X10Y119_SLICE_X12Y119_AQ;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_C1 = CLBLM_R_X7Y106_SLICE_X8Y106_CQ;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_C2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_C3 = CLBLM_L_X8Y114_SLICE_X11Y114_B5Q;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_C4 = CLBLM_L_X10Y104_SLICE_X12Y104_BO6;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_C5 = CLBLM_L_X10Y107_SLICE_X12Y107_BQ;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_C6 = 1'b1;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_D3 = CLBLM_R_X7Y118_SLICE_X8Y118_CQ;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_D4 = CLBLM_R_X7Y114_SLICE_X8Y114_A5Q;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_A1 = CLBLM_R_X7Y118_SLICE_X8Y118_DO6;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_A3 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_A4 = CLBLM_R_X11Y116_SLICE_X14Y116_AQ;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_A5 = CLBLM_R_X7Y111_SLICE_X9Y111_AQ;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_D1 = CLBLM_L_X8Y110_SLICE_X11Y110_DQ;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_A1 = CLBLL_L_X4Y116_SLICE_X4Y116_BO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_A2 = CLBLM_L_X8Y108_SLICE_X10Y108_BQ;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_A3 = CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_D5 = CLBLM_L_X10Y106_SLICE_X13Y106_CQ;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_D6 = CLBLM_L_X8Y113_SLICE_X10Y113_BQ;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_A4 = CLBLL_L_X4Y111_SLICE_X4Y111_BQ;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_A6 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_D2 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_D3 = CLBLM_L_X10Y107_SLICE_X12Y107_BQ;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_A1 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_A2 = CLBLM_L_X12Y112_SLICE_X16Y112_CQ;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_A3 = CLBLM_L_X8Y106_SLICE_X10Y106_AQ;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_A5 = CLBLM_R_X7Y106_SLICE_X9Y106_BQ;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_A6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_B1 = CLBLL_L_X4Y117_SLICE_X4Y117_DQ;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_B2 = CLBLL_L_X4Y112_SLICE_X4Y112_BQ;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_C2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_C3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_C4 = CLBLM_R_X11Y113_SLICE_X14Y113_CQ;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_C5 = CLBLL_L_X4Y114_SLICE_X4Y114_BQ;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_B1 = CLBLM_R_X7Y107_SLICE_X8Y107_DO6;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_B2 = CLBLM_L_X8Y106_SLICE_X10Y106_BQ;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_B3 = CLBLM_L_X8Y110_SLICE_X11Y110_CQ;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_B4 = CLBLM_R_X7Y105_SLICE_X9Y105_CQ;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_B5 = CLBLM_L_X10Y113_SLICE_X13Y113_AQ;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_D3 = CLBLM_R_X7Y118_SLICE_X8Y118_CQ;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_D4 = CLBLM_L_X8Y118_SLICE_X10Y118_AQ;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_D5 = CLBLM_L_X10Y117_SLICE_X13Y117_CO6;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_D6 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_C1 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_D1 = CLBLL_L_X2Y108_SLICE_X1Y108_AO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_D2 = CLBLM_R_X3Y114_SLICE_X2Y114_DO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_D3 = CLBLL_L_X4Y112_SLICE_X5Y112_BO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_D4 = CLBLM_L_X10Y111_SLICE_X12Y111_C5Q;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_D5 = CLBLL_L_X4Y111_SLICE_X5Y111_AQ;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_D6 = CLBLM_R_X3Y112_SLICE_X3Y112_BO5;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_D1 = CLBLM_L_X8Y105_SLICE_X10Y105_BO6;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_D2 = CLBLM_L_X8Y106_SLICE_X10Y106_AQ;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_D3 = CLBLM_L_X8Y110_SLICE_X11Y110_DQ;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_D4 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_D5 = CLBLM_R_X5Y107_SLICE_X7Y107_AQ;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_D6 = CLBLM_L_X8Y113_SLICE_X10Y113_BQ;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_A5 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_A6 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_D6 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_A1 = CLBLL_L_X4Y112_SLICE_X4Y112_CO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_A2 = CLBLM_R_X7Y112_SLICE_X9Y112_AQ;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_A3 = CLBLL_L_X4Y112_SLICE_X5Y112_AQ;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_A5 = CLBLM_R_X11Y110_SLICE_X14Y110_D5Q;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_A6 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_B1 = CLBLL_L_X26Y136_SLICE_X38Y136_AO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_B2 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_B3 = CLBLL_L_X4Y112_SLICE_X5Y112_AQ;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_B4 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_B5 = CLBLM_R_X7Y106_SLICE_X8Y106_BQ;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_B6 = CLBLL_L_X2Y112_SLICE_X0Y112_AO5;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_C1 = CLBLL_L_X2Y112_SLICE_X0Y112_AO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_C2 = CLBLL_L_X2Y112_SLICE_X0Y112_AO5;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_C3 = CLBLL_L_X2Y114_SLICE_X0Y114_AO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_C4 = CLBLM_R_X7Y112_SLICE_X8Y112_DQ;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_C5 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_C6 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_B4 = CLBLM_R_X5Y111_SLICE_X6Y111_CQ;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_B5 = CLBLL_L_X4Y111_SLICE_X4Y111_BQ;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_A1 = CLBLM_R_X7Y115_SLICE_X8Y115_DQ;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_A3 = CLBLM_R_X11Y110_SLICE_X15Y110_AQ;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_A6 = CLBLM_L_X8Y114_SLICE_X10Y114_CQ;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_D1 = CLBLM_R_X7Y108_SLICE_X8Y108_CQ;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_D2 = CLBLM_R_X11Y113_SLICE_X14Y113_CQ;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_D3 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_D4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_D5 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_D6 = CLBLL_L_X4Y114_SLICE_X4Y114_BQ;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_B4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_B6 = CLBLM_L_X10Y111_SLICE_X12Y111_A5Q;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_C1 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_C2 = CLBLM_R_X11Y110_SLICE_X15Y110_CQ;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_C3 = CLBLM_L_X10Y114_SLICE_X13Y114_CQ;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_C4 = CLBLM_R_X5Y115_SLICE_X7Y115_CO6;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_C5 = CLBLM_R_X11Y110_SLICE_X15Y110_AQ;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_D1 = CLBLM_L_X8Y109_SLICE_X10Y109_C5Q;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_D2 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_D3 = CLBLM_L_X10Y114_SLICE_X13Y114_CQ;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_D4 = CLBLM_L_X10Y109_SLICE_X12Y109_AQ;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_D5 = CLBLM_R_X11Y108_SLICE_X15Y108_AQ;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_D6 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_C6 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_A2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_A3 = CLBLM_R_X11Y110_SLICE_X14Y110_AQ;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_A4 = CLBLM_R_X13Y110_SLICE_X18Y110_AQ;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_A5 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_A6 = CLBLM_L_X10Y110_SLICE_X12Y110_B5Q;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_AX = CLBLM_R_X11Y110_SLICE_X14Y110_BO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_B1 = CLBLM_R_X13Y112_SLICE_X18Y112_CQ;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_C6 = CLBLM_R_X7Y110_SLICE_X8Y110_CQ;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_B2 = CLBLM_R_X11Y107_SLICE_X15Y107_BQ;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_B3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_B4 = CLBLM_R_X13Y110_SLICE_X19Y110_BQ;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_B6 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_C4 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_C1 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_C2 = CLBLM_R_X11Y110_SLICE_X14Y110_CQ;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_C3 = CLBLM_L_X8Y115_SLICE_X11Y115_BQ;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_C4 = CLBLM_R_X13Y110_SLICE_X19Y110_BQ;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_C5 = CLBLM_R_X7Y115_SLICE_X9Y115_DO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_C5 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_C6 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_D2 = CLBLM_R_X11Y112_SLICE_X14Y112_C5Q;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_D3 = CLBLM_R_X11Y105_SLICE_X14Y105_AQ;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_D4 = CLBLM_R_X11Y109_SLICE_X14Y109_AQ;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_D5 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_D6 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_D2 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_D3 = 1'b1;
  assign LIOB33_X0Y179_IOB_X0Y180_O = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_D4 = 1'b1;
  assign LIOB33_X0Y179_IOB_X0Y179_O = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_D5 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_D1 = RIOB33_X105Y143_IOB_X1Y144_I;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I0 = LIOB33_X0Y77_IOB_X0Y78_I;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I1 = 1'b1;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_A1 = CLBLM_R_X7Y118_SLICE_X9Y118_BO5;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_A2 = CLBLM_R_X7Y114_SLICE_X8Y114_A5Q;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_A3 = CLBLM_R_X7Y118_SLICE_X8Y118_CQ;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_A4 = CLBLM_L_X8Y118_SLICE_X10Y118_AQ;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_A5 = CLBLM_L_X10Y119_SLICE_X12Y119_AQ;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_A6 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_B3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_B4 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_B1 = CLBLM_L_X10Y116_SLICE_X13Y116_CQ;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_B2 = CLBLM_R_X11Y117_SLICE_X15Y117_CQ;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_B3 = CLBLM_L_X12Y117_SLICE_X17Y117_BQ;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_B4 = CLBLM_L_X10Y117_SLICE_X12Y117_BQ;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_B5 = CLBLM_L_X10Y119_SLICE_X12Y119_CO6;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_B6 = 1'b1;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_A1 = CLBLM_L_X8Y107_SLICE_X11Y107_B5Q;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_A2 = CLBLM_L_X8Y107_SLICE_X11Y107_BQ;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_A3 = CLBLM_L_X8Y107_SLICE_X11Y107_AQ;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_A4 = CLBLM_L_X8Y107_SLICE_X11Y107_DO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_A5 = CLBLM_L_X8Y107_SLICE_X11Y107_A5Q;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_A6 = 1'b1;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_C1 = CLBLM_R_X11Y117_SLICE_X15Y117_DQ;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_C2 = CLBLM_R_X11Y117_SLICE_X15Y117_CQ;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_C3 = CLBLM_R_X7Y118_SLICE_X9Y118_CO5;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_B1 = CLBLM_L_X8Y107_SLICE_X11Y107_B5Q;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_B2 = CLBLM_L_X8Y107_SLICE_X11Y107_BQ;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_B3 = 1'b1;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_B4 = CLBLM_L_X8Y107_SLICE_X11Y107_DO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_B5 = CLBLM_L_X8Y107_SLICE_X11Y107_A5Q;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_B6 = 1'b1;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_D2 = CLBLM_L_X12Y117_SLICE_X17Y117_BQ;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_D3 = 1'b1;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_D4 = CLBLM_R_X11Y117_SLICE_X14Y117_DO6;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_D5 = CLBLM_L_X10Y116_SLICE_X13Y116_CQ;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_D6 = CLBLM_L_X10Y117_SLICE_X12Y117_BQ;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_C4 = CLBLM_R_X5Y115_SLICE_X7Y115_CO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_C2 = CLBLM_L_X8Y107_SLICE_X11Y107_CQ;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_C3 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_A1 = RIOB33_X105Y143_IOB_X1Y144_I;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_A2 = CLBLM_L_X10Y116_SLICE_X13Y116_CQ;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_A4 = CLBLM_R_X3Y114_SLICE_X2Y114_BQ;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_A5 = 1'b1;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_A6 = 1'b1;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_C6 = CLBLM_L_X8Y110_SLICE_X10Y110_BQ;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_C6 = CLBLM_L_X10Y109_SLICE_X12Y109_AQ;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A1 = CLBLM_R_X5Y114_SLICE_X7Y114_AQ;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_B1 = CLBLM_L_X10Y118_SLICE_X13Y118_CO6;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_B2 = CLBLM_L_X10Y117_SLICE_X12Y117_BQ;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_B4 = CLBLM_R_X7Y115_SLICE_X8Y115_DQ;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_B5 = CLBLM_L_X10Y116_SLICE_X12Y116_DO5;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_B6 = CLBLM_L_X10Y117_SLICE_X12Y117_CO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A6 = 1'b1;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_D4 = CLBLM_L_X8Y107_SLICE_X11Y107_A5Q;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B1 = CLBLL_L_X4Y116_SLICE_X5Y116_A5Q;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_C1 = CLBLM_L_X8Y116_SLICE_X11Y116_CO6;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_C2 = CLBLM_L_X8Y116_SLICE_X10Y116_CQ;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_C3 = CLBLM_L_X10Y116_SLICE_X13Y116_CQ;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_C4 = CLBLM_L_X10Y119_SLICE_X12Y119_CO6;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_C5 = CLBLM_L_X10Y117_SLICE_X12Y117_DO6;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_C6 = CLBLM_L_X10Y119_SLICE_X12Y119_BO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_A1 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_A2 = CLBLM_L_X10Y109_SLICE_X12Y109_AQ;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C2 = CLBLM_R_X3Y109_SLICE_X2Y109_A5Q;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C3 = CLBLL_L_X4Y113_SLICE_X5Y113_B5Q;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C4 = CLBLM_L_X12Y113_SLICE_X17Y113_BQ;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_D1 = CLBLM_L_X10Y119_SLICE_X12Y119_AQ;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_D2 = CLBLM_R_X11Y117_SLICE_X15Y117_AQ;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_D3 = CLBLM_R_X7Y118_SLICE_X9Y118_BO5;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_D4 = CLBLM_L_X8Y118_SLICE_X10Y118_AQ;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_D5 = CLBLM_R_X7Y118_SLICE_X8Y118_CQ;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_D6 = CLBLM_R_X7Y114_SLICE_X8Y114_A5Q;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D1 = CLBLM_R_X3Y116_SLICE_X3Y116_AO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D2 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D3 = CLBLL_L_X4Y113_SLICE_X4Y113_AQ;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D4 = CLBLL_L_X2Y110_SLICE_X0Y110_AO5;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D5 = CLBLM_R_X5Y113_SLICE_X6Y113_AQ;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D6 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_C5 = CLBLM_L_X12Y106_SLICE_X16Y106_AQ;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_C6 = CLBLM_R_X3Y108_SLICE_X2Y108_BO6;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_D2 = CLBLM_R_X5Y112_SLICE_X7Y112_CQ;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_D1 = 1'b1;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_D2 = CLBLM_L_X8Y107_SLICE_X10Y107_CQ;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_D3 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_D4 = 1'b1;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_D5 = 1'b1;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_D6 = CLBLM_L_X8Y119_SLICE_X10Y119_AQ;
  assign RIOI3_SING_X105Y150_OLOGIC_X1Y150_T1 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_D5 = CLBLM_R_X11Y114_SLICE_X14Y114_CQ;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A1 = CLBLL_L_X4Y112_SLICE_X4Y112_CO5;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A2 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A3 = CLBLL_L_X4Y113_SLICE_X5Y113_AQ;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A5 = CLBLL_L_X4Y113_SLICE_X4Y113_AQ;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A6 = CLBLM_R_X7Y115_SLICE_X9Y115_A5Q;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_D6 = CLBLM_L_X8Y108_SLICE_X10Y108_BQ;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B1 = CLBLL_L_X4Y111_SLICE_X5Y111_CO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B2 = CLBLL_L_X4Y111_SLICE_X5Y111_BO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B4 = CLBLM_R_X7Y112_SLICE_X9Y112_AQ;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B5 = CLBLM_L_X12Y113_SLICE_X16Y113_AQ;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B6 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C1 = CLBLM_R_X3Y116_SLICE_X3Y116_AO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C3 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C4 = CLBLL_L_X2Y114_SLICE_X0Y114_AO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C5 = CLBLL_L_X2Y110_SLICE_X0Y110_AO5;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C6 = CLBLM_R_X7Y113_SLICE_X8Y113_BQ;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_A1 = CLBLM_R_X11Y112_SLICE_X14Y112_BQ;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_A3 = CLBLM_L_X10Y106_SLICE_X12Y106_AQ;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_A4 = 1'b1;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_A5 = 1'b1;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_A6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D2 = CLBLM_R_X5Y111_SLICE_X6Y111_DO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D3 = CLBLM_R_X5Y115_SLICE_X7Y115_CO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D4 = CLBLM_R_X11Y112_SLICE_X15Y112_CO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D5 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D6 = CLBLL_L_X4Y113_SLICE_X4Y113_CO5;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_B1 = 1'b1;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_B2 = CLBLM_R_X11Y112_SLICE_X15Y112_BQ;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_B3 = CLBLM_R_X5Y106_SLICE_X6Y106_BQ;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_B5 = 1'b1;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_C1 = CLBLM_L_X10Y118_SLICE_X12Y118_AQ;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_C2 = CLBLM_R_X11Y110_SLICE_X14Y110_A5Q;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_C3 = CLBLM_R_X5Y111_SLICE_X6Y111_BQ;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_C5 = CLBLM_R_X11Y110_SLICE_X15Y110_A5Q;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_C6 = 1'b1;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_D1 = CLBLM_R_X11Y110_SLICE_X15Y110_CQ;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_D2 = CLBLM_R_X11Y110_SLICE_X15Y110_DO6;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_D3 = CLBLM_R_X11Y114_SLICE_X14Y114_DQ;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_D4 = CLBLM_R_X7Y107_SLICE_X9Y107_C5Q;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_D5 = 1'b1;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_D6 = CLBLM_R_X11Y115_SLICE_X15Y115_BQ;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_A1 = CLBLM_R_X11Y114_SLICE_X14Y114_BQ;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_A2 = CLBLM_R_X7Y110_SLICE_X8Y110_CQ;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_A3 = CLBLM_R_X11Y109_SLICE_X15Y109_AO6;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_A4 = CLBLM_R_X11Y105_SLICE_X14Y105_CQ;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_A5 = CLBLM_R_X5Y115_SLICE_X7Y115_CO6;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_A6 = CLBLM_R_X11Y115_SLICE_X15Y115_BQ;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_B1 = CLBLL_L_X4Y107_SLICE_X5Y107_BO6;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_B2 = CLBLM_R_X7Y110_SLICE_X8Y110_CQ;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_B3 = CLBLM_R_X11Y115_SLICE_X14Y115_CO6;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_B4 = CLBLM_R_X3Y110_SLICE_X2Y110_BO6;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_B5 = CLBLM_R_X5Y115_SLICE_X7Y115_DO6;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_B6 = CLBLM_R_X11Y111_SLICE_X14Y111_CO6;
  assign LIOI3_X0Y173_OLOGIC_X0Y174_D1 = CLBLM_L_X10Y148_SLICE_X12Y148_AO6;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_C1 = CLBLM_L_X10Y106_SLICE_X13Y106_DO6;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_C2 = CLBLM_L_X10Y110_SLICE_X12Y110_DO6;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_C3 = CLBLM_L_X12Y113_SLICE_X17Y113_BQ;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_C4 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_C5 = CLBLM_R_X11Y111_SLICE_X14Y111_DO6;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_C6 = CLBLM_L_X8Y107_SLICE_X11Y107_BQ;
  assign LIOB33_X0Y181_IOB_X0Y181_O = RIOB33_X105Y133_IOB_X1Y133_I;
  assign LIOB33_X0Y181_IOB_X0Y182_O = RIOB33_X105Y133_IOB_X1Y134_I;
  assign LIOI3_X0Y173_OLOGIC_X0Y174_T1 = 1'b1;
  assign LIOI3_X0Y111_OLOGIC_X0Y112_D1 = CLBLM_R_X11Y110_SLICE_X14Y110_D5Q;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_D1 = CLBLM_R_X11Y113_SLICE_X15Y113_AQ;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_B4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_D2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_D3 = 1'b1;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_D4 = CLBLM_R_X7Y118_SLICE_X8Y118_CQ;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_D5 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_B5 = CLBLM_L_X10Y113_SLICE_X12Y113_DO5;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_D6 = CLBLM_L_X8Y107_SLICE_X11Y107_B5Q;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_B6 = CLBLM_L_X10Y116_SLICE_X12Y116_BQ;
  assign LIOI3_X0Y111_OLOGIC_X0Y112_T1 = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y156_D1 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_A2 = CLBLM_L_X12Y110_SLICE_X16Y110_CO6;
  assign LIOI3_X0Y173_OLOGIC_X0Y173_T1 = 1'b1;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_D1 = 1'b0;
  assign RIOI3_X105Y155_OLOGIC_X1Y156_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_D1 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_T1 = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y155_D1 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_T1 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign RIOI3_X105Y155_OLOGIC_X1Y155_T1 = 1'b1;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_C2 = CLBLM_L_X10Y114_SLICE_X12Y114_CQ;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_AX = CLBLM_L_X12Y110_SLICE_X16Y110_BO6;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_D1 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_C3 = CLBLM_R_X11Y113_SLICE_X15Y113_DQ;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_C4 = CLBLM_R_X5Y115_SLICE_X7Y115_CO6;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_B1 = CLBLM_L_X12Y110_SLICE_X16Y110_AO5;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_C5 = CLBLM_R_X5Y115_SLICE_X6Y115_BQ;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_T1 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_B2 = CLBLM_R_X11Y115_SLICE_X15Y115_AQ;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_C6 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_B5 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_A1 = CLBLM_L_X10Y118_SLICE_X13Y118_DO6;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_A2 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_A3 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_A5 = CLBLM_L_X10Y113_SLICE_X13Y113_DQ;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_A6 = CLBLM_L_X10Y118_SLICE_X13Y118_CO6;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_B1 = CLBLM_L_X10Y119_SLICE_X12Y119_BO6;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_B2 = CLBLM_L_X10Y117_SLICE_X12Y117_DO6;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_B3 = CLBLM_L_X10Y117_SLICE_X12Y117_BQ;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_B4 = CLBLM_R_X7Y118_SLICE_X9Y118_CO5;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_B5 = CLBLM_L_X10Y119_SLICE_X13Y119_AO6;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_B6 = CLBLM_L_X10Y116_SLICE_X12Y116_CQ;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_A1 = CLBLM_L_X8Y108_SLICE_X11Y108_AQ;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_A2 = CLBLM_L_X8Y108_SLICE_X11Y108_BQ;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_C3 = CLBLM_R_X7Y118_SLICE_X8Y118_CQ;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_C4 = CLBLM_L_X10Y117_SLICE_X13Y117_CO6;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_C5 = CLBLM_R_X11Y117_SLICE_X15Y117_AQ;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_A3 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_A5 = 1'b1;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_A6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_C1 = CLBLM_L_X8Y118_SLICE_X10Y118_AQ;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_C2 = CLBLM_L_X10Y119_SLICE_X12Y119_AQ;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_B1 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_B2 = CLBLM_R_X7Y108_SLICE_X9Y108_CO6;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_D1 = CLBLM_L_X8Y116_SLICE_X11Y116_CO6;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_D2 = CLBLM_L_X10Y117_SLICE_X12Y117_DO6;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_D3 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_D4 = CLBLM_L_X10Y118_SLICE_X13Y118_AQ;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_D5 = CLBLM_L_X10Y116_SLICE_X12Y116_DO5;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_D6 = CLBLM_L_X10Y116_SLICE_X13Y116_BQ;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_B4 = CLBLM_R_X11Y110_SLICE_X15Y110_CQ;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_B6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y114_SLICE_X12Y114_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_C1 = CLBLM_L_X8Y108_SLICE_X11Y108_BQ;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_A1 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_A3 = CLBLM_L_X10Y118_SLICE_X13Y118_CO6;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_A4 = CLBLM_L_X10Y116_SLICE_X12Y116_DO5;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_A5 = CLBLM_R_X7Y105_SLICE_X8Y105_AQ;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_A6 = CLBLM_L_X10Y118_SLICE_X12Y118_CO6;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_C6 = CLBLM_R_X13Y112_SLICE_X18Y112_BQ;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_A1 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_A2 = CLBLM_R_X7Y114_SLICE_X8Y114_AQ;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_A4 = CLBLL_L_X4Y108_SLICE_X4Y108_CO6;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_B1 = CLBLM_L_X10Y118_SLICE_X12Y118_DO6;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_B2 = CLBLM_L_X10Y116_SLICE_X12Y116_DO5;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_B6 = CLBLM_R_X11Y113_SLICE_X14Y113_CQ;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_B3 = CLBLM_L_X10Y118_SLICE_X13Y118_CO6;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_B4 = CLBLM_L_X8Y118_SLICE_X10Y118_BQ;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_B5 = CLBLM_L_X10Y118_SLICE_X12Y118_BQ;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_C1 = CLBLM_R_X7Y113_SLICE_X9Y113_A5Q;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_D6 = CLBLM_L_X10Y113_SLICE_X13Y113_BQ;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_C1 = CLBLM_L_X10Y118_SLICE_X13Y118_AQ;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_C2 = CLBLM_L_X10Y118_SLICE_X12Y118_AQ;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_C3 = CLBLM_L_X8Y118_SLICE_X10Y118_CO5;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_C4 = CLBLM_L_X10Y117_SLICE_X12Y117_DO6;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_C5 = CLBLM_L_X8Y117_SLICE_X10Y117_AQ;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_C6 = CLBLM_R_X7Y118_SLICE_X9Y118_CO5;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_A1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_A2 = CLBLM_L_X8Y107_SLICE_X11Y107_CQ;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_A4 = CLBLM_L_X10Y112_SLICE_X12Y112_CQ;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_A6 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_D4 = CLBLL_L_X2Y114_SLICE_X0Y114_AO6;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_D1 = CLBLM_L_X8Y116_SLICE_X11Y116_CO6;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_D2 = CLBLM_L_X10Y118_SLICE_X12Y118_AQ;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_D3 = CLBLM_L_X10Y118_SLICE_X13Y118_AQ;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_D4 = CLBLM_L_X8Y118_SLICE_X10Y118_CO5;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_D5 = CLBLM_L_X8Y116_SLICE_X10Y116_BQ;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_B4 = CLBLM_L_X8Y106_SLICE_X10Y106_CQ;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_B6 = CLBLM_L_X8Y108_SLICE_X10Y108_AO5;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_D6 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_C1 = CLBLM_R_X5Y115_SLICE_X6Y115_AQ;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_C2 = 1'b1;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_C5 = CLBLM_L_X10Y108_SLICE_X12Y108_DO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_C3 = CLBLM_L_X8Y119_SLICE_X10Y119_AQ;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_C4 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_D1 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_D2 = CLBLM_L_X8Y108_SLICE_X10Y108_CQ;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_D3 = CLBLM_L_X8Y108_SLICE_X10Y108_DQ;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_D4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_D6 = CLBLL_L_X4Y110_SLICE_X4Y110_BQ;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_A1 = CLBLM_R_X11Y110_SLICE_X14Y110_CQ;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_A3 = CLBLL_L_X4Y114_SLICE_X5Y114_AQ;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_A4 = CLBLL_L_X4Y113_SLICE_X4Y113_CO6;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_A5 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_A6 = CLBLL_L_X4Y114_SLICE_X5Y114_CO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_A5 = CLBLM_L_X8Y113_SLICE_X11Y113_AQ;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_B1 = CLBLM_R_X3Y113_SLICE_X3Y113_AQ;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_B2 = CLBLM_R_X5Y115_SLICE_X7Y115_CO6;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_B3 = CLBLL_L_X4Y114_SLICE_X5Y114_AQ;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_B4 = CLBLM_R_X5Y111_SLICE_X6Y111_DO6;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_B5 = CLBLM_R_X11Y112_SLICE_X15Y112_CO6;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_B6 = CLBLM_R_X3Y114_SLICE_X2Y114_BQ;
  assign LIOI3_X0Y51_ILOGIC_X0Y52_D = LIOB33_X0Y51_IOB_X0Y52_I;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_C1 = CLBLM_R_X5Y111_SLICE_X6Y111_DO6;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_C2 = CLBLM_R_X3Y114_SLICE_X2Y114_BQ;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_C3 = CLBLM_R_X3Y113_SLICE_X3Y113_AQ;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_C4 = CLBLM_R_X5Y115_SLICE_X7Y115_CO6;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_C5 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_C6 = CLBLM_R_X11Y112_SLICE_X15Y112_CO6;
  assign LIOI3_X0Y51_ILOGIC_X0Y51_D = LIOB33_X0Y51_IOB_X0Y51_I;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOB33_X105Y151_IOB_X1Y151_O = LIOB33_X0Y75_IOB_X0Y76_I;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_A2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_A3 = CLBLM_R_X11Y112_SLICE_X15Y112_AQ;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_A4 = CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_D1 = CLBLL_L_X2Y112_SLICE_X0Y112_AO5;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_D2 = CLBLL_L_X2Y114_SLICE_X0Y114_AO6;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_D3 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_D4 = CLBLL_L_X2Y109_SLICE_X0Y109_AO5;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_D5 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_D6 = CLBLM_L_X10Y113_SLICE_X13Y113_DQ;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_B1 = CLBLM_R_X5Y112_SLICE_X7Y112_DQ;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_B2 = 1'b1;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_A6 = CLBLM_R_X7Y112_SLICE_X9Y112_CO6;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_B1 = 1'b1;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_B2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_B3 = 1'b1;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_B4 = CLBLM_L_X12Y113_SLICE_X17Y113_BQ;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_B6 = CLBLM_R_X13Y112_SLICE_X18Y112_CQ;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_C1 = CLBLM_R_X11Y112_SLICE_X15Y112_DO6;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_C2 = CLBLM_L_X10Y114_SLICE_X12Y114_CQ;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_C3 = CLBLM_R_X11Y111_SLICE_X15Y111_DO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_C4 = CLBLM_R_X13Y112_SLICE_X18Y112_A5Q;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_C5 = CLBLM_L_X12Y109_SLICE_X16Y109_DQ;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_C6 = CLBLM_R_X11Y114_SLICE_X15Y114_BO6;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y57_D = LIOB33_X0Y57_IOB_X0Y57_I;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_D1 = CLBLM_R_X11Y111_SLICE_X15Y111_C5Q;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_D2 = CLBLM_R_X13Y117_SLICE_X18Y117_AQ;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_D3 = CLBLM_R_X11Y113_SLICE_X15Y113_DQ;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_D4 = CLBLM_R_X11Y113_SLICE_X15Y113_CQ;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_D5 = CLBLM_R_X11Y114_SLICE_X15Y114_DO6;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_D6 = 1'b1;
  assign LIOB33_X0Y183_IOB_X0Y184_O = RIOB33_X105Y135_IOB_X1Y136_I;
  assign LIOB33_X0Y183_IOB_X0Y183_O = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_A2 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_A3 = CLBLM_L_X10Y111_SLICE_X12Y111_C5Q;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_A4 = CLBLM_R_X11Y112_SLICE_X14Y112_CQ;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_A5 = CLBLM_R_X11Y112_SLICE_X15Y112_AQ;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_A6 = 1'b1;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_B2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_B3 = CLBLM_L_X12Y111_SLICE_X16Y111_DQ;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_B4 = CLBLM_R_X5Y109_SLICE_X6Y109_DQ;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_B5 = CLBLM_L_X10Y107_SLICE_X13Y107_AQ;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_B6 = 1'b1;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_C1 = CLBLM_L_X10Y117_SLICE_X12Y117_AQ;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_C2 = CLBLM_R_X11Y113_SLICE_X15Y113_CQ;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_C5 = CLBLM_R_X11Y112_SLICE_X14Y112_B5Q;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_C6 = 1'b1;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_D1 = CLBLM_L_X8Y111_SLICE_X11Y111_CQ;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_D2 = 1'b1;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_D3 = CLBLM_L_X8Y114_SLICE_X10Y114_DQ;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_D4 = 1'b1;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_D5 = CLBLM_R_X11Y112_SLICE_X14Y112_B5Q;
  assign CLBLM_R_X11Y112_SLICE_X14Y112_D6 = CLBLM_R_X13Y110_SLICE_X18Y110_BQ;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_A1 = 1'b1;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_A2 = CLBLM_L_X10Y117_SLICE_X12Y117_BQ;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_A3 = CLBLM_L_X10Y119_SLICE_X12Y119_CO6;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_A4 = CLBLM_L_X10Y116_SLICE_X13Y116_CQ;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_A5 = 1'b1;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_A6 = 1'b1;
  assign RIOI3_X105Y171_OLOGIC_X1Y172_T1 = 1'b1;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_B1 = 1'b1;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_B2 = 1'b1;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_B3 = 1'b1;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_B4 = 1'b1;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_B5 = 1'b1;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_B6 = 1'b1;
  assign RIOI3_X105Y161_OLOGIC_X1Y162_T1 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_A1 = CLBLM_L_X8Y104_SLICE_X11Y104_AO5;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_A3 = CLBLM_L_X8Y109_SLICE_X11Y109_AQ;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_A4 = CLBLM_L_X8Y108_SLICE_X10Y108_BQ;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_C5 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_A5 = CLBLM_L_X8Y111_SLICE_X10Y111_CO6;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_A6 = CLBLM_L_X8Y108_SLICE_X11Y108_CO6;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_C1 = 1'b1;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_C2 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_AX = CLBLM_L_X8Y111_SLICE_X10Y111_BO6;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_C3 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_B1 = CLBLM_L_X8Y106_SLICE_X11Y106_A5Q;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_B2 = CLBLM_R_X13Y117_SLICE_X18Y117_AQ;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_B4 = CLBLM_R_X5Y109_SLICE_X6Y109_CQ;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_B6 = CLBLM_L_X8Y109_SLICE_X10Y109_CQ;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_D3 = 1'b1;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_D4 = 1'b1;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_D5 = 1'b1;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_D6 = 1'b1;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_D1 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_C5 = CLBLM_L_X12Y110_SLICE_X17Y110_AQ;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_C6 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_A2 = CLBLM_L_X10Y114_SLICE_X12Y114_AQ;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_A3 = CLBLM_L_X10Y119_SLICE_X12Y119_AQ;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_A4 = CLBLM_L_X8Y118_SLICE_X10Y118_DO6;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_A5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_A6 = CLBLM_L_X10Y117_SLICE_X13Y117_AO5;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_A5 = CLBLM_R_X3Y116_SLICE_X3Y116_AO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_A6 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_B6 = 1'b1;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_B1 = CLBLM_L_X10Y118_SLICE_X12Y118_AQ;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_B2 = CLBLM_L_X10Y116_SLICE_X13Y116_CQ;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_B3 = CLBLM_L_X10Y118_SLICE_X13Y118_AQ;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_C2 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_C3 = 1'b1;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_B4 = CLBLM_L_X10Y118_SLICE_X12Y118_BQ;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_B5 = CLBLM_R_X11Y116_SLICE_X14Y116_BQ;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_B6 = CLBLM_L_X8Y118_SLICE_X10Y118_CO5;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_C1 = 1'b1;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_C1 = CLBLM_R_X11Y116_SLICE_X14Y116_BQ;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_C2 = CLBLM_L_X8Y118_SLICE_X10Y118_CO5;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_C3 = 1'b1;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_C4 = CLBLM_L_X10Y118_SLICE_X12Y118_AQ;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_C5 = CLBLM_L_X10Y118_SLICE_X13Y118_AQ;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_C6 = CLBLM_L_X10Y118_SLICE_X12Y118_BQ;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_A1 = CLBLM_L_X10Y108_SLICE_X12Y108_CQ;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_A2 = CLBLM_R_X11Y111_SLICE_X15Y111_C5Q;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_A3 = CLBLM_L_X8Y109_SLICE_X10Y109_AQ;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_D1 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_B5 = CLBLM_L_X8Y109_SLICE_X10Y109_C5Q;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_B6 = 1'b1;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_D1 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_D3 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_D4 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_D5 = 1'b1;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_D5 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_C2 = CLBLM_L_X8Y109_SLICE_X11Y109_A5Q;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_C3 = CLBLM_R_X7Y109_SLICE_X9Y109_AQ;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_C4 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_C5 = CLBLM_R_X5Y109_SLICE_X6Y109_CQ;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_C6 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_D6 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_D2 = CLBLM_R_X5Y106_SLICE_X6Y106_DQ;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_D3 = CLBLM_L_X8Y109_SLICE_X10Y109_DQ;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_D4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_D5 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_A1 = CLBLM_R_X3Y110_SLICE_X2Y110_DO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_A2 = CLBLM_R_X3Y109_SLICE_X2Y109_CO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_A3 = CLBLM_L_X8Y117_SLICE_X10Y117_AQ;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_A5 = CLBLM_R_X7Y117_SLICE_X9Y117_AQ;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_A6 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_D6 = CLBLM_R_X7Y109_SLICE_X8Y109_DO6;
  assign RIOB33_X105Y153_IOB_X1Y153_O = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_B1 = CLBLL_L_X4Y113_SLICE_X5Y113_DO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_B2 = CLBLL_L_X4Y115_SLICE_X5Y115_BQ;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_B3 = CLBLL_L_X4Y116_SLICE_X4Y116_A5Q;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_B5 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_B6 = CLBLL_L_X4Y115_SLICE_X5Y115_A5Q;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_C1 = CLBLL_L_X4Y116_SLICE_X5Y116_AQ;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_C2 = CLBLL_L_X4Y115_SLICE_X5Y115_CQ;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_C3 = CLBLL_L_X4Y113_SLICE_X5Y113_DO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_C4 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_C6 = CLBLM_R_X5Y110_SLICE_X6Y110_BQ;
  assign RIOI3_X105Y161_OLOGIC_X1Y161_T1 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_D1 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_D2 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_D3 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_D4 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_D5 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_D6 = 1'b1;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_A2 = CLBLM_R_X11Y113_SLICE_X15Y113_BQ;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_A3 = CLBLM_R_X11Y113_SLICE_X15Y113_AQ;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_B2 = CLBLM_R_X11Y113_SLICE_X15Y113_BQ;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_B3 = CLBLM_R_X7Y113_SLICE_X8Y113_CQ;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_B4 = 1'b1;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_B5 = CLBLM_R_X5Y115_SLICE_X7Y115_CO6;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_B6 = CLBLM_L_X10Y114_SLICE_X12Y114_DQ;
  assign LIOB33_X0Y185_IOB_X0Y185_O = RIOB33_X105Y137_IOB_X1Y137_I;
  assign LIOB33_X0Y185_IOB_X0Y186_O = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_C1 = CLBLM_R_X7Y115_SLICE_X9Y115_AQ;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_C2 = CLBLM_R_X11Y113_SLICE_X15Y113_CQ;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_C4 = CLBLM_R_X7Y115_SLICE_X9Y115_DO6;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_C5 = CLBLM_R_X11Y114_SLICE_X15Y114_BO6;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_C6 = 1'b1;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_D2 = CLBLM_R_X11Y113_SLICE_X15Y113_CQ;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_D3 = CLBLM_R_X11Y113_SLICE_X15Y113_DQ;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_D4 = CLBLM_R_X7Y115_SLICE_X9Y115_DO6;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_D5 = CLBLM_R_X11Y107_SLICE_X15Y107_AQ;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_D6 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_D4 = 1'b1;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_A2 = CLBLM_R_X11Y113_SLICE_X14Y113_BQ;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_A3 = CLBLM_R_X11Y113_SLICE_X14Y113_AQ;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_A4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_A5 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_A6 = CLBLM_R_X11Y107_SLICE_X15Y107_AQ;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_B1 = CLBLM_L_X12Y113_SLICE_X17Y113_CQ;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_B2 = CLBLM_R_X11Y113_SLICE_X14Y113_BQ;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_B3 = CLBLM_R_X11Y113_SLICE_X14Y113_DQ;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_B4 = CLBLM_R_X11Y113_SLICE_X14Y113_CQ;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_C1 = CLBLM_L_X10Y112_SLICE_X13Y112_AO6;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_C2 = CLBLM_L_X10Y113_SLICE_X13Y113_BQ;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_C3 = CLBLM_R_X11Y113_SLICE_X14Y113_BQ;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_C6 = CLBLM_R_X13Y112_SLICE_X18Y112_BQ;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_T1 = 1'b1;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_D1 = CLBLM_L_X10Y112_SLICE_X13Y112_AO6;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_D2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_D3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_D4 = CLBLM_R_X13Y112_SLICE_X18Y112_BQ;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_D5 = CLBLM_R_X11Y118_SLICE_X15Y118_A5Q;
  assign CLBLM_R_X11Y113_SLICE_X14Y113_D6 = 1'b1;
  assign RIOB33_X105Y187_IOB_X1Y188_O = CLBLM_L_X12Y117_SLICE_X17Y117_AQ;
  assign RIOB33_X105Y187_IOB_X1Y187_O = CLBLM_R_X11Y115_SLICE_X14Y115_BQ;
  assign LIOI3_X0Y175_OLOGIC_X0Y176_D1 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_D4 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_A1 = CLBLL_L_X4Y116_SLICE_X4Y116_BO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_A3 = CLBLM_L_X8Y110_SLICE_X11Y110_AQ;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_A4 = CLBLM_L_X8Y106_SLICE_X11Y106_BQ;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_A5 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_A6 = CLBLM_L_X8Y115_SLICE_X10Y115_CQ;
  assign LIOI3_X0Y115_OLOGIC_X0Y116_D1 = CLBLM_R_X11Y118_SLICE_X15Y118_AQ;
  assign LIOI3_X0Y175_OLOGIC_X0Y176_T1 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_AX = CLBLM_L_X8Y110_SLICE_X11Y110_BO6;
  assign LIOI3_SING_X0Y199_OLOGIC_X0Y199_D1 = LIOB33_X0Y73_IOB_X0Y74_I;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_B1 = CLBLM_L_X12Y113_SLICE_X17Y113_BQ;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_B2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_B3 = CLBLM_L_X8Y107_SLICE_X11Y107_CQ;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_B5 = CLBLM_L_X8Y110_SLICE_X11Y110_A5Q;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_B6 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_A1 = CLBLM_R_X5Y116_SLICE_X6Y116_DQ;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_A3 = CLBLL_L_X4Y116_SLICE_X4Y116_AQ;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_C1 = CLBLM_L_X8Y112_SLICE_X11Y112_AO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_C2 = CLBLM_L_X8Y110_SLICE_X11Y110_CQ;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_A5 = CLBLL_L_X4Y117_SLICE_X5Y117_BO5;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_A6 = CLBLL_L_X4Y113_SLICE_X5Y113_B5Q;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_C2 = CLBLM_L_X8Y106_SLICE_X10Y106_CQ;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_C3 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_AX = CLBLL_L_X4Y117_SLICE_X5Y117_BO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_C3 = CLBLM_R_X5Y107_SLICE_X7Y107_B5Q;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_C5 = CLBLM_L_X8Y110_SLICE_X10Y110_AQ;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_B1 = CLBLM_R_X5Y116_SLICE_X6Y116_DQ;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_B2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_C4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_B3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_B4 = CLBLM_R_X11Y113_SLICE_X14Y113_CQ;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_B5 = CLBLM_L_X12Y112_SLICE_X16Y112_AQ;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_B6 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_C5 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_D1 = CLBLM_R_X11Y113_SLICE_X14Y113_AQ;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_C1 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_C2 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_C3 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_C4 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_C5 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_C6 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_A1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_D1 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_D2 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_D3 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_D4 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_D5 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X4Y116_D6 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_A3 = CLBLM_L_X8Y110_SLICE_X10Y110_AQ;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_A4 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_A6 = CLBLM_R_X7Y110_SLICE_X9Y110_DO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_B1 = CLBLM_L_X12Y111_SLICE_X16Y111_BQ;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_B2 = CLBLM_L_X8Y110_SLICE_X10Y110_BQ;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_B3 = CLBLM_R_X7Y108_SLICE_X9Y108_BO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_B4 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_B5 = CLBLM_L_X10Y113_SLICE_X13Y113_AQ;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_C1 = CLBLM_R_X7Y110_SLICE_X9Y110_BQ;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_C2 = CLBLM_R_X7Y105_SLICE_X9Y105_AQ;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_C3 = CLBLM_L_X8Y110_SLICE_X10Y110_AQ;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_C4 = CLBLM_R_X7Y105_SLICE_X8Y105_A5Q;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_C5 = CLBLM_L_X10Y113_SLICE_X13Y113_CQ;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_C6 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_T1 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_A1 = CLBLM_R_X5Y116_SLICE_X6Y116_DQ;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_A2 = CLBLM_L_X8Y114_SLICE_X10Y114_BQ;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_D3 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_A3 = CLBLL_L_X4Y116_SLICE_X5Y116_AQ;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_D4 = CLBLM_R_X7Y116_SLICE_X8Y116_CQ;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_D5 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_D6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_A6 = CLBLL_L_X4Y118_SLICE_X4Y118_A5Q;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_D2 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_AX = CLBLM_R_X5Y116_SLICE_X6Y116_AO6;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_B2 = CLBLL_L_X4Y116_SLICE_X5Y116_BQ;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_B3 = RIOB33_X105Y127_IOB_X1Y127_I;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_B4 = CLBLM_R_X7Y117_SLICE_X9Y117_BQ;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_B5 = CLBLL_L_X4Y111_SLICE_X5Y111_AQ;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_B6 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_C1 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_C2 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_C3 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_C4 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_C5 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_C6 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_B3 = 1'b1;
  assign LIOB33_X0Y187_IOB_X0Y187_O = RIOB33_X105Y143_IOB_X1Y144_I;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOB33_X0Y187_IOB_X0Y188_O = RIOB33_X105Y145_IOB_X1Y145_I;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_B5 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_D1 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_D2 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_D3 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_D4 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_D5 = 1'b1;
  assign CLBLL_L_X4Y116_SLICE_X5Y116_D6 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_A1 = CLBLM_R_X11Y114_SLICE_X14Y114_DQ;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_A2 = CLBLM_L_X10Y114_SLICE_X13Y114_CQ;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_A3 = CLBLM_R_X11Y110_SLICE_X15Y110_CQ;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_A4 = CLBLM_L_X12Y113_SLICE_X16Y113_BQ;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_A5 = CLBLM_L_X8Y114_SLICE_X10Y114_BQ;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_A6 = CLBLM_L_X10Y109_SLICE_X12Y109_AQ;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_B1 = CLBLM_L_X12Y109_SLICE_X16Y109_DQ;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_B2 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_B3 = CLBLM_R_X5Y111_SLICE_X6Y111_DO6;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_B4 = CLBLM_R_X11Y115_SLICE_X15Y115_CQ;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_B5 = CLBLM_L_X12Y114_SLICE_X16Y114_BQ;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_B6 = CLBLM_R_X11Y114_SLICE_X15Y114_CO6;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_C1 = CLBLM_R_X11Y114_SLICE_X15Y114_AO6;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_C2 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_C3 = CLBLM_L_X10Y114_SLICE_X12Y114_CQ;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_C4 = CLBLM_L_X10Y114_SLICE_X12Y114_DQ;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_C5 = CLBLM_R_X11Y115_SLICE_X15Y115_DO6;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_C6 = CLBLM_L_X12Y114_SLICE_X16Y114_AQ;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_D1 = CLBLM_L_X12Y113_SLICE_X16Y113_BQ;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_D2 = CLBLM_L_X8Y112_SLICE_X10Y112_AQ;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_D3 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_D4 = CLBLM_L_X8Y114_SLICE_X10Y114_BQ;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_D5 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X15Y114_D6 = CLBLM_R_X11Y111_SLICE_X15Y111_CQ;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_A1 = CLBLM_L_X12Y114_SLICE_X16Y114_CQ;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_A3 = CLBLM_R_X11Y114_SLICE_X14Y114_AQ;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_A4 = CLBLL_L_X4Y116_SLICE_X4Y116_BO6;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_A5 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_A6 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_B1 = CLBLM_L_X8Y119_SLICE_X10Y119_AQ;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_B3 = CLBLM_R_X11Y111_SLICE_X14Y111_AO6;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_B4 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_B5 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_B6 = CLBLM_R_X7Y115_SLICE_X9Y115_BQ;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_C1 = CLBLM_R_X11Y112_SLICE_X15Y112_BQ;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_C2 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_C3 = CLBLM_R_X11Y115_SLICE_X14Y115_BO5;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_C5 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_C6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_D1 = CLBLM_R_X11Y110_SLICE_X15Y110_CQ;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_D2 = 1'b1;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_D3 = CLBLM_R_X11Y114_SLICE_X14Y114_DQ;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_D4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_D5 = CLBLM_L_X10Y115_SLICE_X12Y115_BQ;
  assign CLBLM_R_X11Y114_SLICE_X14Y114_D6 = CLBLM_R_X5Y115_SLICE_X7Y115_CO6;
  assign LIOI3_X0Y53_ILOGIC_X0Y54_D = LIOB33_X0Y53_IOB_X0Y54_I;
  assign LIOI3_X0Y53_ILOGIC_X0Y53_D = LIOB33_X0Y53_IOB_X0Y53_I;
  assign LIOI3_X0Y171_OLOGIC_X0Y172_D1 = CLBLM_R_X103Y138_SLICE_X163Y138_AO6;
  assign LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y70_D = LIOB33_X0Y69_IOB_X0Y70_I;
  assign LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y69_D = LIOB33_X0Y69_IOB_X0Y69_I;
  assign RIOB33_SING_X105Y199_IOB_X1Y199_O = CLBLM_R_X11Y119_SLICE_X14Y119_AQ;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_A1 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_A2 = CLBLM_R_X7Y111_SLICE_X8Y111_CQ;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_A3 = CLBLM_L_X8Y111_SLICE_X11Y111_AQ;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_A4 = CLBLL_L_X4Y116_SLICE_X4Y116_BO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_A5 = CLBLM_L_X12Y110_SLICE_X17Y110_CQ;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_B1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_A1 = CLBLL_L_X4Y116_SLICE_X4Y116_BO5;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_B3 = CLBLM_R_X11Y106_SLICE_X15Y106_AQ;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_A2 = CLBLL_L_X4Y117_SLICE_X4Y117_DQ;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_B4 = CLBLM_L_X8Y112_SLICE_X11Y112_DO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_B5 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_A3 = CLBLL_L_X4Y117_SLICE_X4Y117_AQ;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_A4 = CLBLL_L_X4Y118_SLICE_X4Y118_DO5;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_A5 = CLBLM_R_X5Y111_SLICE_X7Y111_BQ;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_C2 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_C4 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_B1 = CLBLL_L_X4Y116_SLICE_X4Y116_BO5;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_C5 = CLBLM_R_X13Y112_SLICE_X18Y112_BQ;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_B2 = CLBLL_L_X4Y117_SLICE_X4Y117_BQ;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_B3 = CLBLL_L_X4Y116_SLICE_X4Y116_AQ;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_B4 = CLBLM_R_X5Y110_SLICE_X6Y110_BQ;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_B6 = CLBLL_L_X4Y117_SLICE_X5Y117_BO5;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_C2 = CLBLL_L_X4Y116_SLICE_X4Y116_AQ;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_C3 = CLBLL_L_X4Y117_SLICE_X5Y117_BO5;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_C4 = CLBLM_R_X7Y106_SLICE_X9Y106_AQ;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_C5 = CLBLL_L_X4Y117_SLICE_X4Y117_BQ;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_C6 = CLBLM_R_X5Y116_SLICE_X6Y116_DQ;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_D6 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_D3 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_D4 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_D2 = CLBLM_R_X7Y116_SLICE_X8Y116_BQ;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_D3 = CLBLL_L_X4Y117_SLICE_X4Y117_DQ;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_D4 = CLBLM_R_X5Y116_SLICE_X6Y116_DQ;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_D5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_D6 = CLBLL_L_X4Y118_SLICE_X4Y118_DO5;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_A1 = CLBLM_L_X12Y110_SLICE_X17Y110_CQ;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_A3 = CLBLM_L_X8Y111_SLICE_X10Y111_AQ;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_A5 = CLBLM_R_X3Y111_SLICE_X2Y111_CO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_A6 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_B1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_B3 = CLBLM_L_X8Y106_SLICE_X10Y106_AQ;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_B4 = CLBLM_R_X7Y111_SLICE_X9Y111_AQ;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_B5 = CLBLM_R_X5Y109_SLICE_X6Y109_DQ;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_B6 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_C1 = CLBLM_L_X8Y112_SLICE_X10Y112_DO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_C2 = CLBLM_L_X8Y111_SLICE_X10Y111_AQ;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_C3 = CLBLM_L_X8Y111_SLICE_X11Y111_DO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_C4 = CLBLM_L_X12Y106_SLICE_X17Y106_AQ;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_C5 = CLBLM_L_X8Y112_SLICE_X11Y112_AO5;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_C6 = CLBLM_R_X7Y105_SLICE_X8Y105_CQ;
  assign LIOB33_X0Y189_IOB_X0Y190_O = RIOB33_X105Y147_IOB_X1Y147_I;
  assign LIOB33_X0Y189_IOB_X0Y189_O = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_A1 = CLBLL_L_X4Y118_SLICE_X4Y118_DO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_A3 = CLBLL_L_X4Y117_SLICE_X5Y117_AQ;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_A5 = CLBLM_R_X5Y116_SLICE_X6Y116_DQ;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_A6 = CLBLM_L_X8Y115_SLICE_X10Y115_A5Q;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_D3 = CLBLM_L_X10Y112_SLICE_X12Y112_BQ;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_D4 = CLBLM_R_X11Y111_SLICE_X15Y111_BQ;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_D1 = CLBLM_L_X8Y111_SLICE_X11Y111_DO5;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_D5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_D2 = CLBLM_L_X8Y114_SLICE_X10Y114_CQ;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_B1 = CLBLL_L_X4Y118_SLICE_X4Y118_DO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_B3 = CLBLL_L_X4Y117_SLICE_X5Y117_AQ;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_B4 = CLBLL_L_X4Y118_SLICE_X4Y118_BQ;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_B5 = CLBLM_R_X5Y116_SLICE_X7Y116_BQ;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_B6 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_C1 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_C2 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_C3 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_C4 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_C5 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_C6 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_B3 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_B4 = CLBLM_R_X5Y109_SLICE_X7Y109_A5Q;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_D1 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_D2 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_D3 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_D4 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_D5 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_D6 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_B6 = CLBLL_L_X4Y112_SLICE_X4Y112_CO6;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_A1 = CLBLM_R_X11Y115_SLICE_X14Y115_AO5;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_A2 = CLBLM_L_X12Y110_SLICE_X17Y110_CQ;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_A3 = 1'b1;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_A6 = CLBLM_R_X11Y113_SLICE_X14Y113_CQ;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_B1 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_B2 = CLBLM_L_X12Y112_SLICE_X17Y112_A5Q;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_B3 = CLBLM_L_X10Y113_SLICE_X13Y113_AQ;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_B4 = CLBLM_L_X10Y115_SLICE_X13Y115_AQ;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_B6 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_A1 = CLBLM_R_X7Y105_SLICE_X9Y105_DO6;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_A3 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_A4 = CLBLM_R_X5Y113_SLICE_X6Y113_BQ;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_A5 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_A6 = 1'b1;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_C1 = CLBLM_R_X11Y113_SLICE_X15Y113_BQ;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_C2 = CLBLM_R_X11Y115_SLICE_X15Y115_CQ;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_C3 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_B1 = CLBLM_R_X5Y107_SLICE_X6Y107_AQ;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_B2 = CLBLM_R_X7Y105_SLICE_X9Y105_BQ;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_B4 = CLBLM_L_X8Y105_SLICE_X11Y105_AQ;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_B6 = CLBLM_L_X10Y106_SLICE_X12Y106_BO6;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_D1 = CLBLM_R_X11Y113_SLICE_X15Y113_BQ;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_C2 = CLBLM_R_X7Y105_SLICE_X9Y105_CQ;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_C3 = CLBLM_R_X7Y107_SLICE_X8Y107_DO6;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_C4 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_C5 = CLBLM_L_X10Y113_SLICE_X13Y113_AQ;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_C6 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_C6 = CLBLM_L_X8Y105_SLICE_X11Y105_AQ;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_D4 = CLBLM_L_X10Y114_SLICE_X12Y114_AQ;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_A2 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_A3 = CLBLM_L_X10Y111_SLICE_X13Y111_C5Q;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_A4 = CLBLM_R_X11Y116_SLICE_X15Y116_AQ;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_A5 = CLBLM_L_X10Y110_SLICE_X12Y110_AQ;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_D1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_D2 = CLBLM_R_X7Y116_SLICE_X8Y116_CQ;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_D3 = CLBLM_L_X10Y104_SLICE_X12Y104_AQ;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_A2 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_D4 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_D5 = CLBLM_R_X7Y105_SLICE_X9Y105_AQ;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_D6 = CLBLM_R_X3Y110_SLICE_X3Y110_AO6;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_A3 = 1'b1;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_AX = CLBLM_R_X11Y115_SLICE_X15Y115_CQ;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_B1 = CLBLM_R_X7Y115_SLICE_X8Y115_CQ;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_B2 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_A4 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_A1 = CLBLM_R_X7Y115_SLICE_X8Y115_DQ;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_A2 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_A3 = CLBLM_R_X7Y105_SLICE_X8Y105_AQ;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_A4 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_A5 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_A6 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_BX = CLBLM_R_X11Y110_SLICE_X14Y110_DQ;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_AX = CLBLM_R_X7Y105_SLICE_X8Y105_BO6;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_C1 = CLBLM_L_X10Y118_SLICE_X12Y118_AQ;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_B1 = CLBLM_R_X7Y105_SLICE_X8Y105_DO6;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_B2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_B3 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_B5 = CLBLM_L_X8Y104_SLICE_X11Y104_AQ;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_B6 = 1'b1;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_CE = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_D1 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_C2 = CLBLM_R_X7Y105_SLICE_X8Y105_CQ;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_C3 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_C4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_C5 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_C6 = CLBLM_R_X7Y105_SLICE_X9Y105_BQ;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_D3 = 1'b1;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_D4 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_D6 = 1'b1;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_SR = CLBLM_L_X12Y117_SLICE_X16Y117_AO6;
  assign RIOI3_X105Y185_OLOGIC_X1Y186_D1 = CLBLM_L_X12Y111_SLICE_X16Y111_AQ;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_B1 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_D1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_D2 = CLBLM_R_X7Y116_SLICE_X8Y116_CQ;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_D3 = CLBLM_L_X10Y104_SLICE_X12Y104_AQ;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_B2 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_D4 = CLBLM_R_X7Y105_SLICE_X8Y105_A5Q;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_D5 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_D6 = CLBLM_R_X3Y110_SLICE_X2Y110_DO6;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_B3 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_B4 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_B5 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_C1 = 1'b1;
  assign RIOI3_X105Y185_OLOGIC_X1Y186_T1 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_C2 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_C3 = 1'b1;
  assign LIOI3_X0Y151_OLOGIC_X0Y152_T1 = 1'b1;
  assign RIOB33_X105Y159_IOB_X1Y160_O = CLBLM_R_X13Y110_SLICE_X18Y110_DO5;
  assign RIOB33_X105Y159_IOB_X1Y159_O = CLBLM_R_X13Y110_SLICE_X18Y110_DO6;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_A1 = CLBLM_L_X8Y114_SLICE_X10Y114_CQ;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_A2 = CLBLM_L_X8Y114_SLICE_X11Y114_BQ;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_A3 = CLBLM_R_X7Y111_SLICE_X8Y111_CQ;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_A4 = CLBLM_L_X10Y112_SLICE_X12Y112_BQ;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_A5 = CLBLM_R_X7Y117_SLICE_X9Y117_DQ;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_A6 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_A1 = CLBLL_L_X4Y114_SLICE_X4Y114_CQ;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_A2 = CLBLL_L_X4Y118_SLICE_X4Y118_AQ;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_A3 = CLBLL_L_X4Y116_SLICE_X5Y116_AQ;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_A5 = CLBLL_L_X4Y118_SLICE_X4Y118_CO5;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_A6 = CLBLL_L_X4Y118_SLICE_X4Y118_A5Q;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_B1 = CLBLM_R_X7Y112_SLICE_X8Y112_BQ;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_AX = CLBLL_L_X4Y118_SLICE_X4Y118_CO6;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_B5 = CLBLM_L_X10Y111_SLICE_X12Y111_BQ;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_B2 = CLBLL_L_X4Y118_SLICE_X4Y118_BQ;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_B4 = CLBLM_R_X3Y118_SLICE_X3Y118_AO6;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_B5 = CLBLM_L_X10Y117_SLICE_X12Y117_BQ;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_B6 = CLBLM_R_X5Y116_SLICE_X6Y116_DQ;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_C3 = CLBLM_L_X10Y116_SLICE_X13Y116_DO6;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_B6 = CLBLM_L_X8Y109_SLICE_X10Y109_BQ;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_C5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_C2 = CLBLM_R_X5Y116_SLICE_X6Y116_DQ;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_C4 = CLBLL_L_X4Y118_SLICE_X4Y118_A5Q;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_C5 = CLBLM_R_X7Y118_SLICE_X9Y118_AQ;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_C6 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_D1 = CLBLM_R_X7Y117_SLICE_X9Y117_DQ;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_D2 = CLBLM_R_X7Y111_SLICE_X8Y111_CQ;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_D3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_D4 = CLBLM_L_X8Y112_SLICE_X11Y112_AO5;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_D5 = CLBLM_L_X10Y112_SLICE_X12Y112_CQ;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_D1 = CLBLL_L_X4Y116_SLICE_X5Y116_AQ;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_D2 = CLBLL_L_X4Y118_SLICE_X4Y118_AQ;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_D3 = CLBLL_L_X4Y117_SLICE_X4Y117_DQ;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_D4 = CLBLL_L_X4Y118_SLICE_X4Y118_A5Q;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_D5 = CLBLL_L_X4Y117_SLICE_X4Y117_AQ;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_D6 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_D6 = CLBLM_L_X8Y115_SLICE_X10Y115_BQ;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_A1 = CLBLM_L_X8Y115_SLICE_X10Y115_A5Q;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_A3 = CLBLM_R_X7Y112_SLICE_X9Y112_BQ;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_A5 = CLBLM_L_X8Y105_SLICE_X10Y105_AQ;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_A6 = 1'b1;
  assign LIOB33_X0Y191_IOB_X0Y191_O = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_B1 = CLBLM_R_X11Y112_SLICE_X14Y112_CQ;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_B2 = CLBLM_R_X7Y113_SLICE_X8Y113_DQ;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_B3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_B4 = CLBLM_L_X10Y112_SLICE_X12Y112_BQ;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_B5 = CLBLM_L_X8Y111_SLICE_X11Y111_DO5;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_B6 = CLBLM_L_X8Y114_SLICE_X10Y114_CQ;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_C1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_C2 = CLBLM_L_X8Y114_SLICE_X10Y114_CQ;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_C3 = CLBLM_L_X8Y111_SLICE_X11Y111_DO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_C4 = CLBLM_L_X10Y112_SLICE_X12Y112_BQ;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_C5 = CLBLM_R_X7Y115_SLICE_X8Y115_CQ;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_C6 = CLBLM_R_X7Y115_SLICE_X8Y115_BQ;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_A1 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_A2 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_A3 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_A4 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_A5 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_A6 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_B1 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_B2 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_B3 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_B4 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_B5 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_B6 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_D1 = CLBLM_L_X12Y106_SLICE_X17Y106_AQ;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_D2 = CLBLM_L_X10Y110_SLICE_X12Y110_DO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_D3 = CLBLM_R_X7Y113_SLICE_X8Y113_DQ;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_C1 = 1'b1;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_D3 = CLBLM_R_X11Y115_SLICE_X15Y115_AQ;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_C2 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_C3 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_C4 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_C5 = 1'b1;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_D4 = CLBLM_L_X12Y110_SLICE_X17Y110_CQ;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_C6 = 1'b1;
  assign LIOI3_X0Y177_OLOGIC_X0Y178_D1 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_D5 = CLBLM_R_X11Y113_SLICE_X14Y113_CQ;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_D1 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_D2 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_D3 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_D4 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_D5 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_D6 = 1'b1;
  assign CLBLM_L_X10Y115_SLICE_X13Y115_D6 = 1'b1;
  assign LIOI3_X0Y177_OLOGIC_X0Y178_T1 = 1'b1;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_D1 = CLBLM_R_X5Y114_SLICE_X7Y114_CQ;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_A2 = CLBLM_L_X12Y114_SLICE_X17Y114_AQ;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_A3 = CLBLM_R_X11Y116_SLICE_X15Y116_AQ;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_A4 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_A5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_A6 = CLBLM_L_X10Y111_SLICE_X13Y111_DO6;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_T1 = 1'b1;
  assign LIOI3_X0Y177_OLOGIC_X0Y177_D1 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_B1 = 1'b1;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_B2 = 1'b1;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_B3 = 1'b1;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_B4 = 1'b1;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_B5 = 1'b1;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_B6 = 1'b1;
  assign LIOI3_X0Y177_OLOGIC_X0Y177_T1 = 1'b1;
  assign RIOI3_X105Y161_OLOGIC_X1Y162_D1 = CLBLM_L_X12Y114_SLICE_X16Y114_DO5;
  assign LIOI3_X0Y117_OLOGIC_X0Y117_D1 = CLBLL_L_X4Y116_SLICE_X5Y116_BQ;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_A1 = CLBLM_L_X10Y113_SLICE_X13Y113_AQ;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_A2 = CLBLM_L_X12Y109_SLICE_X16Y109_D5Q;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_A3 = CLBLM_R_X7Y106_SLICE_X9Y106_AQ;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_A4 = CLBLM_R_X7Y105_SLICE_X9Y105_AO5;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_A5 = CLBLM_R_X7Y109_SLICE_X9Y109_CQ;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_C1 = 1'b1;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_C2 = 1'b1;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_C3 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_B1 = CLBLM_R_X11Y107_SLICE_X15Y107_BQ;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_B2 = CLBLM_R_X7Y106_SLICE_X9Y106_BQ;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_B3 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_B4 = CLBLL_L_X4Y113_SLICE_X4Y113_BQ;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_B6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_D1 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_C2 = CLBLM_R_X7Y106_SLICE_X9Y106_CQ;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_C3 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_C4 = CLBLM_R_X7Y105_SLICE_X9Y105_CQ;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_C5 = CLBLM_L_X8Y104_SLICE_X10Y104_AO6;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_C6 = CLBLM_R_X7Y112_SLICE_X8Y112_BQ;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_D3 = 1'b1;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_D4 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_A1 = CLBLM_L_X10Y117_SLICE_X13Y117_AO5;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_A3 = CLBLM_R_X11Y116_SLICE_X14Y116_AQ;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_A6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_A4 = CLBLM_L_X12Y114_SLICE_X16Y114_BQ;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_D2 = CLBLM_L_X10Y111_SLICE_X12Y111_CQ;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_D3 = CLBLM_R_X7Y111_SLICE_X8Y111_BQ;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_D4 = CLBLL_L_X4Y107_SLICE_X4Y107_CQ;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_D5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_D6 = 1'b1;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_A5 = CLBLM_L_X8Y116_SLICE_X10Y116_BQ;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_A6 = CLBLM_R_X7Y118_SLICE_X8Y118_DO6;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_AX = CLBLM_R_X11Y117_SLICE_X15Y117_BO6;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_B1 = CLBLM_L_X10Y118_SLICE_X13Y118_CO6;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_B2 = CLBLM_R_X7Y108_SLICE_X9Y108_AQ;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_A1 = CLBLM_L_X12Y107_SLICE_X16Y107_DQ;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_A2 = CLBLM_R_X7Y105_SLICE_X8Y105_CQ;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_A3 = CLBLM_R_X7Y106_SLICE_X8Y106_AQ;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_A5 = CLBLL_L_X4Y110_SLICE_X4Y110_AQ;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_A6 = CLBLM_R_X5Y106_SLICE_X6Y106_CQ;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_C1 = CLBLM_L_X10Y116_SLICE_X12Y116_DO5;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_C2 = CLBLM_L_X10Y117_SLICE_X12Y117_DO6;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_B1 = CLBLM_L_X8Y109_SLICE_X10Y109_CQ;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_B2 = CLBLM_R_X7Y106_SLICE_X8Y106_BQ;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_B1 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_B4 = CLBLM_R_X5Y105_SLICE_X7Y105_BQ;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_B5 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_B6 = CLBLM_L_X8Y104_SLICE_X10Y104_AO6;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_B2 = CLBLM_L_X8Y114_SLICE_X11Y114_CQ;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_D3 = CLBLM_L_X10Y118_SLICE_X13Y118_AQ;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_C2 = CLBLM_R_X7Y106_SLICE_X8Y106_CQ;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_C3 = CLBLM_L_X8Y104_SLICE_X10Y104_AO6;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_C4 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_C5 = CLBLM_R_X7Y109_SLICE_X9Y109_CQ;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_C6 = CLBLM_R_X7Y109_SLICE_X8Y109_AQ;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_B4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_D4 = CLBLM_L_X8Y118_SLICE_X10Y118_AQ;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_D6 = CLBLM_L_X10Y119_SLICE_X12Y119_AQ;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_B5 = CLBLM_R_X11Y112_SLICE_X14Y112_AO5;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE0 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE1 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_D1 = 1'b1;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_B6 = CLBLM_L_X8Y116_SLICE_X11Y116_AQ;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_D2 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_D3 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_D4 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_D5 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_D6 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE0 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE1 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S0 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S1 = 1'b1;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_C2 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_C3 = 1'b1;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign RIOB33_X105Y161_IOB_X1Y162_O = CLBLM_L_X12Y114_SLICE_X16Y114_DO5;
  assign RIOB33_X105Y161_IOB_X1Y161_O = CLBLM_L_X12Y114_SLICE_X16Y114_DO6;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_C5 = 1'b1;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_C6 = CLBLM_L_X10Y114_SLICE_X12Y114_BQ;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_C5 = CLBLM_R_X7Y117_SLICE_X9Y117_AQ;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_A1 = CLBLM_L_X8Y113_SLICE_X11Y113_DO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_A2 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_A4 = CLBLM_L_X8Y114_SLICE_X10Y114_DQ;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_A6 = CLBLM_L_X8Y108_SLICE_X11Y108_CO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_B2 = CLBLM_L_X8Y113_SLICE_X11Y113_BQ;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_B3 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_B4 = CLBLM_L_X8Y113_SLICE_X10Y113_BQ;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_B5 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_B6 = CLBLM_L_X8Y113_SLICE_X11Y113_CO6;
  assign LIOB33_X0Y193_IOB_X0Y193_O = LIOB33_X0Y55_IOB_X0Y56_I;
  assign LIOB33_X0Y193_IOB_X0Y194_O = LIOB33_X0Y59_IOB_X0Y60_I;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_C1 = CLBLM_R_X13Y112_SLICE_X18Y112_CQ;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_C2 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_C3 = CLBLM_L_X12Y113_SLICE_X17Y113_B5Q;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_C4 = CLBLM_L_X8Y114_SLICE_X10Y114_CQ;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_C5 = CLBLM_L_X8Y111_SLICE_X11Y111_DO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_C6 = CLBLM_L_X10Y112_SLICE_X12Y112_BQ;
  assign LIOI3_X0Y55_ILOGIC_X0Y56_D = LIOB33_X0Y55_IOB_X0Y56_I;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_D1 = 1'b1;
  assign LIOI3_X0Y55_ILOGIC_X0Y55_D = LIOB33_X0Y55_IOB_X0Y55_I;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_D2 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_D1 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_D2 = CLBLM_L_X12Y108_SLICE_X16Y108_AQ;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_D3 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_D4 = CLBLM_L_X8Y113_SLICE_X11Y113_AQ;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_D5 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_D6 = CLBLM_R_X7Y115_SLICE_X9Y115_A5Q;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_D3 = 1'b1;
  assign RIOI3_X105Y101_ILOGIC_X1Y102_D = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_D4 = 1'b1;
  assign RIOI3_X105Y101_ILOGIC_X1Y101_D = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_A1 = CLBLL_L_X4Y112_SLICE_X4Y112_CO5;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_A2 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_A3 = CLBLM_L_X8Y113_SLICE_X10Y113_AQ;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_A4 = CLBLM_L_X10Y106_SLICE_X13Y106_AQ;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_A6 = 1'b1;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_D5 = 1'b1;
  assign CLBLM_L_X10Y115_SLICE_X12Y115_D6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y58_D = LIOB33_X0Y57_IOB_X0Y58_I;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_B1 = CLBLM_L_X10Y113_SLICE_X12Y113_CQ;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_B2 = CLBLM_L_X8Y113_SLICE_X10Y113_BQ;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_B3 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_B4 = CLBLM_R_X7Y114_SLICE_X9Y114_BQ;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_B5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_C1 = CLBLM_R_X11Y114_SLICE_X14Y114_AQ;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_C2 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_C4 = CLBLM_L_X8Y112_SLICE_X11Y112_CO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_C5 = CLBLM_R_X5Y113_SLICE_X6Y113_BQ;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_D1 = CLBLM_L_X10Y111_SLICE_X13Y111_C5Q;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_D2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_D3 = RIOB33_X105Y119_IOB_X1Y119_I;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_D4 = CLBLM_R_X5Y111_SLICE_X6Y111_CQ;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_D5 = CLBLM_L_X8Y113_SLICE_X10Y113_D5Q;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_D6 = 1'b1;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_A1 = CLBLM_R_X11Y117_SLICE_X15Y117_BO5;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_A2 = CLBLM_L_X10Y117_SLICE_X13Y117_AO6;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_A3 = CLBLM_R_X11Y117_SLICE_X15Y117_AQ;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_A4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_A6 = CLBLM_L_X12Y112_SLICE_X17Y112_A5Q;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_AX = CLBLM_R_X7Y113_SLICE_X9Y113_BO5;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_B1 = CLBLM_L_X10Y116_SLICE_X13Y116_AQ;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_B2 = CLBLM_L_X10Y117_SLICE_X12Y117_A5Q;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_B3 = 1'b1;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_B5 = CLBLM_R_X7Y118_SLICE_X8Y118_DO6;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_B6 = 1'b1;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_A1 = CLBLM_R_X7Y108_SLICE_X9Y108_DO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_A2 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_A3 = CLBLM_R_X7Y107_SLICE_X9Y107_CQ;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_A4 = 1'b1;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_A6 = CLBLM_L_X8Y119_SLICE_X10Y119_AQ;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_B3 = CLBLM_L_X8Y111_SLICE_X11Y111_BQ;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_C1 = CLBLM_R_X11Y116_SLICE_X15Y116_AQ;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_C2 = CLBLM_R_X11Y117_SLICE_X14Y117_CO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_B1 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_B2 = CLBLM_R_X7Y107_SLICE_X9Y107_BQ;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_B3 = CLBLM_R_X7Y107_SLICE_X9Y107_AQ;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_B4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_B6 = CLBLM_R_X5Y116_SLICE_X6Y116_D5Q;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_D1 = CLBLM_L_X10Y116_SLICE_X12Y116_DO5;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_D2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_C2 = CLBLM_R_X7Y110_SLICE_X9Y110_AQ;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_C3 = CLBLM_L_X8Y108_SLICE_X10Y108_AQ;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_C4 = CLBLM_R_X7Y107_SLICE_X9Y107_AQ;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_C5 = CLBLM_R_X7Y107_SLICE_X9Y107_DO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_C6 = 1'b1;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_D3 = CLBLM_R_X11Y117_SLICE_X15Y117_DQ;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_D4 = CLBLM_R_X11Y117_SLICE_X14Y117_BO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_A1 = CLBLM_R_X11Y117_SLICE_X14Y117_DO6;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_A2 = CLBLM_L_X10Y117_SLICE_X12Y117_DO6;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_A3 = CLBLM_R_X7Y118_SLICE_X9Y118_CO5;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_A4 = CLBLM_L_X10Y119_SLICE_X12Y119_CO6;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_A5 = CLBLM_R_X11Y116_SLICE_X14Y116_BQ;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_D1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_D2 = CLBLM_R_X7Y107_SLICE_X9Y107_CQ;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_D3 = CLBLM_R_X7Y108_SLICE_X8Y108_CQ;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_D4 = 1'b1;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_D5 = CLBLM_L_X10Y108_SLICE_X12Y108_CQ;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_D6 = CLBLM_R_X5Y105_SLICE_X6Y105_BQ;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_A6 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_B1 = CLBLM_L_X10Y116_SLICE_X13Y116_AQ;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_B2 = CLBLM_L_X10Y117_SLICE_X12Y117_DO6;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_B3 = CLBLM_L_X10Y117_SLICE_X13Y117_BO6;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_B4 = CLBLM_L_X10Y117_SLICE_X13Y117_DO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_A1 = CLBLM_R_X7Y105_SLICE_X8Y105_CQ;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_A2 = CLBLM_L_X8Y110_SLICE_X10Y110_BQ;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_A3 = CLBLM_R_X7Y107_SLICE_X8Y107_AQ;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_A4 = CLBLM_L_X12Y106_SLICE_X17Y106_AQ;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_A5 = CLBLL_L_X4Y110_SLICE_X4Y110_AQ;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_C1 = CLBLM_L_X10Y117_SLICE_X13Y117_BO6;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_C2 = CLBLM_L_X10Y116_SLICE_X12Y116_BQ;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_C3 = CLBLM_L_X10Y117_SLICE_X13Y117_DO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_B1 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_B2 = CLBLM_R_X7Y107_SLICE_X8Y107_BQ;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_B4 = CLBLM_R_X7Y107_SLICE_X9Y107_BQ;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_B5 = CLBLM_R_X5Y110_SLICE_X7Y110_AQ;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_B6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_D1 = CLBLM_L_X10Y118_SLICE_X12Y118_AQ;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_D2 = CLBLM_L_X8Y118_SLICE_X10Y118_AQ;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_D3 = CLBLM_L_X10Y118_SLICE_X13Y118_AQ;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_C1 = CLBLM_R_X7Y113_SLICE_X9Y113_AQ;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_C2 = CLBLM_R_X7Y107_SLICE_X8Y107_CQ;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_C3 = CLBLM_L_X8Y107_SLICE_X10Y107_CQ;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_C5 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_C6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_D4 = CLBLM_L_X10Y118_SLICE_X12Y118_BQ;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_D5 = CLBLM_R_X7Y118_SLICE_X8Y118_CQ;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_D6 = CLBLM_L_X10Y119_SLICE_X12Y119_AQ;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_D1 = CLBLM_R_X7Y106_SLICE_X9Y106_AQ;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_D2 = CLBLM_R_X7Y108_SLICE_X9Y108_AQ;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_D3 = CLBLM_L_X8Y110_SLICE_X10Y110_BQ;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_D4 = CLBLM_R_X7Y109_SLICE_X9Y109_CQ;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_D5 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_D6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign RIOB33_X105Y163_IOB_X1Y164_O = CLBLM_L_X8Y110_SLICE_X10Y110_CO5;
  assign RIOB33_X105Y163_IOB_X1Y163_O = CLBLM_L_X8Y110_SLICE_X10Y110_CO6;
  assign LIOB33_X0Y195_IOB_X0Y196_O = LIOB33_X0Y69_IOB_X0Y69_I;
  assign LIOB33_X0Y195_IOB_X0Y195_O = LIOB33_X0Y63_IOB_X0Y64_I;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_A1 = CLBLL_L_X4Y116_SLICE_X4Y116_BO6;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_A2 = CLBLM_L_X8Y111_SLICE_X11Y111_CQ;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_A3 = CLBLM_L_X8Y114_SLICE_X11Y114_AQ;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_A4 = CLBLM_R_X7Y115_SLICE_X9Y115_BQ;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_A5 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_B1 = CLBLM_L_X8Y109_SLICE_X11Y109_BQ;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_B2 = CLBLM_L_X8Y114_SLICE_X11Y114_BQ;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_B4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_B5 = CLBLM_L_X12Y117_SLICE_X17Y117_AQ;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_B6 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_C1 = CLBLM_L_X8Y115_SLICE_X11Y115_AQ;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_C2 = CLBLM_L_X10Y114_SLICE_X12Y114_BQ;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_C3 = CLBLM_L_X8Y111_SLICE_X10Y111_BO5;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_C5 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_C6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_D1 = CLBLM_L_X10Y111_SLICE_X12Y111_BQ;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_D2 = CLBLM_R_X7Y111_SLICE_X8Y111_CQ;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_D3 = CLBLM_R_X7Y117_SLICE_X9Y117_DQ;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_D4 = CLBLM_L_X8Y114_SLICE_X10Y114_CQ;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_D5 = CLBLM_R_X5Y117_SLICE_X7Y117_AQ;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_D6 = CLBLM_L_X10Y112_SLICE_X12Y112_BQ;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_A1 = CLBLM_R_X11Y113_SLICE_X15Y113_DQ;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_A2 = CLBLM_R_X5Y113_SLICE_X6Y113_BQ;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_A3 = CLBLM_L_X8Y114_SLICE_X10Y114_AQ;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_A4 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_A5 = CLBLL_L_X4Y112_SLICE_X4Y112_CO5;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_B1 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_B2 = CLBLM_L_X8Y114_SLICE_X10Y114_BQ;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_B4 = CLBLM_R_X7Y113_SLICE_X9Y113_A5Q;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_B5 = CLBLM_L_X12Y113_SLICE_X16Y113_BQ;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_B6 = CLBLM_R_X5Y115_SLICE_X7Y115_CO6;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_C2 = CLBLM_L_X8Y114_SLICE_X10Y114_CQ;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_C3 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_C4 = CLBLM_R_X7Y112_SLICE_X8Y112_CQ;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_C5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_C6 = CLBLM_L_X8Y115_SLICE_X10Y115_BQ;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_A1 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_A2 = CLBLM_R_X3Y108_SLICE_X2Y108_DO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_A3 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_A4 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_A5 = CLBLM_R_X3Y110_SLICE_X3Y110_DO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_A6 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_D1 = CLBLM_R_X7Y118_SLICE_X8Y118_BQ;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_D2 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_D3 = CLBLM_L_X10Y112_SLICE_X12Y112_CQ;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_D4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_D5 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_D6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_B1 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_B2 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_B3 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_B4 = CLBLM_R_X3Y111_SLICE_X2Y111_CO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_B5 = CLBLL_L_X2Y111_SLICE_X1Y111_DO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_C1 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_C2 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_C3 = CLBLM_R_X3Y109_SLICE_X2Y109_CO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_C4 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_C5 = CLBLM_R_X3Y110_SLICE_X2Y110_DO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_C6 = 1'b1;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_C4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_D1 = 1'b1;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_C5 = CLBLM_L_X10Y107_SLICE_X12Y107_DO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_D2 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_D3 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_D4 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_D5 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_D6 = 1'b1;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_A2 = CLBLL_L_X4Y118_SLICE_X4Y118_AQ;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_A3 = 1'b1;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_A4 = CLBLM_L_X12Y107_SLICE_X16Y107_BQ;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_A5 = RIOB33_X105Y125_IOB_X1Y126_I;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_A6 = 1'b1;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_B5 = CLBLM_R_X11Y106_SLICE_X14Y106_AQ;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_B1 = 1'b1;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_B2 = 1'b1;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_B3 = 1'b1;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_B4 = 1'b1;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_B5 = 1'b1;
  assign CLBLM_R_X11Y118_SLICE_X15Y118_B6 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_A1 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_A2 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_A3 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_A4 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_A5 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_A6 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_A1 = CLBLM_R_X7Y115_SLICE_X8Y115_CQ;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_A2 = CLBLM_L_X8Y110_SLICE_X10Y110_BQ;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_A3 = CLBLM_R_X7Y108_SLICE_X9Y108_AQ;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_B1 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_B2 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_B3 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_B4 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_B5 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_B6 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_B1 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_C1 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_C2 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_C3 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_C4 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_C5 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_C6 = 1'b1;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_D1 = CLBLM_L_X8Y106_SLICE_X11Y106_CO5;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_D2 = CLBLM_R_X5Y110_SLICE_X7Y110_DO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_C1 = CLBLL_L_X4Y107_SLICE_X5Y107_BO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_C2 = CLBLL_L_X4Y108_SLICE_X5Y108_AO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_C3 = CLBLM_L_X10Y112_SLICE_X12Y112_DO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_C4 = CLBLL_L_X2Y110_SLICE_X1Y110_DO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_D3 = CLBLL_L_X4Y107_SLICE_X5Y107_DO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_C6 = CLBLM_R_X3Y110_SLICE_X2Y110_DO6;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_D1 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_D2 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_D3 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_D4 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_D5 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_D6 = 1'b1;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_D5 = CLBLM_L_X10Y107_SLICE_X13Y107_CO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_D1 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_D2 = CLBLM_L_X8Y109_SLICE_X11Y109_CQ;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_D3 = CLBLM_R_X7Y107_SLICE_X9Y107_C5Q;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_D6 = CLBLM_R_X11Y111_SLICE_X14Y111_BO6;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_A1 = CLBLM_L_X8Y113_SLICE_X10Y113_D5Q;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_A2 = CLBLM_R_X5Y106_SLICE_X6Y106_BQ;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_A3 = CLBLM_R_X7Y108_SLICE_X8Y108_AQ;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_A4 = CLBLM_R_X7Y105_SLICE_X8Y105_CQ;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_A5 = CLBLL_L_X4Y110_SLICE_X4Y110_AQ;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_C1 = 1'b1;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_C2 = 1'b1;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_C3 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_B1 = CLBLL_L_X4Y112_SLICE_X4Y112_CO5;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_B2 = CLBLM_R_X7Y107_SLICE_X8Y107_AQ;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_B3 = CLBLM_R_X7Y109_SLICE_X9Y109_DQ;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_B4 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_B5 = CLBLM_R_X7Y108_SLICE_X8Y108_BQ;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_D1 = 1'b1;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_D2 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_C2 = CLBLM_L_X8Y112_SLICE_X10Y112_A5Q;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_C3 = CLBLM_L_X10Y108_SLICE_X12Y108_CQ;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_C5 = CLBLM_R_X7Y108_SLICE_X8Y108_DO6;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_C6 = 1'b1;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_D3 = 1'b1;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_D4 = 1'b1;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_D5 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_D6 = 1'b1;
  assign RIOB33_X105Y165_IOB_X1Y165_O = RIOB33_X105Y125_IOB_X1Y125_I;
  assign LIOI3_X0Y179_OLOGIC_X0Y180_T1 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_D1 = CLBLM_L_X8Y109_SLICE_X11Y109_AQ;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_D2 = CLBLM_R_X11Y111_SLICE_X15Y111_BQ;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_D3 = CLBLM_R_X5Y111_SLICE_X7Y111_CQ;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_D4 = CLBLM_R_X7Y115_SLICE_X8Y115_CQ;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_D5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_D6 = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_D1 = CLBLM_R_X5Y116_SLICE_X7Y116_A5Q;
  assign LIOI3_X0Y179_OLOGIC_X0Y179_D1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_A3 = CLBLM_L_X8Y107_SLICE_X10Y107_AQ;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_T1 = 1'b1;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign RIOI3_X105Y165_OLOGIC_X1Y166_D1 = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_A5 = CLBLM_L_X8Y108_SLICE_X10Y108_DQ;
  assign LIOI3_X0Y179_OLOGIC_X0Y179_T1 = 1'b1;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_A6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_D1 = CLBLM_R_X11Y118_SLICE_X15Y118_A5Q;
  assign RIOI3_X105Y165_OLOGIC_X1Y166_T1 = 1'b1;
  assign LIOB33_X0Y197_IOB_X0Y198_O = LIOB33_X0Y73_IOB_X0Y73_I;
  assign LIOB33_X0Y197_IOB_X0Y197_O = LIOB33_X0Y71_IOB_X0Y72_I;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_T1 = 1'b1;
  assign RIOI3_X105Y165_OLOGIC_X1Y165_D1 = RIOB33_X105Y125_IOB_X1Y125_I;
  assign RIOI3_X105Y165_OLOGIC_X1Y165_T1 = 1'b1;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_B1 = CLBLM_L_X10Y111_SLICE_X12Y111_CQ;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_B2 = CLBLM_L_X8Y107_SLICE_X10Y107_BQ;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_B3 = CLBLM_L_X10Y106_SLICE_X12Y106_BO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_B5 = CLBLM_L_X10Y110_SLICE_X13Y110_BQ;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_A1 = CLBLM_R_X7Y112_SLICE_X9Y112_DO6;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_A2 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_A3 = CLBLM_L_X8Y115_SLICE_X11Y115_AQ;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_A5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_A6 = CLBLM_R_X5Y116_SLICE_X7Y116_A5Q;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_B1 = CLBLM_R_X5Y109_SLICE_X6Y109_CQ;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_B2 = CLBLM_L_X8Y115_SLICE_X11Y115_BQ;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_B4 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_B5 = CLBLM_L_X8Y115_SLICE_X10Y115_AQ;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_B6 = CLBLM_R_X7Y115_SLICE_X9Y115_DO6;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_C1 = CLBLM_L_X10Y114_SLICE_X12Y114_BQ;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_C2 = CLBLM_L_X8Y114_SLICE_X11Y114_CQ;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_C3 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_C4 = CLBLM_L_X8Y115_SLICE_X10Y115_CQ;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_C5 = CLBLM_L_X8Y115_SLICE_X11Y115_DO6;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_C6 = CLBLM_R_X13Y117_SLICE_X18Y117_BQ;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_C1 = CLBLM_L_X8Y107_SLICE_X10Y107_DO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_C2 = CLBLM_L_X10Y107_SLICE_X12Y107_CO6;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_D1 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_D2 = CLBLM_L_X12Y112_SLICE_X17Y112_BQ;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_D3 = CLBLM_L_X12Y112_SLICE_X16Y112_AQ;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_D4 = CLBLM_L_X8Y116_SLICE_X11Y116_BQ;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_D5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y115_SLICE_X11Y115_D6 = CLBLM_R_X7Y115_SLICE_X9Y115_BQ;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_C4 = CLBLM_R_X11Y108_SLICE_X14Y108_BO6;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_A1 = CLBLM_L_X10Y115_SLICE_X13Y115_BQ;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_A2 = CLBLM_R_X11Y118_SLICE_X15Y118_AQ;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_A3 = CLBLM_L_X8Y115_SLICE_X10Y115_AQ;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_A4 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_A6 = CLBLM_R_X7Y115_SLICE_X9Y115_DO6;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_AX = CLBLM_R_X11Y115_SLICE_X14Y115_AO6;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_B1 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_B2 = CLBLM_L_X8Y115_SLICE_X10Y115_BQ;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_B4 = CLBLM_R_X7Y111_SLICE_X9Y111_CQ;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_B6 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_C1 = CLBLM_L_X8Y114_SLICE_X10Y114_AQ;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_A1 = CLBLL_L_X4Y107_SLICE_X5Y107_DO6;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_C5 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_A2 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_A3 = CLBLL_L_X2Y110_SLICE_X1Y110_DO6;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_A4 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_C6 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_A5 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_A6 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_B1 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_B2 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_B3 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_B4 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_B5 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_B6 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_D1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_D2 = CLBLM_L_X10Y115_SLICE_X12Y115_AQ;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_C1 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_C2 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_C3 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_C4 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_C5 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_C6 = 1'b1;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_D5 = CLBLL_L_X4Y114_SLICE_X4Y114_BQ;
  assign CLBLM_L_X8Y115_SLICE_X10Y115_D6 = CLBLM_R_X7Y111_SLICE_X9Y111_CQ;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_D1 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_D2 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_D3 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_D4 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_D5 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_D6 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_A1 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_A2 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_A3 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_A4 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_A5 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_A6 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_B1 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_B2 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_B3 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_B4 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_B5 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_A1 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_A2 = CLBLM_R_X3Y107_SLICE_X3Y107_AQ;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_A3 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_A4 = CLBLL_L_X4Y107_SLICE_X5Y107_DO6;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_A5 = CLBLM_R_X5Y106_SLICE_X7Y106_CO6;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_A6 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_A1 = CLBLM_R_X7Y110_SLICE_X9Y110_BQ;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_A2 = CLBLM_R_X7Y111_SLICE_X8Y111_BQ;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_A3 = CLBLM_R_X7Y109_SLICE_X9Y109_AQ;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_B1 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_B2 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_B3 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_B4 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_B5 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_B6 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_A4 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_A6 = CLBLL_L_X4Y112_SLICE_X4Y112_CO6;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_C1 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_C2 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_C3 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_C4 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_C5 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_C6 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_C2 = CLBLM_R_X7Y109_SLICE_X9Y109_CQ;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_C3 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_C4 = CLBLM_L_X8Y114_SLICE_X11Y114_CQ;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_C5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_C6 = CLBLM_L_X10Y113_SLICE_X13Y113_AQ;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_D1 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_D2 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_D3 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_D4 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_D5 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_D6 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_C3 = CLBLL_L_X2Y114_SLICE_X0Y114_AO5;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_D1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_D2 = CLBLM_L_X8Y109_SLICE_X11Y109_DO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_D3 = CLBLM_L_X12Y112_SLICE_X16Y112_B5Q;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_D4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_D5 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_D6 = CLBLM_R_X5Y106_SLICE_X6Y106_DQ;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_B1 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_A1 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_A3 = CLBLM_R_X7Y109_SLICE_X8Y109_AQ;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_A4 = CLBLL_L_X4Y116_SLICE_X4Y116_BO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_A5 = CLBLM_R_X5Y109_SLICE_X6Y109_DQ;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_A6 = CLBLM_L_X8Y114_SLICE_X11Y114_CQ;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_C1 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_C2 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_C3 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_B1 = CLBLL_L_X4Y112_SLICE_X4Y112_CO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_B2 = CLBLM_R_X7Y109_SLICE_X8Y109_BQ;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_B3 = CLBLM_R_X5Y108_SLICE_X7Y108_AQ;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_C4 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_B4 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_B6 = CLBLM_R_X7Y111_SLICE_X9Y111_BQ;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_D1 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_C1 = CLBLM_R_X7Y113_SLICE_X9Y113_AQ;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_C2 = CLBLM_R_X5Y109_SLICE_X6Y109_DQ;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_C3 = CLBLL_L_X4Y109_SLICE_X5Y109_AQ;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_C4 = CLBLM_L_X8Y112_SLICE_X10Y112_A5Q;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_C5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_C6 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_D2 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_D3 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_D4 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_D6 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_D1 = CLBLM_L_X10Y104_SLICE_X12Y104_AQ;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_C5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_D2 = CLBLL_L_X2Y111_SLICE_X1Y111_DO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_D3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_D4 = CLBLM_R_X7Y109_SLICE_X8Y109_CO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_D5 = CLBLM_R_X7Y116_SLICE_X8Y116_CQ;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_D6 = 1'b1;
  assign LIOI3_X0Y173_OLOGIC_X0Y173_D1 = CLBLM_R_X7Y132_SLICE_X9Y132_AO5;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_A1 = CLBLM_R_X7Y116_SLICE_X8Y116_BQ;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_A2 = CLBLM_L_X12Y108_SLICE_X17Y108_BQ;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_A4 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_A5 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_A6 = CLBLM_L_X10Y116_SLICE_X12Y116_DO6;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_B1 = CLBLM_L_X8Y116_SLICE_X11Y116_DO6;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_B2 = CLBLM_L_X8Y116_SLICE_X11Y116_BQ;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_B3 = CLBLM_L_X10Y117_SLICE_X12Y117_AQ;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_B5 = CLBLM_L_X12Y112_SLICE_X17Y112_BQ;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_C1 = CLBLM_R_X7Y114_SLICE_X8Y114_A5Q;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_C2 = CLBLM_L_X10Y115_SLICE_X13Y115_CQ;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_C3 = CLBLM_R_X7Y118_SLICE_X8Y118_CQ;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_C4 = CLBLM_L_X8Y118_SLICE_X10Y118_AQ;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_C5 = CLBLM_R_X11Y117_SLICE_X15Y117_AQ;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_C6 = CLBLM_L_X10Y119_SLICE_X12Y119_AQ;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A2 = CLBLL_L_X4Y112_SLICE_X4Y112_CO5;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_D1 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_D2 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_D3 = CLBLM_R_X13Y117_SLICE_X18Y117_BQ;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_D4 = CLBLM_R_X5Y112_SLICE_X7Y112_CQ;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A3 = CLBLL_L_X4Y113_SLICE_X4Y113_AQ;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_D5 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_D6 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_A1 = CLBLM_L_X8Y113_SLICE_X10Y113_DQ;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_A2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A5 = CLBLM_R_X5Y105_SLICE_X6Y105_BQ;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_A3 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_A5 = CLBLM_R_X5Y112_SLICE_X7Y112_BQ;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_A6 = RIOB33_X105Y119_IOB_X1Y119_I;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_B1 = CLBLM_R_X7Y118_SLICE_X8Y118_DO6;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_B2 = CLBLM_L_X8Y116_SLICE_X10Y116_BQ;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_B3 = CLBLM_L_X8Y117_SLICE_X10Y117_AQ;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_B4 = CLBLM_R_X5Y112_SLICE_X6Y112_AQ;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_B5 = CLBLM_L_X10Y117_SLICE_X13Y117_AO5;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_A1 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_A2 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_A3 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_C1 = CLBLM_R_X7Y115_SLICE_X9Y115_B5Q;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_C2 = CLBLM_L_X8Y116_SLICE_X10Y116_CQ;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_C3 = CLBLM_L_X10Y117_SLICE_X13Y117_AO5;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_C5 = CLBLM_R_X7Y118_SLICE_X8Y118_DO6;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_C6 = CLBLM_L_X10Y116_SLICE_X12Y116_AQ;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_A4 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_A5 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_A6 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_B5 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_B6 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_B1 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_B2 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_B3 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_B4 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_D1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B3 = CLBLM_R_X5Y112_SLICE_X6Y112_AQ;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_D2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_D3 = CLBLM_L_X8Y116_SLICE_X10Y116_DQ;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_D4 = CLBLM_R_X11Y113_SLICE_X14Y113_CQ;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_D5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B4 = CLBLL_L_X4Y114_SLICE_X4Y114_AQ;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_D6 = CLBLM_L_X10Y115_SLICE_X13Y115_CQ;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_C4 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_C5 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B5 = CLBLM_R_X3Y112_SLICE_X3Y112_AQ;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_D1 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_D2 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_D3 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B6 = CLBLM_R_X11Y113_SLICE_X14Y113_AQ;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_D4 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_D5 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_D6 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C1 = CLBLM_R_X3Y115_SLICE_X2Y115_AQ;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_A1 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_A2 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_A3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_A4 = CLBLL_L_X2Y114_SLICE_X0Y114_AO6;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_A5 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_A6 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_B1 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_B2 = CLBLM_R_X3Y116_SLICE_X3Y116_AO6;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_B3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_B4 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_B5 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_B6 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_A1 = CLBLM_L_X8Y113_SLICE_X10Y113_CQ;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_A2 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C6 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_C1 = CLBLM_R_X3Y111_SLICE_X3Y111_AO6;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_C2 = CLBLL_L_X2Y109_SLICE_X0Y109_AO6;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_C3 = LIOB33_X0Y67_IOB_X0Y67_I;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_C4 = CLBLL_L_X2Y108_SLICE_X1Y108_AO6;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_C5 = CLBLL_L_X2Y108_SLICE_X1Y108_DO6;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_C6 = CLBLM_R_X7Y106_SLICE_X8Y106_AQ;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_B1 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_B2 = CLBLM_R_X7Y110_SLICE_X9Y110_BQ;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_B3 = CLBLM_R_X7Y113_SLICE_X8Y113_C5Q;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_B5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_B6 = CLBLM_R_X7Y110_SLICE_X9Y110_CO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_D1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_D2 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_D3 = CLBLL_L_X2Y114_SLICE_X0Y114_AO5;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_D4 = CLBLL_L_X4Y115_SLICE_X5Y115_BQ;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_D5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_D6 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_C4 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_C4 = CLBLM_L_X8Y110_SLICE_X10Y110_DO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_C6 = CLBLM_R_X7Y111_SLICE_X9Y111_DO5;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_C5 = CLBLM_L_X12Y111_SLICE_X16Y111_BQ;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_D1 = CLBLM_R_X7Y109_SLICE_X8Y109_CO5;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_D2 = CLBLM_L_X10Y104_SLICE_X12Y104_AQ;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_D3 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_C6 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_D4 = CLBLM_R_X7Y116_SLICE_X8Y116_CQ;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_D5 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_D6 = CLBLL_L_X4Y108_SLICE_X5Y108_AO6;
  assign RIOB33_X105Y167_IOB_X1Y167_O = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign RIOB33_X105Y167_IOB_X1Y168_O = CLBLM_L_X10Y148_SLICE_X12Y148_AO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_A1 = CLBLM_R_X11Y110_SLICE_X14Y110_A5Q;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_A2 = CLBLM_R_X7Y105_SLICE_X9Y105_CQ;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_A3 = CLBLM_R_X7Y110_SLICE_X8Y110_AQ;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_A4 = CLBLM_R_X7Y105_SLICE_X8Y105_CQ;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_A5 = CLBLL_L_X4Y110_SLICE_X4Y110_AQ;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_B1 = CLBLM_R_X5Y114_SLICE_X7Y114_BQ;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_B2 = CLBLM_R_X7Y105_SLICE_X8Y105_A5Q;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_B4 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_B6 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_C1 = CLBLM_R_X7Y112_SLICE_X8Y112_AQ;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_C2 = CLBLM_R_X7Y110_SLICE_X8Y110_CQ;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_C3 = CLBLM_R_X5Y115_SLICE_X7Y115_CO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_C5 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_C6 = CLBLM_L_X8Y109_SLICE_X11Y109_CQ;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_A5 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_A6 = LIOB33_X0Y67_IOB_X0Y68_I;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_D2 = CLBLL_L_X2Y110_SLICE_X1Y110_DO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_D3 = CLBLM_L_X8Y106_SLICE_X11Y106_AQ;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_D4 = CLBLM_R_X5Y106_SLICE_X6Y106_CQ;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_D5 = CLBLM_L_X10Y113_SLICE_X13Y113_CQ;
  assign CLBLM_L_X12Y114_SLICE_X17Y114_D1 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_D6 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_A1 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_A2 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_A3 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_A4 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_A5 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_A6 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_B1 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_B2 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_B3 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_B4 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_B5 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_B6 = 1'b1;
  assign LIOI3_X0Y183_OLOGIC_X0Y184_D1 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_C1 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_C2 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_C3 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_C4 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_C5 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_C6 = 1'b1;
  assign LIOI3_X0Y183_OLOGIC_X0Y184_T1 = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_D1 = CLBLM_R_X5Y114_SLICE_X7Y114_C5Q;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_D1 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_D2 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_D3 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_D4 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_D5 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_D6 = 1'b1;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_C4 = CLBLM_L_X10Y118_SLICE_X13Y118_CO6;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_C5 = CLBLM_L_X12Y110_SLICE_X17Y110_DQ;
  assign LIOI3_X0Y183_OLOGIC_X0Y183_D1 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_T1 = 1'b1;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_A1 = CLBLM_R_X7Y118_SLICE_X8Y118_DO6;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_A2 = CLBLM_L_X10Y117_SLICE_X13Y117_AO5;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_A3 = CLBLM_L_X8Y117_SLICE_X10Y117_AQ;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_A4 = CLBLM_R_X5Y116_SLICE_X7Y116_BQ;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_A5 = CLBLM_L_X10Y116_SLICE_X13Y116_BQ;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOI3_X0Y183_OLOGIC_X0Y183_T1 = 1'b1;
  assign RIOI3_X105Y167_OLOGIC_X1Y168_D1 = CLBLM_L_X10Y148_SLICE_X12Y148_AO6;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_D1 = CLBLM_R_X7Y113_SLICE_X8Y113_C5Q;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_B1 = CLBLM_R_X13Y113_SLICE_X18Y113_BQ;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_B2 = CLBLM_L_X10Y117_SLICE_X13Y117_AO5;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_B3 = CLBLM_R_X7Y110_SLICE_X8Y110_DO5;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_B4 = CLBLM_L_X8Y118_SLICE_X10Y118_DO5;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_B6 = CLBLM_L_X8Y117_SLICE_X10Y117_CO6;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_A5 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_A6 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_A1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_A2 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_A3 = CLBLL_L_X2Y114_SLICE_X0Y114_AO5;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_A4 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_C1 = CLBLM_L_X10Y116_SLICE_X12Y116_DO6;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_C2 = CLBLM_R_X11Y117_SLICE_X15Y117_AQ;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_C3 = CLBLM_L_X8Y117_SLICE_X10Y117_BQ;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_C4 = CLBLM_R_X7Y116_SLICE_X8Y116_BQ;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_C5 = CLBLM_L_X8Y117_SLICE_X10Y117_DO6;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_C6 = CLBLM_R_X7Y116_SLICE_X9Y116_CO6;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_B1 = CLBLM_R_X3Y116_SLICE_X3Y116_AO6;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_B2 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_C1 = CLBLL_L_X2Y107_SLICE_X1Y107_AO6;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_C2 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_B5 = CLBLL_L_X2Y109_SLICE_X0Y109_CO6;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_B6 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_C6 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_D1 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_D2 = CLBLM_L_X10Y119_SLICE_X12Y119_AQ;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_D3 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_D4 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_D5 = CLBLM_R_X7Y118_SLICE_X8Y118_CQ;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_D6 = CLBLM_R_X7Y114_SLICE_X8Y114_A5Q;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_D1 = CLBLL_L_X2Y112_SLICE_X0Y112_AO6;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_D2 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_D3 = LIOB33_X0Y67_IOB_X0Y67_I;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_D4 = CLBLL_L_X2Y114_SLICE_X0Y114_AO5;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_D5 = CLBLL_L_X2Y112_SLICE_X0Y112_AO5;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_D6 = CLBLL_L_X4Y115_SLICE_X5Y115_BQ;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_D2 = CLBLM_L_X10Y115_SLICE_X13Y115_CQ;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_D1 = CLBLM_R_X3Y106_SLICE_X2Y106_BO6;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_C4 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_D5 = CLBLM_R_X7Y118_SLICE_X9Y118_BO5;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_T1 = 1'b1;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_C5 = CLBLM_L_X10Y111_SLICE_X13Y111_DO6;
  assign CLBLM_L_X10Y116_SLICE_X13Y116_D6 = CLBLM_L_X8Y118_SLICE_X10Y118_AQ;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign RIOB33_X105Y171_IOB_X1Y172_O = CLBLM_R_X103Y173_SLICE_X163Y173_AO6;
  assign RIOB33_X105Y171_IOB_X1Y171_O = CLBLM_R_X103Y170_SLICE_X163Y170_AO5;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_A1 = CLBLL_L_X2Y108_SLICE_X1Y108_BO5;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_A2 = CLBLL_L_X2Y111_SLICE_X1Y111_BO6;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_A3 = CLBLL_L_X2Y109_SLICE_X0Y109_CO6;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_A4 = CLBLL_L_X2Y108_SLICE_X1Y108_AO5;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_A5 = CLBLL_L_X2Y110_SLICE_X0Y110_BO5;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_A6 = CLBLL_L_X2Y110_SLICE_X1Y110_AO5;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_B1 = CLBLL_L_X2Y108_SLICE_X1Y108_BO5;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_B2 = CLBLL_L_X2Y111_SLICE_X1Y111_BO6;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_B3 = CLBLL_L_X2Y109_SLICE_X0Y109_CO6;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_B4 = CLBLL_L_X2Y110_SLICE_X0Y110_BO5;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_B5 = CLBLL_L_X2Y111_SLICE_X1Y111_AO5;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_B6 = CLBLL_L_X2Y110_SLICE_X1Y110_AO5;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_A1 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_A2 = CLBLM_R_X7Y110_SLICE_X9Y110_DO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_A3 = CLBLM_R_X7Y111_SLICE_X9Y111_AQ;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_C1 = CLBLL_L_X2Y112_SLICE_X1Y112_AO6;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_C2 = CLBLL_L_X2Y109_SLICE_X0Y109_CO6;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_C3 = CLBLL_L_X2Y110_SLICE_X0Y110_BO5;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_C4 = CLBLL_L_X2Y110_SLICE_X1Y110_AO5;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_C5 = CLBLL_L_X2Y108_SLICE_X1Y108_BO5;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_C6 = CLBLL_L_X2Y111_SLICE_X1Y111_BO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_A4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_A6 = CLBLL_L_X4Y113_SLICE_X5Y113_BQ;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_B1 = CLBLM_L_X12Y111_SLICE_X16Y111_CQ;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_B2 = CLBLM_R_X7Y111_SLICE_X9Y111_BQ;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_B4 = CLBLM_R_X7Y110_SLICE_X9Y110_AQ;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_D1 = CLBLL_L_X2Y114_SLICE_X1Y114_AO6;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_D2 = CLBLL_L_X4Y115_SLICE_X5Y115_BQ;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_D3 = LIOB33_X0Y67_IOB_X0Y67_I;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_D4 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_D5 = CLBLL_L_X2Y109_SLICE_X0Y109_AO6;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_D6 = CLBLM_R_X3Y111_SLICE_X3Y111_AO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_C2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_C3 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_C4 = CLBLM_L_X8Y112_SLICE_X10Y112_CO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_C5 = CLBLM_R_X5Y105_SLICE_X6Y105_AQ;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_C6 = CLBLM_R_X7Y110_SLICE_X9Y110_AQ;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_D1 = CLBLM_R_X7Y111_SLICE_X8Y111_AQ;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_D2 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_D3 = CLBLM_R_X5Y114_SLICE_X7Y114_BQ;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_D4 = CLBLM_R_X11Y112_SLICE_X14Y112_CQ;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_D5 = CLBLM_L_X8Y113_SLICE_X11Y113_BQ;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_D6 = 1'b1;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_A6 = CLBLM_L_X10Y117_SLICE_X13Y117_AO5;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_A1 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_A3 = CLBLM_R_X7Y111_SLICE_X8Y111_AQ;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_A4 = CLBLM_L_X8Y112_SLICE_X10Y112_BO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_A5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X12Y114_SLICE_X16Y114_D5 = CLBLM_L_X12Y113_SLICE_X16Y113_AQ;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_A6 = CLBLL_L_X4Y116_SLICE_X4Y116_A5Q;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_B1 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_B2 = CLBLM_R_X7Y107_SLICE_X8Y107_BQ;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_B4 = CLBLM_R_X7Y114_SLICE_X8Y114_CQ;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_B5 = CLBLM_L_X8Y111_SLICE_X10Y111_DO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_A4 = CLBLM_L_X12Y117_SLICE_X16Y117_AQ;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_C2 = CLBLM_R_X7Y111_SLICE_X8Y111_CQ;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_B1 = CLBLM_R_X7Y118_SLICE_X8Y118_DO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_C3 = CLBLM_R_X7Y111_SLICE_X8Y111_DQ;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_C5 = CLBLM_R_X7Y112_SLICE_X8Y112_CQ;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_C6 = 1'b1;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_B2 = CLBLM_L_X10Y116_SLICE_X12Y116_BQ;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_B4 = CLBLM_R_X5Y115_SLICE_X7Y115_BQ;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_D2 = CLBLM_R_X5Y111_SLICE_X6Y111_CQ;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_D3 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_D4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_D5 = CLBLM_R_X7Y109_SLICE_X8Y109_CO5;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_B5 = CLBLM_L_X10Y116_SLICE_X12Y116_CQ;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_D6 = CLBLM_L_X10Y113_SLICE_X13Y113_CQ;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_D3 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_D4 = 1'b1;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_B6 = CLBLM_L_X10Y117_SLICE_X13Y117_AO5;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_D5 = 1'b1;
  assign LIOI3_SING_X0Y50_ILOGIC_X0Y50_D = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign CLBLM_R_X103Y138_SLICE_X163Y138_D6 = 1'b1;
  assign LIOI3_X0Y61_ILOGIC_X0Y62_D = LIOB33_X0Y61_IOB_X0Y62_I;
  assign LIOI3_X0Y61_ILOGIC_X0Y61_D = LIOB33_X0Y61_IOB_X0Y61_I;
  assign CLBLM_R_X11Y112_SLICE_X15Y112_A5 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign RIOI3_X105Y105_ILOGIC_X1Y106_D = RIOB33_X105Y105_IOB_X1Y106_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y105_D = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_C2 = CLBLM_L_X10Y116_SLICE_X12Y116_CQ;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_C3 = CLBLM_R_X7Y118_SLICE_X8Y118_DO6;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_C4 = CLBLM_L_X8Y116_SLICE_X10Y116_CQ;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_A1 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_A2 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_A3 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_A4 = RIOB33_X105Y123_IOB_X1Y124_I;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_A5 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_A6 = 1'b1;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_C5 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_C6 = CLBLM_L_X10Y117_SLICE_X13Y117_AO5;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y114_D = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_B1 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_B2 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_B3 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_B4 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_B5 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_B6 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_D = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_C1 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_C2 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_A1 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_A2 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_A3 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_C6 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_A4 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_A5 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_A6 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_C3 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_C4 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_C5 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_B1 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_B2 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_B3 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_B4 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_D3 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_D4 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_B5 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_B6 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_D1 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_D2 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_C1 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_C2 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_C3 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_C4 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_C5 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_C6 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_D1 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_D2 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_D3 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_D4 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_D5 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_D6 = 1'b1;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_D1 = CLBLM_L_X10Y119_SLICE_X12Y119_AQ;
  assign CLBLM_L_X10Y116_SLICE_X12Y116_D2 = CLBLM_R_X7Y114_SLICE_X8Y114_A5Q;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_B4 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_A1 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_A2 = CLBLM_L_X10Y117_SLICE_X13Y117_CO6;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_A3 = CLBLM_L_X8Y118_SLICE_X10Y118_AQ;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_A4 = CLBLM_L_X8Y116_SLICE_X11Y116_BQ;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_A6 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_A5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_A6 = CLBLM_L_X8Y118_SLICE_X10Y118_CO6;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_A1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_A2 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_A3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_A4 = CLBLL_L_X2Y114_SLICE_X0Y114_AO6;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_A5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_A6 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_B1 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_B2 = CLBLM_L_X8Y118_SLICE_X10Y118_BQ;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_B1 = CLBLM_R_X3Y116_SLICE_X3Y116_AO6;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_B2 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_B3 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_B4 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_B5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_B6 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_B6 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_C1 = CLBLM_R_X7Y114_SLICE_X8Y114_A5Q;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_C1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_C2 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_C3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_C4 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_C4 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_C5 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_C6 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_D1 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_D2 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_D3 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_D4 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_D5 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_D6 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_D1 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_B4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_D2 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_D3 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_D4 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_D5 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_D6 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_B5 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_B6 = CLBLM_R_X7Y117_SLICE_X8Y117_BQ;
  assign RIOB33_X105Y173_IOB_X1Y173_O = CLBLM_R_X103Y173_SLICE_X163Y173_AO5;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_C6 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_A1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_A2 = CLBLM_R_X3Y116_SLICE_X3Y116_AO6;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_A3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_A4 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_A5 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_A6 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_B1 = CLBLL_L_X2Y112_SLICE_X0Y112_CO6;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_B2 = CLBLL_L_X2Y108_SLICE_X1Y108_AO5;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_C2 = CLBLM_L_X10Y119_SLICE_X12Y119_AQ;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_B3 = CLBLL_L_X2Y110_SLICE_X0Y110_AO6;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_B4 = CLBLL_L_X2Y110_SLICE_X0Y110_CO6;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_B5 = CLBLL_L_X2Y109_SLICE_X0Y109_CO6;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_B6 = CLBLL_L_X2Y110_SLICE_X1Y110_AO5;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_C3 = CLBLM_L_X8Y118_SLICE_X10Y118_AQ;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_C1 = CLBLL_L_X2Y111_SLICE_X1Y111_AO6;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_C2 = CLBLL_L_X2Y110_SLICE_X0Y110_CO6;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_C4 = CLBLM_R_X11Y117_SLICE_X15Y117_AQ;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_C3 = CLBLL_L_X2Y110_SLICE_X0Y110_BO6;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_C4 = CLBLL_L_X2Y109_SLICE_X0Y109_CO6;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_C5 = CLBLL_L_X2Y110_SLICE_X1Y110_AO6;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_C6 = CLBLL_L_X2Y111_SLICE_X1Y111_BO6;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_C5 = CLBLM_R_X7Y118_SLICE_X8Y118_CQ;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_A1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_A2 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_A4 = CLBLM_L_X8Y112_SLICE_X11Y112_DO6;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_C6 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_A6 = CLBLM_R_X7Y108_SLICE_X8Y108_CQ;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_D1 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_D2 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_D3 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_D4 = CLBLM_R_X3Y110_SLICE_X2Y110_CO6;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_D5 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_D6 = CLBLL_L_X2Y112_SLICE_X1Y112_BO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_B4 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_B6 = CLBLM_L_X10Y111_SLICE_X13Y111_C5Q;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_C1 = CLBLM_R_X7Y109_SLICE_X8Y109_DO5;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_C2 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_C3 = CLBLM_R_X7Y113_SLICE_X9Y113_CO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_C4 = CLBLM_R_X11Y112_SLICE_X14Y112_CQ;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_C5 = CLBLM_R_X3Y110_SLICE_X2Y110_DO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_C6 = CLBLM_L_X8Y113_SLICE_X11Y113_BQ;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_D1 = CLBLM_R_X7Y109_SLICE_X8Y109_DO5;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_D2 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_D3 = CLBLM_R_X7Y113_SLICE_X9Y113_CO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_D4 = CLBLM_R_X7Y115_SLICE_X8Y115_CQ;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_D5 = CLBLM_R_X5Y111_SLICE_X7Y111_CQ;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_D6 = CLBLM_R_X3Y110_SLICE_X3Y110_AO6;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_A1 = CLBLM_R_X7Y114_SLICE_X8Y114_DO6;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_A3 = CLBLM_R_X7Y112_SLICE_X8Y112_AQ;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_A4 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_A6 = CLBLM_L_X10Y112_SLICE_X12Y112_AQ;
  assign LIOB33_X0Y163_IOB_X0Y163_O = RIOB33_X105Y109_IOB_X1Y110_I;
  assign LIOB33_X0Y163_IOB_X0Y164_O = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_B1 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_B2 = CLBLM_R_X7Y112_SLICE_X8Y112_BQ;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_B4 = CLBLM_R_X7Y113_SLICE_X8Y113_AQ;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_B6 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_D1 = CLBLM_L_X10Y117_SLICE_X13Y117_CO6;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_C1 = CLBLL_L_X4Y107_SLICE_X5Y107_AQ;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_C2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_D2 = CLBLM_L_X8Y118_SLICE_X10Y118_AQ;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_C4 = CLBLM_L_X10Y112_SLICE_X12Y112_AQ;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_C5 = CLBLM_R_X11Y112_SLICE_X14Y112_CQ;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_C6 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_D3 = CLBLM_R_X7Y118_SLICE_X8Y118_CQ;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_D4 = CLBLM_L_X10Y119_SLICE_X12Y119_AQ;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_D1 = CLBLM_L_X10Y104_SLICE_X12Y104_BO6;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_D2 = CLBLM_L_X8Y114_SLICE_X11Y114_B5Q;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_D5 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_D3 = CLBLM_R_X7Y112_SLICE_X8Y112_DQ;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_D4 = CLBLM_R_X5Y106_SLICE_X6Y106_CQ;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_D5 = CLBLM_R_X7Y113_SLICE_X8Y113_DQ;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_D6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_D6 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_A1 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_A2 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_A3 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_A4 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_A5 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_A6 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_B1 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_B2 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_B3 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_B4 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_B5 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_B6 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_C1 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_C2 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_C3 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_C4 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_C5 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_C6 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_D1 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_D2 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_D3 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_D4 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_D5 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_D6 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_A1 = CLBLM_L_X10Y115_SLICE_X13Y115_BQ;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_A3 = CLBLM_L_X8Y119_SLICE_X10Y119_AQ;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_A1 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_A2 = CLBLL_L_X2Y114_SLICE_X0Y114_AO5;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_A3 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_A4 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_A5 = CLBLM_L_X12Y112_SLICE_X16Y112_B5Q;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_A6 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_A4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_B1 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_B1 = CLBLL_L_X2Y112_SLICE_X0Y112_CO6;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_B2 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_B3 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_B4 = CLBLL_L_X2Y114_SLICE_X0Y114_AO6;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_B5 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_B6 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_B3 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_B4 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_B5 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_C1 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_C2 = CLBLM_R_X5Y110_SLICE_X7Y110_AQ;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_C3 = LIOB33_X0Y57_IOB_X0Y58_I;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_C4 = CLBLL_L_X2Y114_SLICE_X0Y114_AO5;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_C5 = CLBLL_L_X2Y112_SLICE_X1Y112_DO6;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_C6 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_C1 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_C2 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_C3 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_C4 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_C5 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_C6 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_D1 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_D2 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_D3 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_D4 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_D5 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_D6 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_D1 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_D2 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_D3 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_D4 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_D5 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_D6 = 1'b1;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_C2 = CLBLM_L_X10Y112_SLICE_X12Y112_DO6;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_C3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_C4 = CLBLM_R_X3Y110_SLICE_X3Y110_DO6;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_A1 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_A2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_A3 = CLBLM_R_X3Y116_SLICE_X3Y116_AO6;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_A4 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_A5 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_A6 = 1'b1;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_C5 = CLBLM_L_X8Y108_SLICE_X11Y108_DO6;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_B1 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_B2 = CLBLL_L_X2Y114_SLICE_X0Y114_AO6;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_B3 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_B4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_B5 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_B6 = 1'b1;
  assign LIOI3_X0Y185_OLOGIC_X0Y186_D1 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_C1 = CLBLL_L_X2Y113_SLICE_X0Y113_AO6;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_C2 = CLBLM_R_X3Y111_SLICE_X2Y111_BO6;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_C3 = CLBLM_R_X3Y113_SLICE_X3Y113_DO6;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_C4 = CLBLM_R_X3Y112_SLICE_X2Y112_CO6;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_C5 = CLBLL_L_X4Y109_SLICE_X4Y109_CO6;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_C6 = CLBLL_L_X2Y110_SLICE_X1Y110_BO6;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_D2 = CLBLM_R_X7Y117_SLICE_X9Y117_A5Q;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_A1 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_A2 = CLBLM_L_X8Y112_SLICE_X10Y112_CO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_A3 = CLBLM_R_X7Y113_SLICE_X9Y113_AQ;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_A5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_A6 = CLBLM_L_X10Y116_SLICE_X12Y116_CQ;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_D1 = CLBLL_L_X2Y109_SLICE_X0Y109_BO6;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_D2 = CLBLM_R_X3Y111_SLICE_X2Y111_BO6;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_D3 = CLBLL_L_X2Y111_SLICE_X0Y111_BO6;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_D4 = CLBLM_R_X3Y112_SLICE_X3Y112_BO6;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_D5 = CLBLM_R_X7Y115_SLICE_X9Y115_AQ;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_D6 = CLBLM_R_X3Y111_SLICE_X2Y111_AO6;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_D5 = CLBLM_R_X5Y116_SLICE_X7Y116_AQ;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_D6 = CLBLM_R_X5Y115_SLICE_X6Y115_BQ;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_B1 = CLBLM_R_X5Y116_SLICE_X6Y116_CQ;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_B2 = CLBLM_L_X10Y111_SLICE_X13Y111_C5Q;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_B5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_B6 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_C2 = CLBLM_L_X10Y104_SLICE_X12Y104_AQ;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_C4 = CLBLM_R_X7Y116_SLICE_X8Y116_CQ;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_C5 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_D1 = CLBLL_L_X4Y107_SLICE_X4Y107_CQ;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_C6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_D1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_D2 = CLBLM_L_X8Y106_SLICE_X10Y106_CQ;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_D2 = CLBLM_L_X8Y109_SLICE_X10Y109_BQ;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_D5 = CLBLM_R_X7Y117_SLICE_X9Y117_DQ;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_D6 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_D3 = CLBLM_R_X7Y114_SLICE_X9Y114_AO5;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_D3 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_D4 = CLBLM_R_X5Y114_SLICE_X7Y114_BQ;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_T1 = 1'b1;
  assign RIOI3_X105Y171_OLOGIC_X1Y171_D1 = CLBLM_R_X103Y170_SLICE_X163Y170_AO5;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_D4 = CLBLM_L_X8Y108_SLICE_X11Y108_AQ;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_A1 = CLBLM_L_X8Y113_SLICE_X10Y113_CQ;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_A2 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_A3 = CLBLM_R_X7Y113_SLICE_X8Y113_AQ;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_A4 = CLBLM_R_X7Y114_SLICE_X8Y114_A5Q;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_D5 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_A6 = CLBLL_L_X4Y112_SLICE_X4Y112_CO5;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_D1 = CLBLM_R_X13Y112_SLICE_X18Y112_AQ;
  assign RIOI3_X105Y171_OLOGIC_X1Y171_T1 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_B1 = CLBLM_R_X5Y109_SLICE_X7Y109_AQ;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_B2 = CLBLM_R_X7Y113_SLICE_X8Y113_BQ;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_B4 = CLBLM_L_X10Y117_SLICE_X12Y117_A5Q;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_B5 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_B6 = CLBLL_L_X4Y112_SLICE_X4Y112_CO5;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_T1 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_C2 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_C3 = CLBLM_R_X7Y107_SLICE_X8Y107_CQ;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_C4 = CLBLM_R_X7Y113_SLICE_X8Y113_BQ;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_C5 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_C6 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_D1 = CLBLM_L_X10Y111_SLICE_X13Y111_CQ;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_T1 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_D2 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_D3 = CLBLM_R_X7Y113_SLICE_X8Y113_DQ;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_D4 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_D5 = CLBLM_L_X8Y113_SLICE_X11Y113_AQ;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_D6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_A3 = CLBLL_L_X4Y114_SLICE_X4Y114_AQ;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_B4 = 1'b1;
  assign LIOI3_X0Y161_OLOGIC_X0Y162_D1 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_B5 = CLBLL_L_X4Y116_SLICE_X4Y116_BO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_B6 = CLBLM_R_X13Y117_SLICE_X18Y117_BQ;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_B2 = 1'b1;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_B3 = CLBLM_R_X11Y110_SLICE_X15Y110_BQ;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_C4 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_C5 = CLBLM_R_X5Y116_SLICE_X6Y116_BQ;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign RIOB33_X105Y177_IOB_X1Y178_O = CLBLM_R_X103Y177_SLICE_X163Y177_AO5;
  assign RIOB33_X105Y177_IOB_X1Y177_O = CLBLM_R_X103Y177_SLICE_X163Y177_AO6;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_A1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_A2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_A3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_A4 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_A5 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_A6 = 1'b1;
  assign LIOI3_X0Y65_ILOGIC_X0Y66_D = LIOB33_X0Y65_IOB_X0Y66_I;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_B1 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_B2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_B3 = CLBLL_L_X4Y109_SLICE_X4Y109_BQ;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_B4 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_B5 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_B6 = CLBLL_L_X2Y114_SLICE_X0Y114_AO6;
  assign LIOI3_X0Y65_ILOGIC_X0Y65_D = LIOB33_X0Y65_IOB_X0Y65_I;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_C1 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_C2 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_C3 = CLBLL_L_X2Y107_SLICE_X1Y107_AO6;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_C4 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_C5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_C6 = CLBLL_L_X2Y110_SLICE_X0Y110_AO5;
  assign RIOI3_X105Y109_ILOGIC_X1Y110_D = RIOB33_X105Y109_IOB_X1Y110_I;
  assign RIOI3_X105Y109_ILOGIC_X1Y109_D = RIOB33_X105Y109_IOB_X1Y109_I;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_D1 = CLBLL_L_X2Y107_SLICE_X0Y107_AO5;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_D1 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_D2 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_D3 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_D4 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_D5 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_D6 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y138_D = RIOB33_X105Y137_IOB_X1Y138_I;
  assign RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y137_D = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_A1 = CLBLL_L_X2Y109_SLICE_X0Y109_AO5;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_A2 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_A3 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_A4 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_A5 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_A6 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_B1 = CLBLL_L_X2Y113_SLICE_X1Y113_DO6;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_B2 = CLBLL_L_X2Y114_SLICE_X1Y114_BO6;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_B3 = CLBLM_R_X3Y113_SLICE_X3Y113_DO6;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_B4 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_B5 = CLBLL_L_X4Y109_SLICE_X4Y109_CO6;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_B6 = CLBLL_L_X2Y112_SLICE_X1Y112_CO6;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_C1 = CLBLL_L_X4Y109_SLICE_X4Y109_BQ;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_C2 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_C3 = CLBLM_L_X10Y114_SLICE_X13Y114_AQ;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_C4 = CLBLM_R_X3Y112_SLICE_X3Y112_BO5;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_C5 = CLBLM_R_X3Y112_SLICE_X2Y112_AO5;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_C6 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_A1 = CLBLM_R_X7Y111_SLICE_X8Y111_CQ;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_A2 = CLBLM_L_X8Y114_SLICE_X10Y114_CQ;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_A3 = CLBLM_R_X7Y117_SLICE_X9Y117_DQ;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_A4 = CLBLM_R_X7Y115_SLICE_X8Y115_BQ;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_D1 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_D2 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_D3 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_D4 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_D5 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_D6 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_A5 = CLBLM_L_X10Y112_SLICE_X12Y112_BQ;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_A6 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_B2 = CLBLM_R_X7Y114_SLICE_X9Y114_BQ;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_B3 = CLBLM_R_X5Y113_SLICE_X7Y113_BQ;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_B4 = CLBLM_R_X11Y115_SLICE_X14Y115_AQ;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_B5 = CLBLL_L_X4Y112_SLICE_X4Y112_CO5;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_B6 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_C1 = CLBLM_R_X7Y114_SLICE_X9Y114_AO6;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_C2 = CLBLM_L_X10Y114_SLICE_X13Y114_BQ;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_C3 = CLBLM_R_X5Y116_SLICE_X6Y116_CQ;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_C4 = CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_C5 = CLBLM_L_X12Y112_SLICE_X17Y112_BQ;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_C6 = CLBLL_L_X4Y116_SLICE_X4Y116_BO6;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_D1 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_D2 = CLBLM_L_X8Y113_SLICE_X10Y113_CQ;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_D3 = CLBLM_R_X7Y111_SLICE_X8Y111_BQ;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_D4 = CLBLM_R_X7Y112_SLICE_X9Y112_AQ;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_D5 = CLBLM_R_X7Y110_SLICE_X9Y110_AQ;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_D6 = CLBLM_R_X5Y113_SLICE_X6Y113_BQ;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_A1 = CLBLM_R_X7Y116_SLICE_X8Y116_DO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_A2 = CLBLM_L_X10Y104_SLICE_X12Y104_AQ;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_A3 = CLBLM_R_X5Y114_SLICE_X6Y114_AQ;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_A4 = CLBLM_R_X3Y110_SLICE_X3Y110_AO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_A6 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_B2 = CLBLM_R_X7Y114_SLICE_X8Y114_BQ;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_B3 = CLBLL_L_X4Y112_SLICE_X4Y112_CO5;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_B4 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_B5 = CLBLM_R_X5Y113_SLICE_X7Y113_BQ;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_B6 = CLBLM_L_X10Y115_SLICE_X12Y115_CQ;
  assign RIOB33_X105Y185_IOB_X1Y186_O = CLBLM_L_X12Y111_SLICE_X16Y111_AQ;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_C2 = CLBLM_R_X7Y111_SLICE_X9Y111_CQ;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_C3 = CLBLM_R_X7Y117_SLICE_X9Y117_BQ;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_C4 = CLBLM_L_X8Y113_SLICE_X11Y113_CO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_C6 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_D1 = CLBLL_L_X4Y110_SLICE_X4Y110_BQ;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_D2 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_D3 = CLBLM_R_X7Y114_SLICE_X9Y114_DO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_D4 = CLBLM_L_X12Y108_SLICE_X16Y108_AQ;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_D5 = CLBLM_L_X8Y115_SLICE_X10Y115_DO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_D6 = CLBLM_R_X5Y113_SLICE_X7Y113_DO6;
  assign RIOB33_X105Y185_IOB_X1Y185_O = CLBLM_L_X8Y110_SLICE_X10Y110_CO5;
  assign CLBLM_L_X10Y114_SLICE_X13Y114_C5 = 1'b1;
  assign RIOB33_X105Y179_IOB_X1Y180_O = CLBLM_R_X13Y110_SLICE_X18Y110_DO6;
  assign RIOB33_X105Y179_IOB_X1Y179_O = CLBLM_R_X13Y117_SLICE_X18Y117_AO5;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_A3 = CLBLL_L_X4Y114_SLICE_X4Y114_AQ;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_A5 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign RIOB33_X105Y169_IOB_X1Y170_O = CLBLM_R_X103Y170_SLICE_X163Y170_AO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_A1 = CLBLL_L_X2Y113_SLICE_X0Y113_DO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_A2 = CLBLM_R_X3Y113_SLICE_X2Y113_BO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_A3 = CLBLL_L_X2Y113_SLICE_X1Y113_CO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_A4 = CLBLL_L_X2Y113_SLICE_X0Y113_BO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_A5 = CLBLL_L_X2Y112_SLICE_X0Y112_BO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_A6 = CLBLL_L_X2Y113_SLICE_X0Y113_CO6;
  assign RIOB33_X105Y169_IOB_X1Y169_O = CLBLM_R_X103Y169_SLICE_X163Y169_AO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_B1 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_B2 = CLBLL_L_X2Y114_SLICE_X0Y114_AO5;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_B3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_B4 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_B5 = LIOB33_X0Y69_IOB_X0Y70_I;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_B6 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_C1 = CLBLL_L_X2Y114_SLICE_X0Y114_AO5;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_C2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_C3 = CLBLL_L_X2Y112_SLICE_X1Y112_DO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_C4 = LIOB33_X0Y53_IOB_X0Y54_I;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_C5 = CLBLM_R_X5Y115_SLICE_X6Y115_CQ;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_C6 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_B2 = CLBLL_L_X4Y114_SLICE_X4Y114_BQ;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_B3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_D1 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_D2 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_D3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_D4 = CLBLM_R_X3Y116_SLICE_X3Y116_AO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_D5 = CLBLM_L_X10Y114_SLICE_X13Y114_AQ;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_D6 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_B4 = CLBLL_L_X4Y111_SLICE_X4Y111_CQ;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_A1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_A2 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_A3 = CLBLL_L_X2Y114_SLICE_X0Y114_AO5;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_A4 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_A5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_A6 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_C2 = CLBLL_L_X4Y114_SLICE_X4Y114_CQ;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_B1 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_B2 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_B3 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_B4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_B5 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_B6 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_C3 = CLBLM_R_X5Y112_SLICE_X7Y112_CQ;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_C1 = CLBLM_R_X3Y115_SLICE_X3Y115_AO6;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_C2 = CLBLL_L_X2Y114_SLICE_X0Y114_AO5;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_C3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_C4 = CLBLL_L_X2Y112_SLICE_X0Y112_AO6;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_C5 = LIOB33_X0Y59_IOB_X0Y59_I;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_C6 = CLBLM_R_X3Y114_SLICE_X2Y114_BQ;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_C5 = CLBLL_L_X4Y113_SLICE_X5Y113_DO6;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_D1 = CLBLL_L_X4Y117_SLICE_X4Y117_CQ;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_C6 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_D1 = CLBLL_L_X2Y113_SLICE_X1Y113_AO6;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_D2 = CLBLL_L_X2Y107_SLICE_X1Y107_AO6;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_D3 = CLBLL_L_X2Y112_SLICE_X0Y112_CO6;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_D4 = CLBLL_L_X2Y113_SLICE_X1Y113_CO6;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_D5 = CLBLL_L_X4Y114_SLICE_X4Y114_AQ;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_D6 = CLBLL_L_X4Y110_SLICE_X5Y110_AQ;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_A2 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_A3 = CLBLM_R_X7Y115_SLICE_X9Y115_AQ;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_A4 = CLBLL_L_X4Y116_SLICE_X4Y116_BO6;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_A5 = CLBLM_R_X7Y115_SLICE_X8Y115_AQ;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_A6 = CLBLM_L_X10Y114_SLICE_X12Y114_BQ;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_AX = CLBLM_R_X7Y115_SLICE_X9Y115_CO5;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_B1 = CLBLM_R_X7Y117_SLICE_X9Y117_A5Q;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_B2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_B3 = CLBLM_R_X7Y109_SLICE_X9Y109_DQ;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_B4 = CLBLM_L_X12Y112_SLICE_X17Y112_BQ;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_B6 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_A1 = CLBLL_L_X4Y112_SLICE_X4Y112_CO5;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_A2 = CLBLL_L_X4Y106_SLICE_X5Y106_BQ;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_A3 = CLBLM_R_X5Y105_SLICE_X7Y105_AQ;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_A4 = CLBLM_R_X7Y105_SLICE_X9Y105_AQ;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_A6 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_C1 = CLBLL_L_X4Y110_SLICE_X4Y110_BQ;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_C2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_B1 = CLBLM_R_X7Y105_SLICE_X8Y105_CQ;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_B2 = CLBLM_R_X5Y105_SLICE_X7Y105_BQ;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_B3 = CLBLM_R_X5Y106_SLICE_X7Y106_BO5;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_B4 = CLBLM_L_X10Y113_SLICE_X13Y113_AQ;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_B6 = CLBLM_R_X5Y107_SLICE_X7Y107_DO6;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_C1 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_C4 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_C2 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_C3 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_C4 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_C5 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_C5 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_C6 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_D1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_D2 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_C6 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_A2 = CLBLM_R_X3Y109_SLICE_X2Y109_AQ;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_D3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_D1 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_D2 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_D3 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_D4 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_D5 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_D6 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_A6 = CLBLM_R_X7Y114_SLICE_X8Y114_A5Q;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_D5 = CLBLM_R_X7Y110_SLICE_X8Y110_AQ;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_B1 = CLBLM_R_X5Y115_SLICE_X7Y115_AQ;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_B2 = CLBLM_R_X7Y115_SLICE_X8Y115_BQ;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_A1 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_A2 = CLBLM_R_X5Y107_SLICE_X7Y107_AQ;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_A3 = CLBLM_R_X5Y105_SLICE_X6Y105_AQ;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_A4 = CLBLL_L_X4Y107_SLICE_X4Y107_DQ;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_A6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_C1 = CLBLM_R_X7Y112_SLICE_X8Y112_C5Q;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_C2 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_B2 = CLBLL_L_X4Y106_SLICE_X5Y106_BQ;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_B4 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_B5 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_B6 = CLBLM_R_X5Y107_SLICE_X6Y107_BQ;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_D1 = CLBLM_R_X11Y114_SLICE_X14Y114_BQ;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_D2 = CLBLM_L_X12Y113_SLICE_X17Y113_AQ;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_C1 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_C2 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_C3 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_C4 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_C5 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_C6 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_D3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_D4 = CLBLM_R_X5Y116_SLICE_X7Y116_AQ;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_D5 = CLBLM_L_X8Y118_SLICE_X10Y118_AQ;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_D6 = 1'b1;
  assign LIOI3_X0Y189_OLOGIC_X0Y190_D1 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_D1 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_D2 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_D3 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_D4 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_D5 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_D6 = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_D1 = CLBLM_R_X11Y115_SLICE_X15Y115_B5Q;
  assign LIOI3_X0Y189_OLOGIC_X0Y190_T1 = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_D1 = CLBLM_R_X3Y115_SLICE_X2Y115_AQ;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_D1 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_D5 = 1'b1;
  assign LIOI3_X0Y189_OLOGIC_X0Y189_D1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X12Y115_SLICE_X17Y115_D6 = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_T1 = 1'b1;
  assign RIOI3_X105Y173_OLOGIC_X1Y174_D1 = CLBLM_R_X103Y174_SLICE_X163Y174_AO6;
  assign LIOI3_X0Y189_OLOGIC_X0Y189_T1 = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_D1 = CLBLL_L_X4Y113_SLICE_X4Y113_BQ;
  assign RIOB33_X105Y181_IOB_X1Y182_O = CLBLM_L_X12Y114_SLICE_X16Y114_DO6;
  assign RIOB33_X105Y181_IOB_X1Y181_O = CLBLM_R_X13Y110_SLICE_X18Y110_DO5;
  assign RIOI3_X105Y173_OLOGIC_X1Y174_T1 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_D2 = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_T1 = 1'b1;
  assign RIOI3_X105Y173_OLOGIC_X1Y173_D1 = CLBLM_R_X103Y173_SLICE_X163Y173_AO5;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_D1 = CLBLM_L_X8Y119_SLICE_X10Y119_AQ;
  assign RIOI3_X105Y173_OLOGIC_X1Y173_T1 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_D3 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_D1 = CLBLM_L_X8Y110_SLICE_X10Y110_CO5;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_D1 = CLBLM_L_X8Y119_SLICE_X10Y119_AO5;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_T1 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_D4 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_D1 = CLBLM_L_X8Y110_SLICE_X10Y110_CO6;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_A1 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_A2 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_A3 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_A4 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_A5 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_A6 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_T1 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_B1 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_B2 = CLBLL_L_X2Y114_SLICE_X0Y114_AO5;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_B3 = CLBLM_R_X3Y115_SLICE_X3Y115_AO6;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_B4 = LIOB33_X0Y71_IOB_X0Y71_I;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_B5 = LIOB33_X0Y55_IOB_X0Y55_I;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_B6 = CLBLL_L_X2Y109_SLICE_X0Y109_AO5;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_C5 = CLBLM_L_X10Y117_SLICE_X13Y117_DO6;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_C4 = CLBLM_L_X10Y119_SLICE_X12Y119_CO6;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_D5 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_C1 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_C2 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_C3 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_C4 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_C5 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_C6 = 1'b1;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_C6 = CLBLM_L_X10Y117_SLICE_X13Y117_BO5;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_D1 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_D2 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_D3 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_D4 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_D5 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X0Y114_D6 = 1'b1;
  assign CLBLM_L_X12Y115_SLICE_X16Y115_B5 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X19Y118_D6 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_A1 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_A2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_A3 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_A4 = CLBLL_L_X2Y114_SLICE_X0Y114_AO5;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_A5 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_A6 = 1'b1;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_D1 = CLBLM_R_X11Y116_SLICE_X14Y116_BQ;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_B1 = LIOB33_X0Y53_IOB_X0Y54_I;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_B2 = CLBLL_L_X2Y114_SLICE_X1Y114_AO5;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_B3 = CLBLM_R_X5Y115_SLICE_X6Y115_CQ;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_B4 = LIOB33_X0Y69_IOB_X0Y70_I;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_B5 = CLBLL_L_X2Y114_SLICE_X1Y114_AO6;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_B6 = CLBLL_L_X2Y113_SLICE_X1Y113_AO5;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_C1 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_C2 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_C3 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_C4 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_C5 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_C6 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_D1 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_D2 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_D3 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_D4 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_D5 = 1'b1;
  assign CLBLL_L_X2Y114_SLICE_X1Y114_D6 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_A1 = CLBLM_R_X7Y116_SLICE_X9Y116_BO5;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_A2 = CLBLM_R_X5Y115_SLICE_X6Y115_BQ;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_A3 = CLBLM_R_X7Y116_SLICE_X9Y116_AQ;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_A5 = CLBLM_R_X7Y132_SLICE_X9Y132_AO6;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_A6 = CLBLM_L_X8Y112_SLICE_X10Y112_AQ;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_B1 = CLBLM_R_X7Y116_SLICE_X9Y116_DO6;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_B2 = CLBLM_R_X7Y117_SLICE_X9Y117_A5Q;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_B3 = CLBLM_R_X7Y117_SLICE_X9Y117_AQ;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_B4 = CLBLM_R_X7Y117_SLICE_X9Y117_BQ;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_B5 = CLBLM_R_X5Y116_SLICE_X7Y116_AQ;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_B6 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_A1 = CLBLM_L_X8Y114_SLICE_X11Y114_B5Q;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_A2 = CLBLM_L_X10Y106_SLICE_X13Y106_CQ;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_A3 = CLBLM_R_X5Y106_SLICE_X7Y106_AQ;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_A5 = CLBLM_R_X7Y106_SLICE_X9Y106_AQ;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_A6 = CLBLM_L_X10Y104_SLICE_X12Y104_BO6;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_C1 = CLBLL_L_X4Y108_SLICE_X5Y108_AO6;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_C2 = CLBLM_R_X7Y114_SLICE_X8Y114_A5Q;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_C3 = CLBLM_L_X8Y118_SLICE_X10Y118_AQ;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_B1 = CLBLM_R_X7Y105_SLICE_X9Y105_CQ;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_B2 = CLBLM_R_X5Y105_SLICE_X7Y105_BQ;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_B3 = CLBLM_R_X7Y107_SLICE_X8Y107_DO6;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_B4 = CLBLM_R_X5Y106_SLICE_X6Y106_BQ;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_B5 = CLBLM_L_X8Y106_SLICE_X10Y106_BQ;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_B6 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_D1 = CLBLM_R_X5Y116_SLICE_X7Y116_BQ;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_C2 = CLBLM_L_X8Y106_SLICE_X11Y106_A5Q;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_C3 = CLBLL_L_X4Y107_SLICE_X4Y107_BO5;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_C4 = CLBLM_R_X3Y108_SLICE_X2Y108_DO6;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_C5 = CLBLM_R_X5Y106_SLICE_X7Y106_DO6;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_C6 = CLBLM_R_X3Y110_SLICE_X2Y110_DO6;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_D3 = CLBLM_R_X5Y115_SLICE_X7Y115_AQ;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_D4 = CLBLM_R_X5Y116_SLICE_X6Y116_CQ;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_A2 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_A3 = CLBLM_L_X8Y115_SLICE_X11Y115_BQ;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_A4 = CLBLM_L_X10Y116_SLICE_X12Y116_DO6;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_A5 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_D1 = CLBLM_L_X8Y104_SLICE_X11Y104_AQ;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_D2 = CLBLM_R_X5Y107_SLICE_X7Y107_CO5;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_D3 = CLBLM_R_X3Y109_SLICE_X2Y109_CO6;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_D4 = CLBLL_L_X4Y117_SLICE_X4Y117_CQ;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_D5 = CLBLL_L_X2Y111_SLICE_X1Y111_DO6;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_D6 = CLBLM_R_X3Y110_SLICE_X3Y110_DO6;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_A6 = CLBLM_R_X7Y117_SLICE_X8Y117_AQ;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_B2 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_B3 = CLBLM_R_X7Y116_SLICE_X8Y116_AQ;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_B4 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_A1 = CLBLM_R_X7Y108_SLICE_X8Y108_CQ;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_A2 = CLBLM_R_X7Y110_SLICE_X8Y110_BQ;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_A3 = CLBLM_R_X5Y106_SLICE_X6Y106_AQ;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_A4 = CLBLL_L_X4Y112_SLICE_X4Y112_CO5;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_A5 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_C1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_C2 = CLBLM_R_X7Y116_SLICE_X8Y116_CQ;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_C3 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_B1 = CLBLM_L_X10Y113_SLICE_X13Y113_AQ;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_B2 = CLBLM_R_X5Y106_SLICE_X6Y106_BQ;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_B3 = CLBLM_R_X7Y109_SLICE_X9Y109_CQ;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_B5 = CLBLM_R_X5Y106_SLICE_X7Y106_BO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_B6 = CLBLM_R_X5Y106_SLICE_X7Y106_BO5;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_D1 = CLBLM_R_X5Y116_SLICE_X6Y116_AO5;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_D2 = CLBLM_R_X11Y117_SLICE_X15Y117_AQ;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_C1 = CLBLM_R_X5Y106_SLICE_X7Y106_BO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_C2 = CLBLM_R_X5Y106_SLICE_X6Y106_CQ;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_C3 = CLBLM_L_X10Y113_SLICE_X13Y113_AQ;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_C5 = CLBLL_L_X4Y111_SLICE_X4Y111_AQ;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_C6 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_D3 = CLBLM_L_X8Y118_SLICE_X10Y118_AQ;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_D4 = CLBLM_R_X7Y114_SLICE_X8Y114_A5Q;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_D5 = CLBLM_R_X7Y118_SLICE_X9Y118_BO5;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_D6 = CLBLM_L_X10Y117_SLICE_X13Y117_CO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_D1 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_D2 = CLBLM_R_X5Y106_SLICE_X6Y106_AQ;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_D3 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_D4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_D6 = CLBLM_R_X7Y107_SLICE_X9Y107_CQ;
  assign RIOB33_X105Y183_IOB_X1Y183_O = CLBLM_L_X12Y114_SLICE_X16Y114_DO5;
  assign RIOB33_X105Y183_IOB_X1Y184_O = CLBLM_L_X8Y110_SLICE_X10Y110_CO6;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_C1 = 1'b1;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_C2 = 1'b1;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_A4 = 1'b1;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_A5 = CLBLM_L_X10Y110_SLICE_X12Y110_AQ;
  assign CLBLM_R_X11Y113_SLICE_X15Y113_A6 = CLBLM_R_X7Y115_SLICE_X9Y115_DO6;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_A1 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_A2 = CLBLM_L_X12Y115_SLICE_X16Y115_AQ;
  assign LIOI3_X0Y185_OLOGIC_X0Y186_T1 = 1'b1;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_A4 = CLBLM_L_X12Y118_SLICE_X16Y118_AQ;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_D1 = RIOB33_X105Y145_IOB_X1Y145_I;
  assign LIOI3_X0Y185_OLOGIC_X0Y185_D1 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_B2 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_B6 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_T1 = 1'b1;
  assign LIOI3_X0Y185_OLOGIC_X0Y185_T1 = 1'b1;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_A1 = CLBLM_L_X10Y112_SLICE_X12Y112_C5Q;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_A3 = CLBLM_R_X7Y117_SLICE_X9Y117_AQ;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_A5 = CLBLM_L_X12Y112_SLICE_X16Y112_B5Q;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_A6 = CLBLM_L_X8Y109_SLICE_X11Y109_BQ;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_AX = CLBLM_R_X7Y117_SLICE_X9Y117_CO6;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_B2 = CLBLM_R_X7Y117_SLICE_X9Y117_BQ;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_B3 = CLBLM_R_X7Y132_SLICE_X9Y132_AO6;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_B4 = CLBLM_R_X5Y116_SLICE_X7Y116_AQ;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_B5 = CLBLM_R_X7Y117_SLICE_X9Y117_CO5;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_B6 = CLBLM_R_X7Y112_SLICE_X8Y112_CQ;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_A1 = CLBLM_R_X7Y107_SLICE_X8Y107_CQ;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_A2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_A3 = CLBLM_R_X5Y107_SLICE_X7Y107_AQ;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_A4 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_A6 = CLBLL_L_X4Y116_SLICE_X5Y116_B5Q;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_C1 = CLBLM_R_X7Y132_SLICE_X9Y132_AO6;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_C2 = CLBLM_L_X8Y110_SLICE_X11Y110_DQ;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_B2 = CLBLM_R_X3Y110_SLICE_X3Y110_DO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_B3 = CLBLM_R_X5Y105_SLICE_X7Y105_AQ;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_B4 = CLBLM_R_X5Y108_SLICE_X7Y108_CO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_B5 = CLBLM_L_X8Y107_SLICE_X10Y107_AQ;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_B6 = 1'b1;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_C1 = CLBLM_L_X8Y106_SLICE_X11Y106_A5Q;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_C2 = CLBLM_L_X8Y109_SLICE_X10Y109_CQ;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_C3 = CLBLM_R_X5Y109_SLICE_X6Y109_CQ;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_C4 = CLBLM_R_X7Y115_SLICE_X8Y115_DQ;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_C5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_C6 = 1'b1;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_D3 = CLBLM_R_X7Y117_SLICE_X9Y117_DQ;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_D4 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_A1 = CLBLM_L_X8Y111_SLICE_X10Y111_A5Q;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_A2 = CLBLM_R_X7Y117_SLICE_X8Y117_BQ;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_A3 = CLBLM_L_X10Y116_SLICE_X12Y116_DO6;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_A4 = 1'b1;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_D1 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_D2 = CLBLM_R_X7Y105_SLICE_X9Y105_CQ;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_D3 = CLBLM_R_X7Y107_SLICE_X8Y107_DO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_D4 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_D5 = CLBLM_L_X8Y106_SLICE_X10Y106_BQ;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_D6 = 1'b1;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_B2 = 1'b1;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_B3 = CLBLM_L_X10Y116_SLICE_X12Y116_DO6;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_B4 = CLBLL_L_X4Y115_SLICE_X5Y115_BQ;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_B5 = CLBLM_L_X8Y116_SLICE_X11Y116_AQ;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_B6 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_A1 = CLBLL_L_X4Y108_SLICE_X5Y108_AO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_A2 = CLBLL_L_X4Y110_SLICE_X4Y110_AQ;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_A3 = CLBLM_R_X5Y107_SLICE_X6Y107_AQ;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_A4 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_A6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_C1 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_C2 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_B1 = CLBLM_R_X7Y105_SLICE_X8Y105_CQ;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_B2 = CLBLM_R_X5Y107_SLICE_X6Y107_BQ;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_B3 = CLBLL_L_X4Y110_SLICE_X4Y110_AQ;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_B4 = CLBLL_L_X4Y109_SLICE_X5Y109_AQ;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_B5 = CLBLM_L_X8Y106_SLICE_X10Y106_BQ;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_C4 = CLBLM_L_X10Y112_SLICE_X12Y112_C5Q;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_C5 = CLBLM_L_X12Y112_SLICE_X16Y112_B5Q;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_C1 = CLBLM_R_X7Y111_SLICE_X9Y111_DO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_C2 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_C3 = CLBLM_R_X7Y111_SLICE_X8Y111_DQ;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_C5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_C6 = CLBLL_L_X4Y107_SLICE_X4Y107_DQ;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_C6 = 1'b1;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_D3 = 1'b1;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_D4 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_D6 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_D1 = CLBLM_L_X8Y106_SLICE_X10Y106_BQ;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_D2 = CLBLM_L_X10Y104_SLICE_X12Y104_BO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_D3 = CLBLM_R_X5Y107_SLICE_X6Y107_DQ;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_D4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_D5 = CLBLM_L_X8Y114_SLICE_X11Y114_B5Q;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_D6 = CLBLM_R_X5Y105_SLICE_X7Y105_BQ;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_D1 = CLBLM_R_X7Y115_SLICE_X8Y115_D5Q;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_D2 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_D3 = CLBLM_R_X7Y115_SLICE_X8Y115_B5Q;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_D4 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_D5 = CLBLM_R_X5Y115_SLICE_X6Y115_DO6;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_D6 = CLBLM_R_X5Y116_SLICE_X6Y116_D5Q;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_B4 = 1'b1;
  assign RIOI3_SING_X105Y149_ILOGIC_X1Y149_D = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_B5 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_A1 = CLBLM_R_X7Y118_SLICE_X8Y118_CQ;
  assign LIOI3_X0Y191_OLOGIC_X0Y192_D1 = LIOB33_X0Y51_IOB_X0Y52_I;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_A3 = CLBLM_L_X8Y118_SLICE_X10Y118_AQ;
  assign CLBLM_R_X13Y118_SLICE_X18Y118_B6 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_A4 = CLBLM_L_X10Y119_SLICE_X12Y119_AQ;
  assign LIOI3_X0Y191_OLOGIC_X0Y192_T1 = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_D1 = CLBLL_L_X52Y126_SLICE_X78Y126_AO6;
  assign LIOI3_X0Y191_OLOGIC_X0Y191_D1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_T1 = 1'b1;
  assign RIOI3_X105Y175_OLOGIC_X1Y176_D1 = CLBLM_R_X103Y174_SLICE_X163Y174_AO5;
  assign LIOI3_X0Y191_OLOGIC_X0Y191_T1 = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_D1 = CLBLM_R_X5Y109_SLICE_X6Y109_CQ;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_C4 = 1'b1;
  assign RIOI3_X105Y175_OLOGIC_X1Y176_T1 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_C5 = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_T1 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_C6 = 1'b1;
  assign RIOI3_X105Y175_OLOGIC_X1Y175_D1 = CLBLM_R_X13Y118_SLICE_X18Y118_AO6;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_B4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_D1 = LIOB33_X0Y57_IOB_X0Y57_I;
  assign RIOI3_X105Y175_OLOGIC_X1Y175_T1 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_B5 = CLBLM_R_X5Y115_SLICE_X6Y115_CQ;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_C2 = CLBLM_L_X8Y109_SLICE_X11Y109_CQ;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_B6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_T1 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_C3 = CLBLM_R_X7Y106_SLICE_X9Y106_CQ;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_D1 = CLBLM_L_X12Y117_SLICE_X17Y117_AQ;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_C4 = CLBLM_R_X5Y115_SLICE_X7Y115_CO6;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_D1 = LIOB33_X0Y55_IOB_X0Y55_I;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_T1 = 1'b1;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_A2 = CLBLM_R_X7Y111_SLICE_X8Y111_BQ;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_A3 = CLBLM_R_X7Y118_SLICE_X9Y118_AQ;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_A4 = 1'b1;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_A5 = CLBLM_L_X10Y117_SLICE_X13Y117_AO5;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_A6 = CLBLM_R_X7Y118_SLICE_X9Y118_CO6;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_D2 = 1'b1;
  assign LIOB33_X0Y101_IOB_X0Y101_O = CLBLL_L_X2Y107_SLICE_X0Y107_AO6;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_B1 = CLBLM_R_X7Y117_SLICE_X8Y117_BQ;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_B2 = CLBLM_R_X7Y118_SLICE_X8Y118_AQ;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_B3 = CLBLM_L_X10Y117_SLICE_X13Y117_AO5;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_B4 = CLBLM_R_X7Y118_SLICE_X8Y118_BQ;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_B5 = CLBLM_R_X7Y118_SLICE_X9Y118_AQ;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_B6 = 1'b1;
  assign LIOB33_X0Y101_IOB_X0Y102_O = CLBLL_L_X2Y106_SLICE_X0Y106_BO5;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_C4 = CLBLM_R_X7Y116_SLICE_X8Y116_AQ;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_T1 = 1'b1;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_A1 = CLBLM_R_X5Y110_SLICE_X6Y110_B5Q;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_A2 = 1'b1;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_A3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_A4 = CLBLM_R_X7Y108_SLICE_X8Y108_DO5;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_A6 = CLBLM_R_X5Y107_SLICE_X6Y107_CQ;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_D5 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_D6 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_B1 = CLBLM_R_X7Y115_SLICE_X8Y115_DQ;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_B2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_B3 = CLBLM_L_X8Y106_SLICE_X11Y106_A5Q;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_B4 = CLBLM_L_X8Y109_SLICE_X10Y109_CQ;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_B6 = CLBLM_R_X5Y109_SLICE_X6Y109_CQ;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_C1 = CLBLM_R_X5Y109_SLICE_X7Y109_BQ;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_D1 = CLBLM_R_X5Y117_SLICE_X7Y117_AQ;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_C2 = CLBLM_R_X5Y109_SLICE_X7Y109_DQ;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_C3 = CLBLM_R_X5Y107_SLICE_X7Y107_B5Q;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_C4 = CLBLM_L_X10Y104_SLICE_X12Y104_BO6;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_C5 = CLBLM_R_X5Y109_SLICE_X7Y109_B5Q;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_D2 = CLBLM_R_X11Y112_SLICE_X14Y112_BQ;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_C6 = CLBLM_R_X5Y108_SLICE_X7Y108_BO6;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_D3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_A2 = CLBLM_R_X7Y118_SLICE_X9Y118_BO6;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_A3 = CLBLM_L_X8Y113_SLICE_X10Y113_AQ;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_D1 = CLBLM_L_X10Y108_SLICE_X12Y108_CQ;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_D4 = CLBLM_L_X8Y107_SLICE_X11Y107_AQ;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_D2 = CLBLM_R_X7Y107_SLICE_X9Y107_CQ;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_D3 = CLBLM_R_X5Y108_SLICE_X6Y108_DO6;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_D4 = CLBLL_L_X4Y112_SLICE_X5Y112_DO6;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_D5 = CLBLM_R_X5Y108_SLICE_X7Y108_AQ;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_D6 = CLBLM_R_X5Y105_SLICE_X6Y105_BQ;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_D5 = 1'b1;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_B2 = CLBLM_R_X7Y118_SLICE_X9Y118_BO6;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_D6 = 1'b1;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_A1 = CLBLM_R_X7Y108_SLICE_X9Y108_BO5;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_A2 = CLBLM_R_X5Y107_SLICE_X7Y107_DO5;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_A3 = CLBLM_L_X8Y110_SLICE_X10Y110_BQ;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_A4 = CLBLM_R_X5Y106_SLICE_X6Y106_BQ;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_A5 = CLBLM_L_X10Y113_SLICE_X13Y113_CQ;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_A6 = CLBLM_R_X5Y106_SLICE_X6Y106_CQ;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_C1 = CLBLM_L_X10Y117_SLICE_X13Y117_CO6;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_C2 = CLBLM_R_X7Y118_SLICE_X8Y118_CQ;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_C3 = CLBLM_L_X10Y119_SLICE_X12Y119_AQ;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_B1 = CLBLL_L_X4Y108_SLICE_X5Y108_AO5;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_B2 = CLBLM_R_X3Y110_SLICE_X3Y110_AO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_B3 = CLBLM_R_X3Y111_SLICE_X2Y111_CO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_B4 = CLBLM_R_X3Y110_SLICE_X2Y110_DO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_B5 = CLBLL_L_X2Y110_SLICE_X1Y110_DO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_B6 = CLBLM_R_X5Y108_SLICE_X6Y108_CO6;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_D1 = CLBLM_R_X7Y117_SLICE_X8Y117_BQ;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_C1 = CLBLM_R_X5Y105_SLICE_X7Y105_BQ;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_C2 = CLBLM_R_X5Y107_SLICE_X7Y107_DO5;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_C3 = CLBLM_R_X5Y106_SLICE_X6Y106_BQ;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_C4 = CLBLM_L_X8Y110_SLICE_X10Y110_BQ;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_C5 = CLBLM_R_X7Y108_SLICE_X9Y108_BO5;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_C6 = CLBLM_R_X7Y108_SLICE_X9Y108_AQ;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_D2 = CLBLM_R_X11Y117_SLICE_X15Y117_AQ;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_D3 = CLBLM_R_X7Y118_SLICE_X8Y118_BQ;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_D4 = CLBLM_R_X7Y118_SLICE_X9Y118_AQ;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_D5 = CLBLM_R_X7Y118_SLICE_X8Y118_AQ;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_D6 = CLBLM_R_X7Y114_SLICE_X8Y114_A5Q;
  assign RIOI3_X105Y111_ILOGIC_X1Y112_D = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_D1 = 1'b1;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_D2 = CLBLM_R_X5Y106_SLICE_X6Y106_DQ;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_D3 = CLBLM_R_X7Y111_SLICE_X8Y111_DQ;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_D4 = CLBLM_R_X5Y107_SLICE_X6Y107_CQ;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_D5 = CLBLM_R_X5Y113_SLICE_X7Y113_BQ;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_D6 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_A5 = CLBLL_L_X4Y112_SLICE_X4Y112_CO5;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_A6 = 1'b1;
  assign LIOI3_X0Y71_ILOGIC_X0Y72_D = LIOB33_X0Y71_IOB_X0Y72_I;
  assign LIOI3_X0Y71_ILOGIC_X0Y71_D = LIOB33_X0Y71_IOB_X0Y71_I;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_B5 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_B6 = 1'b1;
  assign RIOI3_X105Y115_ILOGIC_X1Y116_D = RIOB33_X105Y115_IOB_X1Y116_I;
  assign RIOI3_X105Y115_ILOGIC_X1Y115_D = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_B1 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_B2 = CLBLM_L_X8Y109_SLICE_X10Y109_BQ;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_C4 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_C5 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_C6 = 1'b1;
  assign RIOI3_X105Y111_ILOGIC_X1Y111_D = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_D3 = 1'b1;
  assign LIOB33_X0Y103_IOB_X0Y104_O = CLBLL_L_X2Y106_SLICE_X0Y106_CO6;
  assign LIOB33_X0Y103_IOB_X0Y103_O = CLBLM_R_X3Y107_SLICE_X3Y107_BO6;
  assign RIOB33_X105Y189_IOB_X1Y190_O = CLBLM_R_X13Y113_SLICE_X19Y113_AQ;
  assign RIOB33_X105Y189_IOB_X1Y189_O = CLBLM_L_X10Y112_SLICE_X13Y112_AQ;
  assign RIOI3_X105Y153_OLOGIC_X1Y153_D1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_A1 = CLBLM_R_X7Y109_SLICE_X8Y109_CO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_A4 = CLBLL_L_X4Y106_SLICE_X5Y106_BQ;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_A5 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_A6 = CLBLM_R_X5Y113_SLICE_X7Y113_BQ;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_AX = CLBLM_R_X7Y106_SLICE_X9Y106_DO5;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_B1 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_B2 = CLBLM_R_X5Y109_SLICE_X7Y109_BQ;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_B4 = CLBLM_L_X8Y109_SLICE_X10Y109_BQ;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_B5 = CLBLM_R_X5Y109_SLICE_X7Y109_CO5;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_B6 = CLBLM_R_X5Y107_SLICE_X7Y107_CO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_BX = CLBLM_R_X5Y109_SLICE_X7Y109_CO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_C1 = CLBLM_L_X10Y104_SLICE_X12Y104_BO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_C2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_C3 = CLBLM_R_X5Y114_SLICE_X7Y114_B5Q;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_C4 = CLBLM_R_X5Y108_SLICE_X7Y108_BO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_C5 = CLBLM_R_X5Y109_SLICE_X7Y109_B5Q;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_C6 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_D1 = CLBLM_R_X5Y109_SLICE_X7Y109_CO5;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_D2 = CLBLM_R_X5Y107_SLICE_X7Y107_CO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_D3 = CLBLM_R_X5Y109_SLICE_X7Y109_DQ;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_D4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_D5 = CLBLM_L_X10Y111_SLICE_X13Y111_AQ;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_D6 = CLBLM_R_X5Y109_SLICE_X7Y109_BQ;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_A1 = CLBLM_R_X11Y117_SLICE_X15Y117_DQ;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_A3 = CLBLM_R_X5Y109_SLICE_X6Y109_AQ;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_A4 = CLBLM_R_X7Y109_SLICE_X9Y109_CQ;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_A5 = CLBLL_L_X4Y110_SLICE_X4Y110_AQ;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_A6 = CLBLM_R_X7Y105_SLICE_X8Y105_CQ;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_B1 = CLBLM_R_X5Y106_SLICE_X6Y106_DQ;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_B2 = CLBLM_R_X5Y109_SLICE_X6Y109_BQ;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_B3 = CLBLM_R_X11Y105_SLICE_X14Y105_C5Q;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_B4 = CLBLL_L_X4Y112_SLICE_X4Y112_CO5;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_B6 = 1'b1;
  assign RIOI3_X105Y153_OLOGIC_X1Y153_T1 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_C1 = CLBLM_R_X7Y112_SLICE_X8Y112_C5Q;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_C2 = CLBLM_R_X5Y107_SLICE_X7Y107_B5Q;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_C3 = CLBLM_R_X5Y109_SLICE_X7Y109_B5Q;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_C5 = CLBLM_R_X5Y109_SLICE_X7Y109_DQ;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_C6 = CLBLM_R_X5Y109_SLICE_X7Y109_BQ;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_D1 = CLBLL_L_X4Y108_SLICE_X4Y108_AQ;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_D2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_D3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_D4 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_D5 = CLBLM_R_X7Y110_SLICE_X8Y110_BQ;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_D6 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_C6 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_A1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_A2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_A3 = CLBLM_R_X5Y111_SLICE_X7Y111_BQ;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_A4 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign LIOI3_X0Y115_OLOGIC_X0Y116_T1 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_B1 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_B2 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_B3 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_B4 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_B5 = 1'b1;
  assign LIOB33_X0Y105_IOB_X0Y106_O = CLBLL_L_X2Y106_SLICE_X0Y106_AO5;
  assign LIOB33_X0Y105_IOB_X0Y105_O = CLBLL_L_X2Y106_SLICE_X0Y106_CO5;
  assign LIOI3_X0Y115_OLOGIC_X0Y115_D1 = CLBLM_R_X11Y110_SLICE_X14Y110_DQ;
  assign CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_CE = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_C4 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_C5 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_C6 = 1'b1;
  assign RIOB33_X105Y191_IOB_X1Y192_O = CLBLM_R_X13Y109_SLICE_X19Y109_AQ;
  assign RIOB33_X105Y191_IOB_X1Y191_O = CLBLM_R_X11Y115_SLICE_X14Y115_AQ;
  assign LIOI3_X0Y115_OLOGIC_X0Y115_T1 = 1'b1;
  assign LIOI3_X0Y195_OLOGIC_X0Y196_D1 = LIOB33_X0Y69_IOB_X0Y69_I;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_A1 = CLBLM_R_X5Y114_SLICE_X7Y114_B5Q;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_A2 = CLBLM_R_X11Y111_SLICE_X15Y111_BQ;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_A3 = CLBLM_R_X5Y110_SLICE_X7Y110_AQ;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_A4 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_A6 = CLBLL_L_X4Y113_SLICE_X5Y113_DO6;
  assign LIOI3_X0Y195_OLOGIC_X0Y196_T1 = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_D1 = CLBLL_L_X4Y116_SLICE_X5Y116_AQ;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_B1 = CLBLL_L_X4Y115_SLICE_X5Y115_CQ;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_B2 = CLBLM_R_X5Y111_SLICE_X7Y111_CQ;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_B4 = CLBLL_L_X4Y110_SLICE_X5Y110_AO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_D2 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_B5 = CLBLM_R_X5Y110_SLICE_X7Y110_CO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_B6 = 1'b1;
  assign LIOI3_X0Y195_OLOGIC_X0Y195_D1 = LIOB33_X0Y63_IOB_X0Y64_I;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_C1 = CLBLM_R_X5Y111_SLICE_X7Y111_AQ;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_C2 = CLBLM_R_X5Y115_SLICE_X7Y115_CO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_C3 = CLBLM_R_X5Y110_SLICE_X7Y110_BQ;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_C4 = CLBLM_L_X8Y110_SLICE_X11Y110_BO5;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_C5 = CLBLM_R_X5Y110_SLICE_X7Y110_B5Q;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_C6 = CLBLL_L_X4Y113_SLICE_X5Y113_BQ;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_T1 = 1'b1;
  assign RIOI3_X105Y177_OLOGIC_X1Y178_D1 = CLBLM_R_X103Y177_SLICE_X163Y177_AO5;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y195_OLOGIC_X0Y195_T1 = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_D1 = CLBLL_L_X4Y118_SLICE_X4Y118_A5Q;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_D6 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_D1 = CLBLM_R_X5Y111_SLICE_X7Y111_AQ;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_D2 = CLBLM_R_X3Y107_SLICE_X3Y107_CO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_D3 = CLBLM_R_X5Y115_SLICE_X7Y115_DO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_D4 = CLBLM_R_X5Y110_SLICE_X7Y110_BQ;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_D5 = CLBLM_R_X5Y110_SLICE_X7Y110_B5Q;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_D6 = CLBLL_L_X4Y113_SLICE_X5Y113_BQ;
  assign RIOI3_X105Y177_OLOGIC_X1Y178_T1 = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_T1 = 1'b1;
  assign RIOI3_X105Y177_OLOGIC_X1Y177_D1 = CLBLM_R_X103Y177_SLICE_X163Y177_AO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_A1 = CLBLM_R_X5Y105_SLICE_X7Y105_BQ;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_A2 = CLBLM_R_X5Y110_SLICE_X6Y110_DQ;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_A4 = CLBLM_L_X8Y113_SLICE_X10Y113_D5Q;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_A5 = CLBLM_R_X5Y108_SLICE_X6Y108_AO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_A6 = CLBLM_R_X7Y108_SLICE_X9Y108_AQ;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_D1 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_B1 = CLBLM_R_X5Y110_SLICE_X6Y110_CQ;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_B2 = CLBLM_R_X5Y117_SLICE_X7Y117_AQ;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_B4 = CLBLM_R_X5Y115_SLICE_X6Y115_BQ;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_B5 = CLBLL_L_X4Y107_SLICE_X4Y107_AQ;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_B6 = 1'b1;
  assign RIOI3_X105Y177_OLOGIC_X1Y177_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_T1 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_C1 = CLBLM_L_X10Y104_SLICE_X12Y104_BO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_C2 = CLBLM_R_X5Y110_SLICE_X6Y110_CQ;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_C3 = CLBLM_L_X8Y114_SLICE_X11Y114_B5Q;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_C4 = CLBLM_R_X5Y106_SLICE_X6Y106_BQ;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_C6 = CLBLM_L_X8Y119_SLICE_X10Y119_AQ;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_D1 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_D2 = CLBLM_R_X13Y107_SLICE_X19Y107_BQ;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_D3 = CLBLM_R_X5Y110_SLICE_X6Y110_DQ;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_D4 = CLBLL_L_X4Y113_SLICE_X5Y113_DO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_D5 = CLBLL_L_X4Y116_SLICE_X5Y116_B5Q;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_D6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_T1 = 1'b1;
  assign LIOB33_X0Y107_IOB_X0Y108_O = CLBLL_L_X2Y107_SLICE_X0Y107_AO5;
  assign LIOB33_X0Y107_IOB_X0Y107_O = CLBLM_R_X3Y106_SLICE_X2Y106_BO6;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_C6 = CLBLM_R_X7Y114_SLICE_X8Y114_A5Q;
  assign LIOI3_X0Y73_ILOGIC_X0Y74_D = LIOB33_X0Y73_IOB_X0Y74_I;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y73_ILOGIC_X0Y73_D = LIOB33_X0Y73_IOB_X0Y73_I;
  assign RIOI3_X105Y117_ILOGIC_X1Y118_D = RIOB33_X105Y117_IOB_X1Y118_I;
  assign RIOI3_X105Y117_ILOGIC_X1Y117_D = RIOB33_X105Y117_IOB_X1Y117_I;
  assign RIOB33_X105Y193_IOB_X1Y194_O = CLBLM_R_X11Y119_SLICE_X14Y119_AQ;
  assign RIOB33_X105Y193_IOB_X1Y193_O = CLBLM_L_X12Y118_SLICE_X16Y118_AQ;
  assign LIOB33_X0Y119_IOB_X0Y120_O = CLBLM_R_X13Y112_SLICE_X18Y112_AQ;
  assign LIOB33_X0Y119_IOB_X0Y119_O = CLBLM_L_X10Y111_SLICE_X13Y111_CQ;
  assign CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_I = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_A1 = CLBLM_R_X7Y118_SLICE_X8Y118_AQ;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_A2 = CLBLM_R_X5Y115_SLICE_X7Y115_CO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_A3 = CLBLM_R_X5Y111_SLICE_X7Y111_AQ;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_A5 = CLBLM_L_X8Y110_SLICE_X11Y110_BO5;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_A6 = CLBLM_R_X5Y111_SLICE_X6Y111_DO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_B1 = CLBLM_R_X5Y111_SLICE_X7Y111_DO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_B2 = CLBLM_R_X5Y111_SLICE_X7Y111_BQ;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_B4 = CLBLM_L_X12Y109_SLICE_X16Y109_AQ;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_B6 = CLBLM_R_X5Y108_SLICE_X7Y108_DO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_C1 = CLBLM_L_X8Y111_SLICE_X10Y111_DO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_C2 = CLBLM_R_X5Y111_SLICE_X7Y111_CQ;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_C3 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_C4 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_C6 = CLBLM_R_X5Y106_SLICE_X7Y106_AQ;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_D1 = CLBLM_L_X10Y111_SLICE_X12Y111_AQ;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_D2 = CLBLM_R_X7Y109_SLICE_X9Y109_DQ;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_D3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_D4 = CLBLM_R_X5Y111_SLICE_X6Y111_CQ;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_D5 = CLBLM_R_X5Y109_SLICE_X7Y109_AQ;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_D6 = CLBLL_L_X4Y106_SLICE_X5Y106_BQ;
  assign LIOI3_X0Y175_OLOGIC_X0Y175_D1 = RIOB33_X105Y127_IOB_X1Y127_I;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_A1 = CLBLM_R_X5Y116_SLICE_X6Y116_CQ;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_A2 = CLBLM_R_X7Y108_SLICE_X9Y108_AQ;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_A3 = CLBLM_R_X5Y111_SLICE_X6Y111_AQ;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_A4 = CLBLM_R_X7Y105_SLICE_X8Y105_CQ;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_A6 = CLBLL_L_X4Y110_SLICE_X4Y110_AQ;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_B1 = CLBLM_R_X7Y111_SLICE_X8Y111_DQ;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_B2 = CLBLM_R_X5Y111_SLICE_X6Y111_BQ;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_B4 = CLBLL_L_X4Y112_SLICE_X4Y112_CO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_B5 = CLBLL_L_X4Y116_SLICE_X4Y116_AQ;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_B6 = 1'b1;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_C1 = CLBLM_R_X5Y109_SLICE_X6Y109_AQ;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_C2 = CLBLM_R_X7Y111_SLICE_X9Y111_DO5;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_C4 = CLBLM_L_X10Y111_SLICE_X12Y111_AQ;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_C6 = 1'b1;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_D1 = CLBLM_R_X5Y111_SLICE_X7Y111_AQ;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_D2 = CLBLL_L_X4Y113_SLICE_X5Y113_BQ;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_D3 = 1'b1;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_D4 = CLBLM_R_X5Y110_SLICE_X7Y110_B5Q;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_D5 = 1'b1;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_D6 = CLBLM_R_X5Y110_SLICE_X7Y110_BQ;
  assign LIOI3_SING_X0Y100_OLOGIC_X0Y100_T1 = 1'b1;
  assign LIOI3_X0Y175_OLOGIC_X0Y175_T1 = 1'b1;
  assign LIOB33_X0Y109_IOB_X0Y110_O = CLBLM_R_X3Y106_SLICE_X2Y106_AO6;
  assign LIOB33_X0Y109_IOB_X0Y109_O = CLBLL_L_X2Y107_SLICE_X1Y107_AO5;
  assign RIOI3_SING_X105Y150_OLOGIC_X1Y150_D1 = LIOB33_X0Y75_IOB_X0Y75_I;
  assign RIOB33_X105Y195_IOB_X1Y196_O = CLBLM_L_X12Y117_SLICE_X16Y117_AQ;
  assign RIOB33_X105Y195_IOB_X1Y195_O = CLBLM_L_X12Y110_SLICE_X16Y110_AQ;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_D6 = CLBLM_L_X10Y117_SLICE_X12Y117_DO6;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_B5 = 1'b1;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_C4 = CLBLM_R_X13Y108_SLICE_X19Y108_BQ;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_B6 = 1'b1;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_A1 = CLBLM_R_X7Y105_SLICE_X8Y105_BO5;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_A2 = CLBLM_R_X3Y110_SLICE_X3Y110_AO6;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_A3 = CLBLM_R_X5Y112_SLICE_X7Y112_AQ;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_A4 = CLBLM_L_X10Y119_SLICE_X12Y119_AQ;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_A6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_B1 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_B2 = CLBLM_R_X5Y112_SLICE_X7Y112_BQ;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_B3 = CLBLM_R_X5Y112_SLICE_X7Y112_AQ;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_B4 = CLBLL_L_X4Y112_SLICE_X4Y112_CO6;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_B6 = CLBLM_R_X7Y111_SLICE_X9Y111_CQ;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_C2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_C3 = CLBLM_R_X7Y112_SLICE_X8Y112_DQ;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_C4 = CLBLM_R_X11Y110_SLICE_X14Y110_BO5;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_C5 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_C6 = CLBLM_R_X11Y114_SLICE_X14Y114_CQ;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_D2 = CLBLL_L_X4Y113_SLICE_X5Y113_DO6;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_D3 = CLBLM_R_X5Y112_SLICE_X7Y112_DQ;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_D4 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_D5 = CLBLM_R_X7Y115_SLICE_X8Y115_B5Q;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_D6 = CLBLM_L_X12Y108_SLICE_X16Y108_DQ;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_A1 = CLBLL_L_X4Y108_SLICE_X4Y108_CO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_A2 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_A3 = CLBLM_R_X5Y112_SLICE_X6Y112_AQ;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_A4 = CLBLM_R_X5Y112_SLICE_X6Y112_CQ;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_A6 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_B2 = CLBLM_R_X5Y112_SLICE_X6Y112_BQ;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_B3 = CLBLM_L_X8Y113_SLICE_X11Y113_AQ;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_B4 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_B5 = CLBLM_R_X13Y112_SLICE_X18Y112_AQ;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_B6 = CLBLL_L_X4Y112_SLICE_X4Y112_CO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_C2 = CLBLM_R_X5Y112_SLICE_X6Y112_CQ;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_C3 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_C4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_C5 = CLBLM_R_X11Y114_SLICE_X14Y114_BQ;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_C6 = CLBLL_L_X4Y112_SLICE_X5Y112_AQ;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_C4 = CLBLM_L_X10Y115_SLICE_X13Y115_CQ;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_C5 = CLBLM_R_X7Y118_SLICE_X8Y118_CQ;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_C6 = CLBLM_L_X10Y119_SLICE_X12Y119_AQ;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_D1 = CLBLM_R_X7Y114_SLICE_X9Y114_BQ;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_D2 = CLBLL_L_X2Y109_SLICE_X0Y109_AO5;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_D3 = CLBLL_L_X2Y112_SLICE_X0Y112_AO5;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_D4 = CLBLM_R_X7Y113_SLICE_X8Y113_AQ;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_D5 = CLBLM_R_X3Y116_SLICE_X3Y116_AO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_D6 = 1'b1;
  assign LIOI3_X0Y197_OLOGIC_X0Y198_D1 = LIOB33_X0Y73_IOB_X0Y73_I;
  assign LIOI3_X0Y197_OLOGIC_X0Y198_T1 = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_D1 = CLBLL_L_X4Y117_SLICE_X4Y117_DQ;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_B2 = CLBLM_R_X13Y108_SLICE_X19Y108_BQ;
  assign LIOI3_X0Y197_OLOGIC_X0Y197_D1 = LIOB33_X0Y71_IOB_X0Y72_I;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_T1 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_D2 = 1'b1;
  assign RIOI3_X105Y179_OLOGIC_X1Y180_D1 = CLBLM_R_X13Y110_SLICE_X18Y110_DO6;
  assign LIOI3_X0Y197_OLOGIC_X0Y197_T1 = 1'b1;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_B6 = CLBLM_L_X12Y105_SLICE_X17Y105_BO5;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_D1 = CLBLL_L_X4Y118_SLICE_X4Y118_AQ;
  assign LIOB33_X0Y111_IOB_X0Y112_O = CLBLM_R_X11Y110_SLICE_X14Y110_D5Q;
  assign LIOB33_X0Y111_IOB_X0Y111_O = 1'b0;
  assign RIOI3_X105Y179_OLOGIC_X1Y180_T1 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_D5 = CLBLM_R_X7Y116_SLICE_X9Y116_AQ;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_D6 = CLBLM_R_X5Y115_SLICE_X6Y115_BQ;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_T1 = 1'b1;
  assign RIOI3_X105Y179_OLOGIC_X1Y179_D1 = CLBLM_R_X13Y117_SLICE_X18Y117_AO5;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_D1 = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_C1 = CLBLM_L_X12Y107_SLICE_X16Y107_AQ;
  assign RIOI3_X105Y179_OLOGIC_X1Y179_T1 = 1'b1;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_C2 = CLBLM_L_X12Y106_SLICE_X17Y106_CO6;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_T1 = 1'b1;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_C3 = CLBLM_L_X12Y106_SLICE_X17Y106_DO6;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_C4 = 1'b1;
  assign RIOB33_X105Y197_IOB_X1Y198_O = CLBLL_L_X26Y136_SLICE_X38Y136_AO5;
  assign RIOB33_X105Y197_IOB_X1Y197_O = CLBLL_L_X26Y136_SLICE_X38Y136_AO5;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_D1 = RIOB33_X105Y121_IOB_X1Y122_I;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_T1 = 1'b1;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_C5 = 1'b1;
  assign CLBLM_R_X11Y118_SLICE_X14Y118_C6 = 1'b1;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_B5 = CLBLM_L_X8Y108_SLICE_X11Y108_BQ;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_B5 = CLBLM_L_X10Y113_SLICE_X12Y113_AQ;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_B6 = CLBLM_L_X10Y116_SLICE_X12Y116_DO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_C4 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_A1 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_A2 = CLBLL_L_X4Y112_SLICE_X4Y112_CO5;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_A3 = CLBLM_R_X5Y113_SLICE_X7Y113_AQ;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_A4 = CLBLM_L_X12Y113_SLICE_X17Y113_AQ;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_A6 = CLBLM_R_X7Y114_SLICE_X8Y114_CQ;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_C4 = CLBLL_L_X4Y118_SLICE_X4Y118_A5Q;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_B1 = CLBLM_R_X7Y109_SLICE_X9Y109_DQ;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_B2 = CLBLM_R_X7Y113_SLICE_X9Y113_BO6;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_B3 = CLBLM_R_X5Y113_SLICE_X7Y113_AQ;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_B4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_B6 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_C6 = CLBLM_L_X10Y113_SLICE_X13Y113_AQ;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_C1 = CLBLM_L_X10Y113_SLICE_X12Y113_AQ;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_C2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_C3 = CLBLM_L_X8Y114_SLICE_X11Y114_AQ;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_C4 = CLBLM_R_X5Y114_SLICE_X6Y114_BO6;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_C5 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_C6 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign LIOI3_X0Y75_ILOGIC_X0Y76_D = LIOB33_X0Y75_IOB_X0Y76_I;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y75_ILOGIC_X0Y75_D = LIOB33_X0Y75_IOB_X0Y75_I;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_D1 = CLBLM_R_X7Y115_SLICE_X9Y115_A5Q;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_D2 = CLBLM_L_X12Y108_SLICE_X17Y108_AQ;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_D2 = CLBLM_R_X5Y109_SLICE_X7Y109_A5Q;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_D3 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_D4 = CLBLM_R_X7Y114_SLICE_X8Y114_CQ;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_D5 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_D3 = CLBLM_L_X8Y110_SLICE_X11Y110_DQ;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_D6 = CLBLM_L_X8Y113_SLICE_X11Y113_AQ;
  assign RIOI3_X105Y121_ILOGIC_X1Y122_D = RIOB33_X105Y121_IOB_X1Y122_I;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_D4 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign RIOI3_X105Y121_ILOGIC_X1Y121_D = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_A1 = CLBLM_R_X5Y113_SLICE_X6Y113_AQ;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_A2 = CLBLM_R_X11Y113_SLICE_X14Y113_DQ;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_A3 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_D5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_A4 = CLBLM_L_X10Y111_SLICE_X12Y111_AQ;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_A6 = CLBLL_L_X4Y112_SLICE_X4Y112_CO5;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_D6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_B1 = CLBLM_R_X7Y113_SLICE_X9Y113_DO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_B2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_B4 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_B5 = CLBLM_R_X7Y112_SLICE_X9Y112_AQ;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_B6 = CLBLM_R_X5Y114_SLICE_X7Y114_C5Q;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_C2 = CLBLM_R_X5Y113_SLICE_X6Y113_CQ;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_C3 = CLBLM_L_X8Y110_SLICE_X10Y110_BQ;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_C4 = CLBLM_L_X10Y104_SLICE_X12Y104_BO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_C5 = CLBLM_L_X8Y114_SLICE_X11Y114_B5Q;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_C6 = CLBLL_L_X4Y116_SLICE_X5Y116_A5Q;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_D1 = CLBLL_L_X4Y112_SLICE_X4Y112_AQ;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_D2 = CLBLM_R_X5Y116_SLICE_X6Y116_BQ;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_D3 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_D4 = CLBLM_R_X5Y114_SLICE_X6Y114_BO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_D5 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_D6 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_A5 = CLBLM_R_X11Y105_SLICE_X14Y105_DQ;
  assign LIOB33_X0Y113_IOB_X0Y113_O = RIOB33_X105Y121_IOB_X1Y121_I;
  assign LIOB33_X0Y113_IOB_X0Y114_O = CLBLM_R_X7Y113_SLICE_X8Y113_CQ;
  assign LIOB33_X0Y191_IOB_X0Y192_O = LIOB33_X0Y51_IOB_X0Y52_I;
  assign RIOB33_X105Y173_IOB_X1Y174_O = CLBLM_R_X103Y174_SLICE_X163Y174_AO6;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_A1 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_A2 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_A3 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_A4 = CLBLM_R_X11Y115_SLICE_X14Y115_BQ;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_A5 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_A6 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_B1 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_B2 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_B3 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_B4 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_B5 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_B6 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_C1 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_C2 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_C3 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_C4 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_C5 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_C6 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_D1 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_D2 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_D3 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_D4 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_D5 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_D6 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_A1 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_A2 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_A3 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_A4 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_A5 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_A6 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_B1 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_B2 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_B3 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_B4 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_B5 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_B6 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_D1 = CLBLM_L_X10Y104_SLICE_X12Y104_AQ;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_C1 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_C2 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_C3 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_C4 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_C5 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_C6 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_D1 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_D2 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_D3 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_D4 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_D5 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_D6 = 1'b1;
  assign LIOB33_SING_X0Y100_IOB_X0Y100_O = CLBLL_L_X2Y106_SLICE_X0Y106_BO6;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_A2 = CLBLM_R_X11Y114_SLICE_X14Y114_CQ;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_A3 = CLBLM_R_X5Y114_SLICE_X7Y114_AQ;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_A4 = CLBLM_R_X5Y116_SLICE_X7Y116_AQ;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_A5 = CLBLL_L_X4Y116_SLICE_X4Y116_BO6;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_A6 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_B2 = CLBLM_R_X7Y116_SLICE_X9Y116_AQ;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_B4 = CLBLM_R_X5Y113_SLICE_X6Y113_CQ;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_B5 = CLBLM_L_X8Y114_SLICE_X10Y114_DQ;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_B6 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_C2 = CLBLM_R_X7Y114_SLICE_X8Y114_CQ;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_C3 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_C4 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_C5 = CLBLM_R_X7Y110_SLICE_X8Y110_AQ;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_C6 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_D1 = CLBLM_R_X7Y115_SLICE_X8Y115_D5Q;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_D2 = CLBLL_L_X4Y116_SLICE_X5Y116_B5Q;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_D3 = CLBLM_R_X5Y110_SLICE_X6Y110_BQ;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_D4 = CLBLL_L_X4Y116_SLICE_X4Y116_A5Q;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_D5 = CLBLM_R_X5Y114_SLICE_X7Y114_B5Q;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_D6 = CLBLM_R_X5Y116_SLICE_X6Y116_D5Q;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_A1 = CLBLM_R_X5Y113_SLICE_X6Y113_AQ;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_A2 = CLBLM_R_X7Y115_SLICE_X9Y115_B5Q;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_A3 = CLBLM_R_X5Y114_SLICE_X6Y114_AQ;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_A4 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_A6 = CLBLL_L_X4Y113_SLICE_X5Y113_DO6;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_B1 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_B2 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_B3 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_B4 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_B5 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_B6 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_C1 = CLBLM_L_X8Y114_SLICE_X10Y114_AQ;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_C2 = CLBLL_L_X2Y112_SLICE_X0Y112_AO5;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_C3 = CLBLM_R_X3Y116_SLICE_X3Y116_AO6;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_C4 = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_C5 = CLBLL_L_X2Y114_SLICE_X0Y114_AO6;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_C6 = CLBLL_L_X2Y109_SLICE_X0Y109_AO5;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_D1 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_D2 = CLBLL_L_X4Y116_SLICE_X4Y116_A5Q;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_D3 = CLBLM_R_X5Y114_SLICE_X7Y114_B5Q;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_D4 = CLBLL_L_X4Y116_SLICE_X5Y116_B5Q;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_D5 = CLBLM_R_X5Y110_SLICE_X6Y110_BQ;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_D6 = CLBLM_R_X7Y113_SLICE_X9Y113_A5Q;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_C4 = CLBLM_R_X11Y116_SLICE_X14Y116_BQ;
  assign LIOB33_X0Y115_IOB_X0Y115_O = CLBLM_R_X11Y110_SLICE_X14Y110_DQ;
  assign LIOB33_X0Y115_IOB_X0Y116_O = CLBLM_R_X11Y118_SLICE_X15Y118_AQ;
  assign LIOB33_SING_X0Y149_IOB_X0Y149_O = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X37Y117_SLICE_X57Y117_B4 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X163Y170_A1 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X163Y170_A2 = CLBLM_L_X10Y112_SLICE_X13Y112_AQ;
  assign CLBLM_R_X103Y170_SLICE_X163Y170_A3 = CLBLM_L_X12Y117_SLICE_X17Y117_AQ;
  assign CLBLM_R_X103Y170_SLICE_X163Y170_A4 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X163Y170_A5 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_R_X103Y170_SLICE_X163Y170_A6 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X163Y170_B1 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X163Y170_B2 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X163Y170_B3 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X163Y170_B4 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X163Y170_B5 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X163Y170_B6 = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_D1 = CLBLL_L_X4Y116_SLICE_X4Y116_AQ;
  assign CLBLM_R_X103Y170_SLICE_X163Y170_C1 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X163Y170_C2 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X163Y170_C3 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X163Y170_C4 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X163Y170_C5 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X163Y170_C6 = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_T1 = 1'b1;
  assign RIOI3_X105Y183_OLOGIC_X1Y184_D1 = CLBLM_L_X8Y110_SLICE_X10Y110_CO6;
  assign RIOI3_X105Y159_OLOGIC_X1Y160_T1 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X163Y170_D1 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X163Y170_D2 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X163Y170_D3 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X163Y170_D4 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X163Y170_D5 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X163Y170_D6 = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_D1 = CLBLL_L_X4Y118_SLICE_X4Y118_BQ;
  assign RIOI3_X105Y183_OLOGIC_X1Y184_T1 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X162Y170_A1 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X162Y170_A2 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X162Y170_A3 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X162Y170_A4 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X162Y170_A5 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X162Y170_A6 = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_T1 = 1'b1;
  assign RIOI3_X105Y183_OLOGIC_X1Y183_D1 = CLBLM_L_X12Y114_SLICE_X16Y114_DO5;
  assign LIOB33_SING_X0Y150_IOB_X0Y150_O = LIOB33_X0Y63_IOB_X0Y63_I;
  assign CLBLM_R_X103Y170_SLICE_X162Y170_B1 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X162Y170_B2 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X162Y170_B3 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X162Y170_B4 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X162Y170_B5 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X162Y170_B6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_D1 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign RIOI3_X105Y183_OLOGIC_X1Y183_T1 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X162Y170_C1 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X162Y170_C2 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X162Y170_C3 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X162Y170_C4 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X162Y170_C5 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X162Y170_C6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_T1 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X162Y170_D1 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X162Y170_D2 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X162Y170_D3 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X162Y170_D4 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X162Y170_D5 = 1'b1;
  assign CLBLM_R_X103Y170_SLICE_X162Y170_D6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_D1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_A1 = CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_A3 = CLBLM_R_X5Y115_SLICE_X7Y115_AQ;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_A4 = CLBLM_R_X7Y115_SLICE_X9Y115_CO6;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_A5 = CLBLM_R_X5Y109_SLICE_X7Y109_AQ;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_A6 = CLBLM_R_X5Y116_SLICE_X6Y116_CQ;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_T1 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_B1 = CLBLM_R_X5Y116_SLICE_X6Y116_D5Q;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_B2 = CLBLM_R_X5Y115_SLICE_X7Y115_BQ;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_B4 = CLBLM_L_X8Y117_SLICE_X10Y117_BQ;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_B5 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_B6 = CLBLL_L_X4Y113_SLICE_X5Y113_DO6;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_C1 = CLBLM_R_X5Y115_SLICE_X6Y115_DO5;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_C2 = CLBLM_R_X3Y110_SLICE_X2Y110_BO6;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_C3 = CLBLM_R_X7Y115_SLICE_X8Y115_B5Q;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_C4 = CLBLL_L_X4Y107_SLICE_X5Y107_BO6;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_C5 = CLBLM_R_X5Y114_SLICE_X7Y114_DO6;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_C6 = CLBLM_R_X7Y113_SLICE_X9Y113_A5Q;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_D1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_C3 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_D2 = CLBLM_R_X7Y115_SLICE_X9Y115_B5Q;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_D3 = CLBLM_R_X7Y115_SLICE_X8Y115_B5Q;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_D4 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_D5 = CLBLM_R_X5Y114_SLICE_X7Y114_DO6;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_C4 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_D6 = CLBLM_R_X7Y113_SLICE_X9Y113_A5Q;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_C5 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_A2 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_A3 = CLBLM_R_X5Y115_SLICE_X6Y115_AQ;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_C6 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_A4 = CLBLL_L_X4Y115_SLICE_X5Y115_AQ;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_A5 = CLBLL_L_X4Y116_SLICE_X4Y116_BO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_A6 = CLBLM_L_X8Y116_SLICE_X11Y116_BQ;
  assign LIOB33_X0Y117_IOB_X0Y118_O = CLBLM_R_X5Y114_SLICE_X7Y114_CQ;
  assign LIOB33_X0Y117_IOB_X0Y117_O = CLBLL_L_X4Y116_SLICE_X5Y116_BQ;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_B1 = CLBLM_R_X7Y116_SLICE_X9Y116_BO5;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_B2 = CLBLM_R_X5Y115_SLICE_X6Y115_BQ;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_B4 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_B5 = CLBLL_L_X4Y113_SLICE_X5Y113_AQ;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_B6 = CLBLM_R_X7Y115_SLICE_X9Y115_CO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_C2 = CLBLM_R_X5Y115_SLICE_X6Y115_CQ;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_C3 = CLBLM_R_X13Y117_SLICE_X18Y117_BQ;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_C4 = CLBLM_R_X7Y115_SLICE_X8Y115_D5Q;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_C5 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_C6 = CLBLL_L_X4Y113_SLICE_X5Y113_DO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_D1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_D2 = CLBLM_R_X7Y115_SLICE_X9Y115_B5Q;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_D3 = CLBLL_L_X4Y107_SLICE_X5Y107_BO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_D4 = CLBLM_R_X5Y114_SLICE_X6Y114_DO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_D5 = CLBLM_R_X3Y110_SLICE_X2Y110_BO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_D6 = 1'b1;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_D1 = 1'b1;
  assign LIOB33_SING_X0Y199_IOB_X0Y199_O = LIOB33_X0Y73_IOB_X0Y74_I;
  assign CLBLM_L_X12Y117_SLICE_X17Y117_D2 = 1'b1;
  assign LIOI3_X0Y77_ILOGIC_X0Y78_D = LIOB33_X0Y77_IOB_X0Y78_I;
  assign LIOI3_X0Y77_ILOGIC_X0Y77_D = LIOB33_X0Y77_IOB_X0Y77_I;
  assign RIOI3_X105Y123_ILOGIC_X1Y124_D = RIOB33_X105Y123_IOB_X1Y124_I;
  assign RIOI3_X105Y123_ILOGIC_X1Y123_D = RIOB33_X105Y123_IOB_X1Y123_I;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_D = RIOB33_X105Y107_IOB_X1Y108_I;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_D = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_C4 = 1'b1;
  assign LIOB33_X0Y169_IOB_X0Y170_O = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_C6 = 1'b1;
  assign LIOB33_X0Y169_IOB_X0Y169_O = RIOB33_X105Y121_IOB_X1Y122_I;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_B5 = 1'b1;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_B6 = 1'b1;
  assign RIOB33_X105Y151_IOB_X1Y152_O = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_D2 = 1'b1;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_C4 = 1'b1;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_C5 = 1'b1;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_C6 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_A2 = CLBLM_R_X7Y117_SLICE_X9Y117_A5Q;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_A3 = CLBLM_R_X7Y115_SLICE_X9Y115_CO6;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_A4 = CLBLM_R_X7Y117_SLICE_X9Y117_AQ;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_A5 = CLBLM_R_X5Y111_SLICE_X6Y111_AQ;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_A6 = CLBLM_R_X5Y116_SLICE_X7Y116_AQ;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_AX = CLBLM_R_X5Y116_SLICE_X7Y116_CO6;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_B1 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_B2 = CLBLM_R_X5Y116_SLICE_X7Y116_BQ;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_B4 = CLBLM_R_X7Y115_SLICE_X9Y115_CO6;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_B5 = CLBLM_R_X5Y116_SLICE_X7Y116_CO5;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_B6 = CLBLM_R_X5Y106_SLICE_X6Y106_CQ;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_A1 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_A2 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_A3 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_A4 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_A5 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_A6 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_C1 = CLBLM_R_X5Y115_SLICE_X7Y115_AQ;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_C2 = RIOB33_X105Y127_IOB_X1Y127_I;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_B1 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_B2 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_B3 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_B4 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_B5 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_B6 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_D1 = CLBLM_R_X7Y117_SLICE_X9Y117_AQ;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_C1 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_C2 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_C3 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_C4 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_C5 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_C6 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_D3 = CLBLM_R_X7Y116_SLICE_X9Y116_AQ;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_D4 = CLBLM_R_X7Y117_SLICE_X9Y117_BQ;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_D2 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_A1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_A2 = CLBLL_L_X4Y116_SLICE_X5Y116_A5Q;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_A3 = CLBLL_L_X4Y108_SLICE_X4Y108_CO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_A4 = CLBLM_L_X8Y116_SLICE_X10Y116_CQ;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_D3 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_D1 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_D2 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_D3 = 1'b1;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_D4 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_D4 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_D5 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_D6 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_A6 = 1'b1;
  assign CLBLM_L_X12Y117_SLICE_X16Y117_D5 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_B1 = CLBLM_R_X7Y117_SLICE_X8Y117_AQ;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_B2 = CLBLM_R_X5Y116_SLICE_X6Y116_BQ;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_A1 = CLBLM_R_X3Y109_SLICE_X2Y109_AQ;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_A2 = CLBLM_R_X5Y106_SLICE_X7Y106_CO6;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_A3 = CLBLM_R_X3Y110_SLICE_X3Y110_AO6;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_A4 = CLBLL_L_X4Y113_SLICE_X4Y113_BQ;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_A6 = CLBLM_R_X3Y106_SLICE_X2Y106_CO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_C1 = CLBLM_R_X7Y115_SLICE_X9Y115_CO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_C2 = CLBLM_R_X5Y116_SLICE_X6Y116_CQ;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_C3 = CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_B1 = CLBLM_R_X3Y109_SLICE_X2Y109_AQ;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_B2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_B3 = CLBLM_R_X3Y110_SLICE_X3Y110_AO6;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_B4 = CLBLL_L_X4Y113_SLICE_X4Y113_BQ;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_B5 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_B6 = CLBLM_R_X3Y106_SLICE_X2Y106_CO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_D2 = CLBLM_L_X10Y113_SLICE_X13Y113_AQ;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_C1 = LIOB33_X0Y53_IOB_X0Y53_I;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_C2 = LIOB33_X0Y51_IOB_X0Y51_I;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_C3 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_C4 = CLBLL_L_X2Y110_SLICE_X1Y110_DO6;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_C5 = CLBLM_R_X3Y111_SLICE_X2Y111_CO6;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_C6 = CLBLM_R_X3Y109_SLICE_X2Y109_DO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_D3 = CLBLM_R_X5Y116_SLICE_X6Y116_DQ;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_D4 = CLBLM_R_X7Y117_SLICE_X9Y117_AQ;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_D5 = CLBLM_R_X3Y115_SLICE_X2Y115_AQ;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_D6 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_D1 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_D2 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_D3 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_D4 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_D5 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_D6 = 1'b1;
  assign RIOI3_X105Y167_OLOGIC_X1Y167_D1 = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign RIOI3_X105Y167_OLOGIC_X1Y167_T1 = 1'b1;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_D2 = 1'b1;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_C5 = CLBLM_L_X8Y110_SLICE_X11Y110_AQ;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_D3 = 1'b1;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_C6 = CLBLM_R_X5Y115_SLICE_X7Y115_CO6;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_D4 = 1'b1;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_C1 = CLBLM_R_X11Y108_SLICE_X15Y108_AO6;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_D2 = CLBLM_R_X11Y113_SLICE_X15Y113_CQ;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_D3 = 1'b1;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_C2 = CLBLM_R_X11Y111_SLICE_X15Y111_CQ;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_D5 = CLBLM_R_X11Y113_SLICE_X15Y113_DQ;
  assign CLBLM_R_X11Y115_SLICE_X15Y115_D6 = 1'b1;
  assign LIOB33_X0Y121_IOB_X0Y122_O = CLBLM_R_X5Y116_SLICE_X7Y116_A5Q;
  assign LIOB33_X0Y121_IOB_X0Y121_O = CLBLM_R_X11Y118_SLICE_X15Y118_A5Q;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_A2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_A3 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_A4 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_A5 = CLBLL_L_X4Y117_SLICE_X4Y117_BQ;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_A6 = CLBLM_L_X8Y114_SLICE_X11Y114_DO6;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_B1 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_B2 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_B3 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_B4 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_B5 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_B6 = 1'b1;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_A1 = CLBLL_L_X4Y107_SLICE_X5Y107_DO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_A2 = CLBLM_L_X10Y112_SLICE_X13Y112_AQ;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_A3 = CLBLM_R_X3Y107_SLICE_X3Y107_AQ;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_A4 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_A5 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_C1 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_C2 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_C3 = 1'b1;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_B1 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_B2 = CLBLM_R_X5Y107_SLICE_X7Y107_BQ;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_B3 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_B4 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_B5 = CLBLM_R_X3Y110_SLICE_X3Y110_AO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_B6 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_D1 = 1'b1;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_C1 = CLBLM_R_X3Y108_SLICE_X3Y108_AO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_C2 = CLBLL_L_X2Y111_SLICE_X1Y111_CO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_C3 = CLBLM_R_X3Y110_SLICE_X2Y110_DO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_C4 = CLBLM_R_X3Y109_SLICE_X2Y109_CO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_C5 = CLBLM_R_X3Y111_SLICE_X2Y111_CO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_C6 = CLBLM_R_X3Y110_SLICE_X3Y110_AO6;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_D3 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_D4 = 1'b1;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_A1 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_A2 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_A3 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_A4 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_A5 = 1'b1;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_D1 = 1'b1;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_D2 = 1'b1;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_D3 = 1'b1;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_D4 = 1'b1;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_D5 = 1'b1;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_D6 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_A6 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_B1 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_B2 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_B3 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_B4 = 1'b1;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_A1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_A2 = CLBLL_L_X2Y114_SLICE_X0Y114_AO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_A3 = CLBLM_R_X5Y109_SLICE_X6Y109_AQ;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_A4 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_A5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_A6 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_C1 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_C2 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_C3 = 1'b1;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_B1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_B2 = CLBLL_L_X2Y114_SLICE_X0Y114_AO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_B3 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_B4 = CLBLM_R_X5Y107_SLICE_X6Y107_BQ;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_B5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_B6 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_D1 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_D2 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_D4 = 1'b1;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_C1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_C2 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_C3 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_C4 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_C5 = CLBLM_R_X5Y107_SLICE_X6Y107_DQ;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_C6 = CLBLL_L_X2Y114_SLICE_X0Y114_AO6;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_D5 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_D6 = 1'b1;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_C6 = 1'b1;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_B3 = CLBLM_L_X10Y110_SLICE_X13Y110_BQ;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_T1 = 1'b1;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_B4 = CLBLM_L_X10Y115_SLICE_X13Y115_AQ;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_D1 = 1'b1;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_D2 = 1'b1;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_D3 = CLBLL_L_X2Y108_SLICE_X1Y108_AO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_D4 = CLBLM_R_X7Y106_SLICE_X8Y106_AQ;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_D5 = 1'b1;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_D6 = 1'b1;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_B6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_D1 = LIOB33_X0Y55_IOB_X0Y56_I;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_T1 = 1'b1;
  assign RIOI3_SING_X105Y199_OLOGIC_X1Y199_D1 = CLBLM_R_X11Y119_SLICE_X14Y119_AQ;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_D2 = CLBLM_R_X7Y112_SLICE_X8Y112_CQ;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_C2 = CLBLM_L_X10Y119_SLICE_X12Y119_AQ;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_C3 = CLBLM_L_X10Y118_SLICE_X13Y118_AQ;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_C4 = CLBLM_L_X8Y118_SLICE_X10Y118_AQ;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_D5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_C5 = CLBLM_R_X7Y118_SLICE_X8Y118_CQ;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_D6 = CLBLL_L_X4Y117_SLICE_X4Y117_AQ;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_C6 = CLBLM_L_X10Y117_SLICE_X12Y117_DO6;
  assign RIOI3_SING_X105Y199_OLOGIC_X1Y199_T1 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_A1 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_A2 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_A3 = CLBLM_R_X11Y115_SLICE_X14Y115_AQ;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_A4 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_A5 = CLBLM_R_X13Y113_SLICE_X19Y113_AQ;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_A6 = 1'b1;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_D2 = 1'b1;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_A6 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_B1 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_B2 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_B3 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_B2 = CLBLM_L_X8Y111_SLICE_X11Y111_BQ;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_B4 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_B5 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_B6 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_C1 = 1'b1;
  assign CLBLM_R_X11Y115_SLICE_X14Y115_D5 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_C2 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_C3 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_C4 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_C5 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_C6 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_D1 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_D2 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_D3 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_D4 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_D5 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_D6 = 1'b1;
  assign LIOI3_X0Y79_ILOGIC_X0Y79_D = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_A1 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_A2 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_A3 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_A4 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_A5 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_A6 = 1'b1;
  assign RIOI3_X105Y125_ILOGIC_X1Y126_D = RIOB33_X105Y125_IOB_X1Y126_I;
  assign LIOB33_X0Y123_IOB_X0Y124_O = CLBLM_R_X5Y114_SLICE_X7Y114_C5Q;
  assign LIOB33_X0Y123_IOB_X0Y123_O = CLBLM_R_X7Y113_SLICE_X8Y113_C5Q;
  assign RIOI3_X105Y125_ILOGIC_X1Y125_D = RIOB33_X105Y125_IOB_X1Y125_I;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_B1 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_B2 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_B3 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_B4 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_B5 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_B6 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_C3 = CLBLM_R_X5Y110_SLICE_X7Y110_B5Q;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_C1 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_C2 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_C3 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_C4 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_C5 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_C6 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_D1 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_D2 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_D3 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_D4 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_D5 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_D6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_D = RIOB33_X105Y119_IOB_X1Y119_I;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_C3 = 1'b1;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_C4 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_A1 = CLBLL_L_X2Y109_SLICE_X1Y109_AO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_A2 = CLBLM_R_X3Y109_SLICE_X3Y109_AO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_A3 = CLBLM_R_X3Y108_SLICE_X2Y108_CO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_A4 = CLBLL_L_X4Y108_SLICE_X5Y108_BO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_A5 = CLBLL_L_X4Y109_SLICE_X4Y109_DO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_A6 = CLBLL_L_X2Y109_SLICE_X1Y109_CO6;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_C5 = 1'b1;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_C6 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_B1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_B2 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_B3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_B4 = CLBLL_L_X4Y112_SLICE_X4Y112_BQ;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_B5 = CLBLM_R_X3Y116_SLICE_X3Y116_AO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_B6 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_C1 = CLBLL_L_X4Y108_SLICE_X5Y108_BO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_C2 = CLBLM_R_X3Y108_SLICE_X2Y108_CO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_C3 = CLBLM_R_X5Y107_SLICE_X7Y107_AQ;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_C4 = CLBLM_L_X10Y112_SLICE_X12Y112_DO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_C5 = CLBLL_L_X2Y109_SLICE_X1Y109_AO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_C6 = CLBLM_R_X11Y110_SLICE_X14Y110_AQ;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_D1 = CLBLM_R_X7Y111_SLICE_X8Y111_CQ;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_D2 = CLBLM_R_X7Y117_SLICE_X9Y117_DQ;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_AX = CLBLM_R_X11Y105_SLICE_X15Y105_DO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_D1 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_D2 = CLBLM_R_X5Y109_SLICE_X6Y109_AQ;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_D3 = CLBLM_R_X3Y112_SLICE_X2Y112_AO5;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_D4 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_D5 = CLBLL_L_X2Y110_SLICE_X0Y110_BO5;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_D6 = CLBLM_R_X7Y109_SLICE_X9Y109_AQ;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_D5 = 1'b1;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_B1 = CLBLM_L_X12Y105_SLICE_X16Y105_BO5;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_B2 = CLBLM_R_X11Y105_SLICE_X15Y105_BQ;
  assign RIOB33_X105Y175_IOB_X1Y176_O = CLBLM_R_X103Y174_SLICE_X163Y174_AO5;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_A1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_A2 = CLBLM_R_X7Y109_SLICE_X9Y109_AQ;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_A3 = CLBLM_R_X3Y116_SLICE_X3Y116_AO6;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_A4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_A5 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_A6 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign RIOB33_X105Y175_IOB_X1Y175_O = CLBLM_R_X13Y118_SLICE_X18Y118_AO6;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_B1 = CLBLL_L_X2Y108_SLICE_X1Y108_AO5;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_B2 = CLBLM_R_X3Y108_SLICE_X3Y108_DO6;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_B3 = CLBLL_L_X4Y108_SLICE_X5Y108_BO6;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_B4 = CLBLL_L_X2Y108_SLICE_X1Y108_CO6;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_B5 = CLBLM_L_X10Y112_SLICE_X12Y112_DO6;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_B6 = CLBLL_L_X2Y110_SLICE_X1Y110_CO6;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_D1 = 1'b1;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_B5 = CLBLM_R_X11Y112_SLICE_X15Y112_AQ;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_D2 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_C1 = CLBLM_R_X3Y108_SLICE_X2Y108_AO6;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_C2 = CLBLM_R_X7Y106_SLICE_X8Y106_AQ;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_C3 = CLBLL_L_X2Y109_SLICE_X0Y109_DO6;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_C4 = CLBLM_R_X3Y107_SLICE_X2Y107_AO6;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_C5 = CLBLL_L_X2Y108_SLICE_X1Y108_AO6;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_C6 = CLBLM_R_X3Y111_SLICE_X3Y111_AO6;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_D5 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_D1 = CLBLL_L_X4Y108_SLICE_X5Y108_BO6;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_D2 = CLBLL_L_X2Y110_SLICE_X1Y110_CO6;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_D3 = CLBLL_L_X2Y108_SLICE_X1Y108_AO5;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_D4 = CLBLM_R_X3Y108_SLICE_X3Y108_DO6;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_D5 = CLBLL_L_X2Y109_SLICE_X1Y109_DO6;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_D6 = CLBLM_R_X3Y107_SLICE_X2Y107_DO6;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_C2 = CLBLM_R_X11Y105_SLICE_X15Y105_CQ;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_C5 = CLBLM_R_X7Y105_SLICE_X9Y105_CQ;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_B5 = 1'b1;
  assign CLBLM_R_X37Y117_SLICE_X56Y117_B4 = 1'b1;
  assign CLBLM_R_X103Y138_SLICE_X162Y138_B6 = 1'b1;
  assign CLBLM_R_X37Y117_SLICE_X56Y117_B5 = 1'b1;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_D5 = CLBLM_L_X10Y111_SLICE_X12Y111_BQ;
  assign CLBLM_R_X37Y117_SLICE_X56Y117_B6 = 1'b1;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_D6 = 1'b1;
  assign LIOI3_X0Y67_ILOGIC_X0Y68_D = LIOB33_X0Y67_IOB_X0Y68_I;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_A1 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_A2 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_A3 = CLBLM_R_X11Y119_SLICE_X14Y119_AQ;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_A4 = CLBLM_R_X13Y109_SLICE_X19Y109_AQ;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_A5 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_A6 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_B1 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_B2 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_B3 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_B4 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_B5 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_B6 = 1'b1;
  assign LIOI3_X0Y67_ILOGIC_X0Y67_D = LIOB33_X0Y67_IOB_X0Y67_I;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_C4 = CLBLM_R_X5Y116_SLICE_X6Y116_CQ;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_C1 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_C2 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_C3 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_C4 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_C5 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_C6 = 1'b1;
  assign LIOB33_X0Y125_IOB_X0Y125_O = CLBLM_R_X11Y115_SLICE_X15Y115_B5Q;
  assign LIOB33_X0Y125_IOB_X0Y126_O = CLBLL_L_X4Y117_SLICE_X4Y117_CQ;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_D1 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_D2 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_D3 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_D4 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_D5 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_D6 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_C5 = CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_A1 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_A2 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_A3 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_A4 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_A5 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_A6 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_B1 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_B2 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_B3 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_B4 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_B5 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_B6 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_C6 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_C1 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_C2 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_C3 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_C4 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_C5 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_C6 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_D1 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_D2 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_D3 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_D4 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_D5 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_D6 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_D6 = CLBLM_R_X7Y112_SLICE_X8Y112_BQ;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_A1 = CLBLM_R_X3Y112_SLICE_X3Y112_CO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_A2 = CLBLM_R_X3Y109_SLICE_X2Y109_BO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_A3 = CLBLM_R_X3Y108_SLICE_X3Y108_BO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_A4 = CLBLM_R_X3Y109_SLICE_X3Y109_BO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_A5 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_A6 = CLBLL_L_X2Y111_SLICE_X1Y111_BO5;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_B1 = CLBLM_R_X3Y107_SLICE_X3Y107_BO5;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_B2 = CLBLL_L_X2Y114_SLICE_X0Y114_AO5;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_B3 = CLBLL_L_X2Y112_SLICE_X0Y112_AO5;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_B4 = LIOB33_X0Y65_IOB_X0Y66_I;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_B5 = CLBLL_L_X2Y112_SLICE_X0Y112_AO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_B6 = CLBLM_R_X5Y112_SLICE_X7Y112_DQ;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_C1 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_C2 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_C3 = CLBLL_L_X2Y114_SLICE_X0Y114_AO5;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_C4 = CLBLL_L_X2Y112_SLICE_X0Y112_AO5;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_C5 = CLBLM_R_X5Y112_SLICE_X7Y112_DQ;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_C6 = CLBLM_R_X5Y107_SLICE_X7Y107_BQ;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_D1 = CLBLL_L_X2Y109_SLICE_X0Y109_AO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_D2 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_D3 = CLBLL_L_X4Y112_SLICE_X4Y112_BQ;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_D4 = CLBLM_R_X3Y109_SLICE_X3Y109_CO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_D5 = LIOB33_X0Y65_IOB_X0Y66_I;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_D6 = CLBLL_L_X2Y110_SLICE_X0Y110_BO5;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_A2 = CLBLM_R_X3Y115_SLICE_X2Y115_AQ;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_A3 = CLBLL_L_X4Y109_SLICE_X4Y109_BQ;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_A4 = CLBLL_L_X4Y113_SLICE_X4Y113_BQ;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_A5 = CLBLM_R_X3Y107_SLICE_X3Y107_AQ;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_A6 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_B1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_B2 = CLBLM_R_X5Y115_SLICE_X6Y115_AQ;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_B3 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_B4 = CLBLM_R_X3Y116_SLICE_X3Y116_AO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_B5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_B6 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_C1 = CLBLL_L_X2Y110_SLICE_X1Y110_CO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_C2 = CLBLM_R_X3Y110_SLICE_X3Y110_CO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_C3 = CLBLL_L_X4Y109_SLICE_X5Y109_DO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_C4 = CLBLL_L_X2Y109_SLICE_X0Y109_BO5;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_C5 = CLBLL_L_X4Y112_SLICE_X4Y112_DO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_C6 = CLBLL_L_X2Y112_SLICE_X1Y112_AO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_X105Y191_OLOGIC_X1Y191_D1 = CLBLM_R_X11Y115_SLICE_X14Y115_AQ;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_D1 = CLBLM_R_X3Y109_SLICE_X2Y109_CO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_D2 = CLBLL_L_X4Y113_SLICE_X5Y113_B5Q;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_D3 = CLBLM_R_X3Y110_SLICE_X2Y110_DO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_D4 = CLBLM_R_X3Y109_SLICE_X2Y109_A5Q;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_D5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_D6 = CLBLM_R_X3Y115_SLICE_X2Y115_AQ;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_D1 = LIOB33_X0Y59_IOB_X0Y59_I;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_T1 = 1'b1;
  assign RIOI3_X105Y191_OLOGIC_X1Y191_T1 = 1'b1;
  assign RIOI3_X105Y189_OLOGIC_X1Y190_D1 = CLBLM_R_X13Y113_SLICE_X19Y113_AQ;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_D1 = LIOB33_X0Y57_IOB_X0Y58_I;
  assign RIOI3_X105Y189_OLOGIC_X1Y190_T1 = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_T1 = 1'b1;
  assign RIOI3_X105Y189_OLOGIC_X1Y189_D1 = CLBLM_L_X10Y112_SLICE_X13Y112_AQ;
  assign RIOI3_X105Y189_OLOGIC_X1Y189_T1 = 1'b1;
  assign LIOB33_X0Y127_IOB_X0Y128_O = CLBLM_R_X3Y115_SLICE_X2Y115_AQ;
  assign LIOB33_X0Y127_IOB_X0Y127_O = CLBLL_L_X4Y113_SLICE_X4Y113_BQ;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_A1 = CLBLL_L_X2Y109_SLICE_X1Y109_BO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_A2 = CLBLL_L_X4Y110_SLICE_X5Y110_CO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_A3 = CLBLL_L_X4Y110_SLICE_X4Y110_DO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_A4 = CLBLM_R_X3Y114_SLICE_X3Y114_AO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_A5 = CLBLL_L_X4Y110_SLICE_X5Y110_BO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_A6 = CLBLM_R_X3Y112_SLICE_X2Y112_DO6;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_D1 = LIOB33_X0Y59_IOB_X0Y60_I;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_B1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_B2 = CLBLL_L_X2Y110_SLICE_X0Y110_AO5;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_B3 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_B4 = CLBLM_R_X5Y109_SLICE_X6Y109_BQ;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_B5 = CLBLM_R_X3Y116_SLICE_X3Y116_AO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_B6 = CLBLL_L_X2Y114_SLICE_X0Y114_AO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_C1 = CLBLM_R_X7Y109_SLICE_X8Y109_BQ;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_C2 = CLBLM_R_X3Y112_SLICE_X3Y112_BO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_C3 = CLBLM_R_X3Y111_SLICE_X3Y111_CO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_C4 = CLBLL_L_X2Y110_SLICE_X0Y110_BO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_C5 = CLBLM_R_X5Y114_SLICE_X7Y114_AQ;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_C6 = CLBLM_R_X3Y110_SLICE_X3Y110_BO6;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_C4 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_D1 = CLBLM_R_X5Y115_SLICE_X6Y115_AQ;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_C5 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_D2 = CLBLL_L_X2Y109_SLICE_X1Y109_CO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_D3 = CLBLM_R_X3Y109_SLICE_X3Y109_DO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_D4 = CLBLL_L_X4Y109_SLICE_X4Y109_DO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_D5 = CLBLM_R_X3Y111_SLICE_X3Y111_DO6;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_C6 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_D6 = CLBLL_L_X2Y110_SLICE_X0Y110_CO5;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_A1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_A2 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_A3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_A4 = CLBLL_L_X2Y114_SLICE_X0Y114_AO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_A5 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_A6 = 1'b1;
  assign RIOI3_X105Y127_ILOGIC_X1Y128_D = RIOB33_X105Y127_IOB_X1Y128_I;
  assign RIOI3_X105Y127_ILOGIC_X1Y127_D = RIOB33_X105Y127_IOB_X1Y127_I;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_B1 = CLBLL_L_X2Y111_SLICE_X1Y111_DO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_B2 = CLBLM_R_X3Y108_SLICE_X2Y108_DO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_B3 = CLBLM_R_X3Y110_SLICE_X3Y110_DO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_B4 = CLBLM_R_X3Y110_SLICE_X2Y110_DO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_B5 = CLBLL_L_X2Y112_SLICE_X1Y112_BO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_B6 = CLBLM_R_X3Y109_SLICE_X2Y109_CO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_C1 = CLBLM_R_X3Y110_SLICE_X2Y110_AO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_C2 = CLBLL_L_X2Y110_SLICE_X1Y110_CO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_C3 = CLBLM_R_X3Y112_SLICE_X3Y112_BO5;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_C4 = CLBLL_L_X2Y108_SLICE_X1Y108_AO5;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_C5 = CLBLL_L_X2Y111_SLICE_X1Y111_AO5;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_C6 = CLBLL_L_X2Y112_SLICE_X1Y112_AO6;
  assign RIOB33_X105Y153_IOB_X1Y154_O = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_D1 = CLBLL_L_X4Y109_SLICE_X5Y109_BO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_D2 = CLBLM_R_X3Y111_SLICE_X2Y111_DO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_D3 = CLBLL_L_X2Y111_SLICE_X1Y111_AO5;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_D4 = CLBLL_L_X2Y110_SLICE_X1Y110_CO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_D5 = CLBLM_R_X3Y112_SLICE_X2Y112_DO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_D6 = CLBLL_L_X4Y110_SLICE_X5Y110_DO6;
  assign CLBLM_L_X12Y105_SLICE_X17Y105_A1 = CLBLM_R_X13Y109_SLICE_X19Y109_BQ;
  assign CLBLM_L_X12Y105_SLICE_X17Y105_A2 = CLBLM_L_X12Y107_SLICE_X17Y107_DO5;
  assign CLBLM_L_X12Y105_SLICE_X17Y105_A3 = CLBLM_R_X11Y105_SLICE_X14Y105_DQ;
  assign CLBLM_L_X12Y105_SLICE_X17Y105_A4 = CLBLM_R_X11Y106_SLICE_X15Y106_DO5;
  assign CLBLM_L_X12Y105_SLICE_X17Y105_A5 = CLBLM_R_X13Y113_SLICE_X18Y113_BQ;
  assign CLBLM_L_X12Y105_SLICE_X17Y105_A6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y132_D = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_D3 = 1'b1;
  assign CLBLM_L_X12Y105_SLICE_X17Y105_B1 = CLBLM_R_X13Y109_SLICE_X19Y109_BQ;
  assign CLBLM_L_X12Y105_SLICE_X17Y105_B2 = CLBLM_R_X13Y113_SLICE_X18Y113_BQ;
  assign CLBLM_L_X12Y105_SLICE_X17Y105_B3 = CLBLM_R_X11Y105_SLICE_X15Y105_BQ;
  assign CLBLM_L_X12Y105_SLICE_X17Y105_B4 = CLBLM_L_X12Y107_SLICE_X17Y107_BQ;
  assign CLBLM_L_X12Y105_SLICE_X17Y105_B5 = CLBLM_L_X12Y105_SLICE_X16Y105_AQ;
  assign CLBLM_L_X12Y105_SLICE_X17Y105_B6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y131_D = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X12Y105_SLICE_X17Y105_C1 = CLBLM_L_X12Y105_SLICE_X16Y105_AQ;
  assign CLBLM_L_X12Y105_SLICE_X17Y105_C2 = CLBLM_R_X11Y105_SLICE_X15Y105_BQ;
  assign CLBLM_L_X12Y105_SLICE_X17Y105_C3 = CLBLM_R_X13Y109_SLICE_X19Y109_BQ;
  assign CLBLM_L_X12Y105_SLICE_X17Y105_C4 = CLBLM_R_X13Y113_SLICE_X18Y113_BQ;
  assign CLBLM_L_X12Y105_SLICE_X17Y105_C5 = CLBLM_L_X12Y107_SLICE_X17Y107_BQ;
  assign CLBLM_L_X12Y105_SLICE_X17Y105_C6 = CLBLM_R_X11Y106_SLICE_X15Y106_DO5;
  assign CLBLM_L_X12Y118_SLICE_X17Y118_D6 = 1'b1;
  assign CLBLM_L_X12Y105_SLICE_X17Y105_D1 = 1'b1;
  assign CLBLM_L_X12Y105_SLICE_X17Y105_D2 = 1'b1;
  assign CLBLM_L_X12Y105_SLICE_X17Y105_D3 = 1'b1;
  assign CLBLM_L_X12Y105_SLICE_X17Y105_D4 = 1'b1;
  assign CLBLM_L_X12Y105_SLICE_X17Y105_D5 = 1'b1;
  assign CLBLM_L_X12Y105_SLICE_X17Y105_D6 = 1'b1;
  assign CLBLM_L_X12Y105_SLICE_X16Y105_A1 = CLBLM_L_X12Y107_SLICE_X17Y107_DO6;
  assign CLBLM_L_X12Y105_SLICE_X16Y105_A2 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X12Y105_SLICE_X16Y105_A3 = CLBLM_L_X12Y105_SLICE_X16Y105_AQ;
  assign CLBLM_L_X12Y105_SLICE_X16Y105_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y105_SLICE_X16Y105_A5 = CLBLM_R_X7Y106_SLICE_X8Y106_CQ;
  assign CLBLM_L_X12Y105_SLICE_X16Y105_A6 = CLBLM_L_X12Y105_SLICE_X16Y105_CO6;
  assign CLBLM_L_X12Y105_SLICE_X16Y105_B1 = CLBLM_R_X13Y109_SLICE_X19Y109_BQ;
  assign CLBLM_L_X12Y105_SLICE_X16Y105_B2 = CLBLM_R_X11Y106_SLICE_X15Y106_DO5;
  assign CLBLM_L_X12Y105_SLICE_X16Y105_B3 = CLBLM_L_X12Y105_SLICE_X16Y105_AQ;
  assign CLBLM_L_X12Y105_SLICE_X16Y105_B4 = CLBLM_R_X13Y113_SLICE_X18Y113_BQ;
  assign CLBLM_L_X12Y105_SLICE_X16Y105_B5 = CLBLM_L_X12Y107_SLICE_X17Y107_BQ;
  assign CLBLM_L_X12Y105_SLICE_X16Y105_B6 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_D5 = 1'b1;
  assign CLBLM_L_X12Y105_SLICE_X16Y105_C1 = CLBLM_R_X13Y108_SLICE_X18Y108_BO5;
  assign CLBLM_L_X12Y105_SLICE_X16Y105_C2 = CLBLM_L_X12Y105_SLICE_X16Y105_AQ;
  assign CLBLM_L_X12Y105_SLICE_X16Y105_C3 = CLBLM_R_X11Y106_SLICE_X15Y106_DO5;
  assign CLBLM_L_X12Y105_SLICE_X16Y105_C4 = CLBLM_R_X11Y105_SLICE_X15Y105_BQ;
  assign CLBLM_L_X12Y105_SLICE_X16Y105_C5 = CLBLM_L_X12Y107_SLICE_X17Y107_BQ;
  assign CLBLM_L_X12Y105_SLICE_X16Y105_C6 = 1'b1;
  assign LIOB33_X0Y129_IOB_X0Y129_O = CLBLM_R_X5Y109_SLICE_X6Y109_CQ;
  assign LIOB33_X0Y129_IOB_X0Y130_O = CLBLL_L_X52Y126_SLICE_X78Y126_AO6;
  assign CLBLM_L_X12Y105_SLICE_X16Y105_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_A5 = 1'b1;
  assign CLBLM_L_X12Y105_SLICE_X16Y105_D1 = 1'b1;
  assign CLBLM_L_X12Y105_SLICE_X16Y105_D2 = 1'b1;
  assign CLBLM_L_X12Y105_SLICE_X16Y105_D3 = 1'b1;
  assign CLBLM_L_X12Y105_SLICE_X16Y105_D4 = 1'b1;
  assign CLBLM_L_X12Y105_SLICE_X16Y105_D5 = 1'b1;
  assign CLBLM_L_X12Y105_SLICE_X16Y105_D6 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_A6 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_D6 = 1'b1;
  assign RIOI3_X105Y167_OLOGIC_X1Y168_T1 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_B1 = 1'b1;
  assign RIOI3_SING_X105Y100_ILOGIC_X1Y100_D = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_C3 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_C4 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_C5 = 1'b1;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_C6 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_A1 = CLBLL_L_X2Y114_SLICE_X0Y114_AO5;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_A2 = CLBLL_L_X4Y110_SLICE_X4Y110_CQ;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_A3 = CLBLL_L_X2Y107_SLICE_X1Y107_AO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_A4 = CLBLM_R_X3Y115_SLICE_X3Y115_AO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_A5 = CLBLM_R_X5Y115_SLICE_X7Y115_BQ;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_A6 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_B1 = CLBLL_L_X2Y114_SLICE_X0Y114_AO5;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_B2 = CLBLM_R_X3Y115_SLICE_X3Y115_AO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_B3 = CLBLM_R_X5Y114_SLICE_X6Y114_AQ;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_B4 = CLBLL_L_X4Y110_SLICE_X4Y110_C5Q;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_B5 = CLBLL_L_X2Y107_SLICE_X1Y107_AO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_B6 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_C1 = CLBLM_R_X3Y116_SLICE_X3Y116_AO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_C2 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_C3 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_C4 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_C5 = CLBLM_L_X8Y110_SLICE_X11Y110_AQ;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_C6 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_D1 = CLBLM_R_X3Y110_SLICE_X2Y110_AO5;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_D2 = CLBLL_L_X2Y111_SLICE_X1Y111_BO5;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_D2 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_D3 = CLBLM_R_X5Y112_SLICE_X6Y112_BQ;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_D4 = CLBLM_R_X5Y110_SLICE_X6Y110_CQ;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_D5 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_D6 = CLBLL_L_X2Y111_SLICE_X1Y111_AO6;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_D3 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_A1 = CLBLM_R_X5Y106_SLICE_X7Y106_AQ;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_A2 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_A3 = CLBLL_L_X2Y111_SLICE_X1Y111_BO5;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_A4 = CLBLL_L_X2Y108_SLICE_X1Y108_AO5;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_A5 = CLBLL_L_X2Y110_SLICE_X0Y110_BO6;
  assign CLBLM_L_X12Y118_SLICE_X16Y118_D5 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_A6 = CLBLL_L_X4Y111_SLICE_X4Y111_BQ;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_B1 = CLBLM_R_X3Y112_SLICE_X2Y112_AO5;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_B2 = CLBLM_R_X3Y111_SLICE_X3Y111_BO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_B3 = CLBLM_R_X5Y113_SLICE_X7Y113_AQ;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_B4 = CLBLL_L_X2Y111_SLICE_X0Y111_AO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_B5 = CLBLL_L_X2Y110_SLICE_X0Y110_BO5;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_B6 = CLBLL_L_X4Y108_SLICE_X4Y108_AQ;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_C1 = CLBLM_R_X3Y115_SLICE_X2Y115_CO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_C2 = CLBLL_L_X2Y111_SLICE_X1Y111_AO5;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_C3 = CLBLM_R_X3Y112_SLICE_X2Y112_DO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_C4 = CLBLL_L_X4Y111_SLICE_X5Y111_DO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_C5 = CLBLL_L_X4Y111_SLICE_X4Y111_DO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_C6 = CLBLL_L_X2Y110_SLICE_X1Y110_CO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_D1 = CLBLL_L_X2Y111_SLICE_X0Y111_CO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_D2 = CLBLM_R_X3Y107_SLICE_X2Y107_BO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_D3 = CLBLM_R_X3Y112_SLICE_X2Y112_BO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_D4 = CLBLM_R_X3Y107_SLICE_X2Y107_CO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_D5 = CLBLM_R_X3Y113_SLICE_X2Y113_DO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_D6 = CLBLM_R_X3Y115_SLICE_X2Y115_DO6;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_A1 = 1'b1;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_A3 = CLBLM_L_X12Y106_SLICE_X17Y106_AQ;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_A5 = CLBLM_R_X13Y107_SLICE_X18Y107_AQ;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_A6 = 1'b1;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_B1 = CLBLM_L_X12Y106_SLICE_X17Y106_DO6;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_B2 = CLBLM_L_X12Y107_SLICE_X16Y107_CQ;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_B3 = CLBLM_L_X12Y105_SLICE_X17Y105_AO5;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_B4 = CLBLM_L_X12Y105_SLICE_X17Y105_CO6;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_B5 = CLBLM_L_X12Y107_SLICE_X16Y107_AQ;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_B6 = CLBLM_L_X12Y106_SLICE_X17Y106_CO6;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_A1 = 1'b1;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_A2 = 1'b1;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_A3 = 1'b1;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_A4 = 1'b1;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_C1 = CLBLM_R_X13Y107_SLICE_X19Y107_AQ;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_C2 = CLBLM_L_X12Y105_SLICE_X17Y105_BO5;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_C3 = CLBLM_L_X12Y108_SLICE_X16Y108_BQ;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_A5 = 1'b1;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_C5 = CLBLM_L_X12Y107_SLICE_X16Y107_BQ;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_C6 = CLBLM_R_X13Y107_SLICE_X19Y107_BQ;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_A6 = 1'b1;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_B1 = 1'b1;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_B2 = 1'b1;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_B3 = 1'b1;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_B4 = 1'b1;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_B5 = 1'b1;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_B6 = 1'b1;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_D1 = CLBLM_R_X13Y107_SLICE_X19Y107_AQ;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_D2 = CLBLM_L_X12Y105_SLICE_X17Y105_BO5;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_D3 = CLBLM_L_X12Y108_SLICE_X16Y108_BQ;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_C3 = 1'b1;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_C4 = 1'b1;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_D4 = CLBLM_R_X13Y108_SLICE_X19Y108_BQ;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_D5 = CLBLM_L_X12Y107_SLICE_X16Y107_BQ;
  assign CLBLM_L_X12Y106_SLICE_X17Y106_D6 = CLBLM_R_X13Y107_SLICE_X19Y107_BQ;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_C1 = 1'b1;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_C2 = 1'b1;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_C5 = 1'b1;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_C6 = 1'b1;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_A1 = CLBLM_R_X13Y109_SLICE_X19Y109_BQ;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_A2 = CLBLM_R_X11Y105_SLICE_X15Y105_BQ;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_D1 = 1'b1;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_D2 = 1'b1;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_D3 = 1'b1;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_D4 = 1'b1;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_D5 = 1'b1;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_D6 = 1'b1;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_A3 = CLBLM_L_X12Y105_SLICE_X16Y105_AQ;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_A5 = CLBLM_L_X12Y107_SLICE_X17Y107_BQ;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_A6 = CLBLM_R_X13Y113_SLICE_X18Y113_BQ;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_B1 = CLBLM_L_X12Y108_SLICE_X16Y108_BQ;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_A1 = CLBLM_L_X10Y110_SLICE_X12Y110_B5Q;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_A2 = 1'b1;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_A3 = 1'b1;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_A4 = 1'b1;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_A5 = 1'b1;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_A6 = 1'b1;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_B3 = CLBLM_L_X12Y105_SLICE_X17Y105_CO6;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_B4 = CLBLM_L_X12Y108_SLICE_X17Y108_BQ;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_B5 = CLBLM_L_X12Y105_SLICE_X17Y105_AO5;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_B1 = 1'b1;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_B2 = 1'b1;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_B3 = 1'b1;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_B4 = 1'b1;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_B5 = 1'b1;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_B6 = 1'b1;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_C4 = CLBLM_L_X12Y105_SLICE_X17Y105_AO5;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_C5 = CLBLM_R_X11Y106_SLICE_X14Y106_CQ;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_C6 = CLBLM_L_X12Y105_SLICE_X17Y105_CO6;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_D1 = CLBLM_L_X12Y105_SLICE_X17Y105_AO5;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_D2 = CLBLM_R_X13Y108_SLICE_X19Y108_BQ;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_C3 = 1'b1;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_C4 = 1'b1;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_C5 = 1'b1;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_C6 = 1'b1;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_D6 = CLBLM_R_X11Y105_SLICE_X15Y105_CQ;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_D3 = CLBLM_L_X12Y105_SLICE_X17Y105_CO6;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_D4 = CLBLM_L_X12Y105_SLICE_X17Y105_BO5;
  assign CLBLM_L_X12Y106_SLICE_X16Y106_D5 = CLBLM_L_X12Y108_SLICE_X16Y108_BQ;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_D1 = 1'b1;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_D2 = 1'b1;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_D3 = 1'b1;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_D4 = 1'b1;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_D5 = 1'b1;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_D6 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_A1 = CLBLM_L_X12Y110_SLICE_X16Y110_AQ;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_A2 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_A3 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_A4 = CLBLM_L_X12Y111_SLICE_X16Y111_AQ;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_A5 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_A6 = 1'b1;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_C4 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_B1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_B2 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_B3 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_B4 = 1'b1;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_C5 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_B6 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_B5 = 1'b1;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_C6 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_C1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_C2 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_C3 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_C4 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_C5 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_C6 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_D1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_D2 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_D3 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_D4 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_D5 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_D6 = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_D1 = LIOB33_X0Y61_IOB_X0Y61_I;
  assign LIOI3_X0Y117_OLOGIC_X0Y117_T1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_A1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_A2 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_A3 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_A4 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_A5 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_A6 = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_T1 = 1'b1;
  assign RIOI3_X105Y191_OLOGIC_X1Y192_D1 = CLBLM_R_X13Y109_SLICE_X19Y109_AQ;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_B1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_B2 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_B3 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_B4 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_B5 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_B6 = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_D1 = LIOB33_X0Y71_IOB_X0Y71_I;
  assign RIOI3_X105Y191_OLOGIC_X1Y192_T1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_C1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_C2 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_C3 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_A1 = CLBLM_L_X10Y112_SLICE_X12Y112_C5Q;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_A2 = RIOB33_X105Y139_IOB_X1Y140_I;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_A3 = CLBLM_L_X12Y112_SLICE_X16Y112_B5Q;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_A4 = RIOB33_X105Y141_IOB_X1Y141_I;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_A6 = 1'b1;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_D2 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_C4 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_C5 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_B1 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_B2 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_B3 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_B4 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_B5 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_B6 = 1'b1;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_D5 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_D1 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_C1 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_C2 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_C3 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_C4 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_C5 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_C6 = 1'b1;
  assign CLBLM_R_X11Y116_SLICE_X15Y116_D6 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_D6 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_D1 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_D2 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_D3 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_D4 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_D5 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_A1 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_A3 = CLBLM_R_X3Y112_SLICE_X3Y112_AQ;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_A4 = CLBLM_R_X11Y105_SLICE_X14Y105_CQ;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_A5 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_A6 = CLBLL_L_X4Y108_SLICE_X4Y108_CO6;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_D6 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_A1 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_B1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_B2 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_B3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_B4 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_B5 = CLBLM_R_X3Y116_SLICE_X3Y116_AO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_B6 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_A2 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_A3 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_A4 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_C1 = CLBLM_R_X5Y112_SLICE_X6Y112_BQ;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_C2 = CLBLM_R_X5Y110_SLICE_X6Y110_CQ;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_C3 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_C4 = CLBLL_L_X26Y136_SLICE_X38Y136_AO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_C5 = CLBLL_L_X2Y112_SLICE_X0Y112_AO5;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_C6 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_B1 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_B2 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_C1 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_C2 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_C3 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_C4 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_D1 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_D2 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_D3 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_D4 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_D5 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_D6 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_C5 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_C6 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_D1 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_D2 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_A1 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_A2 = CLBLL_L_X2Y114_SLICE_X0Y114_AO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_A3 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_A4 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_A5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_A6 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_D3 = 1'b1;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_C1 = CLBLM_L_X8Y116_SLICE_X11Y116_CO6;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_D4 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_D5 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_B1 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_B2 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_B3 = CLBLM_L_X8Y109_SLICE_X10Y109_AQ;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_B4 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_B5 = CLBLL_L_X26Y136_SLICE_X38Y136_AO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_B6 = CLBLL_L_X2Y112_SLICE_X0Y112_AO6;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_C2 = CLBLM_R_X7Y118_SLICE_X9Y118_AQ;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_C3 = CLBLM_R_X7Y118_SLICE_X8Y118_AQ;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_C1 = CLBLM_R_X5Y106_SLICE_X7Y106_AQ;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_C2 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_C3 = CLBLM_R_X3Y112_SLICE_X3Y112_BO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_C4 = CLBLM_R_X3Y113_SLICE_X2Y113_AO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_C5 = CLBLM_R_X7Y115_SLICE_X9Y115_AQ;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_C6 = CLBLL_L_X2Y108_SLICE_X1Y108_AO5;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_C4 = CLBLM_R_X7Y117_SLICE_X8Y117_BQ;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_C5 = CLBLM_R_X7Y118_SLICE_X8Y118_BQ;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_C6 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_D1 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_D2 = CLBLL_L_X26Y136_SLICE_X38Y136_AO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_D3 = CLBLM_R_X3Y112_SLICE_X3Y112_BO5;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_D4 = CLBLL_L_X2Y109_SLICE_X0Y109_AO5;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_D5 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_D6 = CLBLL_L_X2Y108_SLICE_X1Y108_AO5;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_B4 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_A1 = CLBLM_L_X12Y107_SLICE_X17Y107_DO6;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_A2 = CLBLM_L_X12Y108_SLICE_X17Y108_CO5;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_A3 = CLBLM_L_X12Y107_SLICE_X17Y107_AQ;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_A4 = CLBLM_L_X8Y109_SLICE_X10Y109_AQ;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_A6 = CLBLM_L_X12Y107_SLICE_X17Y107_CO6;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_B5 = 1'b1;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_B6 = CLBLM_R_X11Y116_SLICE_X14Y116_CO6;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_B2 = CLBLM_L_X12Y105_SLICE_X17Y105_BO6;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_B3 = CLBLM_R_X13Y113_SLICE_X18Y113_AQ;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_B4 = CLBLM_R_X13Y108_SLICE_X18Y108_BO6;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_B5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_B6 = CLBLM_L_X12Y107_SLICE_X17Y107_BQ;
  assign LIOB33_X0Y133_IOB_X0Y133_O = CLBLL_L_X4Y118_SLICE_X4Y118_A5Q;
  assign LIOB33_X0Y133_IOB_X0Y134_O = CLBLL_L_X4Y116_SLICE_X5Y116_AQ;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_C1 = CLBLM_R_X13Y113_SLICE_X18Y113_BQ;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_C2 = CLBLM_R_X11Y105_SLICE_X15Y105_BQ;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_C3 = CLBLM_R_X13Y109_SLICE_X19Y109_BQ;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_C4 = CLBLM_L_X12Y107_SLICE_X17Y107_BQ;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_C5 = CLBLM_L_X12Y105_SLICE_X16Y105_AQ;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_C6 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_D1 = CLBLM_R_X13Y108_SLICE_X18Y108_BO6;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_D2 = CLBLM_R_X11Y105_SLICE_X15Y105_BQ;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_D3 = CLBLM_L_X12Y107_SLICE_X17Y107_BQ;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_D4 = CLBLM_L_X12Y105_SLICE_X16Y105_AQ;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_D5 = CLBLM_L_X12Y107_SLICE_X17Y107_AQ;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_D6 = 1'b1;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_D1 = 1'b1;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_D2 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_A1 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_A2 = CLBLM_L_X12Y106_SLICE_X16Y106_CO6;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_A3 = CLBLM_L_X12Y107_SLICE_X17Y107_CO5;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_A5 = CLBLM_R_X7Y107_SLICE_X9Y107_BQ;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_A6 = CLBLM_L_X12Y108_SLICE_X17Y108_CO5;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_D3 = 1'b1;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_D4 = 1'b1;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_C3 = CLBLM_R_X11Y116_SLICE_X14Y116_AQ;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_D5 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_B1 = CLBLM_L_X10Y118_SLICE_X13Y118_AQ;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_B2 = CLBLM_L_X12Y107_SLICE_X16Y107_BQ;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_B3 = CLBLM_L_X12Y107_SLICE_X17Y107_CO5;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_B4 = CLBLM_L_X12Y106_SLICE_X16Y106_DO6;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_B6 = CLBLM_L_X12Y108_SLICE_X17Y108_CO5;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_D6 = 1'b1;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_C5 = CLBLM_R_X11Y116_SLICE_X14Y116_DO6;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_C6 = CLBLM_L_X8Y116_SLICE_X11Y116_CO6;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_C1 = CLBLM_L_X12Y105_SLICE_X16Y105_CO5;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_C2 = CLBLM_L_X12Y107_SLICE_X16Y107_CQ;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_C4 = CLBLM_L_X8Y113_SLICE_X10Y113_CQ;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_C5 = CLBLM_L_X12Y105_SLICE_X16Y105_BO6;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_C6 = CLBLM_R_X11Y106_SLICE_X14Y106_CQ;
  assign RIOI3_X105Y129_ILOGIC_X1Y130_D = RIOB33_X105Y129_IOB_X1Y130_I;
  assign RIOI3_X105Y129_ILOGIC_X1Y129_D = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_D1 = CLBLM_L_X12Y107_SLICE_X16Y107_DQ;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_D2 = CLBLM_L_X12Y105_SLICE_X16Y105_CO5;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_D3 = CLBLM_L_X12Y105_SLICE_X16Y105_BO6;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_D4 = CLBLM_L_X12Y108_SLICE_X16Y108_CQ;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_D5 = CLBLM_L_X10Y110_SLICE_X13Y110_DQ;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_D6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOI3_SING_X0Y150_OLOGIC_X0Y150_D1 = LIOB33_X0Y63_IOB_X0Y63_I;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_A4 = CLBLM_R_X7Y118_SLICE_X8Y118_AQ;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_D1 = CLBLM_L_X10Y118_SLICE_X12Y118_AQ;
  assign RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y144_D = RIOB33_X105Y143_IOB_X1Y144_I;
  assign RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y143_D = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_A5 = CLBLM_R_X7Y117_SLICE_X8Y117_BQ;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_D2 = CLBLM_L_X10Y118_SLICE_X12Y118_BQ;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_A6 = CLBLM_R_X7Y118_SLICE_X8Y118_BQ;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_B2 = CLBLM_L_X8Y114_SLICE_X11Y114_BQ;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_B3 = CLBLM_L_X12Y113_SLICE_X17Y113_B5Q;
  assign CLBLM_R_X11Y116_SLICE_X14Y116_D5 = CLBLM_R_X7Y118_SLICE_X8Y118_CQ;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_B4 = CLBLM_L_X8Y115_SLICE_X10Y115_BQ;
  assign LIOI3_X0Y79_OLOGIC_X0Y80_D1 = CLBLL_L_X2Y106_SLICE_X0Y106_AO6;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_B3 = CLBLM_R_X7Y114_SLICE_X8Y114_BQ;
  assign LIOI3_SING_X0Y150_OLOGIC_X0Y150_T1 = 1'b1;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_B4 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_C1 = CLBLM_R_X5Y109_SLICE_X6Y109_DQ;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_B5 = CLBLM_R_X7Y117_SLICE_X8Y117_BQ;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_C2 = CLBLM_L_X10Y112_SLICE_X12Y112_BQ;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_B6 = CLBLM_R_X7Y118_SLICE_X8Y118_BQ;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_C3 = CLBLM_L_X8Y118_SLICE_X10Y118_BQ;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_C4 = CLBLM_L_X8Y114_SLICE_X10Y114_CQ;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_C6 = CLBLM_L_X8Y111_SLICE_X11Y111_DO5;
  assign LIOI3_X0Y79_OLOGIC_X0Y80_T1 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_A1 = CLBLM_R_X3Y114_SLICE_X2Y114_BQ;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_A3 = CLBLM_R_X3Y113_SLICE_X3Y113_AQ;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_A4 = CLBLL_L_X4Y113_SLICE_X4Y113_CO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_A5 = CLBLM_R_X3Y112_SLICE_X3Y112_AQ;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_A6 = CLBLL_L_X4Y111_SLICE_X5Y111_BO6;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_C4 = CLBLL_L_X4Y118_SLICE_X4Y118_BQ;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_B1 = CLBLL_L_X2Y112_SLICE_X0Y112_AO5;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_B2 = CLBLM_R_X5Y112_SLICE_X7Y112_BQ;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_B3 = CLBLM_R_X3Y116_SLICE_X3Y116_AO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_B4 = CLBLL_L_X2Y114_SLICE_X0Y114_AO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_B5 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_B6 = CLBLL_L_X2Y109_SLICE_X0Y109_AO5;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_C6 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_A4 = CLBLM_R_X11Y106_SLICE_X14Y106_DQ;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_C1 = CLBLM_R_X3Y115_SLICE_X3Y115_AO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_C2 = CLBLL_L_X2Y114_SLICE_X0Y114_AO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_C3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_C4 = CLBLM_R_X5Y109_SLICE_X7Y109_B5Q;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_C5 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_C6 = CLBLL_L_X2Y112_SLICE_X0Y112_AO6;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_A6 = CLBLM_R_X11Y106_SLICE_X14Y106_BQ;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_D1 = CLBLM_R_X3Y110_SLICE_X2Y110_AO5;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_D2 = CLBLL_L_X4Y113_SLICE_X4Y113_DO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_D3 = CLBLM_R_X5Y113_SLICE_X6Y113_DO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_D4 = CLBLM_R_X3Y113_SLICE_X3Y113_CO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_D5 = CLBLM_R_X5Y113_SLICE_X6Y113_CQ;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_D6 = CLBLM_R_X3Y113_SLICE_X3Y113_BO6;
  assign RIOI3_X105Y161_OLOGIC_X1Y161_D1 = CLBLM_L_X12Y114_SLICE_X16Y114_DO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_A1 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_A2 = CLBLL_L_X26Y136_SLICE_X38Y136_AO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_A3 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_A4 = CLBLL_L_X2Y112_SLICE_X0Y112_AO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_A5 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_A6 = CLBLL_L_X4Y111_SLICE_X4Y111_BQ;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_B1 = CLBLL_L_X2Y114_SLICE_X0Y114_AO5;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_B2 = CLBLL_L_X4Y114_SLICE_X4Y114_AQ;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_B3 = CLBLM_R_X3Y112_SLICE_X2Y112_AO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_B4 = CLBLL_L_X2Y110_SLICE_X0Y110_AO5;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_B5 = CLBLL_L_X2Y113_SLICE_X1Y113_BO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_B6 = CLBLM_R_X3Y114_SLICE_X2Y114_CO6;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_B3 = CLBLM_L_X12Y112_SLICE_X16Y112_CQ;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_B4 = CLBLM_R_X11Y105_SLICE_X15Y105_A5Q;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_C1 = CLBLM_R_X3Y113_SLICE_X3Y113_AQ;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_C2 = CLBLL_L_X2Y114_SLICE_X0Y114_AO5;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_C3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_C4 = CLBLL_L_X2Y112_SLICE_X1Y112_DO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_C5 = CLBLM_R_X5Y110_SLICE_X6Y110_DQ;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_C6 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_B6 = 1'b1;
  assign LIOB33_X0Y135_IOB_X0Y135_O = CLBLL_L_X4Y118_SLICE_X4Y118_AQ;
  assign LIOB33_X0Y135_IOB_X0Y136_O = CLBLL_L_X4Y117_SLICE_X4Y117_DQ;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_D1 = CLBLM_R_X3Y112_SLICE_X3Y112_AQ;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_D2 = CLBLL_L_X2Y114_SLICE_X0Y114_AO5;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_D3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_D4 = CLBLM_R_X3Y115_SLICE_X3Y115_AO5;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_D5 = LIOB33_X0Y63_IOB_X0Y63_I;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_D6 = CLBLL_L_X2Y112_SLICE_X0Y112_AO6;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_A1 = CLBLM_L_X12Y105_SLICE_X16Y105_BO6;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_A2 = CLBLM_R_X7Y109_SLICE_X8Y109_BQ;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_A3 = CLBLM_L_X12Y108_SLICE_X17Y108_AQ;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_A4 = CLBLM_L_X12Y105_SLICE_X16Y105_CO5;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_A5 = CLBLM_L_X12Y107_SLICE_X16Y107_CQ;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_B1 = CLBLM_L_X12Y108_SLICE_X16Y108_DQ;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_B3 = CLBLM_L_X12Y105_SLICE_X16Y105_BO6;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_B4 = CLBLM_L_X12Y105_SLICE_X16Y105_CO5;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_B5 = CLBLM_L_X12Y108_SLICE_X17Y108_BQ;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_B6 = CLBLM_L_X12Y109_SLICE_X17Y109_CQ;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_C6 = 1'b1;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_C1 = CLBLM_L_X12Y107_SLICE_X17Y107_BQ;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_C2 = CLBLM_R_X13Y113_SLICE_X18Y113_BQ;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_C3 = CLBLM_L_X12Y105_SLICE_X16Y105_AQ;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_C4 = CLBLM_R_X13Y108_SLICE_X18Y108_BO5;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_C5 = CLBLM_R_X13Y109_SLICE_X19Y109_BQ;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_C6 = 1'b1;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_D3 = CLBLM_L_X10Y110_SLICE_X12Y110_BQ;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_D4 = CLBLM_L_X8Y110_SLICE_X11Y110_A5Q;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_D1 = CLBLM_R_X11Y105_SLICE_X15Y105_BQ;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_D3 = CLBLM_L_X12Y105_SLICE_X16Y105_AQ;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_D2 = CLBLM_L_X12Y107_SLICE_X17Y107_BQ;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_D5 = CLBLM_R_X13Y109_SLICE_X19Y109_BQ;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_D6 = CLBLM_L_X12Y109_SLICE_X17Y109_BQ;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_D5 = 1'b1;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_D4 = CLBLM_R_X13Y113_SLICE_X18Y113_BQ;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_D6 = CLBLM_L_X10Y109_SLICE_X12Y109_BQ;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_A1 = CLBLM_L_X10Y115_SLICE_X12Y115_CQ;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_A2 = CLBLM_L_X12Y109_SLICE_X17Y109_BQ;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_A3 = CLBLM_R_X7Y115_SLICE_X8Y115_DQ;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_A6 = 1'b1;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_B1 = 1'b1;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_B2 = CLBLM_L_X12Y112_SLICE_X16Y112_AQ;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_B3 = CLBLM_L_X12Y108_SLICE_X17Y108_CO5;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_B5 = CLBLM_L_X12Y106_SLICE_X16Y106_BO6;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_B6 = CLBLM_L_X12Y107_SLICE_X17Y107_CO5;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_C2 = CLBLM_L_X12Y108_SLICE_X16Y108_CQ;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_C3 = CLBLM_L_X12Y105_SLICE_X16Y105_BO6;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_C4 = CLBLM_R_X11Y105_SLICE_X15Y105_CQ;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_C5 = CLBLM_L_X12Y105_SLICE_X16Y105_CO5;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_C6 = CLBLM_R_X7Y109_SLICE_X9Y109_BQ;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_D1 = CLBLM_R_X11Y105_SLICE_X15Y105_A5Q;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_D1 = CLBLM_L_X8Y116_SLICE_X10Y116_DQ;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_D2 = CLBLM_L_X12Y105_SLICE_X16Y105_BO6;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_D3 = CLBLM_L_X12Y108_SLICE_X16Y108_DQ;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_D4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_D5 = CLBLM_L_X12Y105_SLICE_X16Y105_CO5;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_D6 = CLBLM_R_X11Y108_SLICE_X14Y108_AQ;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_D2 = CLBLM_R_X11Y105_SLICE_X15Y105_AQ;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_A4 = CLBLM_R_X7Y108_SLICE_X9Y108_BO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_A6 = CLBLM_L_X10Y113_SLICE_X13Y113_AQ;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_C5 = CLBLM_R_X5Y115_SLICE_X7Y115_DO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_B2 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_B3 = CLBLM_R_X7Y106_SLICE_X9Y106_AQ;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_B4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_B5 = CLBLM_R_X7Y109_SLICE_X9Y109_CQ;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_B6 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_C5 = CLBLM_R_X3Y116_SLICE_X3Y116_AO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_C5 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_D4 = CLBLM_L_X8Y112_SLICE_X11Y112_BO6;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_C6 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_D5 = CLBLM_L_X8Y118_SLICE_X10Y118_BQ;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_D6 = CLBLM_R_X7Y115_SLICE_X8Y115_BQ;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_A1 = CLBLM_R_X3Y114_SLICE_X3Y114_DO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_A2 = CLBLM_R_X3Y115_SLICE_X3Y115_DO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_A3 = CLBLM_R_X3Y115_SLICE_X3Y115_CO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_A4 = CLBLM_R_X3Y114_SLICE_X3Y114_BO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_A5 = CLBLM_R_X3Y114_SLICE_X3Y114_CO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_A6 = CLBLL_L_X4Y114_SLICE_X4Y114_DO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_B1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_B2 = CLBLL_L_X2Y114_SLICE_X0Y114_AO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_B3 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_B4 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_B5 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_B6 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_C1 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_C2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_C3 = CLBLL_L_X2Y114_SLICE_X0Y114_AO5;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_C4 = CLBLL_L_X4Y115_SLICE_X5Y115_CQ;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_C5 = CLBLL_L_X2Y112_SLICE_X0Y112_AO5;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_C6 = CLBLL_L_X2Y112_SLICE_X0Y112_AO6;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_D1 = CLBLL_L_X2Y109_SLICE_X0Y109_AO5;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_D2 = CLBLM_R_X7Y106_SLICE_X9Y106_CQ;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_D3 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_D4 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_D5 = CLBLL_L_X2Y112_SLICE_X0Y112_AO5;
  assign CLBLM_R_X3Y114_SLICE_X3Y114_D6 = CLBLL_L_X2Y114_SLICE_X0Y114_AO6;
  assign LIOB33_X0Y137_IOB_X0Y137_O = CLBLL_L_X4Y117_SLICE_X4Y117_AQ;
  assign LIOB33_X0Y137_IOB_X0Y138_O = CLBLL_L_X4Y117_SLICE_X5Y117_AQ;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_D1 = LIOB33_X0Y53_IOB_X0Y54_I;
  assign LIOI3_X0Y151_OLOGIC_X0Y152_D1 = LIOB33_X0Y65_IOB_X0Y66_I;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_A1 = CLBLM_R_X3Y115_SLICE_X2Y115_AO5;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_A2 = CLBLM_R_X7Y106_SLICE_X9Y106_BQ;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_A3 = CLBLM_R_X3Y114_SLICE_X2Y114_AQ;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_A4 = CLBLL_L_X4Y113_SLICE_X4Y113_CO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_A6 = CLBLL_L_X4Y114_SLICE_X5Y114_BO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_D4 = CLBLM_R_X5Y115_SLICE_X7Y115_CO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_D5 = CLBLM_L_X10Y109_SLICE_X13Y109_BO5;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_B2 = CLBLL_L_X4Y111_SLICE_X5Y111_BO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_B3 = CLBLM_R_X3Y114_SLICE_X2Y114_AQ;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_B4 = CLBLL_L_X4Y113_SLICE_X4Y113_CO6;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_B5 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_B6 = CLBLM_R_X3Y114_SLICE_X2Y114_BQ;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_D6 = CLBLM_R_X7Y107_SLICE_X9Y107_AQ;
  assign LIOI3_X0Y151_OLOGIC_X0Y151_D1 = LIOB33_X0Y65_IOB_X0Y65_I;
  assign RIOI3_X105Y195_OLOGIC_X1Y196_T1 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_C1 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_C2 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_C3 = CLBLL_L_X4Y115_SLICE_X5Y115_A5Q;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_C4 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_C5 = CLBLL_L_X4Y110_SLICE_X5Y110_AQ;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_C6 = 1'b1;
  assign LIOI3_X0Y151_OLOGIC_X0Y151_T1 = 1'b1;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_X105Y195_OLOGIC_X1Y195_D1 = CLBLM_L_X12Y110_SLICE_X16Y110_AQ;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_D1 = CLBLM_R_X3Y114_SLICE_X2Y114_CO5;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_D2 = CLBLL_L_X4Y114_SLICE_X4Y114_CQ;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_D3 = LIOB33_X0Y65_IOB_X0Y65_I;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_D4 = CLBLL_L_X2Y112_SLICE_X0Y112_AO5;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_D5 = CLBLL_L_X2Y114_SLICE_X0Y114_AO5;
  assign CLBLM_R_X3Y114_SLICE_X2Y114_D6 = CLBLL_L_X2Y112_SLICE_X0Y112_AO6;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_A1 = CLBLM_L_X12Y105_SLICE_X16Y105_AQ;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_A2 = CLBLM_R_X13Y113_SLICE_X18Y113_BQ;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_A4 = CLBLM_L_X12Y107_SLICE_X17Y107_BQ;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_A5 = CLBLM_R_X13Y109_SLICE_X19Y109_BQ;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_A6 = CLBLM_L_X12Y109_SLICE_X16Y109_CQ;
  assign RIOI3_X105Y195_OLOGIC_X1Y195_T1 = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_T1 = 1'b1;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_B2 = CLBLM_R_X5Y107_SLICE_X7Y107_BQ;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_B3 = CLBLM_L_X12Y109_SLICE_X17Y109_AQ;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_B4 = 1'b1;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_B5 = CLBLM_L_X12Y108_SLICE_X17Y108_CO6;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_B6 = 1'b1;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_C2 = CLBLM_L_X10Y111_SLICE_X13Y111_BQ;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_C3 = 1'b1;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_C4 = CLBLM_R_X7Y115_SLICE_X8Y115_CQ;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_C6 = 1'b1;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_D1 = CLBLM_R_X37Y117_SLICE_X56Y117_AO6;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_D2 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_D3 = CLBLM_L_X12Y109_SLICE_X17Y109_DQ;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_D4 = CLBLM_R_X7Y109_SLICE_X8Y109_DO6;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_D5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_D6 = CLBLM_R_X11Y112_SLICE_X14Y112_BQ;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_T1 = 1'b1;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_A1 = CLBLM_R_X13Y110_SLICE_X18Y110_AQ;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_A2 = CLBLM_L_X12Y110_SLICE_X17Y110_BQ;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_A3 = CLBLM_L_X12Y109_SLICE_X16Y109_AQ;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_A4 = CLBLM_L_X12Y108_SLICE_X16Y108_AO5;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_A6 = CLBLM_L_X12Y110_SLICE_X16Y110_CO5;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_D1 = RIOB33_X105Y125_IOB_X1Y126_I;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_B1 = CLBLM_L_X12Y117_SLICE_X16Y117_AO6;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_B2 = CLBLM_L_X12Y109_SLICE_X16Y109_BQ;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_B3 = CLBLM_R_X11Y108_SLICE_X14Y108_BO6;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_B4 = CLBLM_R_X11Y109_SLICE_X15Y109_CO6;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_B6 = CLBLM_L_X12Y109_SLICE_X16Y109_DQ;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_T1 = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_D1 = CLBLL_L_X4Y117_SLICE_X4Y117_BQ;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_C1 = CLBLM_L_X8Y106_SLICE_X11Y106_A5Q;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_C2 = CLBLM_L_X12Y108_SLICE_X17Y108_CO6;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_C4 = CLBLM_L_X12Y112_SLICE_X16Y112_CQ;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_C5 = 1'b1;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_C6 = 1'b1;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_D1 = CLBLM_L_X12Y109_SLICE_X16Y109_BQ;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_D2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_D3 = CLBLM_L_X12Y112_SLICE_X17Y112_B5Q;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_D4 = CLBLM_L_X10Y105_SLICE_X12Y105_AQ;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_D5 = CLBLM_R_X13Y109_SLICE_X18Y109_AQ;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_D6 = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_T1 = 1'b1;
  assign LIOB33_X0Y173_IOB_X0Y174_O = CLBLM_L_X10Y148_SLICE_X12Y148_AO6;
  assign LIOB33_X0Y173_IOB_X0Y173_O = CLBLM_R_X7Y132_SLICE_X9Y132_AO5;
  assign RIOB33_X105Y155_IOB_X1Y156_O = RIOB33_X105Y103_IOB_X1Y104_I;
  assign RIOB33_X105Y155_IOB_X1Y155_O = RIOB33_X105Y103_IOB_X1Y103_I;
  assign RIOI3_X105Y133_ILOGIC_X1Y134_D = RIOB33_X105Y133_IOB_X1Y134_I;
  assign RIOI3_X105Y133_ILOGIC_X1Y133_D = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_A1 = 1'b1;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_A2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_A3 = 1'b1;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_A4 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_A5 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_A6 = 1'b1;
  assign LIOB33_X0Y139_IOB_X0Y140_O = CLBLL_L_X4Y116_SLICE_X4Y116_AQ;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_B1 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_B2 = CLBLM_R_X5Y112_SLICE_X6Y112_AQ;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_B3 = CLBLL_L_X2Y114_SLICE_X0Y114_AO5;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_B4 = CLBLL_L_X2Y107_SLICE_X1Y107_AO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_B5 = CLBLM_L_X8Y111_SLICE_X10Y111_A5Q;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_B6 = CLBLM_R_X3Y115_SLICE_X3Y115_AO5;
  assign LIOB33_X0Y139_IOB_X0Y139_O = CLBLL_L_X4Y118_SLICE_X4Y118_BQ;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_C1 = LIOB33_X0Y57_IOB_X0Y57_I;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_C2 = CLBLM_R_X7Y114_SLICE_X8Y114_AQ;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_C3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_C4 = CLBLL_L_X2Y114_SLICE_X0Y114_AO5;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_C5 = CLBLM_R_X3Y115_SLICE_X3Y115_AO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_C6 = CLBLL_L_X2Y107_SLICE_X1Y107_AO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_D1 = CLBLM_R_X3Y115_SLICE_X3Y115_AO6;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_D2 = CLBLL_L_X4Y116_SLICE_X5Y116_A5Q;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_D3 = CLBLL_L_X2Y114_SLICE_X0Y114_AO5;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_D4 = CLBLM_R_X3Y115_SLICE_X3Y115_AO5;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_D5 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y115_SLICE_X3Y115_D6 = CLBLL_L_X4Y114_SLICE_X5Y114_AQ;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_A2 = CLBLM_R_X3Y114_SLICE_X2Y114_BQ;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_A3 = CLBLM_R_X3Y114_SLICE_X2Y114_AQ;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_A4 = CLBLM_R_X3Y113_SLICE_X3Y113_AQ;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_A5 = CLBLL_L_X4Y114_SLICE_X5Y114_AQ;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_A6 = 1'b1;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_B1 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_B2 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_B3 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_B4 = CLBLL_L_X2Y114_SLICE_X0Y114_AO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_B5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_B6 = CLBLL_L_X4Y111_SLICE_X4Y111_CQ;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_C1 = CLBLL_L_X4Y115_SLICE_X4Y115_AO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_C2 = CLBLL_L_X2Y114_SLICE_X0Y114_BO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_C3 = CLBLM_R_X3Y115_SLICE_X3Y115_BO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_C4 = CLBLM_R_X3Y113_SLICE_X2Y113_CO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_C5 = CLBLM_R_X3Y116_SLICE_X2Y116_AO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_C6 = CLBLM_R_X3Y115_SLICE_X2Y115_BO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_D1 = CLBLM_R_X3Y114_SLICE_X2Y114_AQ;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_D2 = CLBLM_R_X3Y115_SLICE_X3Y115_AO6;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_D3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_D4 = CLBLL_L_X2Y114_SLICE_X0Y114_AO5;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_D5 = CLBLL_L_X4Y115_SLICE_X5Y115_AQ;
  assign CLBLM_R_X3Y115_SLICE_X2Y115_D6 = CLBLL_L_X2Y107_SLICE_X1Y107_AO6;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_A1 = CLBLM_R_X5Y115_SLICE_X7Y115_CO6;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_A3 = CLBLM_L_X12Y110_SLICE_X17Y110_AQ;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_A4 = CLBLM_R_X11Y110_SLICE_X14Y110_CQ;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_A5 = 1'b1;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_A6 = CLBLM_L_X8Y115_SLICE_X10Y115_CQ;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_B2 = CLBLM_L_X12Y110_SLICE_X17Y110_BQ;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_B3 = CLBLM_L_X12Y110_SLICE_X16Y110_CO5;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_B5 = CLBLM_R_X7Y115_SLICE_X8Y115_DQ;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_B6 = CLBLM_L_X12Y108_SLICE_X16Y108_AQ;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_C2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_C3 = CLBLM_L_X12Y110_SLICE_X16Y110_BO5;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_C4 = CLBLM_L_X8Y115_SLICE_X10Y115_CQ;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_C5 = 1'b1;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_C6 = CLBLM_L_X12Y108_SLICE_X16Y108_BQ;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_D1 = CLBLM_L_X8Y109_SLICE_X11Y109_CQ;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_D2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_D3 = CLBLM_L_X12Y110_SLICE_X17Y110_DQ;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_D4 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_D5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_D6 = CLBLM_L_X10Y109_SLICE_X13Y109_CO6;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_A1 = CLBLM_L_X8Y109_SLICE_X10Y109_DQ;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_A3 = CLBLM_L_X8Y112_SLICE_X10Y112_A5Q;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_A4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_A5 = CLBLM_L_X12Y110_SLICE_X17Y110_AQ;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_A6 = 1'b1;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_AX = CLBLM_L_X12Y107_SLICE_X16Y107_CQ;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_B1 = CLBLL_L_X4Y117_SLICE_X4Y117_CQ;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_B2 = CLBLM_R_X11Y112_SLICE_X14Y112_BQ;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_B3 = CLBLM_L_X10Y110_SLICE_X13Y110_CQ;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_B4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_B6 = 1'b1;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_C1 = CLBLM_L_X12Y109_SLICE_X16Y109_AQ;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_C2 = CLBLM_L_X12Y110_SLICE_X17Y110_BQ;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_C3 = CLBLM_L_X10Y106_SLICE_X12Y106_BO6;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_C4 = CLBLM_R_X11Y110_SLICE_X15Y110_AQ;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_C5 = CLBLM_R_X13Y110_SLICE_X19Y110_AQ;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_C6 = 1'b1;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_CE = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_D1 = CLBLL_L_X4Y117_SLICE_X5Y117_AQ;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_D1 = CLBLM_L_X12Y109_SLICE_X16Y109_AQ;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_D2 = CLBLM_L_X12Y110_SLICE_X17Y110_BQ;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_D3 = CLBLM_L_X10Y106_SLICE_X12Y106_BO6;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_D4 = CLBLM_R_X11Y110_SLICE_X15Y110_AQ;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_D5 = CLBLM_R_X13Y110_SLICE_X19Y110_AQ;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_D6 = 1'b1;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_SR = CLBLM_L_X12Y117_SLICE_X16Y117_AO6;
  assign CLBLL_L_X26Y136_SLICE_X38Y136_A1 = 1'b1;
  assign CLBLL_L_X26Y136_SLICE_X38Y136_A2 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLL_L_X26Y136_SLICE_X38Y136_A3 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X26Y136_SLICE_X38Y136_A4 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X26Y136_SLICE_X38Y136_A5 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLL_L_X26Y136_SLICE_X38Y136_A6 = 1'b1;
  assign CLBLL_L_X26Y136_SLICE_X38Y136_B1 = 1'b1;
  assign CLBLL_L_X26Y136_SLICE_X38Y136_B2 = 1'b1;
  assign CLBLL_L_X26Y136_SLICE_X38Y136_B3 = 1'b1;
  assign CLBLL_L_X26Y136_SLICE_X38Y136_B4 = 1'b1;
  assign CLBLL_L_X26Y136_SLICE_X38Y136_B5 = 1'b1;
  assign CLBLL_L_X26Y136_SLICE_X38Y136_B6 = 1'b1;
  assign CLBLL_L_X26Y136_SLICE_X38Y136_C1 = 1'b1;
  assign CLBLL_L_X26Y136_SLICE_X38Y136_C2 = 1'b1;
  assign CLBLL_L_X26Y136_SLICE_X38Y136_C3 = 1'b1;
  assign CLBLL_L_X26Y136_SLICE_X38Y136_C4 = 1'b1;
  assign CLBLL_L_X26Y136_SLICE_X38Y136_C5 = 1'b1;
  assign CLBLL_L_X26Y136_SLICE_X38Y136_C6 = 1'b1;
  assign LIOB33_X0Y141_IOB_X0Y141_O = CLBLL_L_X4Y117_SLICE_X4Y117_BQ;
  assign LIOB33_X0Y141_IOB_X0Y142_O = LIOB33_X0Y53_IOB_X0Y54_I;
  assign CLBLL_L_X26Y136_SLICE_X38Y136_D1 = 1'b1;
  assign CLBLL_L_X26Y136_SLICE_X38Y136_D2 = 1'b1;
  assign CLBLL_L_X26Y136_SLICE_X38Y136_D3 = 1'b1;
  assign CLBLL_L_X26Y136_SLICE_X38Y136_D4 = 1'b1;
  assign CLBLL_L_X26Y136_SLICE_X38Y136_D5 = 1'b1;
  assign CLBLL_L_X26Y136_SLICE_X38Y136_D6 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_A1 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_A2 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_A3 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_A4 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_A5 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_A6 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_B1 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_B2 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_B3 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_B4 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_B5 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_B6 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_C1 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_C2 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_C3 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_C4 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_C5 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_C6 = 1'b1;
  assign LIOI3_SING_X0Y100_OLOGIC_X0Y100_D1 = CLBLL_L_X2Y106_SLICE_X0Y106_BO6;
  assign CLBLL_L_X26Y136_SLICE_X39Y136_A1 = 1'b1;
  assign CLBLL_L_X26Y136_SLICE_X39Y136_A2 = 1'b1;
  assign CLBLL_L_X26Y136_SLICE_X39Y136_A3 = 1'b1;
  assign CLBLL_L_X26Y136_SLICE_X39Y136_A4 = 1'b1;
  assign CLBLL_L_X26Y136_SLICE_X39Y136_A5 = 1'b1;
  assign CLBLL_L_X26Y136_SLICE_X39Y136_A6 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_D1 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_D2 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_D3 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_D5 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X3Y116_D6 = 1'b1;
  assign CLBLL_L_X26Y136_SLICE_X39Y136_B1 = 1'b1;
  assign CLBLL_L_X26Y136_SLICE_X39Y136_B2 = 1'b1;
  assign CLBLL_L_X26Y136_SLICE_X39Y136_B3 = 1'b1;
  assign CLBLL_L_X26Y136_SLICE_X39Y136_B4 = 1'b1;
  assign CLBLL_L_X26Y136_SLICE_X39Y136_B5 = 1'b1;
  assign CLBLL_L_X26Y136_SLICE_X39Y136_B6 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_A1 = LIOB33_X0Y61_IOB_X0Y61_I;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_A2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X26Y136_SLICE_X39Y136_C1 = 1'b1;
  assign CLBLL_L_X26Y136_SLICE_X39Y136_C2 = 1'b1;
  assign CLBLL_L_X26Y136_SLICE_X39Y136_C3 = 1'b1;
  assign CLBLL_L_X26Y136_SLICE_X39Y136_C4 = 1'b1;
  assign CLBLL_L_X26Y136_SLICE_X39Y136_C5 = 1'b1;
  assign CLBLL_L_X26Y136_SLICE_X39Y136_C6 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_A3 = CLBLL_L_X2Y114_SLICE_X0Y114_AO5;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_A4 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_A5 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_A6 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_B4 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_B1 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_B2 = 1'b1;
  assign CLBLL_L_X26Y136_SLICE_X39Y136_D1 = 1'b1;
  assign CLBLL_L_X26Y136_SLICE_X39Y136_D2 = 1'b1;
  assign CLBLL_L_X26Y136_SLICE_X39Y136_D3 = 1'b1;
  assign CLBLL_L_X26Y136_SLICE_X39Y136_D4 = 1'b1;
  assign CLBLL_L_X26Y136_SLICE_X39Y136_D5 = 1'b1;
  assign CLBLL_L_X26Y136_SLICE_X39Y136_D6 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_B6 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_C1 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_C2 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_C3 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_C4 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_C5 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_C6 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_D1 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_D2 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_D3 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_D4 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_D5 = 1'b1;
  assign CLBLM_R_X3Y116_SLICE_X2Y116_D6 = 1'b1;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_A1 = 1'b1;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_A2 = 1'b1;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_A3 = 1'b1;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_A4 = 1'b1;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_A5 = 1'b1;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_A6 = 1'b1;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_B1 = 1'b1;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_B2 = 1'b1;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_B3 = 1'b1;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_B4 = 1'b1;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_B5 = 1'b1;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_B6 = 1'b1;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_C1 = 1'b1;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_C2 = 1'b1;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_C3 = 1'b1;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_C4 = 1'b1;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_C5 = 1'b1;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_C6 = 1'b1;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_D1 = 1'b1;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_D2 = 1'b1;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_D3 = 1'b1;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_D4 = 1'b1;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_D5 = 1'b1;
  assign CLBLM_L_X12Y111_SLICE_X17Y111_D6 = 1'b1;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_A1 = 1'b1;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_A2 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_A3 = CLBLM_L_X12Y111_SLICE_X16Y111_AQ;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_A4 = CLBLM_L_X10Y113_SLICE_X12Y113_BQ;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_A6 = CLBLM_L_X8Y119_SLICE_X10Y119_AQ;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_B1 = CLBLM_R_X7Y115_SLICE_X9Y115_DO6;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_B2 = CLBLM_L_X12Y111_SLICE_X16Y111_BQ;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_B4 = CLBLM_L_X12Y108_SLICE_X16Y108_CQ;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_B5 = CLBLM_L_X12Y112_SLICE_X16Y112_DQ;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_B6 = 1'b1;
  assign LIOI3_X0Y153_OLOGIC_X0Y154_D1 = LIOB33_X0Y67_IOB_X0Y68_I;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_C2 = CLBLM_L_X8Y111_SLICE_X11Y111_CQ;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_C3 = CLBLM_R_X11Y107_SLICE_X15Y107_CQ;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_C5 = 1'b1;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_C6 = 1'b1;
  assign LIOI3_X0Y153_OLOGIC_X0Y154_T1 = 1'b1;
  assign RIOI3_X105Y197_OLOGIC_X1Y198_D1 = CLBLL_L_X26Y136_SLICE_X38Y136_AO5;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_D1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_D2 = CLBLM_L_X12Y111_SLICE_X16Y111_CQ;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_D3 = CLBLM_R_X11Y108_SLICE_X15Y108_AQ;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_D4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_D5 = 1'b1;
  assign CLBLM_L_X12Y111_SLICE_X16Y111_D6 = 1'b1;
  assign LIOI3_X0Y153_OLOGIC_X0Y153_D1 = LIOB33_X0Y67_IOB_X0Y67_I;
  assign RIOI3_X105Y197_OLOGIC_X1Y198_T1 = 1'b1;
  assign CLBLM_R_X13Y117_SLICE_X18Y117_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign LIOI3_X0Y153_OLOGIC_X0Y153_T1 = 1'b1;
  assign RIOI3_X105Y197_OLOGIC_X1Y197_D1 = CLBLL_L_X26Y136_SLICE_X38Y136_AO5;
  assign RIOI3_X105Y197_OLOGIC_X1Y197_T1 = 1'b1;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_C3 = CLBLM_L_X10Y118_SLICE_X13Y118_CO6;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_C5 = 1'b1;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_C6 = CLBLM_L_X10Y116_SLICE_X12Y116_DO5;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_D1 = CLBLM_R_X103Y170_SLICE_X163Y170_AO6;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_D1 = CLBLM_R_X103Y169_SLICE_X163Y169_AO6;
  assign LIOB33_X0Y151_IOB_X0Y152_O = LIOB33_X0Y65_IOB_X0Y66_I;
  assign LIOB33_X0Y143_IOB_X0Y143_O = LIOB33_X0Y55_IOB_X0Y55_I;
  assign LIOB33_X0Y151_IOB_X0Y151_O = LIOB33_X0Y65_IOB_X0Y65_I;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_T1 = 1'b1;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_D5 = CLBLM_L_X10Y118_SLICE_X13Y118_CO6;
  assign CLBLM_R_X11Y117_SLICE_X15Y117_D6 = CLBLM_R_X11Y110_SLICE_X15Y110_A5Q;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_T1 = 1'b1;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_D1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign RIOI3_X105Y135_ILOGIC_X1Y136_D = RIOB33_X105Y135_IOB_X1Y136_I;
  assign RIOI3_X105Y135_ILOGIC_X1Y135_D = RIOB33_X105Y135_IOB_X1Y135_I;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_T1 = 1'b1;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_A1 = CLBLM_L_X12Y112_SLICE_X17Y112_B5Q;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_A2 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_A3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_A5 = CLBLM_R_X13Y113_SLICE_X18Y113_DO6;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_A6 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_AX = CLBLM_L_X12Y110_SLICE_X16Y110_AO6;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_B1 = CLBLM_R_X5Y112_SLICE_X7Y112_CQ;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_B2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_B3 = 1'b1;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_B4 = CLBLM_L_X12Y109_SLICE_X16Y109_CQ;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_B5 = CLBLM_L_X12Y112_SLICE_X17Y112_CO5;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_B5 = CLBLM_R_X7Y118_SLICE_X9Y118_CO5;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_BX = CLBLM_L_X12Y112_SLICE_X17Y112_CO6;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_B6 = CLBLM_R_X11Y117_SLICE_X15Y117_CQ;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_C1 = CLBLM_R_X13Y110_SLICE_X18Y110_BQ;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_C2 = CLBLM_R_X11Y111_SLICE_X15Y111_BQ;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_C3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_C5 = CLBLM_L_X12Y110_SLICE_X17Y110_DQ;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_C6 = 1'b1;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_D1 = CLBLM_R_X11Y111_SLICE_X15Y111_BQ;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_D2 = 1'b1;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_D3 = CLBLM_R_X7Y115_SLICE_X8Y115_CQ;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_D4 = CLBLM_L_X12Y111_SLICE_X16Y111_CQ;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_D5 = CLBLM_L_X12Y109_SLICE_X17Y109_CQ;
  assign CLBLM_L_X12Y112_SLICE_X17Y112_D6 = 1'b1;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_A1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_A3 = CLBLM_L_X12Y112_SLICE_X16Y112_AQ;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_A5 = CLBLM_R_X11Y113_SLICE_X15Y113_AQ;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_A6 = CLBLM_R_X11Y113_SLICE_X14Y113_CQ;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_AX = CLBLM_R_X11Y112_SLICE_X14Y112_AO6;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_B1 = CLBLM_R_X11Y116_SLICE_X14Y116_A5Q;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_B2 = CLBLM_L_X10Y112_SLICE_X12Y112_CQ;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_B4 = CLBLM_L_X12Y108_SLICE_X17Y108_CO6;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_B5 = CLBLM_L_X12Y109_SLICE_X17Y109_BQ;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_B6 = 1'b1;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_C4 = CLBLM_R_X11Y117_SLICE_X15Y117_CQ;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_C5 = CLBLM_R_X7Y118_SLICE_X9Y118_CO5;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_C1 = CLBLM_L_X12Y112_SLICE_X16Y112_BQ;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_C2 = 1'b1;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_C3 = 1'b1;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_C5 = CLBLM_R_X11Y114_SLICE_X14Y114_CQ;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_C6 = CLBLM_L_X12Y108_SLICE_X17Y108_CO6;
  assign CLBLM_R_X11Y117_SLICE_X14Y117_C6 = CLBLM_L_X10Y117_SLICE_X12Y117_DO6;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_B6 = 1'b1;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_D1 = 1'b1;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_D2 = CLBLM_L_X12Y113_SLICE_X16Y113_CQ;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_D3 = CLBLM_L_X12Y112_SLICE_X16Y112_DQ;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_D4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_D5 = CLBLM_R_X7Y115_SLICE_X9Y115_DO6;
  assign CLBLM_L_X12Y112_SLICE_X16Y112_D6 = CLBLM_L_X8Y105_SLICE_X11Y105_BQ;
  assign LIOB33_X0Y145_IOB_X0Y146_O = LIOB33_X0Y59_IOB_X0Y59_I;
  assign LIOB33_X0Y145_IOB_X0Y145_O = LIOB33_X0Y57_IOB_X0Y58_I;
  assign CLBLM_R_X13Y106_SLICE_X19Y106_A1 = 1'b1;
  assign CLBLM_R_X13Y106_SLICE_X19Y106_A2 = 1'b1;
  assign CLBLM_R_X13Y106_SLICE_X19Y106_A3 = 1'b1;
  assign CLBLM_R_X13Y106_SLICE_X19Y106_A4 = 1'b1;
  assign CLBLM_R_X13Y106_SLICE_X19Y106_A5 = 1'b1;
  assign CLBLM_R_X13Y106_SLICE_X19Y106_A6 = 1'b1;
  assign CLBLM_R_X13Y106_SLICE_X19Y106_B1 = 1'b1;
  assign CLBLM_R_X13Y106_SLICE_X19Y106_B2 = 1'b1;
  assign CLBLM_R_X13Y106_SLICE_X19Y106_B3 = 1'b1;
  assign CLBLM_R_X13Y106_SLICE_X19Y106_B4 = 1'b1;
  assign CLBLM_R_X13Y106_SLICE_X19Y106_B5 = 1'b1;
  assign CLBLM_R_X13Y106_SLICE_X19Y106_B6 = 1'b1;
  assign CLBLM_R_X13Y106_SLICE_X19Y106_C1 = 1'b1;
  assign CLBLM_R_X13Y106_SLICE_X19Y106_C2 = 1'b1;
  assign CLBLM_R_X13Y106_SLICE_X19Y106_C3 = 1'b1;
  assign CLBLM_R_X13Y106_SLICE_X19Y106_C4 = 1'b1;
  assign CLBLM_R_X13Y106_SLICE_X19Y106_C5 = 1'b1;
  assign CLBLM_R_X13Y106_SLICE_X19Y106_C6 = 1'b1;
  assign RIOI3_X105Y171_OLOGIC_X1Y172_D1 = CLBLM_R_X103Y173_SLICE_X163Y173_AO6;
  assign CLBLM_R_X13Y106_SLICE_X19Y106_D1 = 1'b1;
  assign CLBLM_R_X13Y106_SLICE_X19Y106_D2 = 1'b1;
  assign CLBLM_R_X13Y106_SLICE_X19Y106_D3 = 1'b1;
  assign CLBLM_R_X13Y106_SLICE_X19Y106_D4 = 1'b1;
  assign CLBLM_R_X13Y106_SLICE_X19Y106_D5 = 1'b1;
  assign CLBLM_R_X13Y106_SLICE_X19Y106_D6 = 1'b1;
  assign CLBLM_R_X13Y106_SLICE_X18Y106_A1 = CLBLM_R_X13Y107_SLICE_X19Y107_BQ;
  assign CLBLM_R_X13Y106_SLICE_X18Y106_A2 = CLBLM_L_X12Y105_SLICE_X17Y105_AO5;
  assign CLBLM_R_X13Y106_SLICE_X18Y106_A3 = CLBLM_L_X12Y107_SLICE_X16Y107_DQ;
  assign CLBLM_R_X13Y106_SLICE_X18Y106_A4 = CLBLM_R_X13Y106_SLICE_X18Y106_BO6;
  assign CLBLM_R_X13Y106_SLICE_X18Y106_A5 = CLBLM_L_X12Y105_SLICE_X17Y105_CO6;
  assign CLBLM_R_X13Y106_SLICE_X18Y106_A6 = CLBLM_R_X13Y106_SLICE_X18Y106_CO6;
  assign CLBLM_R_X13Y106_SLICE_X18Y106_B1 = CLBLM_R_X13Y108_SLICE_X19Y108_BQ;
  assign CLBLM_R_X13Y106_SLICE_X18Y106_B2 = CLBLM_R_X13Y109_SLICE_X19Y109_BQ;
  assign CLBLM_R_X13Y106_SLICE_X18Y106_B3 = CLBLM_R_X13Y113_SLICE_X18Y113_BQ;
  assign CLBLM_R_X13Y106_SLICE_X18Y106_B4 = CLBLM_L_X12Y108_SLICE_X16Y108_BQ;
  assign CLBLM_R_X13Y106_SLICE_X18Y106_B5 = CLBLM_L_X12Y107_SLICE_X17Y107_BQ;
  assign CLBLM_R_X13Y106_SLICE_X18Y106_B6 = CLBLM_L_X12Y107_SLICE_X16Y107_BQ;
  assign CLBLM_R_X13Y106_SLICE_X18Y106_C1 = CLBLM_R_X13Y109_SLICE_X19Y109_BQ;
  assign CLBLM_R_X13Y106_SLICE_X18Y106_C2 = CLBLM_L_X12Y107_SLICE_X17Y107_BQ;
  assign CLBLM_R_X13Y106_SLICE_X18Y106_C3 = CLBLM_R_X13Y113_SLICE_X18Y113_BQ;
  assign CLBLM_R_X13Y106_SLICE_X18Y106_C4 = CLBLM_L_X12Y107_SLICE_X16Y107_BQ;
  assign CLBLM_R_X13Y106_SLICE_X18Y106_C5 = CLBLM_R_X13Y108_SLICE_X19Y108_BQ;
  assign CLBLM_R_X13Y106_SLICE_X18Y106_C6 = CLBLM_L_X12Y108_SLICE_X16Y108_BQ;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_A1 = CLBLL_L_X4Y118_SLICE_X4Y118_A5Q;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_A2 = CLBLL_L_X4Y117_SLICE_X4Y117_AQ;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_A3 = CLBLL_L_X4Y118_SLICE_X4Y118_AQ;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_A4 = CLBLL_L_X4Y116_SLICE_X5Y116_AQ;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_A5 = CLBLL_L_X4Y117_SLICE_X4Y117_DQ;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_A6 = CLBLL_L_X4Y117_SLICE_X5Y117_AQ;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_B1 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_B2 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_B3 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_B4 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_B5 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_B6 = 1'b1;
  assign CLBLM_R_X13Y106_SLICE_X18Y106_D1 = CLBLM_R_X13Y107_SLICE_X19Y107_AQ;
  assign CLBLM_R_X13Y106_SLICE_X18Y106_D2 = CLBLM_L_X12Y107_SLICE_X16Y107_AQ;
  assign CLBLM_R_X13Y106_SLICE_X18Y106_D3 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_C1 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_C2 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_C3 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_C4 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_C5 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_C6 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_D1 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_D2 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_D3 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_D4 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_D5 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_D6 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_A1 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_A2 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_A3 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_A4 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_A5 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_A6 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_B1 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_B2 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_B3 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_B4 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_B5 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_B6 = 1'b1;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_B1 = 1'b1;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_B2 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_C1 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_C2 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_C3 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_C4 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_C5 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_C6 = 1'b1;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_B4 = CLBLM_R_X11Y109_SLICE_X15Y109_BO6;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_B5 = CLBLM_L_X10Y105_SLICE_X12Y105_BQ;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_D1 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_D2 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_D3 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_D4 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_D5 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_D6 = 1'b1;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_A2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_A3 = CLBLM_L_X12Y109_SLICE_X17Y109_AQ;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_A4 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_A5 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_A6 = CLBLM_R_X13Y113_SLICE_X18Y113_DO6;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_B1 = CLBLM_L_X12Y113_SLICE_X17Y113_B5Q;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_B2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_B3 = CLBLM_L_X12Y112_SLICE_X17Y112_AQ;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_B5 = CLBLM_R_X11Y115_SLICE_X15Y115_B5Q;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_B6 = 1'b1;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_C1 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_C2 = CLBLM_L_X12Y113_SLICE_X17Y113_CQ;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_C3 = CLBLM_R_X13Y113_SLICE_X19Y113_AQ;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_C4 = CLBLM_R_X7Y110_SLICE_X9Y110_CO6;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_C6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X37Y117_SLICE_X57Y117_A1 = 1'b1;
  assign CLBLM_R_X37Y117_SLICE_X57Y117_A2 = 1'b1;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X37Y117_SLICE_X57Y117_A3 = 1'b1;
  assign CLBLM_R_X37Y117_SLICE_X57Y117_A4 = 1'b1;
  assign CLBLM_R_X37Y117_SLICE_X57Y117_A5 = 1'b1;
  assign CLBLM_R_X37Y117_SLICE_X57Y117_A6 = 1'b1;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_C4 = CLBLM_L_X10Y107_SLICE_X12Y107_DO6;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_D1 = CLBLM_R_X11Y109_SLICE_X15Y109_DO6;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_D2 = 1'b1;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_D3 = CLBLM_L_X12Y114_SLICE_X17Y114_CO6;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_D4 = CLBLM_L_X12Y113_SLICE_X16Y113_DO6;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_D5 = CLBLM_R_X13Y113_SLICE_X18Y113_CQ;
  assign CLBLM_L_X12Y113_SLICE_X17Y113_D6 = CLBLM_L_X12Y114_SLICE_X17Y114_BQ;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_C5 = CLBLM_L_X8Y108_SLICE_X11Y108_AQ;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_C6 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLM_R_X37Y117_SLICE_X57Y117_B1 = 1'b1;
  assign CLBLM_R_X37Y117_SLICE_X57Y117_B2 = 1'b1;
  assign CLBLM_R_X37Y117_SLICE_X57Y117_B3 = 1'b1;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_A2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_A3 = CLBLM_L_X12Y113_SLICE_X16Y113_AQ;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_A4 = CLBLM_L_X12Y113_SLICE_X16Y113_CQ;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_A5 = CLBLM_L_X8Y116_SLICE_X10Y116_AQ;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_A6 = CLBLM_R_X7Y112_SLICE_X9Y112_CO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_D5 = 1'b1;
  assign CLBLM_R_X37Y117_SLICE_X57Y117_C1 = 1'b1;
  assign CLBLM_R_X37Y117_SLICE_X57Y117_C2 = 1'b1;
  assign CLBLM_R_X37Y117_SLICE_X57Y117_C4 = 1'b1;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_B1 = CLBLM_R_X11Y114_SLICE_X14Y114_DQ;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_B2 = CLBLM_L_X12Y113_SLICE_X16Y113_BQ;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_B3 = 1'b1;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_B4 = CLBLM_L_X12Y112_SLICE_X16Y112_DQ;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_B6 = CLBLM_R_X5Y115_SLICE_X7Y115_CO6;
  assign CLBLM_R_X37Y117_SLICE_X57Y117_D1 = 1'b1;
  assign CLBLM_R_X37Y117_SLICE_X57Y117_D2 = 1'b1;
  assign CLBLM_R_X37Y117_SLICE_X57Y117_D3 = 1'b1;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_C2 = CLBLM_L_X12Y113_SLICE_X16Y113_CQ;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_C3 = CLBLM_L_X12Y113_SLICE_X16Y113_BQ;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_C4 = 1'b1;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_C5 = CLBLM_R_X7Y115_SLICE_X9Y115_DO6;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_C6 = CLBLM_R_X11Y113_SLICE_X15Y113_AQ;
  assign CLBLM_R_X37Y117_SLICE_X56Y117_A1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X37Y117_SLICE_X56Y117_A2 = 1'b1;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X37Y117_SLICE_X56Y117_A3 = RIOB33_X105Y119_IOB_X1Y119_I;
  assign CLBLM_R_X37Y117_SLICE_X56Y117_A4 = 1'b1;
  assign CLBLM_R_X37Y117_SLICE_X56Y117_A5 = 1'b1;
  assign CLBLM_R_X37Y117_SLICE_X56Y117_A6 = CLBLM_L_X8Y113_SLICE_X10Y113_DQ;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_D1 = CLBLM_L_X8Y115_SLICE_X10Y115_AQ;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_D2 = CLBLM_L_X12Y113_SLICE_X16Y113_CQ;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_D3 = CLBLM_L_X8Y115_SLICE_X11Y115_BQ;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_D4 = 1'b1;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_D5 = 1'b1;
  assign CLBLM_L_X12Y113_SLICE_X16Y113_D6 = CLBLM_L_X10Y115_SLICE_X13Y115_BQ;
  assign CLBLM_R_X37Y117_SLICE_X56Y117_B1 = 1'b1;
endmodule
